-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 626;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (46,0,76,0,11,0,14,0,219,0,77,0,65,0,38,0,133,0,11,0,248,0,188,0,0,0,125,0,140,0,237,0,90,0,242,0,152,0,220,0,18,0,117,0,173,0,0,0,15,0,0,0,252,0,100,0,74,0,71,0,0,0,211,0,148,0,124,0,233,0,149,0,0,0,114,0,190,0,74,0,136,0,233,0,46,0,123,0,27,0,33,0,216,0,0,0,50,0,133,0,65,0,243,0,5,0,207,0,30,0,53,0,218,0,48,0,152,0,70,0,191,0,73,0,180,0,0,0,0,0,190,0,150,0,26,0,241,0,150,0,0,0,181,0,90,0,0,0,89,0,150,0,211,0,179,0,0,0,95,0,131,0,0,0,26,0,181,0,2,0,0,0,78,0,154,0,63,0,196,0,0,0,0,0,105,0,110,0,46,0,0,0,57,0,0,0,133,0,17,0,223,0,2,0,226,0,95,0,187,0,223,0,212,0,168,0,193,0,95,0,0,0,215,0,17,0,141,0,0,0,0,0,96,0,70,0,210,0,213,0,11,0,101,0,172,0,232,0,219,0,0,0,110,0,243,0,232,0,79,0,0,0,126,0,0,0,220,0,147,0,105,0,176,0,37,0,86,0,0,0,4,0,0,0,0,0,44,0,89,0,13,0,111,0,90,0,144,0,0,0,237,0,222,0,0,0,117,0,171,0,151,0,177,0,140,0,113,0,93,0,72,0,225,0,181,0,0,0,246,0,23,0,28,0,3,0,196,0,0,0,227,0,115,0,115,0,86,0,59,0,222,0,85,0,36,0,176,0,250,0,249,0,0,0,180,0,0,0,243,0,237,0,0,0,231,0,204,0,169,0,0,0,0,0,86,0,72,0,0,0,82,0,166,0,11,0,90,0,0,0,43,0,119,0,168,0,232,0,141,0,93,0,104,0,193,0,168,0,12,0,119,0,76,0,48,0,181,0,176,0,33,0,122,0,13,0,225,0,185,0,239,0,151,0,95,0,0,0,30,0,237,0,152,0,28,0,151,0,4,0,80,0,225,0,244,0,0,0,129,0,238,0,135,0,253,0,0,0,88,0,20,0,193,0,41,0,0,0,43,0,113,0,249,0,70,0,186,0,197,0,163,0,102,0,0,0,203,0,253,0,227,0,27,0,203,0,87,0,0,0,125,0,245,0,70,0,56,0,252,0,126,0,138,0,0,0,130,0,33,0,104,0,65,0,55,0,158,0,60,0,158,0,135,0,188,0,0,0,177,0,109,0,186,0,102,0,237,0,68,0,244,0,131,0,0,0,166,0,178,0,0,0,78,0,182,0,0,0,33,0,0,0,192,0,164,0,247,0,25,0,146,0,0,0,222,0,165,0,134,0,238,0,0,0,11,0,248,0,193,0,183,0,0,0,130,0,189,0,45,0,0,0,0,0,77,0,12,0,243,0,88,0,251,0,133,0,170,0,143,0,160,0,21,0,101,0,0,0,94,0,107,0,36,0,176,0,85,0,145,0,0,0,165,0,217,0,21,0,0,0,0,0,91,0,70,0,54,0,172,0,220,0,137,0,0,0,224,0,224,0,246,0,132,0,37,0,0,0,245,0,217,0,0,0,13,0,0,0,34,0,82,0,0,0,154,0,14,0,247,0,114,0,43,0,27,0,13,0,25,0,74,0,177,0,85,0,0,0,38,0,15,0,141,0,136,0,161,0,47,0,62,0,0,0,163,0,80,0,244,0,147,0,63,0,160,0,4,0,221,0,0,0,28,0,237,0,172,0,0,0,166,0,204,0,170,0,113,0,0,0,180,0,202,0,154,0,52,0,0,0,192,0,171,0,0,0,22,0,50,0,115,0,244,0,28,0,93,0,224,0,159,0,172,0,42,0,65,0,21,0,81,0,114,0,175,0,0,0,0,0,164,0,80,0,249,0,254,0,229,0,229,0,0,0,86,0,0,0,68,0,8,0,80,0,213,0,247,0,15,0,235,0,0,0,50,0,246,0,212,0,131,0,242,0,157,0,182,0,255,0,154,0,147,0,84,0,2,0,126,0,0,0,0,0,0,0,34,0,40,0,24,0,194,0,87,0,0,0,118,0,0,0,101,0,120,0,45,0,0,0,238,0,177,0,154,0,70,0,97,0,62,0,156,0,65,0,171,0,243,0,24,0,149,0,117,0,133,0,111,0,14,0,85,0,0,0,47,0,0,0,118,0,24,0,118,0,83,0,18,0,157,0,0,0,44,0,16,0,79,0,23,0,202,0,238,0,120,0,0,0,46,0,0,0,210,0,179,0,101,0,130,0,157,0,97,0,213,0,22,0,15,0,223,0,220,0,0,0,64,0,38,0,193,0,252,0,62,0,0,0,0,0,155,0,162,0,198,0,17,0,252,0,217,0,149,0,228,0,180,0,75,0,0,0,158,0,249,0,139,0,78,0,211,0,82,0,175,0,59,0,92,0,121,0,4,0,12,0,20,0,54,0,31,0,217,0,153,0,118,0,0,0,11,0,0,0,1,0,0,0,52,0,121,0,0,0,164,0,35,0,0,0,0,0,12,0,0,0,157,0,158,0,156,0,40,0,152,0,100,0,0,0,0,0,177,0,222,0,0,0,63,0,48,0,0,0,0,0,133,0,230,0,0,0,129,0,36,0,44,0,170,0,220,0,168,0,101,0,217,0,148,0,233,0,22,0,131,0,0,0,174,0,0,0,198,0,0,0,0,0,221,0,234,0,62,0,219,0,0,0,137,0,29,0,77,0,93,0,203,0,0,0,228,0,116,0,5,0,65,0,162,0,116,0,222,0,113,0,140,0,173,0);
signal scenario_full  : scenario_type := (46,31,76,31,11,31,14,31,219,31,77,31,65,31,38,31,133,31,11,31,248,31,188,31,188,30,125,31,140,31,237,31,90,31,242,31,152,31,220,31,18,31,117,31,173,31,173,30,15,31,15,30,252,31,100,31,74,31,71,31,71,30,211,31,148,31,124,31,233,31,149,31,149,30,114,31,190,31,74,31,136,31,233,31,46,31,123,31,27,31,33,31,216,31,216,30,50,31,133,31,65,31,243,31,5,31,207,31,30,31,53,31,218,31,48,31,152,31,70,31,191,31,73,31,180,31,180,30,180,29,190,31,150,31,26,31,241,31,150,31,150,30,181,31,90,31,90,30,89,31,150,31,211,31,179,31,179,30,95,31,131,31,131,30,26,31,181,31,2,31,2,30,78,31,154,31,63,31,196,31,196,30,196,29,105,31,110,31,46,31,46,30,57,31,57,30,133,31,17,31,223,31,2,31,226,31,95,31,187,31,223,31,212,31,168,31,193,31,95,31,95,30,215,31,17,31,141,31,141,30,141,29,96,31,70,31,210,31,213,31,11,31,101,31,172,31,232,31,219,31,219,30,110,31,243,31,232,31,79,31,79,30,126,31,126,30,220,31,147,31,105,31,176,31,37,31,86,31,86,30,4,31,4,30,4,29,44,31,89,31,13,31,111,31,90,31,144,31,144,30,237,31,222,31,222,30,117,31,171,31,151,31,177,31,140,31,113,31,93,31,72,31,225,31,181,31,181,30,246,31,23,31,28,31,3,31,196,31,196,30,227,31,115,31,115,31,86,31,59,31,222,31,85,31,36,31,176,31,250,31,249,31,249,30,180,31,180,30,243,31,237,31,237,30,231,31,204,31,169,31,169,30,169,29,86,31,72,31,72,30,82,31,166,31,11,31,90,31,90,30,43,31,119,31,168,31,232,31,141,31,93,31,104,31,193,31,168,31,12,31,119,31,76,31,48,31,181,31,176,31,33,31,122,31,13,31,225,31,185,31,239,31,151,31,95,31,95,30,30,31,237,31,152,31,28,31,151,31,4,31,80,31,225,31,244,31,244,30,129,31,238,31,135,31,253,31,253,30,88,31,20,31,193,31,41,31,41,30,43,31,113,31,249,31,70,31,186,31,197,31,163,31,102,31,102,30,203,31,253,31,227,31,27,31,203,31,87,31,87,30,125,31,245,31,70,31,56,31,252,31,126,31,138,31,138,30,130,31,33,31,104,31,65,31,55,31,158,31,60,31,158,31,135,31,188,31,188,30,177,31,109,31,186,31,102,31,237,31,68,31,244,31,131,31,131,30,166,31,178,31,178,30,78,31,182,31,182,30,33,31,33,30,192,31,164,31,247,31,25,31,146,31,146,30,222,31,165,31,134,31,238,31,238,30,11,31,248,31,193,31,183,31,183,30,130,31,189,31,45,31,45,30,45,29,77,31,12,31,243,31,88,31,251,31,133,31,170,31,143,31,160,31,21,31,101,31,101,30,94,31,107,31,36,31,176,31,85,31,145,31,145,30,165,31,217,31,21,31,21,30,21,29,91,31,70,31,54,31,172,31,220,31,137,31,137,30,224,31,224,31,246,31,132,31,37,31,37,30,245,31,217,31,217,30,13,31,13,30,34,31,82,31,82,30,154,31,14,31,247,31,114,31,43,31,27,31,13,31,25,31,74,31,177,31,85,31,85,30,38,31,15,31,141,31,136,31,161,31,47,31,62,31,62,30,163,31,80,31,244,31,147,31,63,31,160,31,4,31,221,31,221,30,28,31,237,31,172,31,172,30,166,31,204,31,170,31,113,31,113,30,180,31,202,31,154,31,52,31,52,30,192,31,171,31,171,30,22,31,50,31,115,31,244,31,28,31,93,31,224,31,159,31,172,31,42,31,65,31,21,31,81,31,114,31,175,31,175,30,175,29,164,31,80,31,249,31,254,31,229,31,229,31,229,30,86,31,86,30,68,31,8,31,80,31,213,31,247,31,15,31,235,31,235,30,50,31,246,31,212,31,131,31,242,31,157,31,182,31,255,31,154,31,147,31,84,31,2,31,126,31,126,30,126,29,126,28,34,31,40,31,24,31,194,31,87,31,87,30,118,31,118,30,101,31,120,31,45,31,45,30,238,31,177,31,154,31,70,31,97,31,62,31,156,31,65,31,171,31,243,31,24,31,149,31,117,31,133,31,111,31,14,31,85,31,85,30,47,31,47,30,118,31,24,31,118,31,83,31,18,31,157,31,157,30,44,31,16,31,79,31,23,31,202,31,238,31,120,31,120,30,46,31,46,30,210,31,179,31,101,31,130,31,157,31,97,31,213,31,22,31,15,31,223,31,220,31,220,30,64,31,38,31,193,31,252,31,62,31,62,30,62,29,155,31,162,31,198,31,17,31,252,31,217,31,149,31,228,31,180,31,75,31,75,30,158,31,249,31,139,31,78,31,211,31,82,31,175,31,59,31,92,31,121,31,4,31,12,31,20,31,54,31,31,31,217,31,153,31,118,31,118,30,11,31,11,30,1,31,1,30,52,31,121,31,121,30,164,31,35,31,35,30,35,29,12,31,12,30,157,31,158,31,156,31,40,31,152,31,100,31,100,30,100,29,177,31,222,31,222,30,63,31,48,31,48,30,48,29,133,31,230,31,230,30,129,31,36,31,44,31,170,31,220,31,168,31,101,31,217,31,148,31,233,31,22,31,131,31,131,30,174,31,174,30,198,31,198,30,198,29,221,31,234,31,62,31,219,31,219,30,137,31,29,31,77,31,93,31,203,31,203,30,228,31,116,31,5,31,65,31,162,31,116,31,222,31,113,31,140,31,173,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
