-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 212;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,135,0,109,0,0,0,33,0,57,0,223,0,4,0,235,0,0,0,233,0,132,0,226,0,12,0,133,0,51,0,87,0,46,0,112,0,74,0,0,0,123,0,159,0,36,0,0,0,236,0,74,0,150,0,105,0,0,0,0,0,29,0,0,0,0,0,153,0,81,0,143,0,0,0,0,0,122,0,0,0,144,0,172,0,85,0,177,0,7,0,143,0,241,0,0,0,28,0,0,0,171,0,34,0,102,0,18,0,219,0,249,0,196,0,58,0,142,0,124,0,145,0,181,0,88,0,215,0,160,0,237,0,0,0,0,0,247,0,3,0,218,0,77,0,233,0,248,0,143,0,254,0,210,0,0,0,35,0,0,0,73,0,98,0,203,0,0,0,205,0,105,0,71,0,51,0,159,0,64,0,0,0,198,0,0,0,0,0,219,0,0,0,0,0,119,0,255,0,53,0,210,0,198,0,17,0,93,0,235,0,94,0,0,0,159,0,149,0,176,0,188,0,0,0,210,0,58,0,232,0,16,0,0,0,22,0,90,0,109,0,196,0,210,0,249,0,145,0,181,0,19,0,0,0,248,0,55,0,212,0,207,0,197,0,172,0,90,0,132,0,157,0,44,0,76,0,20,0,0,0,19,0,126,0,36,0,42,0,131,0,0,0,207,0,0,0,254,0,0,0,0,0,0,0,18,0,82,0,237,0,104,0,160,0,126,0,191,0,192,0,76,0,0,0,0,0,0,0,135,0,0,0,147,0,0,0,143,0,105,0,103,0,203,0,143,0,211,0,150,0,211,0,167,0,181,0,155,0,173,0,241,0,142,0,100,0,107,0,240,0,201,0,0,0,181,0,0,0,74,0,17,0,0,0,164,0,0,0,0,0,145,0,211,0,32,0,116,0,44,0,202,0,0,0,205,0,44,0,112,0,212,0,248,0,111,0,0,0,63,0,64,0);
signal scenario_full  : scenario_type := (136,31,135,31,109,31,109,30,33,31,57,31,223,31,4,31,235,31,235,30,233,31,132,31,226,31,12,31,133,31,51,31,87,31,46,31,112,31,74,31,74,30,123,31,159,31,36,31,36,30,236,31,74,31,150,31,105,31,105,30,105,29,29,31,29,30,29,29,153,31,81,31,143,31,143,30,143,29,122,31,122,30,144,31,172,31,85,31,177,31,7,31,143,31,241,31,241,30,28,31,28,30,171,31,34,31,102,31,18,31,219,31,249,31,196,31,58,31,142,31,124,31,145,31,181,31,88,31,215,31,160,31,237,31,237,30,237,29,247,31,3,31,218,31,77,31,233,31,248,31,143,31,254,31,210,31,210,30,35,31,35,30,73,31,98,31,203,31,203,30,205,31,105,31,71,31,51,31,159,31,64,31,64,30,198,31,198,30,198,29,219,31,219,30,219,29,119,31,255,31,53,31,210,31,198,31,17,31,93,31,235,31,94,31,94,30,159,31,149,31,176,31,188,31,188,30,210,31,58,31,232,31,16,31,16,30,22,31,90,31,109,31,196,31,210,31,249,31,145,31,181,31,19,31,19,30,248,31,55,31,212,31,207,31,197,31,172,31,90,31,132,31,157,31,44,31,76,31,20,31,20,30,19,31,126,31,36,31,42,31,131,31,131,30,207,31,207,30,254,31,254,30,254,29,254,28,18,31,82,31,237,31,104,31,160,31,126,31,191,31,192,31,76,31,76,30,76,29,76,28,135,31,135,30,147,31,147,30,143,31,105,31,103,31,203,31,143,31,211,31,150,31,211,31,167,31,181,31,155,31,173,31,241,31,142,31,100,31,107,31,240,31,201,31,201,30,181,31,181,30,74,31,17,31,17,30,164,31,164,30,164,29,145,31,211,31,32,31,116,31,44,31,202,31,202,30,205,31,44,31,112,31,212,31,248,31,111,31,111,30,63,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
