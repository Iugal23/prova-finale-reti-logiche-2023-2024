-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 657;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,247,0,0,0,129,0,248,0,89,0,0,0,165,0,0,0,170,0,21,0,0,0,90,0,34,0,196,0,0,0,179,0,0,0,176,0,87,0,139,0,61,0,0,0,14,0,194,0,135,0,86,0,46,0,201,0,252,0,75,0,0,0,131,0,0,0,49,0,228,0,224,0,188,0,0,0,254,0,222,0,69,0,97,0,56,0,198,0,104,0,77,0,0,0,115,0,0,0,140,0,213,0,0,0,49,0,151,0,28,0,153,0,3,0,91,0,14,0,203,0,211,0,53,0,247,0,0,0,0,0,83,0,1,0,3,0,47,0,189,0,0,0,15,0,48,0,0,0,226,0,0,0,0,0,174,0,151,0,105,0,0,0,112,0,0,0,0,0,182,0,0,0,88,0,0,0,203,0,239,0,0,0,0,0,180,0,0,0,133,0,16,0,0,0,82,0,212,0,169,0,40,0,0,0,228,0,0,0,101,0,236,0,99,0,163,0,51,0,148,0,195,0,127,0,247,0,0,0,182,0,224,0,0,0,228,0,179,0,58,0,30,0,0,0,248,0,73,0,29,0,41,0,188,0,147,0,107,0,239,0,247,0,0,0,154,0,174,0,124,0,246,0,179,0,75,0,229,0,65,0,0,0,11,0,0,0,0,0,157,0,203,0,52,0,59,0,82,0,8,0,47,0,180,0,12,0,236,0,69,0,33,0,166,0,172,0,0,0,51,0,83,0,95,0,150,0,253,0,13,0,235,0,104,0,210,0,168,0,0,0,0,0,0,0,0,0,191,0,0,0,231,0,247,0,132,0,115,0,0,0,94,0,0,0,252,0,174,0,148,0,0,0,64,0,0,0,5,0,40,0,205,0,138,0,190,0,111,0,0,0,0,0,0,0,0,0,126,0,242,0,204,0,233,0,0,0,108,0,45,0,215,0,196,0,179,0,192,0,86,0,0,0,117,0,0,0,6,0,128,0,0,0,242,0,0,0,110,0,183,0,210,0,0,0,134,0,172,0,197,0,227,0,134,0,128,0,183,0,191,0,126,0,147,0,0,0,232,0,222,0,245,0,33,0,68,0,0,0,0,0,167,0,0,0,94,0,37,0,0,0,0,0,0,0,0,0,18,0,0,0,102,0,145,0,0,0,43,0,128,0,253,0,184,0,38,0,181,0,89,0,162,0,0,0,169,0,0,0,187,0,139,0,4,0,65,0,152,0,50,0,187,0,160,0,42,0,38,0,182,0,0,0,246,0,48,0,147,0,0,0,125,0,78,0,137,0,18,0,38,0,10,0,206,0,182,0,0,0,204,0,0,0,0,0,167,0,244,0,143,0,0,0,84,0,175,0,146,0,216,0,0,0,191,0,0,0,177,0,131,0,61,0,0,0,100,0,158,0,255,0,0,0,120,0,218,0,0,0,63,0,0,0,4,0,0,0,90,0,0,0,168,0,175,0,161,0,26,0,51,0,151,0,5,0,104,0,0,0,105,0,0,0,42,0,70,0,125,0,236,0,0,0,53,0,99,0,0,0,182,0,224,0,255,0,32,0,0,0,30,0,120,0,234,0,103,0,190,0,101,0,0,0,40,0,229,0,0,0,147,0,206,0,197,0,184,0,0,0,94,0,0,0,70,0,0,0,208,0,112,0,71,0,80,0,208,0,31,0,4,0,252,0,8,0,47,0,5,0,124,0,59,0,164,0,61,0,110,0,0,0,167,0,239,0,60,0,157,0,73,0,0,0,194,0,0,0,10,0,150,0,5,0,70,0,152,0,248,0,192,0,2,0,148,0,150,0,238,0,116,0,148,0,70,0,221,0,0,0,61,0,211,0,207,0,114,0,0,0,206,0,85,0,0,0,111,0,0,0,190,0,100,0,0,0,84,0,178,0,16,0,214,0,65,0,200,0,73,0,0,0,148,0,83,0,0,0,9,0,102,0,0,0,188,0,160,0,69,0,0,0,220,0,215,0,170,0,141,0,110,0,22,0,40,0,133,0,89,0,169,0,68,0,155,0,41,0,0,0,172,0,246,0,134,0,143,0,0,0,243,0,200,0,0,0,18,0,37,0,0,0,0,0,95,0,137,0,141,0,191,0,82,0,123,0,29,0,38,0,0,0,74,0,254,0,38,0,232,0,158,0,44,0,63,0,177,0,34,0,0,0,64,0,135,0,95,0,212,0,223,0,0,0,223,0,0,0,180,0,120,0,182,0,171,0,12,0,41,0,0,0,236,0,67,0,242,0,147,0,226,0,184,0,0,0,0,0,99,0,215,0,224,0,13,0,49,0,0,0,0,0,171,0,219,0,104,0,50,0,217,0,0,0,73,0,3,0,26,0,141,0,220,0,114,0,230,0,28,0,62,0,28,0,98,0,234,0,0,0,104,0,218,0,52,0,39,0,77,0,238,0,132,0,212,0,179,0,184,0,77,0,167,0,189,0,243,0,0,0,1,0,129,0,128,0,15,0,0,0,0,0,67,0,206,0,0,0,117,0,101,0,60,0,6,0,1,0,0,0,162,0,0,0,203,0,177,0,148,0,32,0,89,0,0,0,219,0,121,0,139,0,48,0,82,0,82,0,23,0,98,0,0,0,226,0,14,0,131,0,255,0,0,0,191,0,211,0,232,0,159,0,177,0,67,0,112,0,19,0,250,0,0,0,0,0,0,0,54,0,90,0,0,0,0,0,0,0,191,0,146,0,189,0,103,0,10,0,0,0,43,0,87,0,184,0,56,0,0,0,10,0,13,0,0,0,131,0,44,0,162,0,0,0,112,0,0,0,129,0,23,0,236,0,44,0,213,0,43,0,145,0,0,0,67,0,158,0,179,0,253,0,124,0,236,0,153,0,0,0,207,0,205,0,205,0,220,0,194,0,0,0,0,0,0,0,20,0,125,0,202,0,0,0,108,0,10,0,89,0,0,0,26,0,48,0,179,0,228,0,0,0,108,0);
signal scenario_full  : scenario_type := (0,0,247,31,247,30,129,31,248,31,89,31,89,30,165,31,165,30,170,31,21,31,21,30,90,31,34,31,196,31,196,30,179,31,179,30,176,31,87,31,139,31,61,31,61,30,14,31,194,31,135,31,86,31,46,31,201,31,252,31,75,31,75,30,131,31,131,30,49,31,228,31,224,31,188,31,188,30,254,31,222,31,69,31,97,31,56,31,198,31,104,31,77,31,77,30,115,31,115,30,140,31,213,31,213,30,49,31,151,31,28,31,153,31,3,31,91,31,14,31,203,31,211,31,53,31,247,31,247,30,247,29,83,31,1,31,3,31,47,31,189,31,189,30,15,31,48,31,48,30,226,31,226,30,226,29,174,31,151,31,105,31,105,30,112,31,112,30,112,29,182,31,182,30,88,31,88,30,203,31,239,31,239,30,239,29,180,31,180,30,133,31,16,31,16,30,82,31,212,31,169,31,40,31,40,30,228,31,228,30,101,31,236,31,99,31,163,31,51,31,148,31,195,31,127,31,247,31,247,30,182,31,224,31,224,30,228,31,179,31,58,31,30,31,30,30,248,31,73,31,29,31,41,31,188,31,147,31,107,31,239,31,247,31,247,30,154,31,174,31,124,31,246,31,179,31,75,31,229,31,65,31,65,30,11,31,11,30,11,29,157,31,203,31,52,31,59,31,82,31,8,31,47,31,180,31,12,31,236,31,69,31,33,31,166,31,172,31,172,30,51,31,83,31,95,31,150,31,253,31,13,31,235,31,104,31,210,31,168,31,168,30,168,29,168,28,168,27,191,31,191,30,231,31,247,31,132,31,115,31,115,30,94,31,94,30,252,31,174,31,148,31,148,30,64,31,64,30,5,31,40,31,205,31,138,31,190,31,111,31,111,30,111,29,111,28,111,27,126,31,242,31,204,31,233,31,233,30,108,31,45,31,215,31,196,31,179,31,192,31,86,31,86,30,117,31,117,30,6,31,128,31,128,30,242,31,242,30,110,31,183,31,210,31,210,30,134,31,172,31,197,31,227,31,134,31,128,31,183,31,191,31,126,31,147,31,147,30,232,31,222,31,245,31,33,31,68,31,68,30,68,29,167,31,167,30,94,31,37,31,37,30,37,29,37,28,37,27,18,31,18,30,102,31,145,31,145,30,43,31,128,31,253,31,184,31,38,31,181,31,89,31,162,31,162,30,169,31,169,30,187,31,139,31,4,31,65,31,152,31,50,31,187,31,160,31,42,31,38,31,182,31,182,30,246,31,48,31,147,31,147,30,125,31,78,31,137,31,18,31,38,31,10,31,206,31,182,31,182,30,204,31,204,30,204,29,167,31,244,31,143,31,143,30,84,31,175,31,146,31,216,31,216,30,191,31,191,30,177,31,131,31,61,31,61,30,100,31,158,31,255,31,255,30,120,31,218,31,218,30,63,31,63,30,4,31,4,30,90,31,90,30,168,31,175,31,161,31,26,31,51,31,151,31,5,31,104,31,104,30,105,31,105,30,42,31,70,31,125,31,236,31,236,30,53,31,99,31,99,30,182,31,224,31,255,31,32,31,32,30,30,31,120,31,234,31,103,31,190,31,101,31,101,30,40,31,229,31,229,30,147,31,206,31,197,31,184,31,184,30,94,31,94,30,70,31,70,30,208,31,112,31,71,31,80,31,208,31,31,31,4,31,252,31,8,31,47,31,5,31,124,31,59,31,164,31,61,31,110,31,110,30,167,31,239,31,60,31,157,31,73,31,73,30,194,31,194,30,10,31,150,31,5,31,70,31,152,31,248,31,192,31,2,31,148,31,150,31,238,31,116,31,148,31,70,31,221,31,221,30,61,31,211,31,207,31,114,31,114,30,206,31,85,31,85,30,111,31,111,30,190,31,100,31,100,30,84,31,178,31,16,31,214,31,65,31,200,31,73,31,73,30,148,31,83,31,83,30,9,31,102,31,102,30,188,31,160,31,69,31,69,30,220,31,215,31,170,31,141,31,110,31,22,31,40,31,133,31,89,31,169,31,68,31,155,31,41,31,41,30,172,31,246,31,134,31,143,31,143,30,243,31,200,31,200,30,18,31,37,31,37,30,37,29,95,31,137,31,141,31,191,31,82,31,123,31,29,31,38,31,38,30,74,31,254,31,38,31,232,31,158,31,44,31,63,31,177,31,34,31,34,30,64,31,135,31,95,31,212,31,223,31,223,30,223,31,223,30,180,31,120,31,182,31,171,31,12,31,41,31,41,30,236,31,67,31,242,31,147,31,226,31,184,31,184,30,184,29,99,31,215,31,224,31,13,31,49,31,49,30,49,29,171,31,219,31,104,31,50,31,217,31,217,30,73,31,3,31,26,31,141,31,220,31,114,31,230,31,28,31,62,31,28,31,98,31,234,31,234,30,104,31,218,31,52,31,39,31,77,31,238,31,132,31,212,31,179,31,184,31,77,31,167,31,189,31,243,31,243,30,1,31,129,31,128,31,15,31,15,30,15,29,67,31,206,31,206,30,117,31,101,31,60,31,6,31,1,31,1,30,162,31,162,30,203,31,177,31,148,31,32,31,89,31,89,30,219,31,121,31,139,31,48,31,82,31,82,31,23,31,98,31,98,30,226,31,14,31,131,31,255,31,255,30,191,31,211,31,232,31,159,31,177,31,67,31,112,31,19,31,250,31,250,30,250,29,250,28,54,31,90,31,90,30,90,29,90,28,191,31,146,31,189,31,103,31,10,31,10,30,43,31,87,31,184,31,56,31,56,30,10,31,13,31,13,30,131,31,44,31,162,31,162,30,112,31,112,30,129,31,23,31,236,31,44,31,213,31,43,31,145,31,145,30,67,31,158,31,179,31,253,31,124,31,236,31,153,31,153,30,207,31,205,31,205,31,220,31,194,31,194,30,194,29,194,28,20,31,125,31,202,31,202,30,108,31,10,31,89,31,89,30,26,31,48,31,179,31,228,31,228,30,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
