-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 741;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (194,0,87,0,249,0,45,0,245,0,207,0,99,0,0,0,91,0,174,0,23,0,119,0,85,0,8,0,211,0,0,0,0,0,46,0,0,0,39,0,48,0,59,0,0,0,35,0,131,0,92,0,0,0,0,0,151,0,193,0,21,0,99,0,199,0,190,0,68,0,189,0,75,0,70,0,130,0,169,0,201,0,162,0,214,0,226,0,69,0,183,0,0,0,168,0,110,0,27,0,135,0,102,0,247,0,5,0,202,0,30,0,0,0,154,0,94,0,101,0,0,0,249,0,0,0,0,0,6,0,0,0,179,0,0,0,39,0,255,0,62,0,148,0,24,0,0,0,87,0,0,0,131,0,177,0,0,0,174,0,0,0,192,0,208,0,0,0,73,0,152,0,177,0,0,0,210,0,237,0,26,0,43,0,88,0,48,0,230,0,181,0,27,0,253,0,0,0,0,0,27,0,46,0,0,0,52,0,21,0,122,0,0,0,0,0,176,0,0,0,255,0,0,0,245,0,143,0,0,0,217,0,229,0,103,0,208,0,0,0,137,0,132,0,217,0,53,0,0,0,1,0,232,0,127,0,242,0,158,0,0,0,191,0,16,0,183,0,244,0,39,0,58,0,0,0,227,0,184,0,0,0,123,0,99,0,12,0,110,0,0,0,168,0,0,0,75,0,113,0,18,0,70,0,0,0,166,0,33,0,88,0,71,0,150,0,176,0,5,0,234,0,166,0,147,0,219,0,19,0,234,0,229,0,33,0,154,0,80,0,87,0,131,0,116,0,64,0,228,0,233,0,64,0,165,0,167,0,62,0,0,0,191,0,244,0,180,0,0,0,163,0,52,0,65,0,233,0,0,0,189,0,215,0,79,0,11,0,5,0,88,0,0,0,221,0,82,0,228,0,198,0,127,0,1,0,170,0,12,0,170,0,216,0,73,0,131,0,232,0,214,0,102,0,245,0,237,0,200,0,64,0,223,0,81,0,0,0,184,0,120,0,0,0,0,0,23,0,232,0,254,0,141,0,34,0,0,0,243,0,13,0,0,0,149,0,127,0,150,0,0,0,0,0,22,0,89,0,114,0,152,0,0,0,0,0,54,0,0,0,169,0,0,0,110,0,0,0,241,0,199,0,0,0,0,0,30,0,225,0,172,0,253,0,102,0,0,0,53,0,194,0,0,0,63,0,0,0,2,0,208,0,196,0,0,0,115,0,204,0,123,0,244,0,0,0,124,0,0,0,164,0,196,0,0,0,227,0,138,0,132,0,147,0,0,0,0,0,237,0,153,0,0,0,0,0,0,0,143,0,219,0,15,0,121,0,157,0,174,0,136,0,230,0,30,0,246,0,138,0,0,0,18,0,112,0,107,0,7,0,189,0,31,0,98,0,95,0,232,0,0,0,236,0,89,0,9,0,242,0,81,0,72,0,122,0,85,0,16,0,3,0,247,0,88,0,249,0,202,0,253,0,69,0,74,0,163,0,24,0,102,0,0,0,0,0,242,0,98,0,129,0,181,0,0,0,9,0,104,0,0,0,117,0,60,0,122,0,133,0,28,0,19,0,207,0,251,0,193,0,104,0,113,0,87,0,52,0,10,0,24,0,118,0,0,0,128,0,35,0,255,0,0,0,79,0,42,0,225,0,0,0,115,0,102,0,176,0,118,0,0,0,254,0,209,0,183,0,29,0,95,0,0,0,0,0,62,0,212,0,11,0,0,0,106,0,238,0,0,0,177,0,85,0,212,0,0,0,0,0,0,0,196,0,93,0,191,0,173,0,0,0,0,0,97,0,63,0,224,0,227,0,36,0,220,0,0,0,150,0,90,0,249,0,30,0,172,0,193,0,132,0,76,0,71,0,209,0,179,0,231,0,21,0,129,0,240,0,222,0,73,0,116,0,71,0,55,0,193,0,1,0,179,0,118,0,201,0,0,0,0,0,84,0,184,0,90,0,0,0,76,0,103,0,127,0,0,0,243,0,107,0,127,0,114,0,153,0,43,0,206,0,162,0,0,0,13,0,43,0,66,0,25,0,171,0,117,0,21,0,192,0,204,0,62,0,169,0,0,0,0,0,10,0,0,0,75,0,0,0,171,0,0,0,164,0,167,0,70,0,85,0,163,0,71,0,117,0,0,0,141,0,120,0,241,0,61,0,181,0,250,0,127,0,0,0,134,0,28,0,25,0,32,0,137,0,142,0,48,0,0,0,37,0,160,0,0,0,0,0,220,0,0,0,0,0,135,0,254,0,195,0,149,0,127,0,105,0,254,0,146,0,33,0,192,0,150,0,230,0,0,0,194,0,0,0,40,0,61,0,136,0,165,0,0,0,23,0,127,0,202,0,62,0,135,0,118,0,75,0,139,0,0,0,231,0,215,0,67,0,153,0,145,0,102,0,185,0,109,0,101,0,8,0,201,0,67,0,176,0,0,0,140,0,0,0,221,0,137,0,215,0,0,0,166,0,170,0,0,0,54,0,55,0,16,0,26,0,88,0,0,0,145,0,0,0,84,0,75,0,57,0,0,0,245,0,31,0,233,0,24,0,50,0,0,0,0,0,0,0,93,0,249,0,171,0,177,0,0,0,91,0,128,0,161,0,240,0,11,0,0,0,200,0,35,0,53,0,151,0,145,0,3,0,32,0,76,0,230,0,242,0,227,0,61,0,53,0,117,0,169,0,128,0,89,0,0,0,136,0,0,0,238,0,0,0,92,0,78,0,155,0,0,0,255,0,226,0,0,0,133,0,79,0,25,0,131,0,190,0,169,0,255,0,129,0,58,0,20,0,216,0,0,0,0,0,0,0,251,0,0,0,225,0,6,0,56,0,67,0,52,0,83,0,20,0,101,0,0,0,0,0,133,0,142,0,86,0,244,0,0,0,196,0,0,0,133,0,137,0,107,0,145,0,43,0,0,0,71,0,109,0,73,0,125,0,136,0,0,0,110,0,226,0,0,0,226,0,0,0,2,0,18,0,197,0,44,0,218,0,221,0,116,0,0,0,253,0,24,0,51,0,231,0,0,0,118,0,0,0,0,0,176,0,0,0,165,0,212,0,169,0,164,0,108,0,93,0,229,0,120,0,210,0,143,0,0,0,199,0,33,0,41,0,204,0,0,0,0,0,0,0,232,0,10,0,169,0,164,0,42,0,11,0,205,0,143,0,239,0,93,0,63,0,107,0,2,0,0,0,194,0,101,0,220,0,169,0,184,0,11,0,175,0,192,0,0,0,3,0,238,0,77,0,211,0,0,0,58,0,198,0,159,0,103,0,0,0,0,0,190,0,182,0,30,0,6,0,0,0,174,0,0,0,197,0,195,0,123,0,252,0);
signal scenario_full  : scenario_type := (194,31,87,31,249,31,45,31,245,31,207,31,99,31,99,30,91,31,174,31,23,31,119,31,85,31,8,31,211,31,211,30,211,29,46,31,46,30,39,31,48,31,59,31,59,30,35,31,131,31,92,31,92,30,92,29,151,31,193,31,21,31,99,31,199,31,190,31,68,31,189,31,75,31,70,31,130,31,169,31,201,31,162,31,214,31,226,31,69,31,183,31,183,30,168,31,110,31,27,31,135,31,102,31,247,31,5,31,202,31,30,31,30,30,154,31,94,31,101,31,101,30,249,31,249,30,249,29,6,31,6,30,179,31,179,30,39,31,255,31,62,31,148,31,24,31,24,30,87,31,87,30,131,31,177,31,177,30,174,31,174,30,192,31,208,31,208,30,73,31,152,31,177,31,177,30,210,31,237,31,26,31,43,31,88,31,48,31,230,31,181,31,27,31,253,31,253,30,253,29,27,31,46,31,46,30,52,31,21,31,122,31,122,30,122,29,176,31,176,30,255,31,255,30,245,31,143,31,143,30,217,31,229,31,103,31,208,31,208,30,137,31,132,31,217,31,53,31,53,30,1,31,232,31,127,31,242,31,158,31,158,30,191,31,16,31,183,31,244,31,39,31,58,31,58,30,227,31,184,31,184,30,123,31,99,31,12,31,110,31,110,30,168,31,168,30,75,31,113,31,18,31,70,31,70,30,166,31,33,31,88,31,71,31,150,31,176,31,5,31,234,31,166,31,147,31,219,31,19,31,234,31,229,31,33,31,154,31,80,31,87,31,131,31,116,31,64,31,228,31,233,31,64,31,165,31,167,31,62,31,62,30,191,31,244,31,180,31,180,30,163,31,52,31,65,31,233,31,233,30,189,31,215,31,79,31,11,31,5,31,88,31,88,30,221,31,82,31,228,31,198,31,127,31,1,31,170,31,12,31,170,31,216,31,73,31,131,31,232,31,214,31,102,31,245,31,237,31,200,31,64,31,223,31,81,31,81,30,184,31,120,31,120,30,120,29,23,31,232,31,254,31,141,31,34,31,34,30,243,31,13,31,13,30,149,31,127,31,150,31,150,30,150,29,22,31,89,31,114,31,152,31,152,30,152,29,54,31,54,30,169,31,169,30,110,31,110,30,241,31,199,31,199,30,199,29,30,31,225,31,172,31,253,31,102,31,102,30,53,31,194,31,194,30,63,31,63,30,2,31,208,31,196,31,196,30,115,31,204,31,123,31,244,31,244,30,124,31,124,30,164,31,196,31,196,30,227,31,138,31,132,31,147,31,147,30,147,29,237,31,153,31,153,30,153,29,153,28,143,31,219,31,15,31,121,31,157,31,174,31,136,31,230,31,30,31,246,31,138,31,138,30,18,31,112,31,107,31,7,31,189,31,31,31,98,31,95,31,232,31,232,30,236,31,89,31,9,31,242,31,81,31,72,31,122,31,85,31,16,31,3,31,247,31,88,31,249,31,202,31,253,31,69,31,74,31,163,31,24,31,102,31,102,30,102,29,242,31,98,31,129,31,181,31,181,30,9,31,104,31,104,30,117,31,60,31,122,31,133,31,28,31,19,31,207,31,251,31,193,31,104,31,113,31,87,31,52,31,10,31,24,31,118,31,118,30,128,31,35,31,255,31,255,30,79,31,42,31,225,31,225,30,115,31,102,31,176,31,118,31,118,30,254,31,209,31,183,31,29,31,95,31,95,30,95,29,62,31,212,31,11,31,11,30,106,31,238,31,238,30,177,31,85,31,212,31,212,30,212,29,212,28,196,31,93,31,191,31,173,31,173,30,173,29,97,31,63,31,224,31,227,31,36,31,220,31,220,30,150,31,90,31,249,31,30,31,172,31,193,31,132,31,76,31,71,31,209,31,179,31,231,31,21,31,129,31,240,31,222,31,73,31,116,31,71,31,55,31,193,31,1,31,179,31,118,31,201,31,201,30,201,29,84,31,184,31,90,31,90,30,76,31,103,31,127,31,127,30,243,31,107,31,127,31,114,31,153,31,43,31,206,31,162,31,162,30,13,31,43,31,66,31,25,31,171,31,117,31,21,31,192,31,204,31,62,31,169,31,169,30,169,29,10,31,10,30,75,31,75,30,171,31,171,30,164,31,167,31,70,31,85,31,163,31,71,31,117,31,117,30,141,31,120,31,241,31,61,31,181,31,250,31,127,31,127,30,134,31,28,31,25,31,32,31,137,31,142,31,48,31,48,30,37,31,160,31,160,30,160,29,220,31,220,30,220,29,135,31,254,31,195,31,149,31,127,31,105,31,254,31,146,31,33,31,192,31,150,31,230,31,230,30,194,31,194,30,40,31,61,31,136,31,165,31,165,30,23,31,127,31,202,31,62,31,135,31,118,31,75,31,139,31,139,30,231,31,215,31,67,31,153,31,145,31,102,31,185,31,109,31,101,31,8,31,201,31,67,31,176,31,176,30,140,31,140,30,221,31,137,31,215,31,215,30,166,31,170,31,170,30,54,31,55,31,16,31,26,31,88,31,88,30,145,31,145,30,84,31,75,31,57,31,57,30,245,31,31,31,233,31,24,31,50,31,50,30,50,29,50,28,93,31,249,31,171,31,177,31,177,30,91,31,128,31,161,31,240,31,11,31,11,30,200,31,35,31,53,31,151,31,145,31,3,31,32,31,76,31,230,31,242,31,227,31,61,31,53,31,117,31,169,31,128,31,89,31,89,30,136,31,136,30,238,31,238,30,92,31,78,31,155,31,155,30,255,31,226,31,226,30,133,31,79,31,25,31,131,31,190,31,169,31,255,31,129,31,58,31,20,31,216,31,216,30,216,29,216,28,251,31,251,30,225,31,6,31,56,31,67,31,52,31,83,31,20,31,101,31,101,30,101,29,133,31,142,31,86,31,244,31,244,30,196,31,196,30,133,31,137,31,107,31,145,31,43,31,43,30,71,31,109,31,73,31,125,31,136,31,136,30,110,31,226,31,226,30,226,31,226,30,2,31,18,31,197,31,44,31,218,31,221,31,116,31,116,30,253,31,24,31,51,31,231,31,231,30,118,31,118,30,118,29,176,31,176,30,165,31,212,31,169,31,164,31,108,31,93,31,229,31,120,31,210,31,143,31,143,30,199,31,33,31,41,31,204,31,204,30,204,29,204,28,232,31,10,31,169,31,164,31,42,31,11,31,205,31,143,31,239,31,93,31,63,31,107,31,2,31,2,30,194,31,101,31,220,31,169,31,184,31,11,31,175,31,192,31,192,30,3,31,238,31,77,31,211,31,211,30,58,31,198,31,159,31,103,31,103,30,103,29,190,31,182,31,30,31,6,31,6,30,174,31,174,30,197,31,195,31,123,31,252,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
