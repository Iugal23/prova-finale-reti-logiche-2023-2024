-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 777;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,165,0,83,0,213,0,64,0,207,0,68,0,165,0,184,0,197,0,107,0,0,0,0,0,81,0,184,0,44,0,165,0,99,0,20,0,91,0,46,0,0,0,56,0,231,0,99,0,158,0,133,0,235,0,172,0,0,0,0,0,115,0,0,0,57,0,42,0,0,0,21,0,2,0,191,0,227,0,75,0,0,0,45,0,98,0,0,0,194,0,165,0,49,0,81,0,77,0,209,0,24,0,15,0,23,0,9,0,174,0,0,0,196,0,70,0,12,0,122,0,12,0,0,0,233,0,241,0,0,0,246,0,80,0,0,0,163,0,130,0,15,0,237,0,206,0,88,0,164,0,197,0,126,0,181,0,18,0,0,0,54,0,52,0,0,0,43,0,0,0,46,0,205,0,129,0,217,0,233,0,40,0,0,0,231,0,0,0,85,0,69,0,0,0,35,0,109,0,233,0,8,0,114,0,0,0,37,0,208,0,242,0,230,0,0,0,151,0,50,0,235,0,0,0,17,0,251,0,41,0,0,0,0,0,233,0,3,0,100,0,202,0,0,0,56,0,61,0,0,0,98,0,238,0,235,0,59,0,105,0,0,0,175,0,134,0,209,0,174,0,36,0,112,0,203,0,174,0,27,0,40,0,93,0,70,0,0,0,187,0,121,0,98,0,0,0,110,0,252,0,0,0,235,0,0,0,222,0,0,0,64,0,219,0,37,0,231,0,189,0,87,0,0,0,0,0,204,0,245,0,2,0,247,0,65,0,157,0,0,0,19,0,0,0,4,0,0,0,27,0,186,0,253,0,0,0,0,0,64,0,49,0,0,0,0,0,16,0,212,0,243,0,197,0,250,0,67,0,79,0,78,0,190,0,233,0,9,0,0,0,80,0,13,0,134,0,65,0,71,0,143,0,90,0,130,0,0,0,156,0,23,0,128,0,167,0,254,0,39,0,15,0,179,0,24,0,63,0,74,0,118,0,116,0,124,0,0,0,0,0,174,0,255,0,196,0,0,0,12,0,132,0,0,0,211,0,0,0,191,0,238,0,232,0,53,0,216,0,0,0,36,0,183,0,25,0,40,0,139,0,219,0,154,0,155,0,0,0,22,0,131,0,0,0,130,0,229,0,217,0,70,0,167,0,114,0,0,0,0,0,234,0,63,0,0,0,28,0,202,0,215,0,0,0,26,0,53,0,22,0,168,0,202,0,210,0,195,0,144,0,0,0,219,0,232,0,47,0,100,0,101,0,64,0,0,0,0,0,179,0,239,0,170,0,203,0,0,0,114,0,97,0,0,0,29,0,0,0,82,0,141,0,85,0,172,0,197,0,17,0,0,0,120,0,198,0,198,0,0,0,250,0,0,0,212,0,0,0,165,0,148,0,45,0,74,0,218,0,173,0,74,0,129,0,231,0,0,0,142,0,78,0,164,0,213,0,25,0,0,0,141,0,250,0,229,0,0,0,243,0,46,0,175,0,156,0,137,0,40,0,159,0,78,0,64,0,0,0,0,0,21,0,0,0,108,0,240,0,45,0,113,0,48,0,141,0,0,0,120,0,142,0,0,0,113,0,184,0,27,0,0,0,31,0,234,0,107,0,96,0,19,0,98,0,120,0,130,0,111,0,247,0,187,0,227,0,223,0,41,0,125,0,0,0,129,0,0,0,240,0,185,0,159,0,189,0,96,0,141,0,219,0,166,0,124,0,204,0,167,0,57,0,10,0,168,0,20,0,65,0,142,0,61,0,0,0,129,0,169,0,234,0,127,0,218,0,0,0,0,0,243,0,33,0,182,0,37,0,0,0,15,0,0,0,0,0,250,0,216,0,20,0,0,0,180,0,232,0,221,0,121,0,43,0,141,0,31,0,182,0,212,0,232,0,0,0,246,0,0,0,163,0,0,0,221,0,6,0,166,0,222,0,194,0,0,0,154,0,195,0,34,0,61,0,149,0,52,0,62,0,83,0,49,0,133,0,0,0,233,0,241,0,208,0,147,0,57,0,238,0,33,0,149,0,0,0,196,0,193,0,0,0,243,0,23,0,171,0,88,0,23,0,1,0,46,0,22,0,0,0,75,0,232,0,0,0,250,0,236,0,30,0,0,0,43,0,134,0,111,0,240,0,213,0,47,0,28,0,199,0,128,0,0,0,238,0,123,0,0,0,3,0,164,0,0,0,190,0,190,0,239,0,86,0,0,0,38,0,55,0,130,0,128,0,0,0,167,0,233,0,0,0,221,0,228,0,48,0,175,0,0,0,0,0,159,0,16,0,135,0,177,0,23,0,13,0,248,0,0,0,137,0,108,0,240,0,0,0,231,0,111,0,21,0,141,0,0,0,80,0,0,0,230,0,127,0,0,0,14,0,134,0,156,0,148,0,0,0,133,0,7,0,104,0,63,0,209,0,124,0,79,0,209,0,43,0,115,0,110,0,181,0,66,0,206,0,254,0,0,0,122,0,0,0,0,0,41,0,107,0,221,0,77,0,79,0,65,0,104,0,147,0,58,0,215,0,113,0,225,0,9,0,20,0,226,0,84,0,156,0,69,0,0,0,153,0,0,0,0,0,0,0,6,0,218,0,0,0,103,0,27,0,20,0,14,0,9,0,113,0,0,0,107,0,253,0,165,0,85,0,140,0,197,0,174,0,19,0,0,0,64,0,76,0,107,0,9,0,123,0,24,0,135,0,155,0,21,0,30,0,0,0,0,0,154,0,155,0,15,0,0,0,57,0,192,0,153,0,2,0,54,0,68,0,133,0,193,0,26,0,190,0,140,0,102,0,101,0,28,0,200,0,176,0,163,0,129,0,48,0,62,0,36,0,229,0,134,0,0,0,151,0,164,0,30,0,204,0,106,0,250,0,137,0,255,0,243,0,0,0,92,0,0,0,155,0,201,0,41,0,131,0,88,0,109,0,166,0,160,0,137,0,192,0,15,0,155,0,0,0,0,0,35,0,124,0,249,0,121,0,141,0,0,0,169,0,66,0,135,0,199,0,0,0,244,0,0,0,0,0,136,0,4,0,0,0,0,0,225,0,0,0,164,0,214,0,71,0,87,0,19,0,144,0,243,0,195,0,0,0,0,0,141,0,0,0,245,0,195,0,3,0,199,0,0,0,20,0,103,0,24,0,91,0,0,0,25,0,206,0,0,0,0,0,111,0,0,0,0,0,39,0,0,0,159,0,0,0,246,0,88,0,179,0,0,0,234,0,145,0,86,0,36,0,86,0,0,0,158,0,8,0,0,0,182,0,147,0,94,0,164,0,128,0,52,0,0,0,0,0,0,0,0,0,156,0,145,0,0,0,247,0,0,0,210,0,217,0,236,0,207,0,0,0,30,0,104,0,153,0,0,0,155,0,80,0,151,0,0,0,245,0,220,0,0,0,169,0,0,0,112,0,68,0,23,0,69,0,0,0,0,0,185,0,31,0,0,0,13,0,154,0,36,0,97,0,113,0,130,0,121,0,10,0,39,0,11,0,137,0,0,0);
signal scenario_full  : scenario_type := (0,0,165,31,83,31,213,31,64,31,207,31,68,31,165,31,184,31,197,31,107,31,107,30,107,29,81,31,184,31,44,31,165,31,99,31,20,31,91,31,46,31,46,30,56,31,231,31,99,31,158,31,133,31,235,31,172,31,172,30,172,29,115,31,115,30,57,31,42,31,42,30,21,31,2,31,191,31,227,31,75,31,75,30,45,31,98,31,98,30,194,31,165,31,49,31,81,31,77,31,209,31,24,31,15,31,23,31,9,31,174,31,174,30,196,31,70,31,12,31,122,31,12,31,12,30,233,31,241,31,241,30,246,31,80,31,80,30,163,31,130,31,15,31,237,31,206,31,88,31,164,31,197,31,126,31,181,31,18,31,18,30,54,31,52,31,52,30,43,31,43,30,46,31,205,31,129,31,217,31,233,31,40,31,40,30,231,31,231,30,85,31,69,31,69,30,35,31,109,31,233,31,8,31,114,31,114,30,37,31,208,31,242,31,230,31,230,30,151,31,50,31,235,31,235,30,17,31,251,31,41,31,41,30,41,29,233,31,3,31,100,31,202,31,202,30,56,31,61,31,61,30,98,31,238,31,235,31,59,31,105,31,105,30,175,31,134,31,209,31,174,31,36,31,112,31,203,31,174,31,27,31,40,31,93,31,70,31,70,30,187,31,121,31,98,31,98,30,110,31,252,31,252,30,235,31,235,30,222,31,222,30,64,31,219,31,37,31,231,31,189,31,87,31,87,30,87,29,204,31,245,31,2,31,247,31,65,31,157,31,157,30,19,31,19,30,4,31,4,30,27,31,186,31,253,31,253,30,253,29,64,31,49,31,49,30,49,29,16,31,212,31,243,31,197,31,250,31,67,31,79,31,78,31,190,31,233,31,9,31,9,30,80,31,13,31,134,31,65,31,71,31,143,31,90,31,130,31,130,30,156,31,23,31,128,31,167,31,254,31,39,31,15,31,179,31,24,31,63,31,74,31,118,31,116,31,124,31,124,30,124,29,174,31,255,31,196,31,196,30,12,31,132,31,132,30,211,31,211,30,191,31,238,31,232,31,53,31,216,31,216,30,36,31,183,31,25,31,40,31,139,31,219,31,154,31,155,31,155,30,22,31,131,31,131,30,130,31,229,31,217,31,70,31,167,31,114,31,114,30,114,29,234,31,63,31,63,30,28,31,202,31,215,31,215,30,26,31,53,31,22,31,168,31,202,31,210,31,195,31,144,31,144,30,219,31,232,31,47,31,100,31,101,31,64,31,64,30,64,29,179,31,239,31,170,31,203,31,203,30,114,31,97,31,97,30,29,31,29,30,82,31,141,31,85,31,172,31,197,31,17,31,17,30,120,31,198,31,198,31,198,30,250,31,250,30,212,31,212,30,165,31,148,31,45,31,74,31,218,31,173,31,74,31,129,31,231,31,231,30,142,31,78,31,164,31,213,31,25,31,25,30,141,31,250,31,229,31,229,30,243,31,46,31,175,31,156,31,137,31,40,31,159,31,78,31,64,31,64,30,64,29,21,31,21,30,108,31,240,31,45,31,113,31,48,31,141,31,141,30,120,31,142,31,142,30,113,31,184,31,27,31,27,30,31,31,234,31,107,31,96,31,19,31,98,31,120,31,130,31,111,31,247,31,187,31,227,31,223,31,41,31,125,31,125,30,129,31,129,30,240,31,185,31,159,31,189,31,96,31,141,31,219,31,166,31,124,31,204,31,167,31,57,31,10,31,168,31,20,31,65,31,142,31,61,31,61,30,129,31,169,31,234,31,127,31,218,31,218,30,218,29,243,31,33,31,182,31,37,31,37,30,15,31,15,30,15,29,250,31,216,31,20,31,20,30,180,31,232,31,221,31,121,31,43,31,141,31,31,31,182,31,212,31,232,31,232,30,246,31,246,30,163,31,163,30,221,31,6,31,166,31,222,31,194,31,194,30,154,31,195,31,34,31,61,31,149,31,52,31,62,31,83,31,49,31,133,31,133,30,233,31,241,31,208,31,147,31,57,31,238,31,33,31,149,31,149,30,196,31,193,31,193,30,243,31,23,31,171,31,88,31,23,31,1,31,46,31,22,31,22,30,75,31,232,31,232,30,250,31,236,31,30,31,30,30,43,31,134,31,111,31,240,31,213,31,47,31,28,31,199,31,128,31,128,30,238,31,123,31,123,30,3,31,164,31,164,30,190,31,190,31,239,31,86,31,86,30,38,31,55,31,130,31,128,31,128,30,167,31,233,31,233,30,221,31,228,31,48,31,175,31,175,30,175,29,159,31,16,31,135,31,177,31,23,31,13,31,248,31,248,30,137,31,108,31,240,31,240,30,231,31,111,31,21,31,141,31,141,30,80,31,80,30,230,31,127,31,127,30,14,31,134,31,156,31,148,31,148,30,133,31,7,31,104,31,63,31,209,31,124,31,79,31,209,31,43,31,115,31,110,31,181,31,66,31,206,31,254,31,254,30,122,31,122,30,122,29,41,31,107,31,221,31,77,31,79,31,65,31,104,31,147,31,58,31,215,31,113,31,225,31,9,31,20,31,226,31,84,31,156,31,69,31,69,30,153,31,153,30,153,29,153,28,6,31,218,31,218,30,103,31,27,31,20,31,14,31,9,31,113,31,113,30,107,31,253,31,165,31,85,31,140,31,197,31,174,31,19,31,19,30,64,31,76,31,107,31,9,31,123,31,24,31,135,31,155,31,21,31,30,31,30,30,30,29,154,31,155,31,15,31,15,30,57,31,192,31,153,31,2,31,54,31,68,31,133,31,193,31,26,31,190,31,140,31,102,31,101,31,28,31,200,31,176,31,163,31,129,31,48,31,62,31,36,31,229,31,134,31,134,30,151,31,164,31,30,31,204,31,106,31,250,31,137,31,255,31,243,31,243,30,92,31,92,30,155,31,201,31,41,31,131,31,88,31,109,31,166,31,160,31,137,31,192,31,15,31,155,31,155,30,155,29,35,31,124,31,249,31,121,31,141,31,141,30,169,31,66,31,135,31,199,31,199,30,244,31,244,30,244,29,136,31,4,31,4,30,4,29,225,31,225,30,164,31,214,31,71,31,87,31,19,31,144,31,243,31,195,31,195,30,195,29,141,31,141,30,245,31,195,31,3,31,199,31,199,30,20,31,103,31,24,31,91,31,91,30,25,31,206,31,206,30,206,29,111,31,111,30,111,29,39,31,39,30,159,31,159,30,246,31,88,31,179,31,179,30,234,31,145,31,86,31,36,31,86,31,86,30,158,31,8,31,8,30,182,31,147,31,94,31,164,31,128,31,52,31,52,30,52,29,52,28,52,27,156,31,145,31,145,30,247,31,247,30,210,31,217,31,236,31,207,31,207,30,30,31,104,31,153,31,153,30,155,31,80,31,151,31,151,30,245,31,220,31,220,30,169,31,169,30,112,31,68,31,23,31,69,31,69,30,69,29,185,31,31,31,31,30,13,31,154,31,36,31,97,31,113,31,130,31,121,31,10,31,39,31,11,31,137,31,137,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
