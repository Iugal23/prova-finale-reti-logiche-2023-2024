-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 250;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,28,0,134,0,159,0,39,0,211,0,110,0,146,0,170,0,198,0,105,0,0,0,0,0,217,0,85,0,0,0,16,0,37,0,146,0,0,0,59,0,176,0,113,0,0,0,153,0,238,0,41,0,219,0,11,0,228,0,9,0,149,0,190,0,217,0,205,0,0,0,130,0,0,0,161,0,31,0,0,0,55,0,107,0,70,0,0,0,0,0,243,0,63,0,223,0,0,0,142,0,212,0,251,0,198,0,236,0,32,0,0,0,213,0,199,0,21,0,55,0,68,0,248,0,125,0,45,0,146,0,168,0,188,0,189,0,103,0,86,0,14,0,0,0,0,0,92,0,83,0,38,0,0,0,98,0,127,0,233,0,0,0,223,0,245,0,62,0,195,0,67,0,0,0,68,0,0,0,12,0,53,0,0,0,0,0,135,0,0,0,165,0,217,0,214,0,5,0,98,0,221,0,41,0,12,0,129,0,0,0,119,0,65,0,88,0,0,0,0,0,176,0,17,0,45,0,0,0,224,0,111,0,50,0,61,0,26,0,117,0,156,0,62,0,172,0,200,0,128,0,109,0,55,0,0,0,210,0,96,0,161,0,133,0,199,0,189,0,34,0,69,0,13,0,70,0,4,0,119,0,234,0,0,0,115,0,80,0,0,0,0,0,73,0,228,0,246,0,118,0,0,0,68,0,45,0,215,0,229,0,232,0,3,0,108,0,247,0,46,0,63,0,198,0,29,0,157,0,253,0,150,0,169,0,219,0,237,0,125,0,255,0,92,0,123,0,131,0,0,0,28,0,0,0,0,0,45,0,0,0,153,0,83,0,140,0,158,0,0,0,48,0,195,0,180,0,204,0,0,0,124,0,0,0,105,0,0,0,0,0,146,0,251,0,156,0,179,0,0,0,92,0,95,0,39,0,0,0,97,0,111,0,0,0,0,0,232,0,179,0,0,0,0,0,225,0,69,0,70,0,88,0,224,0,196,0,19,0,122,0,62,0,0,0,204,0,186,0,210,0,7,0,0,0,216,0,0,0,0,0,0,0,133,0,78,0,255,0,169,0,232,0,182,0,93,0,102,0,119,0,99,0,0,0,0,0,183,0,190,0,183,0,199,0,5,0,0,0);
signal scenario_full  : scenario_type := (83,31,28,31,134,31,159,31,39,31,211,31,110,31,146,31,170,31,198,31,105,31,105,30,105,29,217,31,85,31,85,30,16,31,37,31,146,31,146,30,59,31,176,31,113,31,113,30,153,31,238,31,41,31,219,31,11,31,228,31,9,31,149,31,190,31,217,31,205,31,205,30,130,31,130,30,161,31,31,31,31,30,55,31,107,31,70,31,70,30,70,29,243,31,63,31,223,31,223,30,142,31,212,31,251,31,198,31,236,31,32,31,32,30,213,31,199,31,21,31,55,31,68,31,248,31,125,31,45,31,146,31,168,31,188,31,189,31,103,31,86,31,14,31,14,30,14,29,92,31,83,31,38,31,38,30,98,31,127,31,233,31,233,30,223,31,245,31,62,31,195,31,67,31,67,30,68,31,68,30,12,31,53,31,53,30,53,29,135,31,135,30,165,31,217,31,214,31,5,31,98,31,221,31,41,31,12,31,129,31,129,30,119,31,65,31,88,31,88,30,88,29,176,31,17,31,45,31,45,30,224,31,111,31,50,31,61,31,26,31,117,31,156,31,62,31,172,31,200,31,128,31,109,31,55,31,55,30,210,31,96,31,161,31,133,31,199,31,189,31,34,31,69,31,13,31,70,31,4,31,119,31,234,31,234,30,115,31,80,31,80,30,80,29,73,31,228,31,246,31,118,31,118,30,68,31,45,31,215,31,229,31,232,31,3,31,108,31,247,31,46,31,63,31,198,31,29,31,157,31,253,31,150,31,169,31,219,31,237,31,125,31,255,31,92,31,123,31,131,31,131,30,28,31,28,30,28,29,45,31,45,30,153,31,83,31,140,31,158,31,158,30,48,31,195,31,180,31,204,31,204,30,124,31,124,30,105,31,105,30,105,29,146,31,251,31,156,31,179,31,179,30,92,31,95,31,39,31,39,30,97,31,111,31,111,30,111,29,232,31,179,31,179,30,179,29,225,31,69,31,70,31,88,31,224,31,196,31,19,31,122,31,62,31,62,30,204,31,186,31,210,31,7,31,7,30,216,31,216,30,216,29,216,28,133,31,78,31,255,31,169,31,232,31,182,31,93,31,102,31,119,31,99,31,99,30,99,29,183,31,190,31,183,31,199,31,5,31,5,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
