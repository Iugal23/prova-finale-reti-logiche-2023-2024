-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_157 is
end project_tb_157;

architecture project_tb_arch_157 of project_tb_157 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 586;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (76,0,171,0,239,0,82,0,0,0,36,0,30,0,219,0,245,0,205,0,32,0,26,0,234,0,230,0,187,0,56,0,156,0,158,0,126,0,171,0,161,0,171,0,0,0,203,0,166,0,74,0,73,0,65,0,102,0,44,0,0,0,61,0,197,0,158,0,0,0,135,0,15,0,0,0,20,0,0,0,0,0,0,0,28,0,1,0,118,0,190,0,76,0,101,0,0,0,178,0,0,0,0,0,247,0,237,0,217,0,99,0,138,0,147,0,82,0,212,0,150,0,24,0,183,0,239,0,244,0,113,0,136,0,118,0,47,0,139,0,246,0,124,0,118,0,246,0,0,0,57,0,32,0,195,0,106,0,0,0,71,0,125,0,71,0,56,0,183,0,172,0,115,0,190,0,117,0,160,0,216,0,151,0,247,0,0,0,39,0,252,0,16,0,6,0,210,0,0,0,98,0,0,0,145,0,211,0,223,0,3,0,248,0,44,0,213,0,64,0,177,0,0,0,197,0,0,0,203,0,238,0,200,0,102,0,101,0,0,0,0,0,5,0,211,0,37,0,132,0,229,0,0,0,0,0,160,0,119,0,58,0,93,0,189,0,167,0,236,0,71,0,243,0,254,0,48,0,181,0,93,0,137,0,45,0,207,0,0,0,159,0,59,0,103,0,0,0,181,0,150,0,0,0,97,0,172,0,127,0,0,0,226,0,0,0,118,0,232,0,201,0,253,0,113,0,163,0,52,0,0,0,249,0,187,0,233,0,0,0,0,0,0,0,0,0,194,0,64,0,120,0,0,0,216,0,0,0,104,0,19,0,232,0,3,0,15,0,62,0,0,0,0,0,157,0,225,0,123,0,127,0,67,0,76,0,197,0,10,0,246,0,0,0,115,0,97,0,246,0,156,0,176,0,4,0,0,0,99,0,35,0,239,0,172,0,191,0,0,0,0,0,250,0,107,0,116,0,202,0,0,0,85,0,194,0,0,0,221,0,9,0,21,0,0,0,224,0,0,0,177,0,80,0,141,0,140,0,68,0,54,0,69,0,0,0,207,0,95,0,241,0,122,0,7,0,75,0,186,0,133,0,0,0,176,0,0,0,172,0,0,0,129,0,187,0,0,0,143,0,0,0,88,0,30,0,199,0,120,0,232,0,0,0,32,0,45,0,107,0,48,0,17,0,0,0,234,0,91,0,146,0,85,0,0,0,168,0,154,0,0,0,125,0,31,0,197,0,123,0,0,0,61,0,198,0,102,0,90,0,144,0,166,0,135,0,255,0,78,0,53,0,109,0,136,0,56,0,144,0,176,0,0,0,0,0,0,0,92,0,112,0,20,0,52,0,100,0,104,0,11,0,24,0,0,0,158,0,65,0,0,0,189,0,124,0,148,0,245,0,74,0,51,0,184,0,0,0,57,0,44,0,13,0,113,0,36,0,116,0,81,0,0,0,226,0,201,0,199,0,0,0,196,0,232,0,118,0,92,0,0,0,197,0,0,0,134,0,0,0,13,0,54,0,148,0,0,0,91,0,110,0,161,0,169,0,51,0,113,0,0,0,0,0,75,0,85,0,238,0,171,0,152,0,210,0,233,0,135,0,48,0,0,0,0,0,175,0,171,0,103,0,0,0,76,0,204,0,44,0,221,0,111,0,207,0,168,0,48,0,0,0,142,0,0,0,211,0,118,0,252,0,94,0,0,0,0,0,0,0,120,0,199,0,172,0,80,0,235,0,154,0,0,0,251,0,232,0,50,0,0,0,21,0,0,0,0,0,0,0,19,0,0,0,113,0,80,0,0,0,7,0,27,0,193,0,247,0,149,0,0,0,218,0,70,0,117,0,113,0,31,0,186,0,120,0,189,0,67,0,55,0,0,0,0,0,0,0,0,0,90,0,203,0,241,0,14,0,17,0,171,0,93,0,142,0,209,0,62,0,0,0,142,0,247,0,36,0,206,0,151,0,0,0,28,0,120,0,0,0,213,0,188,0,61,0,0,0,60,0,0,0,244,0,197,0,2,0,119,0,147,0,81,0,212,0,0,0,117,0,64,0,0,0,25,0,0,0,54,0,178,0,104,0,40,0,75,0,234,0,0,0,231,0,171,0,203,0,137,0,0,0,80,0,137,0,175,0,200,0,0,0,152,0,0,0,80,0,41,0,88,0,211,0,84,0,222,0,226,0,172,0,0,0,230,0,97,0,185,0,119,0,107,0,225,0,123,0,190,0,0,0,0,0,134,0,0,0,0,0,191,0,93,0,135,0,129,0,215,0,0,0,245,0,41,0,246,0,229,0,197,0,111,0,32,0,12,0,248,0,167,0,224,0,134,0,63,0,145,0,225,0,86,0,225,0,20,0,151,0,0,0,47,0,116,0,0,0,128,0,228,0,113,0,207,0,0,0,40,0,103,0,67,0,81,0,0,0,211,0,0,0,84,0,0,0,178,0,226,0,0,0,68,0,202,0,138,0,9,0,117,0,51,0,234,0,2,0,233,0,0,0,55,0,19,0,47,0,6,0,0,0,168,0,125,0,0,0,47,0,193,0,178,0,91,0,228,0,180,0,169,0,204,0,148,0,0,0,164,0,142,0,74,0,122,0,0,0,253,0,21,0,12,0,1,0,0,0,0,0,155,0);
signal scenario_full  : scenario_type := (76,31,171,31,239,31,82,31,82,30,36,31,30,31,219,31,245,31,205,31,32,31,26,31,234,31,230,31,187,31,56,31,156,31,158,31,126,31,171,31,161,31,171,31,171,30,203,31,166,31,74,31,73,31,65,31,102,31,44,31,44,30,61,31,197,31,158,31,158,30,135,31,15,31,15,30,20,31,20,30,20,29,20,28,28,31,1,31,118,31,190,31,76,31,101,31,101,30,178,31,178,30,178,29,247,31,237,31,217,31,99,31,138,31,147,31,82,31,212,31,150,31,24,31,183,31,239,31,244,31,113,31,136,31,118,31,47,31,139,31,246,31,124,31,118,31,246,31,246,30,57,31,32,31,195,31,106,31,106,30,71,31,125,31,71,31,56,31,183,31,172,31,115,31,190,31,117,31,160,31,216,31,151,31,247,31,247,30,39,31,252,31,16,31,6,31,210,31,210,30,98,31,98,30,145,31,211,31,223,31,3,31,248,31,44,31,213,31,64,31,177,31,177,30,197,31,197,30,203,31,238,31,200,31,102,31,101,31,101,30,101,29,5,31,211,31,37,31,132,31,229,31,229,30,229,29,160,31,119,31,58,31,93,31,189,31,167,31,236,31,71,31,243,31,254,31,48,31,181,31,93,31,137,31,45,31,207,31,207,30,159,31,59,31,103,31,103,30,181,31,150,31,150,30,97,31,172,31,127,31,127,30,226,31,226,30,118,31,232,31,201,31,253,31,113,31,163,31,52,31,52,30,249,31,187,31,233,31,233,30,233,29,233,28,233,27,194,31,64,31,120,31,120,30,216,31,216,30,104,31,19,31,232,31,3,31,15,31,62,31,62,30,62,29,157,31,225,31,123,31,127,31,67,31,76,31,197,31,10,31,246,31,246,30,115,31,97,31,246,31,156,31,176,31,4,31,4,30,99,31,35,31,239,31,172,31,191,31,191,30,191,29,250,31,107,31,116,31,202,31,202,30,85,31,194,31,194,30,221,31,9,31,21,31,21,30,224,31,224,30,177,31,80,31,141,31,140,31,68,31,54,31,69,31,69,30,207,31,95,31,241,31,122,31,7,31,75,31,186,31,133,31,133,30,176,31,176,30,172,31,172,30,129,31,187,31,187,30,143,31,143,30,88,31,30,31,199,31,120,31,232,31,232,30,32,31,45,31,107,31,48,31,17,31,17,30,234,31,91,31,146,31,85,31,85,30,168,31,154,31,154,30,125,31,31,31,197,31,123,31,123,30,61,31,198,31,102,31,90,31,144,31,166,31,135,31,255,31,78,31,53,31,109,31,136,31,56,31,144,31,176,31,176,30,176,29,176,28,92,31,112,31,20,31,52,31,100,31,104,31,11,31,24,31,24,30,158,31,65,31,65,30,189,31,124,31,148,31,245,31,74,31,51,31,184,31,184,30,57,31,44,31,13,31,113,31,36,31,116,31,81,31,81,30,226,31,201,31,199,31,199,30,196,31,232,31,118,31,92,31,92,30,197,31,197,30,134,31,134,30,13,31,54,31,148,31,148,30,91,31,110,31,161,31,169,31,51,31,113,31,113,30,113,29,75,31,85,31,238,31,171,31,152,31,210,31,233,31,135,31,48,31,48,30,48,29,175,31,171,31,103,31,103,30,76,31,204,31,44,31,221,31,111,31,207,31,168,31,48,31,48,30,142,31,142,30,211,31,118,31,252,31,94,31,94,30,94,29,94,28,120,31,199,31,172,31,80,31,235,31,154,31,154,30,251,31,232,31,50,31,50,30,21,31,21,30,21,29,21,28,19,31,19,30,113,31,80,31,80,30,7,31,27,31,193,31,247,31,149,31,149,30,218,31,70,31,117,31,113,31,31,31,186,31,120,31,189,31,67,31,55,31,55,30,55,29,55,28,55,27,90,31,203,31,241,31,14,31,17,31,171,31,93,31,142,31,209,31,62,31,62,30,142,31,247,31,36,31,206,31,151,31,151,30,28,31,120,31,120,30,213,31,188,31,61,31,61,30,60,31,60,30,244,31,197,31,2,31,119,31,147,31,81,31,212,31,212,30,117,31,64,31,64,30,25,31,25,30,54,31,178,31,104,31,40,31,75,31,234,31,234,30,231,31,171,31,203,31,137,31,137,30,80,31,137,31,175,31,200,31,200,30,152,31,152,30,80,31,41,31,88,31,211,31,84,31,222,31,226,31,172,31,172,30,230,31,97,31,185,31,119,31,107,31,225,31,123,31,190,31,190,30,190,29,134,31,134,30,134,29,191,31,93,31,135,31,129,31,215,31,215,30,245,31,41,31,246,31,229,31,197,31,111,31,32,31,12,31,248,31,167,31,224,31,134,31,63,31,145,31,225,31,86,31,225,31,20,31,151,31,151,30,47,31,116,31,116,30,128,31,228,31,113,31,207,31,207,30,40,31,103,31,67,31,81,31,81,30,211,31,211,30,84,31,84,30,178,31,226,31,226,30,68,31,202,31,138,31,9,31,117,31,51,31,234,31,2,31,233,31,233,30,55,31,19,31,47,31,6,31,6,30,168,31,125,31,125,30,47,31,193,31,178,31,91,31,228,31,180,31,169,31,204,31,148,31,148,30,164,31,142,31,74,31,122,31,122,30,253,31,21,31,12,31,1,31,1,30,1,29,155,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
