-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_409 is
end project_tb_409;

architecture project_tb_arch_409 of project_tb_409 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 883;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (116,0,79,0,215,0,159,0,88,0,220,0,139,0,0,0,139,0,0,0,125,0,40,0,122,0,140,0,23,0,213,0,73,0,0,0,148,0,25,0,205,0,0,0,15,0,29,0,10,0,28,0,68,0,73,0,0,0,0,0,0,0,138,0,252,0,4,0,178,0,196,0,175,0,245,0,17,0,130,0,254,0,0,0,213,0,201,0,185,0,243,0,50,0,45,0,164,0,40,0,196,0,100,0,165,0,0,0,0,0,181,0,147,0,144,0,70,0,211,0,129,0,152,0,44,0,203,0,0,0,0,0,130,0,64,0,118,0,94,0,170,0,0,0,0,0,130,0,80,0,202,0,129,0,189,0,71,0,0,0,82,0,48,0,65,0,100,0,144,0,108,0,0,0,0,0,11,0,129,0,126,0,155,0,0,0,0,0,202,0,141,0,91,0,0,0,30,0,7,0,0,0,209,0,46,0,236,0,240,0,0,0,0,0,90,0,0,0,0,0,252,0,0,0,147,0,0,0,19,0,159,0,149,0,168,0,223,0,9,0,0,0,0,0,88,0,86,0,238,0,178,0,185,0,0,0,91,0,193,0,198,0,0,0,192,0,243,0,0,0,34,0,4,0,61,0,193,0,154,0,0,0,0,0,88,0,40,0,53,0,252,0,40,0,0,0,132,0,222,0,56,0,70,0,63,0,102,0,138,0,50,0,95,0,31,0,75,0,9,0,0,0,0,0,0,0,164,0,0,0,0,0,191,0,179,0,248,0,248,0,59,0,85,0,148,0,59,0,0,0,149,0,47,0,77,0,184,0,0,0,112,0,99,0,143,0,212,0,101,0,229,0,180,0,102,0,3,0,101,0,0,0,62,0,9,0,246,0,188,0,157,0,187,0,25,0,108,0,95,0,122,0,0,0,163,0,0,0,60,0,133,0,190,0,0,0,0,0,252,0,175,0,210,0,139,0,0,0,7,0,0,0,31,0,8,0,70,0,0,0,226,0,0,0,187,0,123,0,59,0,0,0,186,0,93,0,0,0,53,0,133,0,193,0,217,0,0,0,210,0,255,0,123,0,185,0,87,0,0,0,96,0,167,0,213,0,110,0,194,0,138,0,233,0,0,0,0,0,171,0,28,0,150,0,10,0,50,0,222,0,127,0,205,0,0,0,13,0,0,0,84,0,82,0,0,0,177,0,176,0,253,0,197,0,224,0,95,0,59,0,241,0,97,0,144,0,48,0,32,0,200,0,18,0,0,0,144,0,156,0,67,0,139,0,39,0,196,0,188,0,217,0,139,0,95,0,188,0,87,0,57,0,235,0,0,0,136,0,124,0,0,0,138,0,212,0,138,0,24,0,217,0,10,0,0,0,229,0,0,0,0,0,82,0,45,0,154,0,132,0,243,0,7,0,208,0,103,0,0,0,133,0,251,0,233,0,109,0,165,0,27,0,123,0,73,0,231,0,224,0,177,0,82,0,20,0,163,0,0,0,181,0,0,0,53,0,87,0,29,0,0,0,171,0,0,0,186,0,0,0,243,0,0,0,0,0,9,0,57,0,86,0,27,0,0,0,190,0,96,0,226,0,99,0,0,0,187,0,255,0,171,0,82,0,0,0,157,0,161,0,197,0,240,0,37,0,0,0,0,0,102,0,255,0,0,0,10,0,1,0,0,0,195,0,97,0,41,0,12,0,0,0,230,0,33,0,0,0,218,0,237,0,0,0,176,0,66,0,187,0,158,0,42,0,148,0,137,0,27,0,191,0,0,0,66,0,0,0,0,0,0,0,191,0,249,0,0,0,194,0,84,0,222,0,17,0,125,0,0,0,218,0,90,0,211,0,53,0,83,0,233,0,162,0,176,0,0,0,30,0,19,0,0,0,96,0,0,0,139,0,27,0,115,0,96,0,0,0,223,0,165,0,0,0,241,0,71,0,0,0,41,0,237,0,0,0,0,0,0,0,48,0,163,0,124,0,0,0,251,0,253,0,67,0,211,0,43,0,67,0,0,0,248,0,197,0,0,0,0,0,16,0,0,0,220,0,253,0,181,0,106,0,167,0,174,0,0,0,53,0,0,0,131,0,24,0,55,0,80,0,36,0,40,0,0,0,0,0,0,0,18,0,250,0,93,0,0,0,125,0,2,0,0,0,105,0,32,0,0,0,226,0,181,0,171,0,203,0,189,0,125,0,150,0,40,0,125,0,53,0,196,0,178,0,88,0,33,0,201,0,10,0,200,0,18,0,0,0,187,0,106,0,0,0,78,0,232,0,41,0,205,0,102,0,0,0,231,0,168,0,242,0,0,0,243,0,155,0,123,0,225,0,0,0,0,0,188,0,0,0,92,0,49,0,118,0,14,0,75,0,147,0,33,0,77,0,136,0,232,0,0,0,4,0,120,0,50,0,129,0,159,0,0,0,176,0,0,0,162,0,203,0,175,0,167,0,83,0,0,0,0,0,110,0,111,0,96,0,92,0,0,0,61,0,0,0,243,0,245,0,165,0,0,0,0,0,74,0,49,0,59,0,201,0,220,0,56,0,196,0,143,0,117,0,174,0,82,0,27,0,201,0,119,0,235,0,207,0,80,0,99,0,105,0,181,0,35,0,192,0,0,0,102,0,14,0,234,0,106,0,0,0,32,0,82,0,116,0,142,0,22,0,182,0,167,0,204,0,169,0,0,0,92,0,56,0,240,0,200,0,162,0,228,0,157,0,237,0,17,0,90,0,21,0,143,0,225,0,171,0,3,0,58,0,0,0,223,0,178,0,148,0,0,0,0,0,0,0,116,0,0,0,124,0,140,0,0,0,23,0,21,0,0,0,188,0,141,0,0,0,177,0,0,0,81,0,215,0,165,0,236,0,251,0,226,0,0,0,119,0,137,0,72,0,127,0,71,0,190,0,220,0,107,0,202,0,18,0,126,0,197,0,118,0,81,0,33,0,24,0,0,0,205,0,0,0,76,0,146,0,161,0,203,0,144,0,0,0,135,0,34,0,139,0,47,0,170,0,153,0,121,0,133,0,228,0,0,0,236,0,18,0,119,0,0,0,54,0,1,0,0,0,141,0,111,0,71,0,67,0,141,0,241,0,93,0,115,0,9,0,186,0,85,0,0,0,59,0,218,0,104,0,199,0,44,0,131,0,0,0,190,0,239,0,55,0,78,0,254,0,88,0,0,0,72,0,171,0,164,0,169,0,66,0,41,0,221,0,0,0,18,0,0,0,30,0,193,0,0,0,0,0,238,0,12,0,121,0,234,0,249,0,7,0,43,0,53,0,0,0,218,0,198,0,0,0,180,0,0,0,155,0,0,0,0,0,162,0,229,0,19,0,249,0,178,0,139,0,14,0,81,0,144,0,227,0,255,0,130,0,0,0,235,0,241,0,77,0,100,0,0,0,89,0,47,0,0,0,161,0,225,0,90,0,163,0,245,0,0,0,183,0,3,0,195,0,214,0,111,0,253,0,0,0,158,0,87,0,96,0,203,0,205,0,89,0,0,0,242,0,12,0,242,0,218,0,146,0,204,0,0,0,27,0,145,0,34,0,158,0,98,0,121,0,191,0,0,0,91,0,97,0,56,0,202,0,0,0,3,0,0,0,115,0,40,0,184,0,54,0,66,0,129,0,24,0,70,0,117,0,0,0,218,0,186,0,180,0,0,0,0,0,0,0,101,0,60,0,189,0,219,0,71,0,60,0,168,0,69,0,40,0,66,0,22,0,130,0,181,0,5,0,0,0,239,0,50,0,224,0,29,0,29,0,0,0,0,0,0,0,14,0,0,0,244,0,241,0,18,0,0,0,255,0,226,0,0,0,0,0,223,0,82,0,83,0,6,0,0,0,195,0,145,0,159,0,252,0,0,0,125,0,144,0,57,0,0,0,129,0,0,0,167,0,0,0,41,0,0,0,90,0,154,0,102,0,99,0,207,0,210,0,184,0,189,0,196,0,199,0,70,0,0,0,182,0);
signal scenario_full  : scenario_type := (116,31,79,31,215,31,159,31,88,31,220,31,139,31,139,30,139,31,139,30,125,31,40,31,122,31,140,31,23,31,213,31,73,31,73,30,148,31,25,31,205,31,205,30,15,31,29,31,10,31,28,31,68,31,73,31,73,30,73,29,73,28,138,31,252,31,4,31,178,31,196,31,175,31,245,31,17,31,130,31,254,31,254,30,213,31,201,31,185,31,243,31,50,31,45,31,164,31,40,31,196,31,100,31,165,31,165,30,165,29,181,31,147,31,144,31,70,31,211,31,129,31,152,31,44,31,203,31,203,30,203,29,130,31,64,31,118,31,94,31,170,31,170,30,170,29,130,31,80,31,202,31,129,31,189,31,71,31,71,30,82,31,48,31,65,31,100,31,144,31,108,31,108,30,108,29,11,31,129,31,126,31,155,31,155,30,155,29,202,31,141,31,91,31,91,30,30,31,7,31,7,30,209,31,46,31,236,31,240,31,240,30,240,29,90,31,90,30,90,29,252,31,252,30,147,31,147,30,19,31,159,31,149,31,168,31,223,31,9,31,9,30,9,29,88,31,86,31,238,31,178,31,185,31,185,30,91,31,193,31,198,31,198,30,192,31,243,31,243,30,34,31,4,31,61,31,193,31,154,31,154,30,154,29,88,31,40,31,53,31,252,31,40,31,40,30,132,31,222,31,56,31,70,31,63,31,102,31,138,31,50,31,95,31,31,31,75,31,9,31,9,30,9,29,9,28,164,31,164,30,164,29,191,31,179,31,248,31,248,31,59,31,85,31,148,31,59,31,59,30,149,31,47,31,77,31,184,31,184,30,112,31,99,31,143,31,212,31,101,31,229,31,180,31,102,31,3,31,101,31,101,30,62,31,9,31,246,31,188,31,157,31,187,31,25,31,108,31,95,31,122,31,122,30,163,31,163,30,60,31,133,31,190,31,190,30,190,29,252,31,175,31,210,31,139,31,139,30,7,31,7,30,31,31,8,31,70,31,70,30,226,31,226,30,187,31,123,31,59,31,59,30,186,31,93,31,93,30,53,31,133,31,193,31,217,31,217,30,210,31,255,31,123,31,185,31,87,31,87,30,96,31,167,31,213,31,110,31,194,31,138,31,233,31,233,30,233,29,171,31,28,31,150,31,10,31,50,31,222,31,127,31,205,31,205,30,13,31,13,30,84,31,82,31,82,30,177,31,176,31,253,31,197,31,224,31,95,31,59,31,241,31,97,31,144,31,48,31,32,31,200,31,18,31,18,30,144,31,156,31,67,31,139,31,39,31,196,31,188,31,217,31,139,31,95,31,188,31,87,31,57,31,235,31,235,30,136,31,124,31,124,30,138,31,212,31,138,31,24,31,217,31,10,31,10,30,229,31,229,30,229,29,82,31,45,31,154,31,132,31,243,31,7,31,208,31,103,31,103,30,133,31,251,31,233,31,109,31,165,31,27,31,123,31,73,31,231,31,224,31,177,31,82,31,20,31,163,31,163,30,181,31,181,30,53,31,87,31,29,31,29,30,171,31,171,30,186,31,186,30,243,31,243,30,243,29,9,31,57,31,86,31,27,31,27,30,190,31,96,31,226,31,99,31,99,30,187,31,255,31,171,31,82,31,82,30,157,31,161,31,197,31,240,31,37,31,37,30,37,29,102,31,255,31,255,30,10,31,1,31,1,30,195,31,97,31,41,31,12,31,12,30,230,31,33,31,33,30,218,31,237,31,237,30,176,31,66,31,187,31,158,31,42,31,148,31,137,31,27,31,191,31,191,30,66,31,66,30,66,29,66,28,191,31,249,31,249,30,194,31,84,31,222,31,17,31,125,31,125,30,218,31,90,31,211,31,53,31,83,31,233,31,162,31,176,31,176,30,30,31,19,31,19,30,96,31,96,30,139,31,27,31,115,31,96,31,96,30,223,31,165,31,165,30,241,31,71,31,71,30,41,31,237,31,237,30,237,29,237,28,48,31,163,31,124,31,124,30,251,31,253,31,67,31,211,31,43,31,67,31,67,30,248,31,197,31,197,30,197,29,16,31,16,30,220,31,253,31,181,31,106,31,167,31,174,31,174,30,53,31,53,30,131,31,24,31,55,31,80,31,36,31,40,31,40,30,40,29,40,28,18,31,250,31,93,31,93,30,125,31,2,31,2,30,105,31,32,31,32,30,226,31,181,31,171,31,203,31,189,31,125,31,150,31,40,31,125,31,53,31,196,31,178,31,88,31,33,31,201,31,10,31,200,31,18,31,18,30,187,31,106,31,106,30,78,31,232,31,41,31,205,31,102,31,102,30,231,31,168,31,242,31,242,30,243,31,155,31,123,31,225,31,225,30,225,29,188,31,188,30,92,31,49,31,118,31,14,31,75,31,147,31,33,31,77,31,136,31,232,31,232,30,4,31,120,31,50,31,129,31,159,31,159,30,176,31,176,30,162,31,203,31,175,31,167,31,83,31,83,30,83,29,110,31,111,31,96,31,92,31,92,30,61,31,61,30,243,31,245,31,165,31,165,30,165,29,74,31,49,31,59,31,201,31,220,31,56,31,196,31,143,31,117,31,174,31,82,31,27,31,201,31,119,31,235,31,207,31,80,31,99,31,105,31,181,31,35,31,192,31,192,30,102,31,14,31,234,31,106,31,106,30,32,31,82,31,116,31,142,31,22,31,182,31,167,31,204,31,169,31,169,30,92,31,56,31,240,31,200,31,162,31,228,31,157,31,237,31,17,31,90,31,21,31,143,31,225,31,171,31,3,31,58,31,58,30,223,31,178,31,148,31,148,30,148,29,148,28,116,31,116,30,124,31,140,31,140,30,23,31,21,31,21,30,188,31,141,31,141,30,177,31,177,30,81,31,215,31,165,31,236,31,251,31,226,31,226,30,119,31,137,31,72,31,127,31,71,31,190,31,220,31,107,31,202,31,18,31,126,31,197,31,118,31,81,31,33,31,24,31,24,30,205,31,205,30,76,31,146,31,161,31,203,31,144,31,144,30,135,31,34,31,139,31,47,31,170,31,153,31,121,31,133,31,228,31,228,30,236,31,18,31,119,31,119,30,54,31,1,31,1,30,141,31,111,31,71,31,67,31,141,31,241,31,93,31,115,31,9,31,186,31,85,31,85,30,59,31,218,31,104,31,199,31,44,31,131,31,131,30,190,31,239,31,55,31,78,31,254,31,88,31,88,30,72,31,171,31,164,31,169,31,66,31,41,31,221,31,221,30,18,31,18,30,30,31,193,31,193,30,193,29,238,31,12,31,121,31,234,31,249,31,7,31,43,31,53,31,53,30,218,31,198,31,198,30,180,31,180,30,155,31,155,30,155,29,162,31,229,31,19,31,249,31,178,31,139,31,14,31,81,31,144,31,227,31,255,31,130,31,130,30,235,31,241,31,77,31,100,31,100,30,89,31,47,31,47,30,161,31,225,31,90,31,163,31,245,31,245,30,183,31,3,31,195,31,214,31,111,31,253,31,253,30,158,31,87,31,96,31,203,31,205,31,89,31,89,30,242,31,12,31,242,31,218,31,146,31,204,31,204,30,27,31,145,31,34,31,158,31,98,31,121,31,191,31,191,30,91,31,97,31,56,31,202,31,202,30,3,31,3,30,115,31,40,31,184,31,54,31,66,31,129,31,24,31,70,31,117,31,117,30,218,31,186,31,180,31,180,30,180,29,180,28,101,31,60,31,189,31,219,31,71,31,60,31,168,31,69,31,40,31,66,31,22,31,130,31,181,31,5,31,5,30,239,31,50,31,224,31,29,31,29,31,29,30,29,29,29,28,14,31,14,30,244,31,241,31,18,31,18,30,255,31,226,31,226,30,226,29,223,31,82,31,83,31,6,31,6,30,195,31,145,31,159,31,252,31,252,30,125,31,144,31,57,31,57,30,129,31,129,30,167,31,167,30,41,31,41,30,90,31,154,31,102,31,99,31,207,31,210,31,184,31,189,31,196,31,199,31,70,31,70,30,182,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
