-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 427;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,0,0,217,0,57,0,70,0,112,0,24,0,52,0,180,0,163,0,80,0,0,0,224,0,178,0,87,0,96,0,0,0,48,0,154,0,141,0,206,0,5,0,192,0,226,0,0,0,131,0,164,0,195,0,196,0,0,0,14,0,0,0,65,0,77,0,2,0,0,0,25,0,39,0,97,0,0,0,162,0,65,0,33,0,22,0,121,0,26,0,65,0,0,0,145,0,158,0,118,0,199,0,131,0,250,0,18,0,213,0,182,0,16,0,181,0,233,0,166,0,100,0,68,0,98,0,144,0,0,0,178,0,117,0,62,0,0,0,0,0,0,0,0,0,155,0,55,0,254,0,116,0,26,0,221,0,34,0,93,0,155,0,165,0,172,0,39,0,214,0,124,0,150,0,226,0,233,0,0,0,22,0,72,0,0,0,1,0,0,0,248,0,0,0,220,0,0,0,173,0,0,0,0,0,23,0,0,0,104,0,60,0,93,0,0,0,201,0,84,0,182,0,1,0,105,0,230,0,42,0,109,0,209,0,0,0,112,0,171,0,0,0,161,0,0,0,12,0,25,0,0,0,124,0,51,0,0,0,222,0,124,0,78,0,0,0,88,0,0,0,121,0,0,0,144,0,20,0,36,0,0,0,0,0,171,0,0,0,105,0,3,0,231,0,202,0,0,0,213,0,78,0,0,0,24,0,0,0,242,0,81,0,201,0,40,0,0,0,243,0,155,0,171,0,13,0,173,0,131,0,158,0,96,0,0,0,234,0,183,0,136,0,30,0,145,0,24,0,0,0,121,0,170,0,186,0,0,0,222,0,1,0,0,0,142,0,144,0,86,0,127,0,170,0,26,0,33,0,172,0,16,0,110,0,123,0,24,0,74,0,201,0,182,0,207,0,115,0,184,0,230,0,43,0,194,0,220,0,0,0,76,0,242,0,189,0,252,0,87,0,163,0,0,0,160,0,22,0,17,0,0,0,34,0,0,0,16,0,74,0,128,0,151,0,205,0,245,0,122,0,230,0,252,0,164,0,73,0,188,0,235,0,127,0,201,0,0,0,237,0,0,0,136,0,4,0,0,0,227,0,138,0,0,0,194,0,0,0,119,0,164,0,0,0,92,0,0,0,0,0,3,0,234,0,66,0,204,0,9,0,81,0,149,0,251,0,34,0,162,0,202,0,115,0,6,0,148,0,213,0,0,0,0,0,216,0,203,0,61,0,0,0,0,0,58,0,8,0,91,0,145,0,50,0,95,0,98,0,238,0,35,0,0,0,227,0,157,0,0,0,0,0,200,0,4,0,0,0,63,0,156,0,177,0,177,0,121,0,61,0,241,0,234,0,166,0,0,0,186,0,0,0,78,0,138,0,102,0,114,0,0,0,89,0,237,0,165,0,0,0,176,0,0,0,40,0,0,0,0,0,0,0,119,0,1,0,204,0,124,0,32,0,210,0,62,0,0,0,0,0,0,0,17,0,10,0,0,0,155,0,159,0,0,0,0,0,121,0,0,0,203,0,113,0,156,0,0,0,219,0,42,0,214,0,0,0,36,0,0,0,171,0,171,0,251,0,40,0,232,0,179,0,199,0,73,0,226,0,193,0,203,0,0,0,250,0,138,0,231,0,195,0,143,0,123,0,79,0,207,0,52,0,198,0,190,0,0,0,98,0,254,0,64,0,194,0,22,0,178,0,173,0,0,0,164,0,168,0,72,0,101,0,158,0,196,0,0,0,175,0,162,0,0,0,32,0,190,0,187,0,142,0,164,0,0,0,163,0,148,0,94,0,97,0,0,0,168,0,12,0,67,0,160,0,115,0,215,0,66,0,120,0,116,0,81,0,178,0,0,0,160,0,135,0,215,0,35,0,155,0,85,0,230,0,115,0,0,0,246,0,0,0,0,0,22,0,0,0,55,0,43,0);
signal scenario_full  : scenario_type := (134,31,134,30,217,31,57,31,70,31,112,31,24,31,52,31,180,31,163,31,80,31,80,30,224,31,178,31,87,31,96,31,96,30,48,31,154,31,141,31,206,31,5,31,192,31,226,31,226,30,131,31,164,31,195,31,196,31,196,30,14,31,14,30,65,31,77,31,2,31,2,30,25,31,39,31,97,31,97,30,162,31,65,31,33,31,22,31,121,31,26,31,65,31,65,30,145,31,158,31,118,31,199,31,131,31,250,31,18,31,213,31,182,31,16,31,181,31,233,31,166,31,100,31,68,31,98,31,144,31,144,30,178,31,117,31,62,31,62,30,62,29,62,28,62,27,155,31,55,31,254,31,116,31,26,31,221,31,34,31,93,31,155,31,165,31,172,31,39,31,214,31,124,31,150,31,226,31,233,31,233,30,22,31,72,31,72,30,1,31,1,30,248,31,248,30,220,31,220,30,173,31,173,30,173,29,23,31,23,30,104,31,60,31,93,31,93,30,201,31,84,31,182,31,1,31,105,31,230,31,42,31,109,31,209,31,209,30,112,31,171,31,171,30,161,31,161,30,12,31,25,31,25,30,124,31,51,31,51,30,222,31,124,31,78,31,78,30,88,31,88,30,121,31,121,30,144,31,20,31,36,31,36,30,36,29,171,31,171,30,105,31,3,31,231,31,202,31,202,30,213,31,78,31,78,30,24,31,24,30,242,31,81,31,201,31,40,31,40,30,243,31,155,31,171,31,13,31,173,31,131,31,158,31,96,31,96,30,234,31,183,31,136,31,30,31,145,31,24,31,24,30,121,31,170,31,186,31,186,30,222,31,1,31,1,30,142,31,144,31,86,31,127,31,170,31,26,31,33,31,172,31,16,31,110,31,123,31,24,31,74,31,201,31,182,31,207,31,115,31,184,31,230,31,43,31,194,31,220,31,220,30,76,31,242,31,189,31,252,31,87,31,163,31,163,30,160,31,22,31,17,31,17,30,34,31,34,30,16,31,74,31,128,31,151,31,205,31,245,31,122,31,230,31,252,31,164,31,73,31,188,31,235,31,127,31,201,31,201,30,237,31,237,30,136,31,4,31,4,30,227,31,138,31,138,30,194,31,194,30,119,31,164,31,164,30,92,31,92,30,92,29,3,31,234,31,66,31,204,31,9,31,81,31,149,31,251,31,34,31,162,31,202,31,115,31,6,31,148,31,213,31,213,30,213,29,216,31,203,31,61,31,61,30,61,29,58,31,8,31,91,31,145,31,50,31,95,31,98,31,238,31,35,31,35,30,227,31,157,31,157,30,157,29,200,31,4,31,4,30,63,31,156,31,177,31,177,31,121,31,61,31,241,31,234,31,166,31,166,30,186,31,186,30,78,31,138,31,102,31,114,31,114,30,89,31,237,31,165,31,165,30,176,31,176,30,40,31,40,30,40,29,40,28,119,31,1,31,204,31,124,31,32,31,210,31,62,31,62,30,62,29,62,28,17,31,10,31,10,30,155,31,159,31,159,30,159,29,121,31,121,30,203,31,113,31,156,31,156,30,219,31,42,31,214,31,214,30,36,31,36,30,171,31,171,31,251,31,40,31,232,31,179,31,199,31,73,31,226,31,193,31,203,31,203,30,250,31,138,31,231,31,195,31,143,31,123,31,79,31,207,31,52,31,198,31,190,31,190,30,98,31,254,31,64,31,194,31,22,31,178,31,173,31,173,30,164,31,168,31,72,31,101,31,158,31,196,31,196,30,175,31,162,31,162,30,32,31,190,31,187,31,142,31,164,31,164,30,163,31,148,31,94,31,97,31,97,30,168,31,12,31,67,31,160,31,115,31,215,31,66,31,120,31,116,31,81,31,178,31,178,30,160,31,135,31,215,31,35,31,155,31,85,31,230,31,115,31,115,30,246,31,246,30,246,29,22,31,22,30,55,31,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
