-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_613 is
end project_tb_613;

architecture project_tb_arch_613 of project_tb_613 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 424;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (50,0,112,0,120,0,65,0,255,0,0,0,63,0,95,0,0,0,0,0,0,0,166,0,37,0,28,0,0,0,0,0,221,0,202,0,94,0,129,0,228,0,212,0,206,0,152,0,0,0,0,0,245,0,122,0,61,0,169,0,0,0,213,0,147,0,0,0,180,0,0,0,131,0,0,0,78,0,3,0,159,0,0,0,154,0,0,0,137,0,0,0,121,0,149,0,80,0,222,0,140,0,43,0,243,0,250,0,105,0,55,0,30,0,0,0,69,0,136,0,240,0,181,0,0,0,202,0,0,0,24,0,241,0,18,0,92,0,0,0,223,0,115,0,8,0,216,0,228,0,136,0,191,0,179,0,184,0,167,0,221,0,0,0,6,0,233,0,133,0,232,0,105,0,141,0,199,0,51,0,158,0,31,0,252,0,28,0,3,0,255,0,0,0,64,0,220,0,196,0,0,0,19,0,31,0,106,0,172,0,32,0,0,0,182,0,188,0,101,0,235,0,87,0,140,0,111,0,130,0,51,0,0,0,0,0,167,0,174,0,2,0,49,0,0,0,0,0,36,0,123,0,224,0,179,0,187,0,29,0,228,0,0,0,171,0,60,0,228,0,223,0,127,0,108,0,0,0,0,0,127,0,240,0,0,0,57,0,41,0,79,0,153,0,0,0,3,0,0,0,43,0,52,0,123,0,68,0,117,0,0,0,140,0,215,0,190,0,0,0,155,0,0,0,160,0,167,0,13,0,173,0,121,0,117,0,17,0,108,0,0,0,0,0,59,0,155,0,0,0,34,0,199,0,0,0,140,0,109,0,87,0,12,0,0,0,61,0,123,0,153,0,119,0,5,0,0,0,80,0,181,0,187,0,250,0,0,0,0,0,150,0,27,0,237,0,39,0,0,0,16,0,255,0,0,0,38,0,0,0,0,0,89,0,226,0,17,0,38,0,132,0,195,0,158,0,0,0,225,0,37,0,0,0,136,0,34,0,228,0,34,0,0,0,245,0,122,0,13,0,32,0,43,0,0,0,0,0,25,0,0,0,181,0,189,0,154,0,16,0,171,0,241,0,115,0,117,0,36,0,194,0,228,0,0,0,55,0,0,0,213,0,195,0,122,0,126,0,62,0,70,0,51,0,134,0,95,0,55,0,0,0,44,0,64,0,0,0,168,0,175,0,111,0,128,0,73,0,83,0,162,0,248,0,0,0,7,0,248,0,39,0,226,0,175,0,168,0,14,0,242,0,0,0,28,0,211,0,0,0,128,0,125,0,252,0,59,0,227,0,150,0,0,0,0,0,151,0,0,0,12,0,154,0,201,0,213,0,17,0,0,0,109,0,205,0,29,0,60,0,86,0,128,0,0,0,124,0,0,0,140,0,0,0,145,0,235,0,0,0,223,0,79,0,228,0,210,0,118,0,0,0,140,0,178,0,226,0,0,0,47,0,215,0,62,0,81,0,0,0,16,0,50,0,199,0,145,0,0,0,161,0,31,0,210,0,101,0,83,0,107,0,110,0,123,0,187,0,0,0,141,0,0,0,150,0,174,0,174,0,0,0,232,0,248,0,115,0,213,0,60,0,0,0,210,0,99,0,193,0,228,0,104,0,156,0,32,0,248,0,23,0,26,0,213,0,11,0,0,0,187,0,40,0,0,0,214,0,7,0,195,0,0,0,100,0,179,0,6,0,85,0,0,0,31,0,208,0,200,0,108,0,55,0,0,0,22,0,8,0,169,0,249,0,199,0,19,0,0,0,150,0,227,0,60,0,0,0,132,0,49,0,208,0,33,0,152,0,93,0,106,0,0,0,0,0,176,0,204,0,250,0,1,0,97,0,31,0,0,0,237,0,133,0,221,0,100,0,8,0,214,0,172,0,252,0,0,0,0,0,130,0,0,0,0,0,59,0);
signal scenario_full  : scenario_type := (50,31,112,31,120,31,65,31,255,31,255,30,63,31,95,31,95,30,95,29,95,28,166,31,37,31,28,31,28,30,28,29,221,31,202,31,94,31,129,31,228,31,212,31,206,31,152,31,152,30,152,29,245,31,122,31,61,31,169,31,169,30,213,31,147,31,147,30,180,31,180,30,131,31,131,30,78,31,3,31,159,31,159,30,154,31,154,30,137,31,137,30,121,31,149,31,80,31,222,31,140,31,43,31,243,31,250,31,105,31,55,31,30,31,30,30,69,31,136,31,240,31,181,31,181,30,202,31,202,30,24,31,241,31,18,31,92,31,92,30,223,31,115,31,8,31,216,31,228,31,136,31,191,31,179,31,184,31,167,31,221,31,221,30,6,31,233,31,133,31,232,31,105,31,141,31,199,31,51,31,158,31,31,31,252,31,28,31,3,31,255,31,255,30,64,31,220,31,196,31,196,30,19,31,31,31,106,31,172,31,32,31,32,30,182,31,188,31,101,31,235,31,87,31,140,31,111,31,130,31,51,31,51,30,51,29,167,31,174,31,2,31,49,31,49,30,49,29,36,31,123,31,224,31,179,31,187,31,29,31,228,31,228,30,171,31,60,31,228,31,223,31,127,31,108,31,108,30,108,29,127,31,240,31,240,30,57,31,41,31,79,31,153,31,153,30,3,31,3,30,43,31,52,31,123,31,68,31,117,31,117,30,140,31,215,31,190,31,190,30,155,31,155,30,160,31,167,31,13,31,173,31,121,31,117,31,17,31,108,31,108,30,108,29,59,31,155,31,155,30,34,31,199,31,199,30,140,31,109,31,87,31,12,31,12,30,61,31,123,31,153,31,119,31,5,31,5,30,80,31,181,31,187,31,250,31,250,30,250,29,150,31,27,31,237,31,39,31,39,30,16,31,255,31,255,30,38,31,38,30,38,29,89,31,226,31,17,31,38,31,132,31,195,31,158,31,158,30,225,31,37,31,37,30,136,31,34,31,228,31,34,31,34,30,245,31,122,31,13,31,32,31,43,31,43,30,43,29,25,31,25,30,181,31,189,31,154,31,16,31,171,31,241,31,115,31,117,31,36,31,194,31,228,31,228,30,55,31,55,30,213,31,195,31,122,31,126,31,62,31,70,31,51,31,134,31,95,31,55,31,55,30,44,31,64,31,64,30,168,31,175,31,111,31,128,31,73,31,83,31,162,31,248,31,248,30,7,31,248,31,39,31,226,31,175,31,168,31,14,31,242,31,242,30,28,31,211,31,211,30,128,31,125,31,252,31,59,31,227,31,150,31,150,30,150,29,151,31,151,30,12,31,154,31,201,31,213,31,17,31,17,30,109,31,205,31,29,31,60,31,86,31,128,31,128,30,124,31,124,30,140,31,140,30,145,31,235,31,235,30,223,31,79,31,228,31,210,31,118,31,118,30,140,31,178,31,226,31,226,30,47,31,215,31,62,31,81,31,81,30,16,31,50,31,199,31,145,31,145,30,161,31,31,31,210,31,101,31,83,31,107,31,110,31,123,31,187,31,187,30,141,31,141,30,150,31,174,31,174,31,174,30,232,31,248,31,115,31,213,31,60,31,60,30,210,31,99,31,193,31,228,31,104,31,156,31,32,31,248,31,23,31,26,31,213,31,11,31,11,30,187,31,40,31,40,30,214,31,7,31,195,31,195,30,100,31,179,31,6,31,85,31,85,30,31,31,208,31,200,31,108,31,55,31,55,30,22,31,8,31,169,31,249,31,199,31,19,31,19,30,150,31,227,31,60,31,60,30,132,31,49,31,208,31,33,31,152,31,93,31,106,31,106,30,106,29,176,31,204,31,250,31,1,31,97,31,31,31,31,30,237,31,133,31,221,31,100,31,8,31,214,31,172,31,252,31,252,30,252,29,130,31,130,30,130,29,59,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
