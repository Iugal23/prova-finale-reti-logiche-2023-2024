-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_991 is
end project_tb_991;

architecture project_tb_arch_991 of project_tb_991 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 158;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (110,0,118,0,75,0,117,0,243,0,83,0,0,0,194,0,195,0,186,0,248,0,118,0,131,0,228,0,205,0,0,0,191,0,5,0,227,0,57,0,34,0,5,0,246,0,219,0,0,0,182,0,240,0,182,0,208,0,0,0,0,0,0,0,197,0,242,0,0,0,253,0,0,0,41,0,130,0,0,0,8,0,3,0,188,0,234,0,153,0,237,0,0,0,132,0,231,0,42,0,210,0,130,0,150,0,106,0,171,0,0,0,101,0,58,0,0,0,206,0,0,0,221,0,0,0,183,0,67,0,234,0,117,0,151,0,107,0,53,0,230,0,9,0,128,0,90,0,0,0,164,0,168,0,235,0,233,0,0,0,38,0,126,0,94,0,162,0,87,0,24,0,190,0,74,0,0,0,0,0,138,0,0,0,114,0,0,0,0,0,132,0,0,0,120,0,95,0,0,0,0,0,7,0,181,0,148,0,240,0,150,0,0,0,0,0,78,0,190,0,33,0,79,0,29,0,199,0,209,0,129,0,214,0,137,0,177,0,54,0,188,0,219,0,158,0,76,0,250,0,203,0,0,0,28,0,241,0,156,0,0,0,90,0,221,0,0,0,11,0,235,0,180,0,209,0,181,0,12,0,0,0,245,0,175,0,152,0,107,0,187,0,222,0,254,0,111,0,92,0,206,0,0,0,244,0,59,0,43,0,25,0,71,0,59,0);
signal scenario_full  : scenario_type := (110,31,118,31,75,31,117,31,243,31,83,31,83,30,194,31,195,31,186,31,248,31,118,31,131,31,228,31,205,31,205,30,191,31,5,31,227,31,57,31,34,31,5,31,246,31,219,31,219,30,182,31,240,31,182,31,208,31,208,30,208,29,208,28,197,31,242,31,242,30,253,31,253,30,41,31,130,31,130,30,8,31,3,31,188,31,234,31,153,31,237,31,237,30,132,31,231,31,42,31,210,31,130,31,150,31,106,31,171,31,171,30,101,31,58,31,58,30,206,31,206,30,221,31,221,30,183,31,67,31,234,31,117,31,151,31,107,31,53,31,230,31,9,31,128,31,90,31,90,30,164,31,168,31,235,31,233,31,233,30,38,31,126,31,94,31,162,31,87,31,24,31,190,31,74,31,74,30,74,29,138,31,138,30,114,31,114,30,114,29,132,31,132,30,120,31,95,31,95,30,95,29,7,31,181,31,148,31,240,31,150,31,150,30,150,29,78,31,190,31,33,31,79,31,29,31,199,31,209,31,129,31,214,31,137,31,177,31,54,31,188,31,219,31,158,31,76,31,250,31,203,31,203,30,28,31,241,31,156,31,156,30,90,31,221,31,221,30,11,31,235,31,180,31,209,31,181,31,12,31,12,30,245,31,175,31,152,31,107,31,187,31,222,31,254,31,111,31,92,31,206,31,206,30,244,31,59,31,43,31,25,31,71,31,59,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
