-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 684;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (215,0,0,0,169,0,141,0,0,0,206,0,0,0,63,0,6,0,196,0,167,0,202,0,229,0,46,0,197,0,92,0,217,0,227,0,204,0,0,0,0,0,30,0,140,0,125,0,0,0,115,0,196,0,112,0,133,0,0,0,126,0,0,0,121,0,186,0,147,0,135,0,130,0,7,0,0,0,78,0,71,0,169,0,16,0,157,0,82,0,55,0,180,0,133,0,197,0,0,0,240,0,36,0,26,0,0,0,159,0,226,0,162,0,13,0,178,0,202,0,39,0,35,0,207,0,118,0,145,0,188,0,93,0,0,0,192,0,14,0,161,0,145,0,201,0,166,0,96,0,135,0,0,0,0,0,246,0,213,0,0,0,234,0,0,0,1,0,0,0,6,0,147,0,194,0,223,0,106,0,0,0,243,0,20,0,214,0,0,0,145,0,101,0,0,0,11,0,122,0,107,0,0,0,97,0,9,0,20,0,108,0,17,0,236,0,19,0,171,0,62,0,39,0,0,0,94,0,124,0,220,0,84,0,224,0,128,0,169,0,100,0,239,0,174,0,51,0,0,0,0,0,213,0,80,0,33,0,0,0,48,0,188,0,0,0,182,0,172,0,217,0,0,0,0,0,0,0,151,0,37,0,227,0,91,0,76,0,0,0,216,0,65,0,52,0,0,0,94,0,149,0,27,0,67,0,60,0,254,0,228,0,20,0,17,0,244,0,73,0,0,0,0,0,25,0,79,0,181,0,204,0,32,0,188,0,135,0,183,0,0,0,60,0,38,0,0,0,128,0,0,0,149,0,254,0,193,0,241,0,17,0,0,0,212,0,98,0,84,0,133,0,227,0,92,0,136,0,76,0,89,0,156,0,0,0,93,0,166,0,223,0,116,0,117,0,137,0,0,0,137,0,16,0,111,0,49,0,223,0,61,0,162,0,0,0,190,0,158,0,70,0,71,0,39,0,69,0,0,0,175,0,0,0,57,0,87,0,34,0,194,0,22,0,153,0,204,0,28,0,0,0,95,0,85,0,12,0,147,0,0,0,66,0,95,0,0,0,153,0,175,0,143,0,0,0,0,0,39,0,169,0,125,0,95,0,138,0,5,0,44,0,117,0,0,0,247,0,62,0,49,0,0,0,0,0,74,0,171,0,175,0,135,0,87,0,72,0,0,0,0,0,29,0,57,0,102,0,127,0,188,0,25,0,104,0,180,0,199,0,0,0,95,0,100,0,3,0,164,0,205,0,123,0,122,0,51,0,251,0,0,0,78,0,4,0,144,0,109,0,17,0,104,0,0,0,63,0,235,0,0,0,205,0,0,0,51,0,175,0,3,0,0,0,179,0,0,0,110,0,226,0,0,0,143,0,121,0,191,0,172,0,173,0,0,0,211,0,214,0,136,0,192,0,237,0,10,0,235,0,15,0,0,0,172,0,158,0,103,0,0,0,163,0,174,0,167,0,79,0,197,0,26,0,47,0,0,0,141,0,252,0,70,0,81,0,2,0,113,0,103,0,0,0,0,0,0,0,59,0,13,0,0,0,12,0,235,0,69,0,0,0,96,0,136,0,0,0,67,0,55,0,0,0,96,0,25,0,202,0,120,0,0,0,199,0,29,0,0,0,221,0,108,0,253,0,25,0,18,0,128,0,0,0,84,0,234,0,47,0,108,0,135,0,55,0,43,0,150,0,82,0,1,0,143,0,255,0,206,0,42,0,235,0,0,0,253,0,216,0,115,0,115,0,212,0,0,0,214,0,71,0,75,0,3,0,175,0,0,0,163,0,0,0,0,0,234,0,235,0,0,0,167,0,0,0,152,0,191,0,45,0,129,0,207,0,210,0,0,0,176,0,187,0,0,0,79,0,28,0,124,0,105,0,208,0,168,0,118,0,0,0,126,0,34,0,178,0,34,0,232,0,20,0,111,0,0,0,101,0,0,0,19,0,243,0,0,0,8,0,0,0,231,0,0,0,85,0,46,0,0,0,235,0,74,0,246,0,131,0,83,0,61,0,198,0,143,0,222,0,6,0,99,0,146,0,59,0,143,0,64,0,194,0,0,0,172,0,209,0,0,0,69,0,141,0,2,0,111,0,38,0,0,0,222,0,25,0,146,0,228,0,0,0,51,0,38,0,68,0,84,0,0,0,120,0,0,0,155,0,86,0,159,0,224,0,0,0,153,0,0,0,198,0,182,0,233,0,10,0,21,0,130,0,40,0,29,0,245,0,0,0,76,0,245,0,54,0,166,0,131,0,101,0,212,0,53,0,60,0,198,0,0,0,0,0,167,0,182,0,67,0,134,0,91,0,74,0,168,0,252,0,82,0,44,0,0,0,140,0,121,0,0,0,247,0,205,0,243,0,0,0,190,0,34,0,25,0,0,0,149,0,111,0,13,0,25,0,0,0,140,0,18,0,198,0,91,0,142,0,180,0,0,0,94,0,140,0,200,0,72,0,198,0,0,0,246,0,98,0,0,0,9,0,101,0,250,0,84,0,89,0,6,0,124,0,236,0,108,0,61,0,215,0,77,0,171,0,181,0,146,0,0,0,73,0,0,0,101,0,168,0,35,0,156,0,18,0,0,0,0,0,236,0,0,0,0,0,0,0,44,0,212,0,0,0,28,0,171,0,11,0,26,0,136,0,75,0,153,0,75,0,0,0,149,0,253,0,245,0,0,0,121,0,127,0,0,0,229,0,157,0,115,0,211,0,52,0,182,0,248,0,109,0,121,0,113,0,219,0,23,0,88,0,134,0,167,0,69,0,53,0,149,0,93,0,18,0,254,0,0,0,192,0,223,0,0,0,179,0,57,0,16,0,61,0,102,0,254,0,207,0,189,0,154,0,0,0,251,0,214,0,176,0,3,0,0,0,180,0,89,0,12,0,160,0,183,0,172,0,226,0,134,0,255,0,110,0,108,0,187,0,208,0,150,0,30,0,194,0,193,0,90,0,49,0,28,0,250,0,71,0,44,0,0,0,209,0,0,0,182,0,0,0,0,0,0,0,3,0,113,0,115,0,213,0,115,0,158,0,243,0,68,0,13,0,80,0,175,0,126,0,136,0,15,0,220,0);
signal scenario_full  : scenario_type := (215,31,215,30,169,31,141,31,141,30,206,31,206,30,63,31,6,31,196,31,167,31,202,31,229,31,46,31,197,31,92,31,217,31,227,31,204,31,204,30,204,29,30,31,140,31,125,31,125,30,115,31,196,31,112,31,133,31,133,30,126,31,126,30,121,31,186,31,147,31,135,31,130,31,7,31,7,30,78,31,71,31,169,31,16,31,157,31,82,31,55,31,180,31,133,31,197,31,197,30,240,31,36,31,26,31,26,30,159,31,226,31,162,31,13,31,178,31,202,31,39,31,35,31,207,31,118,31,145,31,188,31,93,31,93,30,192,31,14,31,161,31,145,31,201,31,166,31,96,31,135,31,135,30,135,29,246,31,213,31,213,30,234,31,234,30,1,31,1,30,6,31,147,31,194,31,223,31,106,31,106,30,243,31,20,31,214,31,214,30,145,31,101,31,101,30,11,31,122,31,107,31,107,30,97,31,9,31,20,31,108,31,17,31,236,31,19,31,171,31,62,31,39,31,39,30,94,31,124,31,220,31,84,31,224,31,128,31,169,31,100,31,239,31,174,31,51,31,51,30,51,29,213,31,80,31,33,31,33,30,48,31,188,31,188,30,182,31,172,31,217,31,217,30,217,29,217,28,151,31,37,31,227,31,91,31,76,31,76,30,216,31,65,31,52,31,52,30,94,31,149,31,27,31,67,31,60,31,254,31,228,31,20,31,17,31,244,31,73,31,73,30,73,29,25,31,79,31,181,31,204,31,32,31,188,31,135,31,183,31,183,30,60,31,38,31,38,30,128,31,128,30,149,31,254,31,193,31,241,31,17,31,17,30,212,31,98,31,84,31,133,31,227,31,92,31,136,31,76,31,89,31,156,31,156,30,93,31,166,31,223,31,116,31,117,31,137,31,137,30,137,31,16,31,111,31,49,31,223,31,61,31,162,31,162,30,190,31,158,31,70,31,71,31,39,31,69,31,69,30,175,31,175,30,57,31,87,31,34,31,194,31,22,31,153,31,204,31,28,31,28,30,95,31,85,31,12,31,147,31,147,30,66,31,95,31,95,30,153,31,175,31,143,31,143,30,143,29,39,31,169,31,125,31,95,31,138,31,5,31,44,31,117,31,117,30,247,31,62,31,49,31,49,30,49,29,74,31,171,31,175,31,135,31,87,31,72,31,72,30,72,29,29,31,57,31,102,31,127,31,188,31,25,31,104,31,180,31,199,31,199,30,95,31,100,31,3,31,164,31,205,31,123,31,122,31,51,31,251,31,251,30,78,31,4,31,144,31,109,31,17,31,104,31,104,30,63,31,235,31,235,30,205,31,205,30,51,31,175,31,3,31,3,30,179,31,179,30,110,31,226,31,226,30,143,31,121,31,191,31,172,31,173,31,173,30,211,31,214,31,136,31,192,31,237,31,10,31,235,31,15,31,15,30,172,31,158,31,103,31,103,30,163,31,174,31,167,31,79,31,197,31,26,31,47,31,47,30,141,31,252,31,70,31,81,31,2,31,113,31,103,31,103,30,103,29,103,28,59,31,13,31,13,30,12,31,235,31,69,31,69,30,96,31,136,31,136,30,67,31,55,31,55,30,96,31,25,31,202,31,120,31,120,30,199,31,29,31,29,30,221,31,108,31,253,31,25,31,18,31,128,31,128,30,84,31,234,31,47,31,108,31,135,31,55,31,43,31,150,31,82,31,1,31,143,31,255,31,206,31,42,31,235,31,235,30,253,31,216,31,115,31,115,31,212,31,212,30,214,31,71,31,75,31,3,31,175,31,175,30,163,31,163,30,163,29,234,31,235,31,235,30,167,31,167,30,152,31,191,31,45,31,129,31,207,31,210,31,210,30,176,31,187,31,187,30,79,31,28,31,124,31,105,31,208,31,168,31,118,31,118,30,126,31,34,31,178,31,34,31,232,31,20,31,111,31,111,30,101,31,101,30,19,31,243,31,243,30,8,31,8,30,231,31,231,30,85,31,46,31,46,30,235,31,74,31,246,31,131,31,83,31,61,31,198,31,143,31,222,31,6,31,99,31,146,31,59,31,143,31,64,31,194,31,194,30,172,31,209,31,209,30,69,31,141,31,2,31,111,31,38,31,38,30,222,31,25,31,146,31,228,31,228,30,51,31,38,31,68,31,84,31,84,30,120,31,120,30,155,31,86,31,159,31,224,31,224,30,153,31,153,30,198,31,182,31,233,31,10,31,21,31,130,31,40,31,29,31,245,31,245,30,76,31,245,31,54,31,166,31,131,31,101,31,212,31,53,31,60,31,198,31,198,30,198,29,167,31,182,31,67,31,134,31,91,31,74,31,168,31,252,31,82,31,44,31,44,30,140,31,121,31,121,30,247,31,205,31,243,31,243,30,190,31,34,31,25,31,25,30,149,31,111,31,13,31,25,31,25,30,140,31,18,31,198,31,91,31,142,31,180,31,180,30,94,31,140,31,200,31,72,31,198,31,198,30,246,31,98,31,98,30,9,31,101,31,250,31,84,31,89,31,6,31,124,31,236,31,108,31,61,31,215,31,77,31,171,31,181,31,146,31,146,30,73,31,73,30,101,31,168,31,35,31,156,31,18,31,18,30,18,29,236,31,236,30,236,29,236,28,44,31,212,31,212,30,28,31,171,31,11,31,26,31,136,31,75,31,153,31,75,31,75,30,149,31,253,31,245,31,245,30,121,31,127,31,127,30,229,31,157,31,115,31,211,31,52,31,182,31,248,31,109,31,121,31,113,31,219,31,23,31,88,31,134,31,167,31,69,31,53,31,149,31,93,31,18,31,254,31,254,30,192,31,223,31,223,30,179,31,57,31,16,31,61,31,102,31,254,31,207,31,189,31,154,31,154,30,251,31,214,31,176,31,3,31,3,30,180,31,89,31,12,31,160,31,183,31,172,31,226,31,134,31,255,31,110,31,108,31,187,31,208,31,150,31,30,31,194,31,193,31,90,31,49,31,28,31,250,31,71,31,44,31,44,30,209,31,209,30,182,31,182,30,182,29,182,28,3,31,113,31,115,31,213,31,115,31,158,31,243,31,68,31,13,31,80,31,175,31,126,31,136,31,15,31,220,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
