-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 475;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,255,0,236,0,0,0,0,0,0,0,139,0,168,0,152,0,179,0,0,0,0,0,0,0,123,0,179,0,23,0,9,0,63,0,247,0,75,0,31,0,236,0,30,0,158,0,109,0,37,0,4,0,105,0,101,0,71,0,155,0,76,0,8,0,101,0,0,0,143,0,235,0,0,0,0,0,13,0,81,0,0,0,128,0,135,0,0,0,148,0,237,0,70,0,228,0,115,0,56,0,0,0,108,0,27,0,37,0,207,0,121,0,233,0,199,0,99,0,192,0,232,0,0,0,0,0,13,0,0,0,223,0,161,0,242,0,120,0,210,0,112,0,155,0,178,0,0,0,183,0,11,0,63,0,91,0,0,0,0,0,0,0,191,0,68,0,77,0,169,0,135,0,57,0,123,0,0,0,200,0,0,0,214,0,0,0,20,0,139,0,9,0,195,0,226,0,11,0,201,0,193,0,92,0,0,0,0,0,84,0,105,0,0,0,0,0,230,0,144,0,180,0,163,0,17,0,47,0,0,0,29,0,0,0,127,0,18,0,212,0,241,0,104,0,121,0,32,0,8,0,250,0,0,0,199,0,38,0,165,0,136,0,18,0,31,0,158,0,17,0,84,0,0,0,76,0,183,0,70,0,0,0,178,0,209,0,0,0,0,0,117,0,214,0,0,0,58,0,95,0,0,0,201,0,96,0,254,0,149,0,92,0,195,0,100,0,233,0,239,0,213,0,0,0,164,0,60,0,71,0,150,0,0,0,89,0,189,0,127,0,13,0,103,0,93,0,234,0,247,0,106,0,163,0,152,0,252,0,43,0,201,0,0,0,122,0,0,0,41,0,95,0,96,0,12,0,101,0,0,0,139,0,237,0,126,0,203,0,0,0,121,0,247,0,197,0,77,0,205,0,0,0,61,0,0,0,154,0,49,0,171,0,246,0,179,0,110,0,100,0,237,0,219,0,80,0,0,0,177,0,176,0,137,0,14,0,179,0,0,0,255,0,98,0,105,0,194,0,0,0,0,0,216,0,154,0,6,0,22,0,171,0,0,0,218,0,216,0,48,0,100,0,165,0,0,0,119,0,219,0,138,0,107,0,173,0,88,0,61,0,168,0,181,0,16,0,29,0,0,0,238,0,0,0,162,0,54,0,206,0,205,0,189,0,100,0,30,0,138,0,0,0,0,0,190,0,111,0,41,0,247,0,137,0,31,0,61,0,179,0,85,0,142,0,0,0,203,0,141,0,185,0,87,0,190,0,145,0,63,0,215,0,39,0,37,0,250,0,97,0,0,0,211,0,0,0,16,0,182,0,165,0,226,0,121,0,214,0,178,0,108,0,252,0,21,0,24,0,111,0,64,0,163,0,247,0,0,0,93,0,88,0,216,0,173,0,41,0,100,0,56,0,0,0,93,0,51,0,168,0,66,0,150,0,0,0,0,0,77,0,227,0,98,0,0,0,202,0,52,0,89,0,114,0,228,0,62,0,190,0,0,0,176,0,0,0,0,0,194,0,0,0,166,0,0,0,99,0,0,0,92,0,97,0,177,0,85,0,166,0,171,0,146,0,112,0,125,0,176,0,179,0,190,0,63,0,108,0,21,0,70,0,135,0,219,0,250,0,49,0,194,0,0,0,26,0,206,0,0,0,224,0,224,0,218,0,82,0,218,0,3,0,77,0,0,0,182,0,222,0,133,0,154,0,242,0,0,0,0,0,44,0,161,0,233,0,184,0,195,0,179,0,152,0,0,0,186,0,0,0,62,0,106,0,77,0,120,0,90,0,0,0,192,0,20,0,67,0,0,0,38,0,109,0,83,0,16,0,104,0,74,0,130,0,30,0,0,0,222,0,250,0,191,0,165,0,54,0,213,0,193,0,85,0,13,0,106,0,0,0,0,0,143,0,20,0,123,0,200,0,112,0,111,0,250,0,78,0,73,0,118,0,247,0,0,0,0,0,0,0,170,0,43,0,184,0,182,0,202,0,42,0,59,0,69,0,118,0,6,0,0,0,0,0,93,0,182,0,127,0,149,0,87,0,10,0,67,0,0,0,5,0,117,0,180,0,213,0,77,0,167,0,0,0,116,0,0,0,0,0,171,0,240,0,37,0,88,0,70,0,127,0,163,0,154,0,0,0);
signal scenario_full  : scenario_type := (139,31,255,31,236,31,236,30,236,29,236,28,139,31,168,31,152,31,179,31,179,30,179,29,179,28,123,31,179,31,23,31,9,31,63,31,247,31,75,31,31,31,236,31,30,31,158,31,109,31,37,31,4,31,105,31,101,31,71,31,155,31,76,31,8,31,101,31,101,30,143,31,235,31,235,30,235,29,13,31,81,31,81,30,128,31,135,31,135,30,148,31,237,31,70,31,228,31,115,31,56,31,56,30,108,31,27,31,37,31,207,31,121,31,233,31,199,31,99,31,192,31,232,31,232,30,232,29,13,31,13,30,223,31,161,31,242,31,120,31,210,31,112,31,155,31,178,31,178,30,183,31,11,31,63,31,91,31,91,30,91,29,91,28,191,31,68,31,77,31,169,31,135,31,57,31,123,31,123,30,200,31,200,30,214,31,214,30,20,31,139,31,9,31,195,31,226,31,11,31,201,31,193,31,92,31,92,30,92,29,84,31,105,31,105,30,105,29,230,31,144,31,180,31,163,31,17,31,47,31,47,30,29,31,29,30,127,31,18,31,212,31,241,31,104,31,121,31,32,31,8,31,250,31,250,30,199,31,38,31,165,31,136,31,18,31,31,31,158,31,17,31,84,31,84,30,76,31,183,31,70,31,70,30,178,31,209,31,209,30,209,29,117,31,214,31,214,30,58,31,95,31,95,30,201,31,96,31,254,31,149,31,92,31,195,31,100,31,233,31,239,31,213,31,213,30,164,31,60,31,71,31,150,31,150,30,89,31,189,31,127,31,13,31,103,31,93,31,234,31,247,31,106,31,163,31,152,31,252,31,43,31,201,31,201,30,122,31,122,30,41,31,95,31,96,31,12,31,101,31,101,30,139,31,237,31,126,31,203,31,203,30,121,31,247,31,197,31,77,31,205,31,205,30,61,31,61,30,154,31,49,31,171,31,246,31,179,31,110,31,100,31,237,31,219,31,80,31,80,30,177,31,176,31,137,31,14,31,179,31,179,30,255,31,98,31,105,31,194,31,194,30,194,29,216,31,154,31,6,31,22,31,171,31,171,30,218,31,216,31,48,31,100,31,165,31,165,30,119,31,219,31,138,31,107,31,173,31,88,31,61,31,168,31,181,31,16,31,29,31,29,30,238,31,238,30,162,31,54,31,206,31,205,31,189,31,100,31,30,31,138,31,138,30,138,29,190,31,111,31,41,31,247,31,137,31,31,31,61,31,179,31,85,31,142,31,142,30,203,31,141,31,185,31,87,31,190,31,145,31,63,31,215,31,39,31,37,31,250,31,97,31,97,30,211,31,211,30,16,31,182,31,165,31,226,31,121,31,214,31,178,31,108,31,252,31,21,31,24,31,111,31,64,31,163,31,247,31,247,30,93,31,88,31,216,31,173,31,41,31,100,31,56,31,56,30,93,31,51,31,168,31,66,31,150,31,150,30,150,29,77,31,227,31,98,31,98,30,202,31,52,31,89,31,114,31,228,31,62,31,190,31,190,30,176,31,176,30,176,29,194,31,194,30,166,31,166,30,99,31,99,30,92,31,97,31,177,31,85,31,166,31,171,31,146,31,112,31,125,31,176,31,179,31,190,31,63,31,108,31,21,31,70,31,135,31,219,31,250,31,49,31,194,31,194,30,26,31,206,31,206,30,224,31,224,31,218,31,82,31,218,31,3,31,77,31,77,30,182,31,222,31,133,31,154,31,242,31,242,30,242,29,44,31,161,31,233,31,184,31,195,31,179,31,152,31,152,30,186,31,186,30,62,31,106,31,77,31,120,31,90,31,90,30,192,31,20,31,67,31,67,30,38,31,109,31,83,31,16,31,104,31,74,31,130,31,30,31,30,30,222,31,250,31,191,31,165,31,54,31,213,31,193,31,85,31,13,31,106,31,106,30,106,29,143,31,20,31,123,31,200,31,112,31,111,31,250,31,78,31,73,31,118,31,247,31,247,30,247,29,247,28,170,31,43,31,184,31,182,31,202,31,42,31,59,31,69,31,118,31,6,31,6,30,6,29,93,31,182,31,127,31,149,31,87,31,10,31,67,31,67,30,5,31,117,31,180,31,213,31,77,31,167,31,167,30,116,31,116,30,116,29,171,31,240,31,37,31,88,31,70,31,127,31,163,31,154,31,154,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
