-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_440 is
end project_tb_440;

architecture project_tb_arch_440 of project_tb_440 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 971;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,140,0,106,0,123,0,242,0,205,0,37,0,130,0,165,0,156,0,196,0,22,0,156,0,135,0,49,0,0,0,0,0,44,0,83,0,118,0,0,0,17,0,96,0,222,0,102,0,0,0,122,0,0,0,252,0,245,0,58,0,0,0,163,0,127,0,158,0,75,0,173,0,221,0,233,0,56,0,168,0,17,0,119,0,203,0,235,0,136,0,45,0,206,0,142,0,157,0,0,0,4,0,182,0,0,0,95,0,136,0,247,0,251,0,225,0,0,0,103,0,0,0,57,0,184,0,0,0,178,0,0,0,180,0,160,0,92,0,0,0,7,0,0,0,176,0,94,0,111,0,118,0,197,0,114,0,0,0,199,0,245,0,0,0,193,0,24,0,113,0,84,0,114,0,58,0,248,0,68,0,13,0,0,0,239,0,147,0,47,0,56,0,17,0,148,0,0,0,78,0,125,0,37,0,232,0,165,0,0,0,243,0,196,0,71,0,242,0,156,0,103,0,229,0,54,0,52,0,32,0,249,0,203,0,0,0,0,0,25,0,153,0,75,0,44,0,130,0,23,0,85,0,0,0,42,0,202,0,43,0,51,0,2,0,230,0,40,0,229,0,248,0,246,0,76,0,10,0,43,0,112,0,138,0,164,0,36,0,200,0,84,0,30,0,80,0,38,0,0,0,128,0,39,0,211,0,0,0,219,0,102,0,90,0,91,0,50,0,219,0,149,0,72,0,0,0,145,0,15,0,0,0,0,0,216,0,199,0,244,0,90,0,82,0,123,0,106,0,0,0,0,0,0,0,46,0,238,0,0,0,35,0,202,0,0,0,98,0,248,0,176,0,0,0,59,0,0,0,185,0,65,0,239,0,212,0,179,0,100,0,163,0,0,0,235,0,91,0,251,0,204,0,218,0,64,0,196,0,9,0,143,0,12,0,156,0,0,0,44,0,0,0,129,0,0,0,65,0,165,0,37,0,24,0,227,0,100,0,188,0,165,0,241,0,0,0,0,0,0,0,99,0,0,0,227,0,0,0,14,0,0,0,213,0,202,0,156,0,130,0,93,0,233,0,29,0,138,0,154,0,0,0,0,0,227,0,0,0,49,0,125,0,148,0,165,0,0,0,122,0,38,0,39,0,92,0,196,0,149,0,70,0,60,0,237,0,157,0,0,0,249,0,44,0,0,0,51,0,101,0,67,0,243,0,0,0,181,0,0,0,187,0,113,0,57,0,216,0,207,0,157,0,77,0,0,0,48,0,139,0,0,0,0,0,92,0,163,0,173,0,239,0,0,0,10,0,195,0,17,0,158,0,120,0,150,0,3,0,242,0,0,0,0,0,15,0,47,0,0,0,42,0,22,0,0,0,79,0,105,0,131,0,34,0,0,0,197,0,51,0,174,0,0,0,253,0,140,0,0,0,202,0,36,0,228,0,0,0,98,0,0,0,207,0,0,0,0,0,149,0,0,0,242,0,64,0,13,0,173,0,172,0,12,0,185,0,143,0,113,0,199,0,177,0,116,0,44,0,69,0,112,0,240,0,209,0,0,0,0,0,210,0,121,0,99,0,59,0,105,0,136,0,0,0,217,0,87,0,0,0,37,0,0,0,79,0,125,0,154,0,52,0,0,0,39,0,0,0,94,0,0,0,61,0,37,0,72,0,109,0,184,0,8,0,204,0,239,0,168,0,0,0,0,0,158,0,130,0,131,0,239,0,46,0,62,0,209,0,35,0,250,0,77,0,106,0,224,0,37,0,140,0,188,0,0,0,26,0,115,0,59,0,113,0,131,0,0,0,179,0,141,0,15,0,0,0,232,0,0,0,0,0,78,0,0,0,5,0,221,0,35,0,0,0,29,0,109,0,81,0,244,0,197,0,246,0,128,0,84,0,176,0,80,0,22,0,0,0,176,0,0,0,22,0,16,0,242,0,101,0,231,0,248,0,0,0,145,0,199,0,0,0,76,0,0,0,127,0,0,0,188,0,185,0,233,0,204,0,147,0,211,0,98,0,90,0,39,0,138,0,125,0,0,0,15,0,176,0,0,0,0,0,156,0,177,0,19,0,128,0,100,0,90,0,254,0,0,0,118,0,142,0,0,0,233,0,58,0,145,0,28,0,153,0,209,0,0,0,225,0,214,0,73,0,192,0,206,0,96,0,205,0,197,0,43,0,0,0,233,0,94,0,134,0,0,0,40,0,108,0,193,0,119,0,33,0,244,0,0,0,22,0,240,0,32,0,193,0,212,0,37,0,49,0,46,0,241,0,151,0,173,0,0,0,31,0,106,0,159,0,191,0,201,0,0,0,111,0,0,0,0,0,242,0,127,0,145,0,219,0,0,0,71,0,171,0,222,0,0,0,208,0,102,0,189,0,78,0,34,0,196,0,0,0,137,0,233,0,5,0,225,0,0,0,0,0,90,0,0,0,213,0,0,0,0,0,203,0,26,0,162,0,0,0,0,0,0,0,0,0,179,0,118,0,0,0,130,0,0,0,0,0,0,0,203,0,143,0,42,0,90,0,195,0,214,0,0,0,236,0,0,0,52,0,225,0,229,0,91,0,216,0,148,0,11,0,0,0,30,0,154,0,0,0,143,0,0,0,48,0,158,0,0,0,98,0,156,0,204,0,70,0,160,0,249,0,154,0,0,0,0,0,246,0,108,0,217,0,67,0,203,0,0,0,118,0,52,0,183,0,86,0,72,0,195,0,75,0,166,0,7,0,225,0,146,0,72,0,191,0,78,0,0,0,248,0,244,0,33,0,30,0,97,0,157,0,117,0,246,0,97,0,39,0,141,0,0,0,229,0,128,0,211,0,183,0,93,0,61,0,80,0,135,0,4,0,180,0,0,0,104,0,15,0,56,0,86,0,13,0,210,0,0,0,0,0,30,0,111,0,78,0,0,0,67,0,0,0,93,0,193,0,61,0,38,0,85,0,87,0,97,0,189,0,193,0,13,0,167,0,0,0,253,0,19,0,96,0,210,0,72,0,86,0,107,0,204,0,202,0,253,0,0,0,0,0,0,0,235,0,136,0,235,0,137,0,2,0,0,0,249,0,0,0,246,0,65,0,0,0,246,0,100,0,0,0,81,0,11,0,130,0,0,0,198,0,127,0,204,0,107,0,107,0,183,0,128,0,3,0,173,0,119,0,164,0,138,0,123,0,250,0,175,0,1,0,159,0,193,0,76,0,206,0,67,0,20,0,171,0,20,0,158,0,184,0,147,0,191,0,254,0,114,0,116,0,73,0,197,0,140,0,160,0,17,0,180,0,215,0,163,0,191,0,0,0,156,0,20,0,142,0,158,0,167,0,162,0,0,0,23,0,144,0,48,0,192,0,9,0,92,0,32,0,97,0,132,0,0,0,105,0,0,0,0,0,0,0,18,0,217,0,150,0,84,0,125,0,91,0,164,0,245,0,40,0,173,0,236,0,47,0,104,0,182,0,38,0,198,0,34,0,174,0,111,0,0,0,0,0,226,0,121,0,0,0,5,0,73,0,255,0,101,0,116,0,0,0,20,0,228,0,118,0,240,0,153,0,122,0,0,0,49,0,93,0,0,0,151,0,0,0,119,0,220,0,250,0,179,0,67,0,214,0,145,0,44,0,0,0,86,0,0,0,95,0,0,0,71,0,141,0,206,0,216,0,0,0,76,0,0,0,9,0,210,0,102,0,69,0,154,0,241,0,0,0,86,0,60,0,232,0,150,0,99,0,121,0,98,0,172,0,207,0,100,0,0,0,128,0,195,0,98,0,163,0,112,0,64,0,140,0,96,0,156,0,234,0,123,0,151,0,0,0,0,0,165,0,183,0,4,0,202,0,44,0,168,0,245,0,0,0,55,0,12,0,193,0,215,0,67,0,32,0,62,0,172,0,58,0,17,0,0,0,65,0,0,0,187,0,102,0,88,0,115,0,61,0,17,0,0,0,184,0,0,0,181,0,92,0,56,0,0,0,0,0,192,0,0,0,209,0,0,0,100,0,83,0,223,0,40,0,221,0,62,0,173,0,43,0,0,0,54,0,210,0,73,0,15,0,146,0,14,0,100,0,164,0,146,0,0,0,83,0,0,0,233,0,0,0,22,0,211,0,109,0,0,0,195,0,151,0,92,0,0,0,199,0,0,0,71,0,145,0,195,0,212,0,0,0,11,0,159,0,175,0,183,0,0,0,166,0,69,0,13,0,0,0,48,0,66,0,69,0,8,0,204,0,62,0,0,0,237,0,107,0,120,0,120,0,3,0,0,0,0,0,40,0,179,0,133,0,29,0,240,0,163,0,172,0,193,0,65,0,239,0,164,0,196,0,237,0,0,0,188,0,0,0,71,0,0,0,105,0,172,0,223,0,0,0);
signal scenario_full  : scenario_type := (219,31,140,31,106,31,123,31,242,31,205,31,37,31,130,31,165,31,156,31,196,31,22,31,156,31,135,31,49,31,49,30,49,29,44,31,83,31,118,31,118,30,17,31,96,31,222,31,102,31,102,30,122,31,122,30,252,31,245,31,58,31,58,30,163,31,127,31,158,31,75,31,173,31,221,31,233,31,56,31,168,31,17,31,119,31,203,31,235,31,136,31,45,31,206,31,142,31,157,31,157,30,4,31,182,31,182,30,95,31,136,31,247,31,251,31,225,31,225,30,103,31,103,30,57,31,184,31,184,30,178,31,178,30,180,31,160,31,92,31,92,30,7,31,7,30,176,31,94,31,111,31,118,31,197,31,114,31,114,30,199,31,245,31,245,30,193,31,24,31,113,31,84,31,114,31,58,31,248,31,68,31,13,31,13,30,239,31,147,31,47,31,56,31,17,31,148,31,148,30,78,31,125,31,37,31,232,31,165,31,165,30,243,31,196,31,71,31,242,31,156,31,103,31,229,31,54,31,52,31,32,31,249,31,203,31,203,30,203,29,25,31,153,31,75,31,44,31,130,31,23,31,85,31,85,30,42,31,202,31,43,31,51,31,2,31,230,31,40,31,229,31,248,31,246,31,76,31,10,31,43,31,112,31,138,31,164,31,36,31,200,31,84,31,30,31,80,31,38,31,38,30,128,31,39,31,211,31,211,30,219,31,102,31,90,31,91,31,50,31,219,31,149,31,72,31,72,30,145,31,15,31,15,30,15,29,216,31,199,31,244,31,90,31,82,31,123,31,106,31,106,30,106,29,106,28,46,31,238,31,238,30,35,31,202,31,202,30,98,31,248,31,176,31,176,30,59,31,59,30,185,31,65,31,239,31,212,31,179,31,100,31,163,31,163,30,235,31,91,31,251,31,204,31,218,31,64,31,196,31,9,31,143,31,12,31,156,31,156,30,44,31,44,30,129,31,129,30,65,31,165,31,37,31,24,31,227,31,100,31,188,31,165,31,241,31,241,30,241,29,241,28,99,31,99,30,227,31,227,30,14,31,14,30,213,31,202,31,156,31,130,31,93,31,233,31,29,31,138,31,154,31,154,30,154,29,227,31,227,30,49,31,125,31,148,31,165,31,165,30,122,31,38,31,39,31,92,31,196,31,149,31,70,31,60,31,237,31,157,31,157,30,249,31,44,31,44,30,51,31,101,31,67,31,243,31,243,30,181,31,181,30,187,31,113,31,57,31,216,31,207,31,157,31,77,31,77,30,48,31,139,31,139,30,139,29,92,31,163,31,173,31,239,31,239,30,10,31,195,31,17,31,158,31,120,31,150,31,3,31,242,31,242,30,242,29,15,31,47,31,47,30,42,31,22,31,22,30,79,31,105,31,131,31,34,31,34,30,197,31,51,31,174,31,174,30,253,31,140,31,140,30,202,31,36,31,228,31,228,30,98,31,98,30,207,31,207,30,207,29,149,31,149,30,242,31,64,31,13,31,173,31,172,31,12,31,185,31,143,31,113,31,199,31,177,31,116,31,44,31,69,31,112,31,240,31,209,31,209,30,209,29,210,31,121,31,99,31,59,31,105,31,136,31,136,30,217,31,87,31,87,30,37,31,37,30,79,31,125,31,154,31,52,31,52,30,39,31,39,30,94,31,94,30,61,31,37,31,72,31,109,31,184,31,8,31,204,31,239,31,168,31,168,30,168,29,158,31,130,31,131,31,239,31,46,31,62,31,209,31,35,31,250,31,77,31,106,31,224,31,37,31,140,31,188,31,188,30,26,31,115,31,59,31,113,31,131,31,131,30,179,31,141,31,15,31,15,30,232,31,232,30,232,29,78,31,78,30,5,31,221,31,35,31,35,30,29,31,109,31,81,31,244,31,197,31,246,31,128,31,84,31,176,31,80,31,22,31,22,30,176,31,176,30,22,31,16,31,242,31,101,31,231,31,248,31,248,30,145,31,199,31,199,30,76,31,76,30,127,31,127,30,188,31,185,31,233,31,204,31,147,31,211,31,98,31,90,31,39,31,138,31,125,31,125,30,15,31,176,31,176,30,176,29,156,31,177,31,19,31,128,31,100,31,90,31,254,31,254,30,118,31,142,31,142,30,233,31,58,31,145,31,28,31,153,31,209,31,209,30,225,31,214,31,73,31,192,31,206,31,96,31,205,31,197,31,43,31,43,30,233,31,94,31,134,31,134,30,40,31,108,31,193,31,119,31,33,31,244,31,244,30,22,31,240,31,32,31,193,31,212,31,37,31,49,31,46,31,241,31,151,31,173,31,173,30,31,31,106,31,159,31,191,31,201,31,201,30,111,31,111,30,111,29,242,31,127,31,145,31,219,31,219,30,71,31,171,31,222,31,222,30,208,31,102,31,189,31,78,31,34,31,196,31,196,30,137,31,233,31,5,31,225,31,225,30,225,29,90,31,90,30,213,31,213,30,213,29,203,31,26,31,162,31,162,30,162,29,162,28,162,27,179,31,118,31,118,30,130,31,130,30,130,29,130,28,203,31,143,31,42,31,90,31,195,31,214,31,214,30,236,31,236,30,52,31,225,31,229,31,91,31,216,31,148,31,11,31,11,30,30,31,154,31,154,30,143,31,143,30,48,31,158,31,158,30,98,31,156,31,204,31,70,31,160,31,249,31,154,31,154,30,154,29,246,31,108,31,217,31,67,31,203,31,203,30,118,31,52,31,183,31,86,31,72,31,195,31,75,31,166,31,7,31,225,31,146,31,72,31,191,31,78,31,78,30,248,31,244,31,33,31,30,31,97,31,157,31,117,31,246,31,97,31,39,31,141,31,141,30,229,31,128,31,211,31,183,31,93,31,61,31,80,31,135,31,4,31,180,31,180,30,104,31,15,31,56,31,86,31,13,31,210,31,210,30,210,29,30,31,111,31,78,31,78,30,67,31,67,30,93,31,193,31,61,31,38,31,85,31,87,31,97,31,189,31,193,31,13,31,167,31,167,30,253,31,19,31,96,31,210,31,72,31,86,31,107,31,204,31,202,31,253,31,253,30,253,29,253,28,235,31,136,31,235,31,137,31,2,31,2,30,249,31,249,30,246,31,65,31,65,30,246,31,100,31,100,30,81,31,11,31,130,31,130,30,198,31,127,31,204,31,107,31,107,31,183,31,128,31,3,31,173,31,119,31,164,31,138,31,123,31,250,31,175,31,1,31,159,31,193,31,76,31,206,31,67,31,20,31,171,31,20,31,158,31,184,31,147,31,191,31,254,31,114,31,116,31,73,31,197,31,140,31,160,31,17,31,180,31,215,31,163,31,191,31,191,30,156,31,20,31,142,31,158,31,167,31,162,31,162,30,23,31,144,31,48,31,192,31,9,31,92,31,32,31,97,31,132,31,132,30,105,31,105,30,105,29,105,28,18,31,217,31,150,31,84,31,125,31,91,31,164,31,245,31,40,31,173,31,236,31,47,31,104,31,182,31,38,31,198,31,34,31,174,31,111,31,111,30,111,29,226,31,121,31,121,30,5,31,73,31,255,31,101,31,116,31,116,30,20,31,228,31,118,31,240,31,153,31,122,31,122,30,49,31,93,31,93,30,151,31,151,30,119,31,220,31,250,31,179,31,67,31,214,31,145,31,44,31,44,30,86,31,86,30,95,31,95,30,71,31,141,31,206,31,216,31,216,30,76,31,76,30,9,31,210,31,102,31,69,31,154,31,241,31,241,30,86,31,60,31,232,31,150,31,99,31,121,31,98,31,172,31,207,31,100,31,100,30,128,31,195,31,98,31,163,31,112,31,64,31,140,31,96,31,156,31,234,31,123,31,151,31,151,30,151,29,165,31,183,31,4,31,202,31,44,31,168,31,245,31,245,30,55,31,12,31,193,31,215,31,67,31,32,31,62,31,172,31,58,31,17,31,17,30,65,31,65,30,187,31,102,31,88,31,115,31,61,31,17,31,17,30,184,31,184,30,181,31,92,31,56,31,56,30,56,29,192,31,192,30,209,31,209,30,100,31,83,31,223,31,40,31,221,31,62,31,173,31,43,31,43,30,54,31,210,31,73,31,15,31,146,31,14,31,100,31,164,31,146,31,146,30,83,31,83,30,233,31,233,30,22,31,211,31,109,31,109,30,195,31,151,31,92,31,92,30,199,31,199,30,71,31,145,31,195,31,212,31,212,30,11,31,159,31,175,31,183,31,183,30,166,31,69,31,13,31,13,30,48,31,66,31,69,31,8,31,204,31,62,31,62,30,237,31,107,31,120,31,120,31,3,31,3,30,3,29,40,31,179,31,133,31,29,31,240,31,163,31,172,31,193,31,65,31,239,31,164,31,196,31,237,31,237,30,188,31,188,30,71,31,71,30,105,31,172,31,223,31,223,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
