-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 655;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (224,0,109,0,110,0,209,0,71,0,211,0,117,0,0,0,58,0,96,0,202,0,50,0,129,0,173,0,104,0,0,0,236,0,0,0,0,0,85,0,0,0,210,0,13,0,204,0,136,0,188,0,177,0,39,0,63,0,168,0,109,0,0,0,0,0,9,0,93,0,55,0,141,0,0,0,0,0,27,0,56,0,128,0,199,0,0,0,201,0,15,0,64,0,182,0,31,0,53,0,108,0,137,0,98,0,220,0,207,0,149,0,179,0,116,0,151,0,7,0,93,0,0,0,124,0,1,0,187,0,127,0,0,0,0,0,168,0,4,0,140,0,0,0,13,0,48,0,82,0,31,0,137,0,64,0,73,0,241,0,238,0,60,0,62,0,18,0,172,0,157,0,0,0,6,0,151,0,80,0,49,0,228,0,18,0,0,0,211,0,247,0,84,0,232,0,20,0,226,0,0,0,0,0,38,0,252,0,166,0,137,0,114,0,166,0,233,0,210,0,72,0,52,0,1,0,181,0,34,0,81,0,14,0,51,0,195,0,214,0,172,0,200,0,185,0,168,0,81,0,11,0,242,0,46,0,230,0,253,0,114,0,165,0,57,0,70,0,0,0,86,0,198,0,157,0,52,0,0,0,249,0,62,0,94,0,57,0,19,0,69,0,110,0,89,0,63,0,114,0,46,0,112,0,126,0,123,0,224,0,4,0,86,0,209,0,15,0,80,0,0,0,99,0,149,0,67,0,174,0,239,0,173,0,2,0,0,0,0,0,108,0,0,0,0,0,203,0,141,0,87,0,176,0,183,0,144,0,0,0,244,0,0,0,146,0,37,0,0,0,150,0,42,0,0,0,233,0,0,0,62,0,47,0,76,0,24,0,141,0,248,0,255,0,0,0,0,0,185,0,159,0,212,0,114,0,79,0,13,0,120,0,190,0,85,0,0,0,101,0,153,0,231,0,254,0,131,0,119,0,0,0,205,0,0,0,168,0,0,0,106,0,133,0,0,0,0,0,237,0,86,0,38,0,76,0,111,0,180,0,0,0,0,0,202,0,136,0,183,0,0,0,102,0,214,0,0,0,53,0,178,0,154,0,80,0,55,0,236,0,0,0,26,0,26,0,211,0,0,0,149,0,0,0,253,0,0,0,159,0,91,0,183,0,120,0,31,0,152,0,206,0,0,0,177,0,142,0,120,0,100,0,140,0,241,0,84,0,75,0,128,0,0,0,160,0,172,0,0,0,85,0,222,0,127,0,45,0,0,0,0,0,0,0,121,0,200,0,116,0,0,0,51,0,162,0,0,0,0,0,52,0,100,0,91,0,169,0,36,0,77,0,59,0,204,0,0,0,211,0,0,0,174,0,128,0,68,0,44,0,131,0,13,0,101,0,0,0,0,0,237,0,0,0,79,0,0,0,67,0,174,0,66,0,0,0,19,0,224,0,144,0,97,0,0,0,56,0,228,0,78,0,0,0,122,0,180,0,180,0,192,0,141,0,0,0,249,0,105,0,5,0,221,0,164,0,0,0,174,0,229,0,20,0,99,0,226,0,0,0,241,0,245,0,127,0,230,0,211,0,250,0,98,0,0,0,70,0,0,0,37,0,25,0,0,0,81,0,100,0,115,0,0,0,218,0,96,0,141,0,0,0,25,0,93,0,3,0,25,0,197,0,164,0,12,0,217,0,24,0,72,0,125,0,7,0,188,0,56,0,0,0,7,0,0,0,84,0,0,0,32,0,0,0,202,0,89,0,3,0,194,0,61,0,164,0,0,0,0,0,246,0,124,0,215,0,76,0,41,0,21,0,0,0,226,0,195,0,96,0,0,0,145,0,122,0,82,0,12,0,0,0,146,0,0,0,63,0,139,0,8,0,75,0,0,0,0,0,176,0,56,0,64,0,215,0,107,0,42,0,9,0,120,0,175,0,193,0,252,0,128,0,0,0,84,0,0,0,193,0,0,0,24,0,0,0,0,0,254,0,211,0,160,0,0,0,179,0,53,0,16,0,49,0,118,0,78,0,135,0,171,0,104,0,117,0,5,0,151,0,0,0,186,0,0,0,227,0,130,0,20,0,190,0,35,0,47,0,56,0,73,0,167,0,25,0,234,0,151,0,97,0,15,0,0,0,144,0,143,0,196,0,10,0,164,0,50,0,116,0,43,0,122,0,87,0,57,0,128,0,127,0,166,0,55,0,116,0,253,0,248,0,247,0,33,0,159,0,21,0,1,0,180,0,192,0,39,0,149,0,0,0,250,0,235,0,220,0,0,0,0,0,107,0,210,0,0,0,23,0,164,0,0,0,52,0,0,0,0,0,218,0,29,0,55,0,8,0,147,0,209,0,107,0,235,0,253,0,25,0,210,0,21,0,239,0,169,0,186,0,216,0,62,0,84,0,129,0,51,0,253,0,255,0,5,0,0,0,83,0,5,0,247,0,206,0,114,0,0,0,170,0,0,0,115,0,225,0,179,0,19,0,0,0,236,0,53,0,103,0,0,0,0,0,252,0,228,0,172,0,255,0,208,0,10,0,16,0,52,0,100,0,170,0,5,0,196,0,79,0,182,0,161,0,0,0,253,0,37,0,239,0,143,0,0,0,30,0,226,0,29,0,233,0,0,0,131,0,103,0,125,0,153,0,0,0,0,0,198,0,47,0,24,0,25,0,77,0,161,0,118,0,130,0,245,0,190,0,32,0,17,0,227,0,226,0,0,0,188,0,0,0,103,0,147,0,22,0,0,0,52,0,22,0,165,0,254,0,55,0,205,0,201,0,0,0,0,0,0,0,241,0,165,0,188,0,0,0,147,0,134,0,18,0,0,0,82,0,69,0,113,0,0,0,116,0,131,0,153,0,224,0,104,0,32,0,27,0,20,0,199,0,172,0,0,0,143,0,230,0,158,0,0,0,114,0,69,0,0,0,49,0,6,0,0,0,231,0,206,0);
signal scenario_full  : scenario_type := (224,31,109,31,110,31,209,31,71,31,211,31,117,31,117,30,58,31,96,31,202,31,50,31,129,31,173,31,104,31,104,30,236,31,236,30,236,29,85,31,85,30,210,31,13,31,204,31,136,31,188,31,177,31,39,31,63,31,168,31,109,31,109,30,109,29,9,31,93,31,55,31,141,31,141,30,141,29,27,31,56,31,128,31,199,31,199,30,201,31,15,31,64,31,182,31,31,31,53,31,108,31,137,31,98,31,220,31,207,31,149,31,179,31,116,31,151,31,7,31,93,31,93,30,124,31,1,31,187,31,127,31,127,30,127,29,168,31,4,31,140,31,140,30,13,31,48,31,82,31,31,31,137,31,64,31,73,31,241,31,238,31,60,31,62,31,18,31,172,31,157,31,157,30,6,31,151,31,80,31,49,31,228,31,18,31,18,30,211,31,247,31,84,31,232,31,20,31,226,31,226,30,226,29,38,31,252,31,166,31,137,31,114,31,166,31,233,31,210,31,72,31,52,31,1,31,181,31,34,31,81,31,14,31,51,31,195,31,214,31,172,31,200,31,185,31,168,31,81,31,11,31,242,31,46,31,230,31,253,31,114,31,165,31,57,31,70,31,70,30,86,31,198,31,157,31,52,31,52,30,249,31,62,31,94,31,57,31,19,31,69,31,110,31,89,31,63,31,114,31,46,31,112,31,126,31,123,31,224,31,4,31,86,31,209,31,15,31,80,31,80,30,99,31,149,31,67,31,174,31,239,31,173,31,2,31,2,30,2,29,108,31,108,30,108,29,203,31,141,31,87,31,176,31,183,31,144,31,144,30,244,31,244,30,146,31,37,31,37,30,150,31,42,31,42,30,233,31,233,30,62,31,47,31,76,31,24,31,141,31,248,31,255,31,255,30,255,29,185,31,159,31,212,31,114,31,79,31,13,31,120,31,190,31,85,31,85,30,101,31,153,31,231,31,254,31,131,31,119,31,119,30,205,31,205,30,168,31,168,30,106,31,133,31,133,30,133,29,237,31,86,31,38,31,76,31,111,31,180,31,180,30,180,29,202,31,136,31,183,31,183,30,102,31,214,31,214,30,53,31,178,31,154,31,80,31,55,31,236,31,236,30,26,31,26,31,211,31,211,30,149,31,149,30,253,31,253,30,159,31,91,31,183,31,120,31,31,31,152,31,206,31,206,30,177,31,142,31,120,31,100,31,140,31,241,31,84,31,75,31,128,31,128,30,160,31,172,31,172,30,85,31,222,31,127,31,45,31,45,30,45,29,45,28,121,31,200,31,116,31,116,30,51,31,162,31,162,30,162,29,52,31,100,31,91,31,169,31,36,31,77,31,59,31,204,31,204,30,211,31,211,30,174,31,128,31,68,31,44,31,131,31,13,31,101,31,101,30,101,29,237,31,237,30,79,31,79,30,67,31,174,31,66,31,66,30,19,31,224,31,144,31,97,31,97,30,56,31,228,31,78,31,78,30,122,31,180,31,180,31,192,31,141,31,141,30,249,31,105,31,5,31,221,31,164,31,164,30,174,31,229,31,20,31,99,31,226,31,226,30,241,31,245,31,127,31,230,31,211,31,250,31,98,31,98,30,70,31,70,30,37,31,25,31,25,30,81,31,100,31,115,31,115,30,218,31,96,31,141,31,141,30,25,31,93,31,3,31,25,31,197,31,164,31,12,31,217,31,24,31,72,31,125,31,7,31,188,31,56,31,56,30,7,31,7,30,84,31,84,30,32,31,32,30,202,31,89,31,3,31,194,31,61,31,164,31,164,30,164,29,246,31,124,31,215,31,76,31,41,31,21,31,21,30,226,31,195,31,96,31,96,30,145,31,122,31,82,31,12,31,12,30,146,31,146,30,63,31,139,31,8,31,75,31,75,30,75,29,176,31,56,31,64,31,215,31,107,31,42,31,9,31,120,31,175,31,193,31,252,31,128,31,128,30,84,31,84,30,193,31,193,30,24,31,24,30,24,29,254,31,211,31,160,31,160,30,179,31,53,31,16,31,49,31,118,31,78,31,135,31,171,31,104,31,117,31,5,31,151,31,151,30,186,31,186,30,227,31,130,31,20,31,190,31,35,31,47,31,56,31,73,31,167,31,25,31,234,31,151,31,97,31,15,31,15,30,144,31,143,31,196,31,10,31,164,31,50,31,116,31,43,31,122,31,87,31,57,31,128,31,127,31,166,31,55,31,116,31,253,31,248,31,247,31,33,31,159,31,21,31,1,31,180,31,192,31,39,31,149,31,149,30,250,31,235,31,220,31,220,30,220,29,107,31,210,31,210,30,23,31,164,31,164,30,52,31,52,30,52,29,218,31,29,31,55,31,8,31,147,31,209,31,107,31,235,31,253,31,25,31,210,31,21,31,239,31,169,31,186,31,216,31,62,31,84,31,129,31,51,31,253,31,255,31,5,31,5,30,83,31,5,31,247,31,206,31,114,31,114,30,170,31,170,30,115,31,225,31,179,31,19,31,19,30,236,31,53,31,103,31,103,30,103,29,252,31,228,31,172,31,255,31,208,31,10,31,16,31,52,31,100,31,170,31,5,31,196,31,79,31,182,31,161,31,161,30,253,31,37,31,239,31,143,31,143,30,30,31,226,31,29,31,233,31,233,30,131,31,103,31,125,31,153,31,153,30,153,29,198,31,47,31,24,31,25,31,77,31,161,31,118,31,130,31,245,31,190,31,32,31,17,31,227,31,226,31,226,30,188,31,188,30,103,31,147,31,22,31,22,30,52,31,22,31,165,31,254,31,55,31,205,31,201,31,201,30,201,29,201,28,241,31,165,31,188,31,188,30,147,31,134,31,18,31,18,30,82,31,69,31,113,31,113,30,116,31,131,31,153,31,224,31,104,31,32,31,27,31,20,31,199,31,172,31,172,30,143,31,230,31,158,31,158,30,114,31,69,31,69,30,49,31,6,31,6,30,231,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
