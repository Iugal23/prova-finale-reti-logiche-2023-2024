-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 613;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (191,0,3,0,129,0,57,0,38,0,0,0,41,0,1,0,249,0,0,0,0,0,138,0,240,0,123,0,247,0,0,0,253,0,98,0,131,0,43,0,192,0,71,0,96,0,238,0,0,0,134,0,232,0,85,0,0,0,116,0,36,0,0,0,243,0,167,0,1,0,0,0,150,0,50,0,0,0,251,0,46,0,225,0,162,0,25,0,157,0,176,0,164,0,230,0,132,0,238,0,64,0,213,0,153,0,79,0,247,0,255,0,38,0,108,0,77,0,36,0,79,0,248,0,51,0,0,0,178,0,160,0,106,0,182,0,254,0,0,0,137,0,48,0,37,0,0,0,11,0,0,0,213,0,75,0,125,0,46,0,220,0,0,0,63,0,115,0,207,0,154,0,39,0,97,0,30,0,189,0,174,0,0,0,0,0,0,0,246,0,1,0,113,0,42,0,217,0,0,0,203,0,0,0,0,0,186,0,33,0,243,0,194,0,150,0,2,0,79,0,27,0,72,0,147,0,0,0,163,0,0,0,86,0,0,0,161,0,55,0,0,0,34,0,226,0,192,0,170,0,40,0,214,0,215,0,235,0,72,0,24,0,249,0,60,0,4,0,236,0,0,0,230,0,79,0,204,0,79,0,78,0,0,0,109,0,149,0,57,0,4,0,93,0,251,0,118,0,59,0,86,0,105,0,18,0,103,0,61,0,229,0,0,0,249,0,155,0,42,0,246,0,232,0,237,0,78,0,162,0,55,0,179,0,0,0,0,0,249,0,103,0,0,0,67,0,44,0,194,0,220,0,9,0,0,0,207,0,87,0,0,0,213,0,0,0,179,0,0,0,228,0,242,0,74,0,255,0,52,0,0,0,206,0,230,0,0,0,41,0,35,0,188,0,140,0,89,0,0,0,23,0,7,0,117,0,106,0,230,0,0,0,35,0,199,0,95,0,0,0,162,0,0,0,19,0,0,0,0,0,0,0,167,0,23,0,248,0,83,0,148,0,151,0,0,0,234,0,68,0,23,0,0,0,35,0,126,0,0,0,231,0,0,0,161,0,164,0,0,0,0,0,152,0,0,0,119,0,244,0,38,0,89,0,0,0,0,0,166,0,0,0,34,0,48,0,5,0,35,0,121,0,201,0,0,0,183,0,200,0,91,0,0,0,67,0,7,0,0,0,0,0,230,0,191,0,194,0,143,0,250,0,152,0,0,0,74,0,0,0,0,0,228,0,208,0,0,0,73,0,114,0,0,0,153,0,39,0,48,0,0,0,71,0,212,0,106,0,82,0,119,0,253,0,57,0,76,0,255,0,188,0,0,0,62,0,1,0,16,0,175,0,0,0,33,0,0,0,168,0,192,0,121,0,11,0,166,0,0,0,101,0,230,0,75,0,136,0,181,0,189,0,91,0,0,0,90,0,14,0,0,0,131,0,249,0,88,0,34,0,95,0,122,0,44,0,0,0,138,0,44,0,191,0,110,0,248,0,180,0,0,0,1,0,242,0,216,0,176,0,49,0,8,0,252,0,151,0,97,0,41,0,0,0,38,0,1,0,162,0,112,0,0,0,56,0,130,0,220,0,4,0,113,0,129,0,202,0,78,0,110,0,167,0,180,0,151,0,237,0,0,0,114,0,227,0,212,0,35,0,0,0,36,0,240,0,64,0,181,0,221,0,48,0,249,0,166,0,0,0,0,0,12,0,0,0,148,0,177,0,16,0,156,0,65,0,232,0,0,0,0,0,141,0,49,0,215,0,209,0,0,0,1,0,122,0,135,0,0,0,128,0,144,0,83,0,0,0,108,0,0,0,0,0,145,0,0,0,10,0,172,0,0,0,0,0,50,0,0,0,32,0,253,0,12,0,213,0,38,0,0,0,156,0,165,0,129,0,43,0,250,0,194,0,0,0,0,0,192,0,131,0,89,0,0,0,89,0,161,0,187,0,78,0,177,0,118,0,71,0,159,0,114,0,241,0,130,0,152,0,187,0,125,0,230,0,174,0,73,0,49,0,87,0,119,0,206,0,129,0,243,0,0,0,9,0,0,0,216,0,162,0,87,0,114,0,0,0,202,0,196,0,69,0,227,0,0,0,80,0,0,0,94,0,158,0,0,0,187,0,0,0,212,0,129,0,0,0,161,0,134,0,12,0,0,0,4,0,16,0,110,0,47,0,66,0,252,0,0,0,149,0,11,0,163,0,0,0,253,0,93,0,185,0,0,0,156,0,218,0,212,0,43,0,92,0,59,0,0,0,9,0,35,0,140,0,238,0,0,0,0,0,106,0,237,0,140,0,80,0,0,0,26,0,206,0,19,0,139,0,0,0,55,0,255,0,11,0,104,0,172,0,208,0,156,0,203,0,1,0,121,0,191,0,177,0,115,0,219,0,132,0,203,0,0,0,223,0,0,0,151,0,247,0,0,0,170,0,107,0,62,0,144,0,142,0,37,0,137,0,160,0,11,0,0,0,35,0,66,0,0,0,243,0,0,0,174,0,167,0,120,0,0,0,114,0,20,0,194,0,169,0,192,0,0,0,222,0,0,0,108,0,0,0,0,0,83,0,47,0,243,0,34,0,117,0,195,0,107,0,72,0,53,0,73,0,119,0,133,0,143,0,45,0,162,0,88,0,128,0,159,0,0,0,224,0,31,0,175,0,247,0,23,0,31,0,0,0,241,0,44,0,0,0,211,0,128,0,127,0,0,0,99,0,66,0,60,0,204,0,82,0,178,0,217,0,0,0,173,0,115,0,14,0,103,0);
signal scenario_full  : scenario_type := (191,31,3,31,129,31,57,31,38,31,38,30,41,31,1,31,249,31,249,30,249,29,138,31,240,31,123,31,247,31,247,30,253,31,98,31,131,31,43,31,192,31,71,31,96,31,238,31,238,30,134,31,232,31,85,31,85,30,116,31,36,31,36,30,243,31,167,31,1,31,1,30,150,31,50,31,50,30,251,31,46,31,225,31,162,31,25,31,157,31,176,31,164,31,230,31,132,31,238,31,64,31,213,31,153,31,79,31,247,31,255,31,38,31,108,31,77,31,36,31,79,31,248,31,51,31,51,30,178,31,160,31,106,31,182,31,254,31,254,30,137,31,48,31,37,31,37,30,11,31,11,30,213,31,75,31,125,31,46,31,220,31,220,30,63,31,115,31,207,31,154,31,39,31,97,31,30,31,189,31,174,31,174,30,174,29,174,28,246,31,1,31,113,31,42,31,217,31,217,30,203,31,203,30,203,29,186,31,33,31,243,31,194,31,150,31,2,31,79,31,27,31,72,31,147,31,147,30,163,31,163,30,86,31,86,30,161,31,55,31,55,30,34,31,226,31,192,31,170,31,40,31,214,31,215,31,235,31,72,31,24,31,249,31,60,31,4,31,236,31,236,30,230,31,79,31,204,31,79,31,78,31,78,30,109,31,149,31,57,31,4,31,93,31,251,31,118,31,59,31,86,31,105,31,18,31,103,31,61,31,229,31,229,30,249,31,155,31,42,31,246,31,232,31,237,31,78,31,162,31,55,31,179,31,179,30,179,29,249,31,103,31,103,30,67,31,44,31,194,31,220,31,9,31,9,30,207,31,87,31,87,30,213,31,213,30,179,31,179,30,228,31,242,31,74,31,255,31,52,31,52,30,206,31,230,31,230,30,41,31,35,31,188,31,140,31,89,31,89,30,23,31,7,31,117,31,106,31,230,31,230,30,35,31,199,31,95,31,95,30,162,31,162,30,19,31,19,30,19,29,19,28,167,31,23,31,248,31,83,31,148,31,151,31,151,30,234,31,68,31,23,31,23,30,35,31,126,31,126,30,231,31,231,30,161,31,164,31,164,30,164,29,152,31,152,30,119,31,244,31,38,31,89,31,89,30,89,29,166,31,166,30,34,31,48,31,5,31,35,31,121,31,201,31,201,30,183,31,200,31,91,31,91,30,67,31,7,31,7,30,7,29,230,31,191,31,194,31,143,31,250,31,152,31,152,30,74,31,74,30,74,29,228,31,208,31,208,30,73,31,114,31,114,30,153,31,39,31,48,31,48,30,71,31,212,31,106,31,82,31,119,31,253,31,57,31,76,31,255,31,188,31,188,30,62,31,1,31,16,31,175,31,175,30,33,31,33,30,168,31,192,31,121,31,11,31,166,31,166,30,101,31,230,31,75,31,136,31,181,31,189,31,91,31,91,30,90,31,14,31,14,30,131,31,249,31,88,31,34,31,95,31,122,31,44,31,44,30,138,31,44,31,191,31,110,31,248,31,180,31,180,30,1,31,242,31,216,31,176,31,49,31,8,31,252,31,151,31,97,31,41,31,41,30,38,31,1,31,162,31,112,31,112,30,56,31,130,31,220,31,4,31,113,31,129,31,202,31,78,31,110,31,167,31,180,31,151,31,237,31,237,30,114,31,227,31,212,31,35,31,35,30,36,31,240,31,64,31,181,31,221,31,48,31,249,31,166,31,166,30,166,29,12,31,12,30,148,31,177,31,16,31,156,31,65,31,232,31,232,30,232,29,141,31,49,31,215,31,209,31,209,30,1,31,122,31,135,31,135,30,128,31,144,31,83,31,83,30,108,31,108,30,108,29,145,31,145,30,10,31,172,31,172,30,172,29,50,31,50,30,32,31,253,31,12,31,213,31,38,31,38,30,156,31,165,31,129,31,43,31,250,31,194,31,194,30,194,29,192,31,131,31,89,31,89,30,89,31,161,31,187,31,78,31,177,31,118,31,71,31,159,31,114,31,241,31,130,31,152,31,187,31,125,31,230,31,174,31,73,31,49,31,87,31,119,31,206,31,129,31,243,31,243,30,9,31,9,30,216,31,162,31,87,31,114,31,114,30,202,31,196,31,69,31,227,31,227,30,80,31,80,30,94,31,158,31,158,30,187,31,187,30,212,31,129,31,129,30,161,31,134,31,12,31,12,30,4,31,16,31,110,31,47,31,66,31,252,31,252,30,149,31,11,31,163,31,163,30,253,31,93,31,185,31,185,30,156,31,218,31,212,31,43,31,92,31,59,31,59,30,9,31,35,31,140,31,238,31,238,30,238,29,106,31,237,31,140,31,80,31,80,30,26,31,206,31,19,31,139,31,139,30,55,31,255,31,11,31,104,31,172,31,208,31,156,31,203,31,1,31,121,31,191,31,177,31,115,31,219,31,132,31,203,31,203,30,223,31,223,30,151,31,247,31,247,30,170,31,107,31,62,31,144,31,142,31,37,31,137,31,160,31,11,31,11,30,35,31,66,31,66,30,243,31,243,30,174,31,167,31,120,31,120,30,114,31,20,31,194,31,169,31,192,31,192,30,222,31,222,30,108,31,108,30,108,29,83,31,47,31,243,31,34,31,117,31,195,31,107,31,72,31,53,31,73,31,119,31,133,31,143,31,45,31,162,31,88,31,128,31,159,31,159,30,224,31,31,31,175,31,247,31,23,31,31,31,31,30,241,31,44,31,44,30,211,31,128,31,127,31,127,30,99,31,66,31,60,31,204,31,82,31,178,31,217,31,217,30,173,31,115,31,14,31,103,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
