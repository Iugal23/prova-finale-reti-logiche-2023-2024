-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 293;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,0,0,2,0,165,0,0,0,21,0,1,0,42,0,199,0,77,0,233,0,241,0,0,0,77,0,89,0,180,0,187,0,0,0,47,0,47,0,0,0,97,0,249,0,0,0,116,0,177,0,56,0,0,0,254,0,0,0,141,0,177,0,55,0,198,0,0,0,76,0,71,0,107,0,141,0,0,0,0,0,197,0,0,0,186,0,0,0,62,0,163,0,0,0,242,0,103,0,0,0,20,0,25,0,0,0,0,0,94,0,254,0,0,0,72,0,207,0,151,0,220,0,64,0,12,0,222,0,0,0,214,0,101,0,147,0,0,0,241,0,102,0,197,0,0,0,0,0,129,0,154,0,211,0,91,0,42,0,0,0,0,0,108,0,121,0,0,0,212,0,56,0,69,0,25,0,67,0,184,0,199,0,247,0,185,0,126,0,104,0,58,0,0,0,133,0,0,0,86,0,0,0,0,0,250,0,60,0,6,0,150,0,15,0,73,0,0,0,172,0,0,0,56,0,207,0,136,0,141,0,193,0,43,0,0,0,197,0,113,0,0,0,97,0,0,0,107,0,36,0,85,0,0,0,98,0,0,0,36,0,90,0,239,0,151,0,26,0,134,0,48,0,45,0,0,0,40,0,252,0,0,0,7,0,245,0,177,0,0,0,86,0,40,0,0,0,0,0,22,0,114,0,58,0,0,0,95,0,210,0,166,0,0,0,0,0,190,0,144,0,152,0,62,0,14,0,59,0,0,0,214,0,86,0,112,0,0,0,0,0,57,0,126,0,198,0,3,0,0,0,65,0,147,0,28,0,0,0,192,0,6,0,170,0,52,0,201,0,0,0,0,0,151,0,19,0,54,0,0,0,173,0,0,0,0,0,23,0,182,0,93,0,243,0,240,0,217,0,189,0,0,0,118,0,0,0,215,0,0,0,92,0,95,0,0,0,53,0,0,0,109,0,40,0,179,0,195,0,36,0,0,0,198,0,0,0,0,0,33,0,24,0,9,0,0,0,117,0,151,0,179,0,71,0,133,0,26,0,177,0,153,0,44,0,109,0,58,0,0,0,228,0,94,0,88,0,0,0,9,0,68,0,95,0,229,0,4,0,193,0,254,0,0,0,167,0,0,0,252,0,9,0,226,0,184,0,204,0,212,0,74,0,95,0,50,0,4,0,16,0,121,0,203,0,0,0,0,0,109,0,220,0,15,0,61,0,171,0,35,0,0,0,107,0,203,0,139,0,123,0,142,0,171,0,0,0,153,0,13,0,247,0,252,0,98,0,100,0,175,0,12,0,101,0,7,0,240,0,197,0,84,0,107,0);
signal scenario_full  : scenario_type := (214,31,214,30,2,31,165,31,165,30,21,31,1,31,42,31,199,31,77,31,233,31,241,31,241,30,77,31,89,31,180,31,187,31,187,30,47,31,47,31,47,30,97,31,249,31,249,30,116,31,177,31,56,31,56,30,254,31,254,30,141,31,177,31,55,31,198,31,198,30,76,31,71,31,107,31,141,31,141,30,141,29,197,31,197,30,186,31,186,30,62,31,163,31,163,30,242,31,103,31,103,30,20,31,25,31,25,30,25,29,94,31,254,31,254,30,72,31,207,31,151,31,220,31,64,31,12,31,222,31,222,30,214,31,101,31,147,31,147,30,241,31,102,31,197,31,197,30,197,29,129,31,154,31,211,31,91,31,42,31,42,30,42,29,108,31,121,31,121,30,212,31,56,31,69,31,25,31,67,31,184,31,199,31,247,31,185,31,126,31,104,31,58,31,58,30,133,31,133,30,86,31,86,30,86,29,250,31,60,31,6,31,150,31,15,31,73,31,73,30,172,31,172,30,56,31,207,31,136,31,141,31,193,31,43,31,43,30,197,31,113,31,113,30,97,31,97,30,107,31,36,31,85,31,85,30,98,31,98,30,36,31,90,31,239,31,151,31,26,31,134,31,48,31,45,31,45,30,40,31,252,31,252,30,7,31,245,31,177,31,177,30,86,31,40,31,40,30,40,29,22,31,114,31,58,31,58,30,95,31,210,31,166,31,166,30,166,29,190,31,144,31,152,31,62,31,14,31,59,31,59,30,214,31,86,31,112,31,112,30,112,29,57,31,126,31,198,31,3,31,3,30,65,31,147,31,28,31,28,30,192,31,6,31,170,31,52,31,201,31,201,30,201,29,151,31,19,31,54,31,54,30,173,31,173,30,173,29,23,31,182,31,93,31,243,31,240,31,217,31,189,31,189,30,118,31,118,30,215,31,215,30,92,31,95,31,95,30,53,31,53,30,109,31,40,31,179,31,195,31,36,31,36,30,198,31,198,30,198,29,33,31,24,31,9,31,9,30,117,31,151,31,179,31,71,31,133,31,26,31,177,31,153,31,44,31,109,31,58,31,58,30,228,31,94,31,88,31,88,30,9,31,68,31,95,31,229,31,4,31,193,31,254,31,254,30,167,31,167,30,252,31,9,31,226,31,184,31,204,31,212,31,74,31,95,31,50,31,4,31,16,31,121,31,203,31,203,30,203,29,109,31,220,31,15,31,61,31,171,31,35,31,35,30,107,31,203,31,139,31,123,31,142,31,171,31,171,30,153,31,13,31,247,31,252,31,98,31,100,31,175,31,12,31,101,31,7,31,240,31,197,31,84,31,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
