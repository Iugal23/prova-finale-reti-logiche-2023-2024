-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 510;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,237,0,131,0,0,0,155,0,136,0,0,0,0,0,0,0,42,0,185,0,0,0,93,0,211,0,0,0,0,0,113,0,154,0,0,0,0,0,211,0,252,0,0,0,226,0,237,0,165,0,0,0,214,0,211,0,0,0,0,0,59,0,83,0,249,0,157,0,96,0,255,0,86,0,58,0,30,0,211,0,211,0,138,0,0,0,188,0,129,0,45,0,108,0,0,0,130,0,148,0,148,0,36,0,0,0,66,0,0,0,0,0,104,0,170,0,227,0,37,0,0,0,0,0,0,0,137,0,17,0,184,0,197,0,36,0,91,0,169,0,128,0,0,0,102,0,203,0,118,0,0,0,154,0,146,0,226,0,117,0,0,0,238,0,43,0,153,0,215,0,69,0,252,0,0,0,110,0,105,0,83,0,0,0,254,0,0,0,164,0,69,0,121,0,30,0,136,0,127,0,221,0,96,0,132,0,165,0,0,0,0,0,0,0,65,0,225,0,4,0,0,0,152,0,53,0,62,0,169,0,155,0,231,0,237,0,252,0,0,0,201,0,172,0,115,0,253,0,0,0,91,0,37,0,9,0,0,0,0,0,86,0,57,0,172,0,0,0,93,0,0,0,68,0,230,0,0,0,0,0,96,0,116,0,0,0,254,0,0,0,155,0,0,0,215,0,0,0,97,0,83,0,29,0,138,0,196,0,129,0,182,0,152,0,0,0,245,0,0,0,123,0,105,0,235,0,0,0,133,0,0,0,75,0,135,0,104,0,130,0,146,0,67,0,0,0,223,0,26,0,242,0,168,0,94,0,0,0,142,0,248,0,40,0,61,0,133,0,246,0,43,0,128,0,158,0,218,0,166,0,248,0,10,0,113,0,132,0,0,0,0,0,0,0,225,0,130,0,170,0,156,0,17,0,197,0,250,0,6,0,228,0,228,0,210,0,65,0,190,0,71,0,154,0,219,0,241,0,60,0,228,0,51,0,40,0,221,0,177,0,223,0,122,0,67,0,0,0,0,0,204,0,231,0,128,0,116,0,234,0,33,0,104,0,0,0,0,0,218,0,42,0,70,0,30,0,0,0,3,0,185,0,167,0,141,0,0,0,251,0,233,0,0,0,116,0,51,0,146,0,147,0,132,0,199,0,0,0,0,0,0,0,6,0,0,0,123,0,84,0,47,0,217,0,144,0,103,0,151,0,133,0,229,0,137,0,0,0,255,0,215,0,151,0,169,0,216,0,89,0,0,0,94,0,0,0,235,0,0,0,133,0,0,0,190,0,30,0,0,0,228,0,0,0,80,0,51,0,40,0,98,0,151,0,101,0,60,0,37,0,27,0,189,0,0,0,199,0,112,0,35,0,240,0,0,0,213,0,97,0,211,0,167,0,172,0,0,0,244,0,92,0,124,0,152,0,190,0,180,0,8,0,137,0,53,0,80,0,4,0,189,0,217,0,0,0,103,0,23,0,45,0,0,0,245,0,127,0,214,0,58,0,245,0,0,0,112,0,200,0,37,0,0,0,248,0,0,0,119,0,121,0,0,0,182,0,241,0,226,0,8,0,158,0,138,0,0,0,192,0,65,0,208,0,228,0,247,0,0,0,2,0,193,0,162,0,19,0,97,0,122,0,179,0,17,0,44,0,22,0,142,0,184,0,113,0,130,0,184,0,165,0,39,0,243,0,223,0,63,0,162,0,197,0,214,0,215,0,97,0,247,0,207,0,62,0,105,0,48,0,97,0,75,0,119,0,66,0,103,0,45,0,0,0,120,0,0,0,0,0,160,0,162,0,153,0,113,0,75,0,122,0,0,0,213,0,3,0,92,0,12,0,64,0,140,0,219,0,209,0,0,0,53,0,197,0,85,0,96,0,131,0,34,0,127,0,216,0,0,0,190,0,26,0,67,0,246,0,83,0,0,0,158,0,9,0,162,0,184,0,234,0,205,0,86,0,218,0,92,0,180,0,0,0,0,0,0,0,93,0,205,0,0,0,200,0,0,0,0,0,222,0,140,0,0,0,28,0,33,0,170,0,59,0,0,0,245,0,198,0,0,0,108,0,120,0,10,0,36,0,122,0,57,0,89,0,108,0,0,0,168,0,17,0,47,0,26,0,183,0,133,0,38,0,0,0,172,0,223,0,189,0,154,0,172,0,32,0,205,0,0,0,126,0,43,0,213,0,0,0,192,0,80,0,142,0,7,0,139,0,0,0,248,0,65,0,193,0,57,0,219,0,227,0,29,0,110,0,36,0,130,0,32,0,90,0,209,0,82,0,70,0,0,0,20,0,0,0);
signal scenario_full  : scenario_type := (154,31,237,31,131,31,131,30,155,31,136,31,136,30,136,29,136,28,42,31,185,31,185,30,93,31,211,31,211,30,211,29,113,31,154,31,154,30,154,29,211,31,252,31,252,30,226,31,237,31,165,31,165,30,214,31,211,31,211,30,211,29,59,31,83,31,249,31,157,31,96,31,255,31,86,31,58,31,30,31,211,31,211,31,138,31,138,30,188,31,129,31,45,31,108,31,108,30,130,31,148,31,148,31,36,31,36,30,66,31,66,30,66,29,104,31,170,31,227,31,37,31,37,30,37,29,37,28,137,31,17,31,184,31,197,31,36,31,91,31,169,31,128,31,128,30,102,31,203,31,118,31,118,30,154,31,146,31,226,31,117,31,117,30,238,31,43,31,153,31,215,31,69,31,252,31,252,30,110,31,105,31,83,31,83,30,254,31,254,30,164,31,69,31,121,31,30,31,136,31,127,31,221,31,96,31,132,31,165,31,165,30,165,29,165,28,65,31,225,31,4,31,4,30,152,31,53,31,62,31,169,31,155,31,231,31,237,31,252,31,252,30,201,31,172,31,115,31,253,31,253,30,91,31,37,31,9,31,9,30,9,29,86,31,57,31,172,31,172,30,93,31,93,30,68,31,230,31,230,30,230,29,96,31,116,31,116,30,254,31,254,30,155,31,155,30,215,31,215,30,97,31,83,31,29,31,138,31,196,31,129,31,182,31,152,31,152,30,245,31,245,30,123,31,105,31,235,31,235,30,133,31,133,30,75,31,135,31,104,31,130,31,146,31,67,31,67,30,223,31,26,31,242,31,168,31,94,31,94,30,142,31,248,31,40,31,61,31,133,31,246,31,43,31,128,31,158,31,218,31,166,31,248,31,10,31,113,31,132,31,132,30,132,29,132,28,225,31,130,31,170,31,156,31,17,31,197,31,250,31,6,31,228,31,228,31,210,31,65,31,190,31,71,31,154,31,219,31,241,31,60,31,228,31,51,31,40,31,221,31,177,31,223,31,122,31,67,31,67,30,67,29,204,31,231,31,128,31,116,31,234,31,33,31,104,31,104,30,104,29,218,31,42,31,70,31,30,31,30,30,3,31,185,31,167,31,141,31,141,30,251,31,233,31,233,30,116,31,51,31,146,31,147,31,132,31,199,31,199,30,199,29,199,28,6,31,6,30,123,31,84,31,47,31,217,31,144,31,103,31,151,31,133,31,229,31,137,31,137,30,255,31,215,31,151,31,169,31,216,31,89,31,89,30,94,31,94,30,235,31,235,30,133,31,133,30,190,31,30,31,30,30,228,31,228,30,80,31,51,31,40,31,98,31,151,31,101,31,60,31,37,31,27,31,189,31,189,30,199,31,112,31,35,31,240,31,240,30,213,31,97,31,211,31,167,31,172,31,172,30,244,31,92,31,124,31,152,31,190,31,180,31,8,31,137,31,53,31,80,31,4,31,189,31,217,31,217,30,103,31,23,31,45,31,45,30,245,31,127,31,214,31,58,31,245,31,245,30,112,31,200,31,37,31,37,30,248,31,248,30,119,31,121,31,121,30,182,31,241,31,226,31,8,31,158,31,138,31,138,30,192,31,65,31,208,31,228,31,247,31,247,30,2,31,193,31,162,31,19,31,97,31,122,31,179,31,17,31,44,31,22,31,142,31,184,31,113,31,130,31,184,31,165,31,39,31,243,31,223,31,63,31,162,31,197,31,214,31,215,31,97,31,247,31,207,31,62,31,105,31,48,31,97,31,75,31,119,31,66,31,103,31,45,31,45,30,120,31,120,30,120,29,160,31,162,31,153,31,113,31,75,31,122,31,122,30,213,31,3,31,92,31,12,31,64,31,140,31,219,31,209,31,209,30,53,31,197,31,85,31,96,31,131,31,34,31,127,31,216,31,216,30,190,31,26,31,67,31,246,31,83,31,83,30,158,31,9,31,162,31,184,31,234,31,205,31,86,31,218,31,92,31,180,31,180,30,180,29,180,28,93,31,205,31,205,30,200,31,200,30,200,29,222,31,140,31,140,30,28,31,33,31,170,31,59,31,59,30,245,31,198,31,198,30,108,31,120,31,10,31,36,31,122,31,57,31,89,31,108,31,108,30,168,31,17,31,47,31,26,31,183,31,133,31,38,31,38,30,172,31,223,31,189,31,154,31,172,31,32,31,205,31,205,30,126,31,43,31,213,31,213,30,192,31,80,31,142,31,7,31,139,31,139,30,248,31,65,31,193,31,57,31,219,31,227,31,29,31,110,31,36,31,130,31,32,31,90,31,209,31,82,31,70,31,70,30,20,31,20,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
