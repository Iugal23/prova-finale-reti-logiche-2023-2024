-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_564 is
end project_tb_564;

architecture project_tb_arch_564 of project_tb_564 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 517;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,95,0,100,0,84,0,150,0,146,0,140,0,168,0,167,0,0,0,88,0,58,0,184,0,125,0,152,0,214,0,0,0,80,0,67,0,62,0,0,0,170,0,221,0,49,0,0,0,68,0,150,0,87,0,242,0,113,0,142,0,68,0,249,0,169,0,213,0,211,0,175,0,161,0,0,0,50,0,49,0,113,0,111,0,0,0,204,0,173,0,0,0,57,0,238,0,0,0,0,0,144,0,212,0,140,0,250,0,63,0,26,0,70,0,222,0,138,0,219,0,44,0,0,0,186,0,0,0,74,0,63,0,22,0,43,0,198,0,75,0,0,0,0,0,214,0,70,0,79,0,44,0,220,0,244,0,70,0,122,0,1,0,158,0,0,0,254,0,0,0,161,0,0,0,0,0,193,0,17,0,82,0,2,0,125,0,89,0,95,0,33,0,195,0,242,0,17,0,85,0,42,0,53,0,48,0,0,0,0,0,140,0,165,0,201,0,68,0,169,0,146,0,109,0,219,0,0,0,35,0,253,0,219,0,86,0,88,0,248,0,31,0,3,0,99,0,19,0,207,0,155,0,76,0,228,0,96,0,73,0,168,0,66,0,224,0,147,0,235,0,237,0,51,0,18,0,41,0,51,0,189,0,0,0,37,0,198,0,90,0,55,0,213,0,49,0,239,0,40,0,101,0,96,0,236,0,110,0,249,0,13,0,13,0,55,0,164,0,188,0,236,0,97,0,3,0,89,0,0,0,198,0,136,0,190,0,62,0,250,0,84,0,72,0,102,0,129,0,237,0,115,0,159,0,159,0,249,0,236,0,41,0,0,0,32,0,104,0,162,0,34,0,224,0,38,0,227,0,0,0,84,0,225,0,179,0,227,0,184,0,142,0,111,0,253,0,152,0,98,0,0,0,67,0,95,0,84,0,0,0,134,0,0,0,193,0,0,0,134,0,0,0,173,0,237,0,0,0,166,0,118,0,61,0,214,0,229,0,18,0,0,0,110,0,162,0,189,0,142,0,37,0,118,0,148,0,189,0,47,0,3,0,0,0,120,0,189,0,32,0,124,0,27,0,9,0,0,0,39,0,227,0,249,0,194,0,97,0,139,0,227,0,14,0,218,0,192,0,216,0,59,0,128,0,29,0,0,0,126,0,134,0,250,0,112,0,193,0,27,0,183,0,0,0,216,0,239,0,0,0,82,0,205,0,229,0,0,0,39,0,252,0,17,0,246,0,135,0,0,0,91,0,205,0,0,0,22,0,23,0,83,0,253,0,45,0,0,0,11,0,66,0,229,0,96,0,0,0,69,0,149,0,252,0,6,0,189,0,104,0,116,0,0,0,0,0,80,0,163,0,69,0,0,0,223,0,233,0,102,0,0,0,0,0,228,0,192,0,0,0,37,0,0,0,60,0,233,0,157,0,98,0,96,0,0,0,132,0,133,0,32,0,193,0,86,0,1,0,0,0,252,0,56,0,226,0,128,0,0,0,230,0,143,0,169,0,139,0,164,0,54,0,0,0,21,0,166,0,32,0,246,0,238,0,38,0,114,0,165,0,190,0,0,0,213,0,39,0,151,0,0,0,0,0,81,0,0,0,0,0,204,0,112,0,135,0,35,0,0,0,0,0,107,0,95,0,155,0,124,0,189,0,215,0,0,0,217,0,241,0,40,0,0,0,0,0,234,0,208,0,40,0,0,0,72,0,141,0,223,0,101,0,59,0,218,0,0,0,226,0,91,0,0,0,37,0,199,0,138,0,0,0,21,0,222,0,212,0,218,0,100,0,190,0,215,0,109,0,0,0,23,0,118,0,185,0,186,0,0,0,103,0,0,0,0,0,119,0,232,0,0,0,108,0,187,0,31,0,80,0,0,0,203,0,123,0,253,0,117,0,0,0,16,0,218,0,186,0,71,0,178,0,63,0,0,0,0,0,154,0,168,0,137,0,191,0,0,0,102,0,162,0,0,0,45,0,0,0,70,0,86,0,170,0,157,0,0,0,134,0,120,0,84,0,71,0,191,0,154,0,137,0,97,0,250,0,121,0,0,0,197,0,40,0,210,0,126,0,62,0,140,0,248,0,99,0,0,0,69,0,0,0,45,0,48,0,0,0,95,0,0,0,253,0,0,0,3,0,0,0,178,0,197,0,31,0,167,0,47,0,0,0,145,0,0,0,163,0,0,0,139,0,74,0,125,0,168,0,123,0,162,0,219,0,106,0,137,0,104,0,209,0,0,0,88,0,106,0,200,0,83,0,0,0,0,0,0,0,49,0,175,0,0,0,234,0,0,0,213,0,239,0,185,0,211,0,61,0,108,0,118,0);
signal scenario_full  : scenario_type := (35,31,95,31,100,31,84,31,150,31,146,31,140,31,168,31,167,31,167,30,88,31,58,31,184,31,125,31,152,31,214,31,214,30,80,31,67,31,62,31,62,30,170,31,221,31,49,31,49,30,68,31,150,31,87,31,242,31,113,31,142,31,68,31,249,31,169,31,213,31,211,31,175,31,161,31,161,30,50,31,49,31,113,31,111,31,111,30,204,31,173,31,173,30,57,31,238,31,238,30,238,29,144,31,212,31,140,31,250,31,63,31,26,31,70,31,222,31,138,31,219,31,44,31,44,30,186,31,186,30,74,31,63,31,22,31,43,31,198,31,75,31,75,30,75,29,214,31,70,31,79,31,44,31,220,31,244,31,70,31,122,31,1,31,158,31,158,30,254,31,254,30,161,31,161,30,161,29,193,31,17,31,82,31,2,31,125,31,89,31,95,31,33,31,195,31,242,31,17,31,85,31,42,31,53,31,48,31,48,30,48,29,140,31,165,31,201,31,68,31,169,31,146,31,109,31,219,31,219,30,35,31,253,31,219,31,86,31,88,31,248,31,31,31,3,31,99,31,19,31,207,31,155,31,76,31,228,31,96,31,73,31,168,31,66,31,224,31,147,31,235,31,237,31,51,31,18,31,41,31,51,31,189,31,189,30,37,31,198,31,90,31,55,31,213,31,49,31,239,31,40,31,101,31,96,31,236,31,110,31,249,31,13,31,13,31,55,31,164,31,188,31,236,31,97,31,3,31,89,31,89,30,198,31,136,31,190,31,62,31,250,31,84,31,72,31,102,31,129,31,237,31,115,31,159,31,159,31,249,31,236,31,41,31,41,30,32,31,104,31,162,31,34,31,224,31,38,31,227,31,227,30,84,31,225,31,179,31,227,31,184,31,142,31,111,31,253,31,152,31,98,31,98,30,67,31,95,31,84,31,84,30,134,31,134,30,193,31,193,30,134,31,134,30,173,31,237,31,237,30,166,31,118,31,61,31,214,31,229,31,18,31,18,30,110,31,162,31,189,31,142,31,37,31,118,31,148,31,189,31,47,31,3,31,3,30,120,31,189,31,32,31,124,31,27,31,9,31,9,30,39,31,227,31,249,31,194,31,97,31,139,31,227,31,14,31,218,31,192,31,216,31,59,31,128,31,29,31,29,30,126,31,134,31,250,31,112,31,193,31,27,31,183,31,183,30,216,31,239,31,239,30,82,31,205,31,229,31,229,30,39,31,252,31,17,31,246,31,135,31,135,30,91,31,205,31,205,30,22,31,23,31,83,31,253,31,45,31,45,30,11,31,66,31,229,31,96,31,96,30,69,31,149,31,252,31,6,31,189,31,104,31,116,31,116,30,116,29,80,31,163,31,69,31,69,30,223,31,233,31,102,31,102,30,102,29,228,31,192,31,192,30,37,31,37,30,60,31,233,31,157,31,98,31,96,31,96,30,132,31,133,31,32,31,193,31,86,31,1,31,1,30,252,31,56,31,226,31,128,31,128,30,230,31,143,31,169,31,139,31,164,31,54,31,54,30,21,31,166,31,32,31,246,31,238,31,38,31,114,31,165,31,190,31,190,30,213,31,39,31,151,31,151,30,151,29,81,31,81,30,81,29,204,31,112,31,135,31,35,31,35,30,35,29,107,31,95,31,155,31,124,31,189,31,215,31,215,30,217,31,241,31,40,31,40,30,40,29,234,31,208,31,40,31,40,30,72,31,141,31,223,31,101,31,59,31,218,31,218,30,226,31,91,31,91,30,37,31,199,31,138,31,138,30,21,31,222,31,212,31,218,31,100,31,190,31,215,31,109,31,109,30,23,31,118,31,185,31,186,31,186,30,103,31,103,30,103,29,119,31,232,31,232,30,108,31,187,31,31,31,80,31,80,30,203,31,123,31,253,31,117,31,117,30,16,31,218,31,186,31,71,31,178,31,63,31,63,30,63,29,154,31,168,31,137,31,191,31,191,30,102,31,162,31,162,30,45,31,45,30,70,31,86,31,170,31,157,31,157,30,134,31,120,31,84,31,71,31,191,31,154,31,137,31,97,31,250,31,121,31,121,30,197,31,40,31,210,31,126,31,62,31,140,31,248,31,99,31,99,30,69,31,69,30,45,31,48,31,48,30,95,31,95,30,253,31,253,30,3,31,3,30,178,31,197,31,31,31,167,31,47,31,47,30,145,31,145,30,163,31,163,30,139,31,74,31,125,31,168,31,123,31,162,31,219,31,106,31,137,31,104,31,209,31,209,30,88,31,106,31,200,31,83,31,83,30,83,29,83,28,49,31,175,31,175,30,234,31,234,30,213,31,239,31,185,31,211,31,61,31,108,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
