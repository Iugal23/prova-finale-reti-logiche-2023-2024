-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 671;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (163,0,0,0,240,0,57,0,115,0,155,0,196,0,5,0,192,0,161,0,119,0,64,0,226,0,0,0,18,0,249,0,104,0,0,0,69,0,94,0,0,0,0,0,154,0,71,0,185,0,118,0,153,0,190,0,223,0,98,0,0,0,0,0,0,0,0,0,45,0,115,0,77,0,0,0,0,0,231,0,90,0,133,0,135,0,219,0,221,0,155,0,0,0,213,0,0,0,159,0,0,0,174,0,0,0,31,0,137,0,140,0,55,0,202,0,24,0,95,0,38,0,12,0,179,0,69,0,243,0,221,0,205,0,75,0,233,0,226,0,14,0,125,0,67,0,49,0,130,0,36,0,90,0,85,0,201,0,0,0,5,0,218,0,241,0,215,0,193,0,231,0,83,0,242,0,53,0,50,0,202,0,0,0,203,0,225,0,27,0,179,0,0,0,84,0,99,0,27,0,139,0,0,0,0,0,109,0,224,0,233,0,210,0,29,0,223,0,92,0,37,0,188,0,27,0,29,0,44,0,0,0,132,0,0,0,0,0,0,0,137,0,0,0,207,0,0,0,0,0,174,0,109,0,223,0,179,0,78,0,74,0,49,0,162,0,75,0,122,0,253,0,196,0,188,0,100,0,0,0,135,0,176,0,0,0,30,0,0,0,0,0,66,0,10,0,182,0,106,0,216,0,111,0,188,0,0,0,52,0,245,0,203,0,10,0,114,0,184,0,157,0,31,0,0,0,88,0,66,0,0,0,29,0,128,0,0,0,128,0,0,0,31,0,200,0,102,0,157,0,97,0,191,0,172,0,0,0,60,0,75,0,137,0,141,0,125,0,252,0,165,0,0,0,111,0,9,0,0,0,225,0,203,0,199,0,2,0,85,0,217,0,0,0,186,0,0,0,230,0,160,0,114,0,0,0,0,0,35,0,167,0,0,0,0,0,67,0,0,0,163,0,178,0,121,0,0,0,219,0,148,0,96,0,0,0,186,0,54,0,70,0,207,0,228,0,0,0,152,0,0,0,0,0,0,0,0,0,129,0,107,0,131,0,209,0,237,0,0,0,50,0,0,0,44,0,200,0,181,0,75,0,0,0,126,0,57,0,142,0,140,0,178,0,231,0,226,0,172,0,219,0,95,0,6,0,23,0,149,0,0,0,17,0,215,0,119,0,0,0,15,0,191,0,54,0,237,0,96,0,0,0,209,0,93,0,0,0,74,0,0,0,0,0,115,0,0,0,135,0,0,0,0,0,193,0,12,0,147,0,103,0,25,0,206,0,4,0,0,0,140,0,143,0,50,0,194,0,214,0,191,0,75,0,77,0,251,0,0,0,2,0,231,0,90,0,30,0,0,0,11,0,100,0,30,0,153,0,172,0,37,0,101,0,55,0,0,0,6,0,47,0,141,0,189,0,227,0,0,0,240,0,73,0,137,0,201,0,248,0,225,0,167,0,87,0,0,0,196,0,249,0,23,0,184,0,135,0,132,0,0,0,0,0,248,0,142,0,5,0,116,0,161,0,90,0,0,0,21,0,163,0,252,0,130,0,110,0,0,0,140,0,235,0,49,0,140,0,46,0,195,0,0,0,35,0,208,0,129,0,195,0,188,0,246,0,185,0,33,0,87,0,163,0,240,0,239,0,0,0,201,0,158,0,238,0,76,0,65,0,0,0,17,0,73,0,16,0,226,0,220,0,57,0,90,0,107,0,0,0,213,0,132,0,141,0,182,0,252,0,187,0,85,0,0,0,182,0,28,0,126,0,51,0,122,0,212,0,0,0,0,0,65,0,226,0,96,0,225,0,151,0,0,0,0,0,46,0,145,0,130,0,176,0,0,0,69,0,153,0,227,0,250,0,135,0,121,0,0,0,25,0,235,0,121,0,246,0,175,0,122,0,192,0,138,0,90,0,8,0,238,0,38,0,6,0,19,0,236,0,33,0,64,0,179,0,0,0,199,0,0,0,40,0,5,0,177,0,78,0,226,0,0,0,34,0,16,0,0,0,94,0,0,0,164,0,0,0,253,0,100,0,0,0,140,0,134,0,125,0,11,0,204,0,155,0,121,0,0,0,194,0,157,0,2,0,118,0,212,0,62,0,0,0,162,0,21,0,252,0,210,0,122,0,152,0,165,0,40,0,39,0,3,0,205,0,173,0,182,0,181,0,0,0,86,0,59,0,94,0,181,0,109,0,0,0,106,0,8,0,203,0,235,0,225,0,193,0,145,0,153,0,0,0,32,0,37,0,171,0,42,0,161,0,109,0,79,0,184,0,0,0,23,0,247,0,0,0,0,0,183,0,0,0,0,0,0,0,224,0,96,0,238,0,153,0,167,0,218,0,178,0,50,0,128,0,36,0,196,0,208,0,89,0,63,0,61,0,97,0,0,0,244,0,161,0,45,0,137,0,25,0,13,0,134,0,134,0,241,0,131,0,185,0,0,0,0,0,211,0,175,0,82,0,179,0,0,0,201,0,95,0,0,0,206,0,0,0,19,0,0,0,31,0,107,0,70,0,0,0,2,0,120,0,83,0,46,0,143,0,73,0,204,0,107,0,0,0,0,0,55,0,145,0,0,0,0,0,0,0,42,0,133,0,0,0,202,0,0,0,0,0,0,0,0,0,0,0,120,0,0,0,240,0,195,0,245,0,31,0,184,0,228,0,0,0,229,0,0,0,0,0,119,0,128,0,155,0,196,0,32,0,174,0,0,0,0,0,55,0,246,0,227,0,105,0,89,0,110,0,69,0,0,0,44,0,137,0,221,0,74,0,135,0,42,0,144,0,154,0,0,0,203,0,50,0,11,0,91,0,172,0,15,0,208,0,157,0,249,0,219,0,0,0,189,0,134,0,195,0,182,0,11,0,0,0,199,0,0,0,0,0,76,0,21,0,0,0,177,0,132,0,41,0,228,0,4,0,77,0,119,0,78,0,0,0,140,0,245,0,144,0,125,0,0,0,93,0,74,0,0,0,247,0,130,0,255,0,79,0,223,0,109,0,118,0,48,0,242,0,209,0);
signal scenario_full  : scenario_type := (163,31,163,30,240,31,57,31,115,31,155,31,196,31,5,31,192,31,161,31,119,31,64,31,226,31,226,30,18,31,249,31,104,31,104,30,69,31,94,31,94,30,94,29,154,31,71,31,185,31,118,31,153,31,190,31,223,31,98,31,98,30,98,29,98,28,98,27,45,31,115,31,77,31,77,30,77,29,231,31,90,31,133,31,135,31,219,31,221,31,155,31,155,30,213,31,213,30,159,31,159,30,174,31,174,30,31,31,137,31,140,31,55,31,202,31,24,31,95,31,38,31,12,31,179,31,69,31,243,31,221,31,205,31,75,31,233,31,226,31,14,31,125,31,67,31,49,31,130,31,36,31,90,31,85,31,201,31,201,30,5,31,218,31,241,31,215,31,193,31,231,31,83,31,242,31,53,31,50,31,202,31,202,30,203,31,225,31,27,31,179,31,179,30,84,31,99,31,27,31,139,31,139,30,139,29,109,31,224,31,233,31,210,31,29,31,223,31,92,31,37,31,188,31,27,31,29,31,44,31,44,30,132,31,132,30,132,29,132,28,137,31,137,30,207,31,207,30,207,29,174,31,109,31,223,31,179,31,78,31,74,31,49,31,162,31,75,31,122,31,253,31,196,31,188,31,100,31,100,30,135,31,176,31,176,30,30,31,30,30,30,29,66,31,10,31,182,31,106,31,216,31,111,31,188,31,188,30,52,31,245,31,203,31,10,31,114,31,184,31,157,31,31,31,31,30,88,31,66,31,66,30,29,31,128,31,128,30,128,31,128,30,31,31,200,31,102,31,157,31,97,31,191,31,172,31,172,30,60,31,75,31,137,31,141,31,125,31,252,31,165,31,165,30,111,31,9,31,9,30,225,31,203,31,199,31,2,31,85,31,217,31,217,30,186,31,186,30,230,31,160,31,114,31,114,30,114,29,35,31,167,31,167,30,167,29,67,31,67,30,163,31,178,31,121,31,121,30,219,31,148,31,96,31,96,30,186,31,54,31,70,31,207,31,228,31,228,30,152,31,152,30,152,29,152,28,152,27,129,31,107,31,131,31,209,31,237,31,237,30,50,31,50,30,44,31,200,31,181,31,75,31,75,30,126,31,57,31,142,31,140,31,178,31,231,31,226,31,172,31,219,31,95,31,6,31,23,31,149,31,149,30,17,31,215,31,119,31,119,30,15,31,191,31,54,31,237,31,96,31,96,30,209,31,93,31,93,30,74,31,74,30,74,29,115,31,115,30,135,31,135,30,135,29,193,31,12,31,147,31,103,31,25,31,206,31,4,31,4,30,140,31,143,31,50,31,194,31,214,31,191,31,75,31,77,31,251,31,251,30,2,31,231,31,90,31,30,31,30,30,11,31,100,31,30,31,153,31,172,31,37,31,101,31,55,31,55,30,6,31,47,31,141,31,189,31,227,31,227,30,240,31,73,31,137,31,201,31,248,31,225,31,167,31,87,31,87,30,196,31,249,31,23,31,184,31,135,31,132,31,132,30,132,29,248,31,142,31,5,31,116,31,161,31,90,31,90,30,21,31,163,31,252,31,130,31,110,31,110,30,140,31,235,31,49,31,140,31,46,31,195,31,195,30,35,31,208,31,129,31,195,31,188,31,246,31,185,31,33,31,87,31,163,31,240,31,239,31,239,30,201,31,158,31,238,31,76,31,65,31,65,30,17,31,73,31,16,31,226,31,220,31,57,31,90,31,107,31,107,30,213,31,132,31,141,31,182,31,252,31,187,31,85,31,85,30,182,31,28,31,126,31,51,31,122,31,212,31,212,30,212,29,65,31,226,31,96,31,225,31,151,31,151,30,151,29,46,31,145,31,130,31,176,31,176,30,69,31,153,31,227,31,250,31,135,31,121,31,121,30,25,31,235,31,121,31,246,31,175,31,122,31,192,31,138,31,90,31,8,31,238,31,38,31,6,31,19,31,236,31,33,31,64,31,179,31,179,30,199,31,199,30,40,31,5,31,177,31,78,31,226,31,226,30,34,31,16,31,16,30,94,31,94,30,164,31,164,30,253,31,100,31,100,30,140,31,134,31,125,31,11,31,204,31,155,31,121,31,121,30,194,31,157,31,2,31,118,31,212,31,62,31,62,30,162,31,21,31,252,31,210,31,122,31,152,31,165,31,40,31,39,31,3,31,205,31,173,31,182,31,181,31,181,30,86,31,59,31,94,31,181,31,109,31,109,30,106,31,8,31,203,31,235,31,225,31,193,31,145,31,153,31,153,30,32,31,37,31,171,31,42,31,161,31,109,31,79,31,184,31,184,30,23,31,247,31,247,30,247,29,183,31,183,30,183,29,183,28,224,31,96,31,238,31,153,31,167,31,218,31,178,31,50,31,128,31,36,31,196,31,208,31,89,31,63,31,61,31,97,31,97,30,244,31,161,31,45,31,137,31,25,31,13,31,134,31,134,31,241,31,131,31,185,31,185,30,185,29,211,31,175,31,82,31,179,31,179,30,201,31,95,31,95,30,206,31,206,30,19,31,19,30,31,31,107,31,70,31,70,30,2,31,120,31,83,31,46,31,143,31,73,31,204,31,107,31,107,30,107,29,55,31,145,31,145,30,145,29,145,28,42,31,133,31,133,30,202,31,202,30,202,29,202,28,202,27,202,26,120,31,120,30,240,31,195,31,245,31,31,31,184,31,228,31,228,30,229,31,229,30,229,29,119,31,128,31,155,31,196,31,32,31,174,31,174,30,174,29,55,31,246,31,227,31,105,31,89,31,110,31,69,31,69,30,44,31,137,31,221,31,74,31,135,31,42,31,144,31,154,31,154,30,203,31,50,31,11,31,91,31,172,31,15,31,208,31,157,31,249,31,219,31,219,30,189,31,134,31,195,31,182,31,11,31,11,30,199,31,199,30,199,29,76,31,21,31,21,30,177,31,132,31,41,31,228,31,4,31,77,31,119,31,78,31,78,30,140,31,245,31,144,31,125,31,125,30,93,31,74,31,74,30,247,31,130,31,255,31,79,31,223,31,109,31,118,31,48,31,242,31,209,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
