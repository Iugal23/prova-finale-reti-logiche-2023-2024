-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_239 is
end project_tb_239;

architecture project_tb_arch_239 of project_tb_239 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 739;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (27,0,225,0,214,0,0,0,209,0,32,0,56,0,247,0,143,0,17,0,4,0,95,0,4,0,0,0,247,0,0,0,0,0,0,0,0,0,30,0,167,0,60,0,0,0,108,0,0,0,199,0,188,0,118,0,0,0,0,0,0,0,149,0,0,0,0,0,96,0,0,0,182,0,254,0,0,0,250,0,72,0,0,0,198,0,212,0,0,0,67,0,142,0,203,0,0,0,218,0,150,0,176,0,83,0,245,0,116,0,0,0,10,0,152,0,131,0,187,0,105,0,33,0,138,0,91,0,109,0,215,0,0,0,178,0,84,0,84,0,182,0,85,0,0,0,125,0,151,0,0,0,69,0,239,0,224,0,37,0,110,0,93,0,86,0,50,0,0,0,233,0,228,0,144,0,230,0,100,0,195,0,0,0,0,0,137,0,231,0,0,0,118,0,200,0,204,0,67,0,64,0,202,0,134,0,98,0,15,0,90,0,197,0,44,0,135,0,108,0,0,0,140,0,62,0,62,0,86,0,0,0,201,0,0,0,33,0,0,0,202,0,0,0,242,0,131,0,212,0,79,0,230,0,78,0,228,0,18,0,174,0,116,0,232,0,177,0,173,0,0,0,160,0,152,0,151,0,0,0,81,0,5,0,214,0,105,0,223,0,149,0,0,0,27,0,37,0,44,0,254,0,0,0,63,0,250,0,0,0,121,0,199,0,0,0,2,0,111,0,102,0,0,0,244,0,14,0,36,0,200,0,186,0,25,0,64,0,67,0,29,0,226,0,0,0,0,0,118,0,5,0,0,0,15,0,0,0,0,0,42,0,0,0,65,0,142,0,187,0,0,0,0,0,202,0,171,0,16,0,120,0,64,0,175,0,97,0,116,0,134,0,29,0,184,0,74,0,238,0,193,0,77,0,0,0,166,0,0,0,51,0,54,0,114,0,108,0,0,0,0,0,176,0,139,0,65,0,246,0,68,0,76,0,107,0,176,0,0,0,37,0,210,0,163,0,233,0,54,0,233,0,189,0,250,0,134,0,127,0,0,0,228,0,0,0,39,0,244,0,201,0,177,0,81,0,90,0,0,0,177,0,106,0,212,0,159,0,142,0,87,0,0,0,173,0,147,0,177,0,4,0,181,0,0,0,82,0,120,0,0,0,75,0,0,0,58,0,87,0,108,0,102,0,162,0,222,0,80,0,3,0,163,0,17,0,0,0,175,0,58,0,49,0,0,0,113,0,185,0,65,0,18,0,25,0,17,0,0,0,47,0,14,0,74,0,211,0,88,0,0,0,70,0,133,0,120,0,197,0,160,0,33,0,0,0,0,0,0,0,0,0,142,0,0,0,173,0,17,0,26,0,137,0,42,0,242,0,96,0,236,0,182,0,116,0,0,0,0,0,37,0,204,0,238,0,184,0,252,0,0,0,231,0,251,0,52,0,79,0,0,0,170,0,0,0,27,0,42,0,161,0,40,0,77,0,0,0,24,0,141,0,124,0,157,0,48,0,103,0,177,0,0,0,40,0,198,0,127,0,9,0,125,0,50,0,200,0,0,0,172,0,54,0,140,0,1,0,0,0,98,0,197,0,2,0,153,0,0,0,242,0,224,0,105,0,205,0,0,0,152,0,0,0,151,0,167,0,64,0,136,0,238,0,0,0,233,0,157,0,140,0,165,0,28,0,126,0,189,0,226,0,225,0,0,0,0,0,50,0,169,0,251,0,165,0,0,0,203,0,50,0,46,0,0,0,58,0,0,0,157,0,210,0,176,0,0,0,129,0,49,0,214,0,213,0,0,0,233,0,112,0,104,0,175,0,72,0,66,0,139,0,49,0,49,0,0,0,227,0,0,0,96,0,94,0,144,0,252,0,167,0,76,0,62,0,87,0,103,0,147,0,178,0,181,0,0,0,139,0,150,0,219,0,153,0,42,0,79,0,234,0,237,0,0,0,51,0,27,0,180,0,42,0,0,0,203,0,0,0,221,0,3,0,195,0,40,0,165,0,24,0,142,0,79,0,60,0,180,0,0,0,245,0,212,0,22,0,9,0,0,0,237,0,249,0,31,0,2,0,0,0,88,0,0,0,0,0,14,0,213,0,36,0,118,0,135,0,57,0,18,0,106,0,130,0,82,0,249,0,0,0,191,0,156,0,13,0,164,0,205,0,217,0,73,0,133,0,0,0,210,0,103,0,133,0,135,0,162,0,230,0,156,0,149,0,235,0,70,0,28,0,141,0,182,0,215,0,212,0,215,0,167,0,0,0,60,0,41,0,240,0,134,0,28,0,125,0,202,0,0,0,195,0,67,0,0,0,116,0,57,0,20,0,116,0,89,0,56,0,0,0,0,0,150,0,0,0,199,0,109,0,0,0,0,0,239,0,237,0,16,0,197,0,47,0,102,0,0,0,0,0,27,0,92,0,252,0,0,0,0,0,8,0,165,0,232,0,171,0,127,0,0,0,9,0,43,0,55,0,22,0,185,0,0,0,79,0,239,0,0,0,180,0,132,0,0,0,44,0,0,0,131,0,134,0,0,0,255,0,242,0,121,0,101,0,0,0,149,0,0,0,0,0,0,0,199,0,77,0,44,0,7,0,201,0,128,0,242,0,0,0,255,0,118,0,58,0,193,0,45,0,0,0,0,0,241,0,139,0,253,0,115,0,219,0,57,0,116,0,82,0,0,0,10,0,1,0,0,0,217,0,38,0,136,0,19,0,144,0,29,0,222,0,146,0,212,0,0,0,0,0,116,0,108,0,162,0,25,0,168,0,188,0,243,0,211,0,35,0,68,0,0,0,115,0,30,0,179,0,253,0,156,0,0,0,98,0,179,0,164,0,188,0,106,0,120,0,107,0,183,0,0,0,109,0,0,0,3,0,176,0,124,0,99,0,132,0,73,0,181,0,148,0,210,0,0,0,116,0,115,0,92,0,0,0,52,0,84,0,95,0,41,0,105,0,242,0,70,0,115,0,49,0,69,0,0,0,169,0,164,0,3,0,83,0,0,0,0,0,82,0,0,0,50,0,212,0,2,0,176,0,0,0,6,0,172,0,80,0,47,0,202,0,178,0,213,0,178,0,250,0,224,0,35,0,96,0,48,0,0,0,0,0,117,0,0,0,215,0,0,0,29,0,42,0,11,0,0,0,230,0,10,0,219,0,219,0,134,0,7,0,0,0,200,0,61,0,78,0,121,0,177,0,60,0,245,0,252,0,0,0,226,0,15,0,151,0,9,0,0,0,166,0,233,0,66,0,74,0,67,0,41,0,22,0,108,0,229,0,189,0,38,0,0,0,240,0,19,0,0,0,146,0,97,0,110,0);
signal scenario_full  : scenario_type := (27,31,225,31,214,31,214,30,209,31,32,31,56,31,247,31,143,31,17,31,4,31,95,31,4,31,4,30,247,31,247,30,247,29,247,28,247,27,30,31,167,31,60,31,60,30,108,31,108,30,199,31,188,31,118,31,118,30,118,29,118,28,149,31,149,30,149,29,96,31,96,30,182,31,254,31,254,30,250,31,72,31,72,30,198,31,212,31,212,30,67,31,142,31,203,31,203,30,218,31,150,31,176,31,83,31,245,31,116,31,116,30,10,31,152,31,131,31,187,31,105,31,33,31,138,31,91,31,109,31,215,31,215,30,178,31,84,31,84,31,182,31,85,31,85,30,125,31,151,31,151,30,69,31,239,31,224,31,37,31,110,31,93,31,86,31,50,31,50,30,233,31,228,31,144,31,230,31,100,31,195,31,195,30,195,29,137,31,231,31,231,30,118,31,200,31,204,31,67,31,64,31,202,31,134,31,98,31,15,31,90,31,197,31,44,31,135,31,108,31,108,30,140,31,62,31,62,31,86,31,86,30,201,31,201,30,33,31,33,30,202,31,202,30,242,31,131,31,212,31,79,31,230,31,78,31,228,31,18,31,174,31,116,31,232,31,177,31,173,31,173,30,160,31,152,31,151,31,151,30,81,31,5,31,214,31,105,31,223,31,149,31,149,30,27,31,37,31,44,31,254,31,254,30,63,31,250,31,250,30,121,31,199,31,199,30,2,31,111,31,102,31,102,30,244,31,14,31,36,31,200,31,186,31,25,31,64,31,67,31,29,31,226,31,226,30,226,29,118,31,5,31,5,30,15,31,15,30,15,29,42,31,42,30,65,31,142,31,187,31,187,30,187,29,202,31,171,31,16,31,120,31,64,31,175,31,97,31,116,31,134,31,29,31,184,31,74,31,238,31,193,31,77,31,77,30,166,31,166,30,51,31,54,31,114,31,108,31,108,30,108,29,176,31,139,31,65,31,246,31,68,31,76,31,107,31,176,31,176,30,37,31,210,31,163,31,233,31,54,31,233,31,189,31,250,31,134,31,127,31,127,30,228,31,228,30,39,31,244,31,201,31,177,31,81,31,90,31,90,30,177,31,106,31,212,31,159,31,142,31,87,31,87,30,173,31,147,31,177,31,4,31,181,31,181,30,82,31,120,31,120,30,75,31,75,30,58,31,87,31,108,31,102,31,162,31,222,31,80,31,3,31,163,31,17,31,17,30,175,31,58,31,49,31,49,30,113,31,185,31,65,31,18,31,25,31,17,31,17,30,47,31,14,31,74,31,211,31,88,31,88,30,70,31,133,31,120,31,197,31,160,31,33,31,33,30,33,29,33,28,33,27,142,31,142,30,173,31,17,31,26,31,137,31,42,31,242,31,96,31,236,31,182,31,116,31,116,30,116,29,37,31,204,31,238,31,184,31,252,31,252,30,231,31,251,31,52,31,79,31,79,30,170,31,170,30,27,31,42,31,161,31,40,31,77,31,77,30,24,31,141,31,124,31,157,31,48,31,103,31,177,31,177,30,40,31,198,31,127,31,9,31,125,31,50,31,200,31,200,30,172,31,54,31,140,31,1,31,1,30,98,31,197,31,2,31,153,31,153,30,242,31,224,31,105,31,205,31,205,30,152,31,152,30,151,31,167,31,64,31,136,31,238,31,238,30,233,31,157,31,140,31,165,31,28,31,126,31,189,31,226,31,225,31,225,30,225,29,50,31,169,31,251,31,165,31,165,30,203,31,50,31,46,31,46,30,58,31,58,30,157,31,210,31,176,31,176,30,129,31,49,31,214,31,213,31,213,30,233,31,112,31,104,31,175,31,72,31,66,31,139,31,49,31,49,31,49,30,227,31,227,30,96,31,94,31,144,31,252,31,167,31,76,31,62,31,87,31,103,31,147,31,178,31,181,31,181,30,139,31,150,31,219,31,153,31,42,31,79,31,234,31,237,31,237,30,51,31,27,31,180,31,42,31,42,30,203,31,203,30,221,31,3,31,195,31,40,31,165,31,24,31,142,31,79,31,60,31,180,31,180,30,245,31,212,31,22,31,9,31,9,30,237,31,249,31,31,31,2,31,2,30,88,31,88,30,88,29,14,31,213,31,36,31,118,31,135,31,57,31,18,31,106,31,130,31,82,31,249,31,249,30,191,31,156,31,13,31,164,31,205,31,217,31,73,31,133,31,133,30,210,31,103,31,133,31,135,31,162,31,230,31,156,31,149,31,235,31,70,31,28,31,141,31,182,31,215,31,212,31,215,31,167,31,167,30,60,31,41,31,240,31,134,31,28,31,125,31,202,31,202,30,195,31,67,31,67,30,116,31,57,31,20,31,116,31,89,31,56,31,56,30,56,29,150,31,150,30,199,31,109,31,109,30,109,29,239,31,237,31,16,31,197,31,47,31,102,31,102,30,102,29,27,31,92,31,252,31,252,30,252,29,8,31,165,31,232,31,171,31,127,31,127,30,9,31,43,31,55,31,22,31,185,31,185,30,79,31,239,31,239,30,180,31,132,31,132,30,44,31,44,30,131,31,134,31,134,30,255,31,242,31,121,31,101,31,101,30,149,31,149,30,149,29,149,28,199,31,77,31,44,31,7,31,201,31,128,31,242,31,242,30,255,31,118,31,58,31,193,31,45,31,45,30,45,29,241,31,139,31,253,31,115,31,219,31,57,31,116,31,82,31,82,30,10,31,1,31,1,30,217,31,38,31,136,31,19,31,144,31,29,31,222,31,146,31,212,31,212,30,212,29,116,31,108,31,162,31,25,31,168,31,188,31,243,31,211,31,35,31,68,31,68,30,115,31,30,31,179,31,253,31,156,31,156,30,98,31,179,31,164,31,188,31,106,31,120,31,107,31,183,31,183,30,109,31,109,30,3,31,176,31,124,31,99,31,132,31,73,31,181,31,148,31,210,31,210,30,116,31,115,31,92,31,92,30,52,31,84,31,95,31,41,31,105,31,242,31,70,31,115,31,49,31,69,31,69,30,169,31,164,31,3,31,83,31,83,30,83,29,82,31,82,30,50,31,212,31,2,31,176,31,176,30,6,31,172,31,80,31,47,31,202,31,178,31,213,31,178,31,250,31,224,31,35,31,96,31,48,31,48,30,48,29,117,31,117,30,215,31,215,30,29,31,42,31,11,31,11,30,230,31,10,31,219,31,219,31,134,31,7,31,7,30,200,31,61,31,78,31,121,31,177,31,60,31,245,31,252,31,252,30,226,31,15,31,151,31,9,31,9,30,166,31,233,31,66,31,74,31,67,31,41,31,22,31,108,31,229,31,189,31,38,31,38,30,240,31,19,31,19,30,146,31,97,31,110,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
