-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 468;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (152,0,175,0,239,0,59,0,96,0,170,0,211,0,0,0,0,0,143,0,0,0,0,0,0,0,110,0,47,0,179,0,253,0,212,0,152,0,20,0,162,0,0,0,0,0,251,0,129,0,173,0,3,0,95,0,200,0,103,0,169,0,65,0,166,0,152,0,0,0,9,0,121,0,22,0,205,0,134,0,191,0,72,0,0,0,186,0,234,0,102,0,208,0,33,0,232,0,102,0,0,0,154,0,42,0,43,0,140,0,75,0,95,0,0,0,75,0,230,0,84,0,67,0,31,0,0,0,107,0,205,0,132,0,1,0,239,0,3,0,196,0,101,0,48,0,219,0,55,0,35,0,0,0,108,0,0,0,185,0,85,0,73,0,49,0,189,0,147,0,10,0,0,0,0,0,117,0,82,0,0,0,0,0,0,0,187,0,5,0,0,0,237,0,9,0,213,0,140,0,52,0,182,0,147,0,0,0,23,0,0,0,142,0,217,0,46,0,10,0,0,0,254,0,114,0,231,0,66,0,0,0,222,0,42,0,20,0,0,0,29,0,9,0,8,0,0,0,0,0,54,0,174,0,48,0,0,0,52,0,0,0,107,0,32,0,202,0,90,0,47,0,123,0,210,0,101,0,171,0,182,0,135,0,17,0,163,0,0,0,0,0,113,0,39,0,118,0,103,0,64,0,112,0,98,0,161,0,63,0,79,0,207,0,175,0,205,0,204,0,63,0,109,0,57,0,165,0,23,0,124,0,61,0,0,0,125,0,187,0,0,0,101,0,80,0,82,0,240,0,122,0,0,0,234,0,0,0,81,0,222,0,99,0,225,0,31,0,238,0,17,0,131,0,3,0,0,0,203,0,189,0,33,0,36,0,2,0,228,0,25,0,139,0,112,0,240,0,163,0,65,0,147,0,0,0,84,0,201,0,65,0,0,0,176,0,176,0,177,0,0,0,60,0,0,0,130,0,197,0,80,0,251,0,0,0,223,0,118,0,83,0,110,0,237,0,16,0,165,0,205,0,20,0,0,0,161,0,158,0,195,0,0,0,24,0,86,0,0,0,19,0,0,0,118,0,0,0,204,0,102,0,0,0,199,0,217,0,88,0,35,0,108,0,62,0,226,0,0,0,0,0,42,0,36,0,135,0,119,0,58,0,0,0,166,0,244,0,95,0,233,0,227,0,0,0,196,0,0,0,138,0,38,0,92,0,135,0,89,0,168,0,0,0,227,0,132,0,112,0,0,0,163,0,53,0,246,0,0,0,153,0,88,0,52,0,216,0,249,0,245,0,131,0,148,0,179,0,128,0,49,0,161,0,139,0,158,0,231,0,80,0,30,0,0,0,166,0,214,0,118,0,107,0,223,0,8,0,209,0,143,0,0,0,131,0,252,0,59,0,134,0,215,0,0,0,0,0,85,0,100,0,0,0,35,0,123,0,0,0,92,0,89,0,0,0,0,0,143,0,166,0,76,0,210,0,236,0,68,0,44,0,3,0,150,0,51,0,219,0,181,0,130,0,81,0,137,0,202,0,216,0,129,0,242,0,138,0,246,0,0,0,140,0,0,0,209,0,114,0,198,0,255,0,193,0,108,0,64,0,53,0,119,0,167,0,117,0,161,0,4,0,195,0,109,0,0,0,0,0,17,0,82,0,82,0,192,0,233,0,0,0,31,0,243,0,17,0,187,0,106,0,0,0,0,0,128,0,117,0,216,0,31,0,200,0,0,0,48,0,0,0,113,0,3,0,190,0,5,0,124,0,97,0,126,0,0,0,207,0,0,0,0,0,52,0,0,0,97,0,168,0,5,0,29,0,18,0,255,0,103,0,37,0,71,0,64,0,84,0,0,0,101,0,126,0,221,0,144,0,156,0,225,0,215,0,93,0,201,0,57,0,12,0,65,0,195,0,127,0,168,0,223,0,13,0,54,0,0,0,155,0,243,0,157,0,0,0,100,0,248,0,96,0,138,0,0,0,44,0,188,0,90,0,180,0,128,0,0,0,73,0,171,0,177,0,35,0,233,0,69,0,209,0,140,0,0,0,113,0,0,0,44,0,84,0,227,0,143,0,81,0,123,0,255,0,94,0,54,0,163,0,111,0,0,0);
signal scenario_full  : scenario_type := (152,31,175,31,239,31,59,31,96,31,170,31,211,31,211,30,211,29,143,31,143,30,143,29,143,28,110,31,47,31,179,31,253,31,212,31,152,31,20,31,162,31,162,30,162,29,251,31,129,31,173,31,3,31,95,31,200,31,103,31,169,31,65,31,166,31,152,31,152,30,9,31,121,31,22,31,205,31,134,31,191,31,72,31,72,30,186,31,234,31,102,31,208,31,33,31,232,31,102,31,102,30,154,31,42,31,43,31,140,31,75,31,95,31,95,30,75,31,230,31,84,31,67,31,31,31,31,30,107,31,205,31,132,31,1,31,239,31,3,31,196,31,101,31,48,31,219,31,55,31,35,31,35,30,108,31,108,30,185,31,85,31,73,31,49,31,189,31,147,31,10,31,10,30,10,29,117,31,82,31,82,30,82,29,82,28,187,31,5,31,5,30,237,31,9,31,213,31,140,31,52,31,182,31,147,31,147,30,23,31,23,30,142,31,217,31,46,31,10,31,10,30,254,31,114,31,231,31,66,31,66,30,222,31,42,31,20,31,20,30,29,31,9,31,8,31,8,30,8,29,54,31,174,31,48,31,48,30,52,31,52,30,107,31,32,31,202,31,90,31,47,31,123,31,210,31,101,31,171,31,182,31,135,31,17,31,163,31,163,30,163,29,113,31,39,31,118,31,103,31,64,31,112,31,98,31,161,31,63,31,79,31,207,31,175,31,205,31,204,31,63,31,109,31,57,31,165,31,23,31,124,31,61,31,61,30,125,31,187,31,187,30,101,31,80,31,82,31,240,31,122,31,122,30,234,31,234,30,81,31,222,31,99,31,225,31,31,31,238,31,17,31,131,31,3,31,3,30,203,31,189,31,33,31,36,31,2,31,228,31,25,31,139,31,112,31,240,31,163,31,65,31,147,31,147,30,84,31,201,31,65,31,65,30,176,31,176,31,177,31,177,30,60,31,60,30,130,31,197,31,80,31,251,31,251,30,223,31,118,31,83,31,110,31,237,31,16,31,165,31,205,31,20,31,20,30,161,31,158,31,195,31,195,30,24,31,86,31,86,30,19,31,19,30,118,31,118,30,204,31,102,31,102,30,199,31,217,31,88,31,35,31,108,31,62,31,226,31,226,30,226,29,42,31,36,31,135,31,119,31,58,31,58,30,166,31,244,31,95,31,233,31,227,31,227,30,196,31,196,30,138,31,38,31,92,31,135,31,89,31,168,31,168,30,227,31,132,31,112,31,112,30,163,31,53,31,246,31,246,30,153,31,88,31,52,31,216,31,249,31,245,31,131,31,148,31,179,31,128,31,49,31,161,31,139,31,158,31,231,31,80,31,30,31,30,30,166,31,214,31,118,31,107,31,223,31,8,31,209,31,143,31,143,30,131,31,252,31,59,31,134,31,215,31,215,30,215,29,85,31,100,31,100,30,35,31,123,31,123,30,92,31,89,31,89,30,89,29,143,31,166,31,76,31,210,31,236,31,68,31,44,31,3,31,150,31,51,31,219,31,181,31,130,31,81,31,137,31,202,31,216,31,129,31,242,31,138,31,246,31,246,30,140,31,140,30,209,31,114,31,198,31,255,31,193,31,108,31,64,31,53,31,119,31,167,31,117,31,161,31,4,31,195,31,109,31,109,30,109,29,17,31,82,31,82,31,192,31,233,31,233,30,31,31,243,31,17,31,187,31,106,31,106,30,106,29,128,31,117,31,216,31,31,31,200,31,200,30,48,31,48,30,113,31,3,31,190,31,5,31,124,31,97,31,126,31,126,30,207,31,207,30,207,29,52,31,52,30,97,31,168,31,5,31,29,31,18,31,255,31,103,31,37,31,71,31,64,31,84,31,84,30,101,31,126,31,221,31,144,31,156,31,225,31,215,31,93,31,201,31,57,31,12,31,65,31,195,31,127,31,168,31,223,31,13,31,54,31,54,30,155,31,243,31,157,31,157,30,100,31,248,31,96,31,138,31,138,30,44,31,188,31,90,31,180,31,128,31,128,30,73,31,171,31,177,31,35,31,233,31,69,31,209,31,140,31,140,30,113,31,113,30,44,31,84,31,227,31,143,31,81,31,123,31,255,31,94,31,54,31,163,31,111,31,111,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
