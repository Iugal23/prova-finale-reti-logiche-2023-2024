-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 432;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (112,0,244,0,0,0,149,0,120,0,121,0,158,0,215,0,158,0,161,0,220,0,36,0,164,0,0,0,145,0,0,0,62,0,0,0,65,0,93,0,155,0,0,0,10,0,128,0,212,0,18,0,0,0,222,0,21,0,0,0,101,0,100,0,102,0,98,0,0,0,77,0,0,0,0,0,227,0,140,0,49,0,172,0,108,0,174,0,238,0,194,0,13,0,63,0,202,0,232,0,0,0,0,0,249,0,12,0,0,0,156,0,254,0,246,0,234,0,147,0,220,0,64,0,1,0,53,0,91,0,0,0,0,0,0,0,79,0,185,0,105,0,214,0,236,0,168,0,24,0,100,0,65,0,82,0,0,0,230,0,244,0,240,0,75,0,73,0,43,0,243,0,182,0,0,0,55,0,0,0,227,0,0,0,56,0,33,0,40,0,172,0,136,0,148,0,239,0,0,0,214,0,90,0,0,0,201,0,184,0,104,0,40,0,159,0,87,0,11,0,200,0,174,0,66,0,168,0,0,0,57,0,155,0,12,0,0,0,0,0,247,0,149,0,253,0,98,0,97,0,28,0,130,0,127,0,134,0,225,0,61,0,0,0,157,0,206,0,204,0,147,0,0,0,223,0,175,0,96,0,36,0,59,0,69,0,99,0,222,0,173,0,61,0,56,0,237,0,0,0,222,0,154,0,0,0,0,0,70,0,0,0,139,0,8,0,29,0,18,0,148,0,198,0,0,0,27,0,59,0,198,0,45,0,4,0,0,0,0,0,28,0,131,0,147,0,0,0,176,0,253,0,0,0,145,0,39,0,128,0,98,0,39,0,148,0,82,0,27,0,0,0,111,0,128,0,0,0,0,0,24,0,2,0,123,0,0,0,0,0,243,0,194,0,66,0,0,0,250,0,216,0,0,0,0,0,10,0,26,0,0,0,0,0,50,0,116,0,106,0,114,0,153,0,251,0,29,0,43,0,0,0,191,0,40,0,0,0,2,0,0,0,48,0,0,0,161,0,227,0,0,0,0,0,17,0,44,0,230,0,0,0,0,0,83,0,122,0,42,0,147,0,0,0,5,0,3,0,225,0,116,0,224,0,82,0,37,0,36,0,220,0,121,0,126,0,0,0,0,0,47,0,61,0,254,0,0,0,19,0,188,0,140,0,173,0,0,0,28,0,0,0,109,0,34,0,0,0,0,0,210,0,0,0,0,0,0,0,162,0,51,0,65,0,205,0,194,0,220,0,0,0,0,0,0,0,212,0,1,0,0,0,245,0,0,0,116,0,108,0,161,0,133,0,253,0,27,0,0,0,155,0,71,0,53,0,248,0,69,0,228,0,5,0,113,0,103,0,164,0,192,0,211,0,93,0,0,0,102,0,0,0,251,0,0,0,254,0,0,0,111,0,180,0,93,0,0,0,29,0,35,0,129,0,0,0,216,0,81,0,43,0,135,0,199,0,212,0,56,0,208,0,253,0,99,0,120,0,0,0,65,0,0,0,0,0,0,0,0,0,56,0,88,0,130,0,157,0,244,0,156,0,200,0,38,0,44,0,238,0,134,0,169,0,0,0,247,0,134,0,228,0,125,0,230,0,0,0,25,0,0,0,178,0,137,0,217,0,160,0,142,0,7,0,178,0,139,0,5,0,62,0,94,0,78,0,73,0,79,0,162,0,77,0,252,0,23,0,105,0,0,0,125,0,97,0,0,0,0,0,232,0,212,0,157,0,30,0,215,0,133,0,0,0,206,0,182,0,217,0,229,0,137,0,230,0,101,0,213,0,141,0,192,0,81,0,40,0,133,0,231,0,39,0,16,0,1,0,133,0,165,0,233,0,159,0,172,0,162,0,0,0,187,0,62,0,0,0,19,0,3,0,182,0,134,0,115,0,252,0,219,0,9,0,235,0,124,0,0,0,0,0,239,0,222,0,100,0,98,0,78,0,63,0);
signal scenario_full  : scenario_type := (112,31,244,31,244,30,149,31,120,31,121,31,158,31,215,31,158,31,161,31,220,31,36,31,164,31,164,30,145,31,145,30,62,31,62,30,65,31,93,31,155,31,155,30,10,31,128,31,212,31,18,31,18,30,222,31,21,31,21,30,101,31,100,31,102,31,98,31,98,30,77,31,77,30,77,29,227,31,140,31,49,31,172,31,108,31,174,31,238,31,194,31,13,31,63,31,202,31,232,31,232,30,232,29,249,31,12,31,12,30,156,31,254,31,246,31,234,31,147,31,220,31,64,31,1,31,53,31,91,31,91,30,91,29,91,28,79,31,185,31,105,31,214,31,236,31,168,31,24,31,100,31,65,31,82,31,82,30,230,31,244,31,240,31,75,31,73,31,43,31,243,31,182,31,182,30,55,31,55,30,227,31,227,30,56,31,33,31,40,31,172,31,136,31,148,31,239,31,239,30,214,31,90,31,90,30,201,31,184,31,104,31,40,31,159,31,87,31,11,31,200,31,174,31,66,31,168,31,168,30,57,31,155,31,12,31,12,30,12,29,247,31,149,31,253,31,98,31,97,31,28,31,130,31,127,31,134,31,225,31,61,31,61,30,157,31,206,31,204,31,147,31,147,30,223,31,175,31,96,31,36,31,59,31,69,31,99,31,222,31,173,31,61,31,56,31,237,31,237,30,222,31,154,31,154,30,154,29,70,31,70,30,139,31,8,31,29,31,18,31,148,31,198,31,198,30,27,31,59,31,198,31,45,31,4,31,4,30,4,29,28,31,131,31,147,31,147,30,176,31,253,31,253,30,145,31,39,31,128,31,98,31,39,31,148,31,82,31,27,31,27,30,111,31,128,31,128,30,128,29,24,31,2,31,123,31,123,30,123,29,243,31,194,31,66,31,66,30,250,31,216,31,216,30,216,29,10,31,26,31,26,30,26,29,50,31,116,31,106,31,114,31,153,31,251,31,29,31,43,31,43,30,191,31,40,31,40,30,2,31,2,30,48,31,48,30,161,31,227,31,227,30,227,29,17,31,44,31,230,31,230,30,230,29,83,31,122,31,42,31,147,31,147,30,5,31,3,31,225,31,116,31,224,31,82,31,37,31,36,31,220,31,121,31,126,31,126,30,126,29,47,31,61,31,254,31,254,30,19,31,188,31,140,31,173,31,173,30,28,31,28,30,109,31,34,31,34,30,34,29,210,31,210,30,210,29,210,28,162,31,51,31,65,31,205,31,194,31,220,31,220,30,220,29,220,28,212,31,1,31,1,30,245,31,245,30,116,31,108,31,161,31,133,31,253,31,27,31,27,30,155,31,71,31,53,31,248,31,69,31,228,31,5,31,113,31,103,31,164,31,192,31,211,31,93,31,93,30,102,31,102,30,251,31,251,30,254,31,254,30,111,31,180,31,93,31,93,30,29,31,35,31,129,31,129,30,216,31,81,31,43,31,135,31,199,31,212,31,56,31,208,31,253,31,99,31,120,31,120,30,65,31,65,30,65,29,65,28,65,27,56,31,88,31,130,31,157,31,244,31,156,31,200,31,38,31,44,31,238,31,134,31,169,31,169,30,247,31,134,31,228,31,125,31,230,31,230,30,25,31,25,30,178,31,137,31,217,31,160,31,142,31,7,31,178,31,139,31,5,31,62,31,94,31,78,31,73,31,79,31,162,31,77,31,252,31,23,31,105,31,105,30,125,31,97,31,97,30,97,29,232,31,212,31,157,31,30,31,215,31,133,31,133,30,206,31,182,31,217,31,229,31,137,31,230,31,101,31,213,31,141,31,192,31,81,31,40,31,133,31,231,31,39,31,16,31,1,31,133,31,165,31,233,31,159,31,172,31,162,31,162,30,187,31,62,31,62,30,19,31,3,31,182,31,134,31,115,31,252,31,219,31,9,31,235,31,124,31,124,30,124,29,239,31,222,31,100,31,98,31,78,31,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
