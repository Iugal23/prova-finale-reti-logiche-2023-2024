-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 639;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (177,0,144,0,56,0,0,0,220,0,142,0,105,0,120,0,248,0,187,0,0,0,0,0,0,0,0,0,212,0,129,0,0,0,0,0,2,0,0,0,52,0,0,0,147,0,154,0,123,0,13,0,64,0,0,0,45,0,114,0,0,0,0,0,121,0,0,0,0,0,167,0,211,0,26,0,0,0,226,0,243,0,168,0,86,0,255,0,229,0,129,0,96,0,216,0,144,0,0,0,83,0,132,0,195,0,78,0,0,0,0,0,129,0,118,0,75,0,176,0,0,0,185,0,39,0,43,0,21,0,107,0,2,0,109,0,128,0,138,0,78,0,159,0,158,0,50,0,49,0,19,0,143,0,109,0,101,0,241,0,14,0,184,0,182,0,243,0,0,0,153,0,133,0,50,0,172,0,65,0,0,0,0,0,0,0,0,0,189,0,31,0,0,0,161,0,202,0,0,0,0,0,0,0,224,0,231,0,28,0,205,0,226,0,82,0,44,0,65,0,38,0,0,0,223,0,195,0,38,0,167,0,254,0,190,0,155,0,73,0,0,0,233,0,141,0,203,0,93,0,74,0,197,0,130,0,197,0,207,0,0,0,230,0,184,0,0,0,215,0,148,0,0,0,0,0,0,0,18,0,0,0,70,0,122,0,204,0,64,0,117,0,192,0,32,0,53,0,141,0,66,0,0,0,57,0,76,0,0,0,145,0,111,0,0,0,0,0,172,0,173,0,148,0,184,0,222,0,125,0,63,0,133,0,0,0,187,0,244,0,64,0,13,0,33,0,48,0,47,0,186,0,86,0,67,0,42,0,116,0,147,0,7,0,175,0,21,0,0,0,43,0,66,0,119,0,223,0,228,0,42,0,0,0,116,0,81,0,180,0,14,0,108,0,57,0,253,0,0,0,0,0,106,0,221,0,0,0,219,0,248,0,80,0,63,0,126,0,80,0,95,0,0,0,0,0,236,0,152,0,63,0,167,0,21,0,16,0,166,0,173,0,135,0,219,0,129,0,220,0,136,0,75,0,0,0,91,0,78,0,0,0,58,0,41,0,82,0,58,0,0,0,126,0,206,0,90,0,139,0,52,0,0,0,144,0,226,0,211,0,0,0,59,0,49,0,0,0,80,0,0,0,0,0,30,0,24,0,0,0,236,0,190,0,19,0,116,0,174,0,129,0,203,0,243,0,239,0,7,0,0,0,101,0,88,0,205,0,101,0,0,0,183,0,165,0,0,0,89,0,210,0,189,0,1,0,150,0,85,0,243,0,175,0,252,0,19,0,137,0,206,0,0,0,148,0,200,0,1,0,48,0,1,0,148,0,86,0,9,0,237,0,175,0,148,0,0,0,129,0,0,0,199,0,147,0,154,0,49,0,7,0,87,0,160,0,0,0,135,0,207,0,21,0,231,0,46,0,220,0,165,0,0,0,110,0,132,0,245,0,90,0,97,0,0,0,78,0,247,0,4,0,0,0,250,0,33,0,1,0,20,0,255,0,4,0,128,0,0,0,0,0,53,0,0,0,0,0,154,0,0,0,44,0,160,0,0,0,58,0,21,0,191,0,3,0,231,0,54,0,208,0,250,0,133,0,43,0,222,0,239,0,14,0,33,0,167,0,42,0,252,0,26,0,0,0,0,0,124,0,0,0,13,0,0,0,0,0,227,0,61,0,0,0,174,0,0,0,226,0,111,0,102,0,236,0,71,0,0,0,60,0,0,0,141,0,16,0,24,0,68,0,49,0,159,0,71,0,0,0,180,0,0,0,178,0,226,0,0,0,233,0,8,0,0,0,90,0,15,0,235,0,121,0,0,0,36,0,97,0,0,0,7,0,96,0,183,0,6,0,0,0,0,0,0,0,20,0,49,0,47,0,0,0,115,0,0,0,255,0,175,0,218,0,51,0,0,0,100,0,68,0,57,0,152,0,0,0,225,0,215,0,62,0,15,0,160,0,114,0,173,0,0,0,6,0,116,0,168,0,100,0,147,0,76,0,242,0,137,0,139,0,159,0,38,0,32,0,168,0,38,0,0,0,243,0,71,0,180,0,114,0,62,0,230,0,0,0,65,0,161,0,0,0,140,0,121,0,87,0,0,0,143,0,0,0,10,0,0,0,213,0,242,0,69,0,65,0,151,0,210,0,0,0,165,0,141,0,202,0,29,0,218,0,136,0,0,0,102,0,9,0,32,0,102,0,14,0,87,0,154,0,203,0,40,0,192,0,0,0,124,0,255,0,148,0,0,0,137,0,114,0,128,0,23,0,123,0,15,0,53,0,145,0,212,0,153,0,250,0,58,0,14,0,178,0,0,0,180,0,160,0,116,0,37,0,101,0,102,0,0,0,166,0,203,0,63,0,41,0,243,0,187,0,37,0,137,0,181,0,0,0,12,0,252,0,0,0,103,0,7,0,90,0,177,0,121,0,82,0,183,0,93,0,62,0,107,0,173,0,0,0,0,0,169,0,225,0,141,0,0,0,0,0,0,0,129,0,5,0,0,0,12,0,38,0,133,0,0,0,5,0,36,0,41,0,41,0,161,0,88,0,0,0,132,0,248,0,0,0,209,0,11,0,0,0,142,0,227,0,220,0,165,0,90,0,23,0,123,0,164,0,212,0,95,0,20,0,0,0,115,0,34,0,0,0,133,0,139,0,139,0,50,0,133,0,0,0,48,0,236,0,250,0,0,0,249,0,0,0,0,0,56,0,217,0,195,0,207,0,210,0,168,0,204,0,44,0,219,0,159,0,0,0,34,0,0,0,190,0,0,0,0,0,58,0,0,0,141,0,38,0,0,0,39,0,99,0,52,0,81,0,198,0,50,0,134,0,0,0,44,0,0,0,175,0,220,0,83,0,172,0,12,0,235,0,218,0);
signal scenario_full  : scenario_type := (177,31,144,31,56,31,56,30,220,31,142,31,105,31,120,31,248,31,187,31,187,30,187,29,187,28,187,27,212,31,129,31,129,30,129,29,2,31,2,30,52,31,52,30,147,31,154,31,123,31,13,31,64,31,64,30,45,31,114,31,114,30,114,29,121,31,121,30,121,29,167,31,211,31,26,31,26,30,226,31,243,31,168,31,86,31,255,31,229,31,129,31,96,31,216,31,144,31,144,30,83,31,132,31,195,31,78,31,78,30,78,29,129,31,118,31,75,31,176,31,176,30,185,31,39,31,43,31,21,31,107,31,2,31,109,31,128,31,138,31,78,31,159,31,158,31,50,31,49,31,19,31,143,31,109,31,101,31,241,31,14,31,184,31,182,31,243,31,243,30,153,31,133,31,50,31,172,31,65,31,65,30,65,29,65,28,65,27,189,31,31,31,31,30,161,31,202,31,202,30,202,29,202,28,224,31,231,31,28,31,205,31,226,31,82,31,44,31,65,31,38,31,38,30,223,31,195,31,38,31,167,31,254,31,190,31,155,31,73,31,73,30,233,31,141,31,203,31,93,31,74,31,197,31,130,31,197,31,207,31,207,30,230,31,184,31,184,30,215,31,148,31,148,30,148,29,148,28,18,31,18,30,70,31,122,31,204,31,64,31,117,31,192,31,32,31,53,31,141,31,66,31,66,30,57,31,76,31,76,30,145,31,111,31,111,30,111,29,172,31,173,31,148,31,184,31,222,31,125,31,63,31,133,31,133,30,187,31,244,31,64,31,13,31,33,31,48,31,47,31,186,31,86,31,67,31,42,31,116,31,147,31,7,31,175,31,21,31,21,30,43,31,66,31,119,31,223,31,228,31,42,31,42,30,116,31,81,31,180,31,14,31,108,31,57,31,253,31,253,30,253,29,106,31,221,31,221,30,219,31,248,31,80,31,63,31,126,31,80,31,95,31,95,30,95,29,236,31,152,31,63,31,167,31,21,31,16,31,166,31,173,31,135,31,219,31,129,31,220,31,136,31,75,31,75,30,91,31,78,31,78,30,58,31,41,31,82,31,58,31,58,30,126,31,206,31,90,31,139,31,52,31,52,30,144,31,226,31,211,31,211,30,59,31,49,31,49,30,80,31,80,30,80,29,30,31,24,31,24,30,236,31,190,31,19,31,116,31,174,31,129,31,203,31,243,31,239,31,7,31,7,30,101,31,88,31,205,31,101,31,101,30,183,31,165,31,165,30,89,31,210,31,189,31,1,31,150,31,85,31,243,31,175,31,252,31,19,31,137,31,206,31,206,30,148,31,200,31,1,31,48,31,1,31,148,31,86,31,9,31,237,31,175,31,148,31,148,30,129,31,129,30,199,31,147,31,154,31,49,31,7,31,87,31,160,31,160,30,135,31,207,31,21,31,231,31,46,31,220,31,165,31,165,30,110,31,132,31,245,31,90,31,97,31,97,30,78,31,247,31,4,31,4,30,250,31,33,31,1,31,20,31,255,31,4,31,128,31,128,30,128,29,53,31,53,30,53,29,154,31,154,30,44,31,160,31,160,30,58,31,21,31,191,31,3,31,231,31,54,31,208,31,250,31,133,31,43,31,222,31,239,31,14,31,33,31,167,31,42,31,252,31,26,31,26,30,26,29,124,31,124,30,13,31,13,30,13,29,227,31,61,31,61,30,174,31,174,30,226,31,111,31,102,31,236,31,71,31,71,30,60,31,60,30,141,31,16,31,24,31,68,31,49,31,159,31,71,31,71,30,180,31,180,30,178,31,226,31,226,30,233,31,8,31,8,30,90,31,15,31,235,31,121,31,121,30,36,31,97,31,97,30,7,31,96,31,183,31,6,31,6,30,6,29,6,28,20,31,49,31,47,31,47,30,115,31,115,30,255,31,175,31,218,31,51,31,51,30,100,31,68,31,57,31,152,31,152,30,225,31,215,31,62,31,15,31,160,31,114,31,173,31,173,30,6,31,116,31,168,31,100,31,147,31,76,31,242,31,137,31,139,31,159,31,38,31,32,31,168,31,38,31,38,30,243,31,71,31,180,31,114,31,62,31,230,31,230,30,65,31,161,31,161,30,140,31,121,31,87,31,87,30,143,31,143,30,10,31,10,30,213,31,242,31,69,31,65,31,151,31,210,31,210,30,165,31,141,31,202,31,29,31,218,31,136,31,136,30,102,31,9,31,32,31,102,31,14,31,87,31,154,31,203,31,40,31,192,31,192,30,124,31,255,31,148,31,148,30,137,31,114,31,128,31,23,31,123,31,15,31,53,31,145,31,212,31,153,31,250,31,58,31,14,31,178,31,178,30,180,31,160,31,116,31,37,31,101,31,102,31,102,30,166,31,203,31,63,31,41,31,243,31,187,31,37,31,137,31,181,31,181,30,12,31,252,31,252,30,103,31,7,31,90,31,177,31,121,31,82,31,183,31,93,31,62,31,107,31,173,31,173,30,173,29,169,31,225,31,141,31,141,30,141,29,141,28,129,31,5,31,5,30,12,31,38,31,133,31,133,30,5,31,36,31,41,31,41,31,161,31,88,31,88,30,132,31,248,31,248,30,209,31,11,31,11,30,142,31,227,31,220,31,165,31,90,31,23,31,123,31,164,31,212,31,95,31,20,31,20,30,115,31,34,31,34,30,133,31,139,31,139,31,50,31,133,31,133,30,48,31,236,31,250,31,250,30,249,31,249,30,249,29,56,31,217,31,195,31,207,31,210,31,168,31,204,31,44,31,219,31,159,31,159,30,34,31,34,30,190,31,190,30,190,29,58,31,58,30,141,31,38,31,38,30,39,31,99,31,52,31,81,31,198,31,50,31,134,31,134,30,44,31,44,30,175,31,220,31,83,31,172,31,12,31,235,31,218,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
