-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 999;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (121,0,49,0,76,0,41,0,7,0,0,0,106,0,174,0,10,0,226,0,173,0,163,0,141,0,0,0,0,0,0,0,146,0,216,0,0,0,153,0,157,0,76,0,37,0,0,0,255,0,116,0,5,0,0,0,0,0,35,0,115,0,4,0,1,0,69,0,204,0,56,0,226,0,60,0,14,0,0,0,66,0,118,0,0,0,28,0,249,0,0,0,0,0,169,0,119,0,145,0,160,0,101,0,212,0,243,0,57,0,25,0,164,0,219,0,104,0,143,0,0,0,23,0,0,0,0,0,154,0,0,0,245,0,57,0,167,0,78,0,217,0,100,0,0,0,0,0,140,0,199,0,113,0,104,0,38,0,17,0,251,0,0,0,156,0,0,0,0,0,251,0,3,0,156,0,45,0,59,0,175,0,237,0,236,0,156,0,167,0,207,0,213,0,0,0,159,0,212,0,119,0,225,0,217,0,70,0,221,0,218,0,123,0,0,0,28,0,194,0,28,0,121,0,1,0,189,0,227,0,254,0,144,0,215,0,238,0,115,0,187,0,230,0,227,0,131,0,36,0,253,0,245,0,170,0,247,0,115,0,202,0,92,0,56,0,3,0,221,0,90,0,50,0,0,0,235,0,97,0,69,0,92,0,0,0,0,0,219,0,139,0,91,0,204,0,58,0,232,0,151,0,74,0,0,0,146,0,228,0,177,0,210,0,39,0,240,0,154,0,175,0,236,0,153,0,93,0,29,0,6,0,227,0,203,0,9,0,182,0,110,0,12,0,157,0,85,0,201,0,0,0,0,0,16,0,68,0,87,0,149,0,214,0,0,0,17,0,112,0,12,0,32,0,26,0,230,0,169,0,119,0,126,0,187,0,221,0,66,0,179,0,92,0,59,0,175,0,87,0,131,0,46,0,208,0,34,0,35,0,31,0,66,0,224,0,0,0,69,0,43,0,153,0,165,0,66,0,62,0,0,0,33,0,218,0,125,0,0,0,208,0,239,0,19,0,76,0,0,0,234,0,63,0,79,0,169,0,94,0,74,0,32,0,188,0,196,0,232,0,246,0,0,0,118,0,18,0,0,0,169,0,7,0,76,0,82,0,161,0,113,0,66,0,8,0,188,0,0,0,218,0,162,0,165,0,0,0,68,0,0,0,186,0,255,0,0,0,0,0,19,0,125,0,251,0,103,0,22,0,247,0,29,0,185,0,233,0,191,0,252,0,65,0,0,0,112,0,0,0,211,0,1,0,24,0,210,0,229,0,244,0,143,0,155,0,126,0,86,0,0,0,242,0,124,0,4,0,201,0,244,0,67,0,0,0,177,0,106,0,229,0,252,0,228,0,188,0,55,0,186,0,171,0,252,0,201,0,73,0,7,0,23,0,204,0,0,0,0,0,36,0,249,0,181,0,242,0,185,0,0,0,0,0,143,0,68,0,0,0,0,0,129,0,0,0,39,0,0,0,28,0,16,0,160,0,143,0,88,0,40,0,141,0,75,0,22,0,4,0,253,0,0,0,0,0,0,0,200,0,163,0,214,0,183,0,244,0,41,0,0,0,0,0,110,0,52,0,151,0,97,0,6,0,184,0,30,0,107,0,57,0,0,0,0,0,140,0,59,0,14,0,227,0,0,0,178,0,0,0,162,0,0,0,79,0,226,0,117,0,85,0,217,0,206,0,195,0,244,0,133,0,63,0,106,0,42,0,101,0,232,0,82,0,0,0,54,0,221,0,151,0,0,0,120,0,71,0,186,0,159,0,122,0,233,0,115,0,61,0,2,0,143,0,0,0,178,0,107,0,123,0,118,0,227,0,149,0,0,0,0,0,177,0,200,0,202,0,58,0,143,0,143,0,122,0,55,0,0,0,156,0,61,0,196,0,0,0,76,0,41,0,0,0,35,0,138,0,244,0,10,0,0,0,45,0,0,0,0,0,135,0,0,0,0,0,0,0,36,0,0,0,154,0,17,0,26,0,86,0,108,0,51,0,213,0,83,0,122,0,129,0,253,0,194,0,218,0,0,0,161,0,248,0,234,0,0,0,0,0,37,0,77,0,160,0,0,0,127,0,253,0,18,0,174,0,45,0,114,0,65,0,162,0,114,0,170,0,115,0,86,0,99,0,0,0,0,0,0,0,0,0,2,0,14,0,0,0,38,0,220,0,151,0,247,0,109,0,0,0,231,0,32,0,158,0,0,0,145,0,253,0,210,0,0,0,0,0,60,0,69,0,91,0,81,0,0,0,212,0,46,0,87,0,162,0,161,0,227,0,166,0,145,0,0,0,98,0,23,0,99,0,0,0,0,0,0,0,24,0,207,0,125,0,187,0,0,0,42,0,0,0,57,0,152,0,96,0,249,0,103,0,3,0,237,0,7,0,70,0,182,0,191,0,0,0,60,0,220,0,221,0,11,0,133,0,250,0,222,0,123,0,191,0,195,0,144,0,69,0,183,0,0,0,98,0,228,0,119,0,241,0,12,0,44,0,80,0,142,0,101,0,0,0,232,0,160,0,139,0,0,0,136,0,14,0,65,0,195,0,0,0,177,0,61,0,95,0,129,0,45,0,0,0,0,0,133,0,0,0,204,0,134,0,237,0,0,0,18,0,0,0,152,0,0,0,93,0,0,0,188,0,147,0,169,0,201,0,96,0,166,0,34,0,247,0,0,0,196,0,17,0,85,0,34,0,230,0,207,0,32,0,0,0,0,0,133,0,16,0,0,0,126,0,0,0,0,0,0,0,0,0,205,0,196,0,85,0,164,0,101,0,178,0,160,0,72,0,25,0,53,0,163,0,183,0,73,0,203,0,127,0,117,0,27,0,77,0,0,0,22,0,157,0,152,0,55,0,219,0,240,0,254,0,229,0,0,0,254,0,0,0,172,0,0,0,0,0,0,0,116,0,13,0,0,0,30,0,232,0,117,0,139,0,168,0,217,0,0,0,0,0,14,0,252,0,0,0,0,0,137,0,16,0,192,0,21,0,116,0,151,0,15,0,36,0,223,0,130,0,222,0,0,0,0,0,150,0,167,0,22,0,0,0,124,0,110,0,232,0,18,0,8,0,234,0,217,0,95,0,148,0,8,0,204,0,105,0,246,0,165,0,43,0,0,0,78,0,139,0,0,0,5,0,163,0,166,0,88,0,49,0,207,0,107,0,67,0,0,0,33,0,0,0,93,0,0,0,162,0,13,0,0,0,113,0,156,0,0,0,109,0,164,0,160,0,82,0,106,0,181,0,0,0,80,0,109,0,7,0,144,0,253,0,138,0,0,0,127,0,103,0,91,0,40,0,0,0,163,0,130,0,69,0,129,0,105,0,196,0,31,0,176,0,8,0,0,0,64,0,35,0,70,0,22,0,224,0,202,0,197,0,57,0,203,0,202,0,235,0,117,0,128,0,0,0,0,0,167,0,24,0,35,0,132,0,0,0,117,0,145,0,166,0,45,0,215,0,133,0,0,0,65,0,111,0,86,0,31,0,109,0,242,0,252,0,134,0,127,0,86,0,221,0,85,0,0,0,216,0,239,0,88,0,0,0,215,0,112,0,120,0,155,0,159,0,0,0,168,0,150,0,78,0,237,0,42,0,192,0,184,0,236,0,247,0,0,0,89,0,157,0,102,0,9,0,0,0,87,0,161,0,0,0,217,0,99,0,0,0,0,0,0,0,0,0,0,0,55,0,0,0,101,0,132,0,93,0,199,0,140,0,0,0,231,0,20,0,18,0,254,0,0,0,36,0,173,0,0,0,250,0,38,0,133,0,207,0,133,0,36,0,0,0,116,0,53,0,106,0,217,0,0,0,30,0,250,0,71,0,31,0,0,0,0,0,217,0,0,0,0,0,137,0,198,0,0,0,168,0,0,0,0,0,200,0,112,0,121,0,0,0,0,0,4,0,149,0,198,0,221,0,0,0,111,0,0,0,13,0,0,0,0,0,237,0,245,0,63,0,204,0,49,0,240,0,22,0,25,0,103,0,93,0,60,0,128,0,125,0,0,0,58,0,183,0,231,0,0,0,193,0,213,0,129,0,0,0,37,0,11,0,176,0,139,0,0,0,100,0,27,0,175,0,188,0,101,0,171,0,69,0,188,0,138,0,0,0,149,0,81,0,134,0,42,0,0,0,211,0,148,0,21,0,0,0,93,0,24,0,0,0,69,0,115,0,78,0,30,0,87,0,102,0,0,0,0,0,169,0,54,0,67,0,156,0,129,0,167,0,0,0,57,0,0,0,13,0,0,0,46,0,221,0,203,0,37,0,0,0,93,0,204,0,0,0,1,0,63,0,209,0,0,0,72,0,0,0,72,0,92,0,106,0,0,0,201,0,0,0,174,0,0,0,0,0,0,0,109,0,18,0,128,0,0,0,59,0,40,0,158,0,44,0,213,0,217,0,223,0,0,0,233,0,214,0,192,0,74,0,84,0,105,0,251,0,0,0,24,0,218,0,205,0,91,0,61,0,215,0,0,0,27,0,195,0,201,0);
signal scenario_full  : scenario_type := (121,31,49,31,76,31,41,31,7,31,7,30,106,31,174,31,10,31,226,31,173,31,163,31,141,31,141,30,141,29,141,28,146,31,216,31,216,30,153,31,157,31,76,31,37,31,37,30,255,31,116,31,5,31,5,30,5,29,35,31,115,31,4,31,1,31,69,31,204,31,56,31,226,31,60,31,14,31,14,30,66,31,118,31,118,30,28,31,249,31,249,30,249,29,169,31,119,31,145,31,160,31,101,31,212,31,243,31,57,31,25,31,164,31,219,31,104,31,143,31,143,30,23,31,23,30,23,29,154,31,154,30,245,31,57,31,167,31,78,31,217,31,100,31,100,30,100,29,140,31,199,31,113,31,104,31,38,31,17,31,251,31,251,30,156,31,156,30,156,29,251,31,3,31,156,31,45,31,59,31,175,31,237,31,236,31,156,31,167,31,207,31,213,31,213,30,159,31,212,31,119,31,225,31,217,31,70,31,221,31,218,31,123,31,123,30,28,31,194,31,28,31,121,31,1,31,189,31,227,31,254,31,144,31,215,31,238,31,115,31,187,31,230,31,227,31,131,31,36,31,253,31,245,31,170,31,247,31,115,31,202,31,92,31,56,31,3,31,221,31,90,31,50,31,50,30,235,31,97,31,69,31,92,31,92,30,92,29,219,31,139,31,91,31,204,31,58,31,232,31,151,31,74,31,74,30,146,31,228,31,177,31,210,31,39,31,240,31,154,31,175,31,236,31,153,31,93,31,29,31,6,31,227,31,203,31,9,31,182,31,110,31,12,31,157,31,85,31,201,31,201,30,201,29,16,31,68,31,87,31,149,31,214,31,214,30,17,31,112,31,12,31,32,31,26,31,230,31,169,31,119,31,126,31,187,31,221,31,66,31,179,31,92,31,59,31,175,31,87,31,131,31,46,31,208,31,34,31,35,31,31,31,66,31,224,31,224,30,69,31,43,31,153,31,165,31,66,31,62,31,62,30,33,31,218,31,125,31,125,30,208,31,239,31,19,31,76,31,76,30,234,31,63,31,79,31,169,31,94,31,74,31,32,31,188,31,196,31,232,31,246,31,246,30,118,31,18,31,18,30,169,31,7,31,76,31,82,31,161,31,113,31,66,31,8,31,188,31,188,30,218,31,162,31,165,31,165,30,68,31,68,30,186,31,255,31,255,30,255,29,19,31,125,31,251,31,103,31,22,31,247,31,29,31,185,31,233,31,191,31,252,31,65,31,65,30,112,31,112,30,211,31,1,31,24,31,210,31,229,31,244,31,143,31,155,31,126,31,86,31,86,30,242,31,124,31,4,31,201,31,244,31,67,31,67,30,177,31,106,31,229,31,252,31,228,31,188,31,55,31,186,31,171,31,252,31,201,31,73,31,7,31,23,31,204,31,204,30,204,29,36,31,249,31,181,31,242,31,185,31,185,30,185,29,143,31,68,31,68,30,68,29,129,31,129,30,39,31,39,30,28,31,16,31,160,31,143,31,88,31,40,31,141,31,75,31,22,31,4,31,253,31,253,30,253,29,253,28,200,31,163,31,214,31,183,31,244,31,41,31,41,30,41,29,110,31,52,31,151,31,97,31,6,31,184,31,30,31,107,31,57,31,57,30,57,29,140,31,59,31,14,31,227,31,227,30,178,31,178,30,162,31,162,30,79,31,226,31,117,31,85,31,217,31,206,31,195,31,244,31,133,31,63,31,106,31,42,31,101,31,232,31,82,31,82,30,54,31,221,31,151,31,151,30,120,31,71,31,186,31,159,31,122,31,233,31,115,31,61,31,2,31,143,31,143,30,178,31,107,31,123,31,118,31,227,31,149,31,149,30,149,29,177,31,200,31,202,31,58,31,143,31,143,31,122,31,55,31,55,30,156,31,61,31,196,31,196,30,76,31,41,31,41,30,35,31,138,31,244,31,10,31,10,30,45,31,45,30,45,29,135,31,135,30,135,29,135,28,36,31,36,30,154,31,17,31,26,31,86,31,108,31,51,31,213,31,83,31,122,31,129,31,253,31,194,31,218,31,218,30,161,31,248,31,234,31,234,30,234,29,37,31,77,31,160,31,160,30,127,31,253,31,18,31,174,31,45,31,114,31,65,31,162,31,114,31,170,31,115,31,86,31,99,31,99,30,99,29,99,28,99,27,2,31,14,31,14,30,38,31,220,31,151,31,247,31,109,31,109,30,231,31,32,31,158,31,158,30,145,31,253,31,210,31,210,30,210,29,60,31,69,31,91,31,81,31,81,30,212,31,46,31,87,31,162,31,161,31,227,31,166,31,145,31,145,30,98,31,23,31,99,31,99,30,99,29,99,28,24,31,207,31,125,31,187,31,187,30,42,31,42,30,57,31,152,31,96,31,249,31,103,31,3,31,237,31,7,31,70,31,182,31,191,31,191,30,60,31,220,31,221,31,11,31,133,31,250,31,222,31,123,31,191,31,195,31,144,31,69,31,183,31,183,30,98,31,228,31,119,31,241,31,12,31,44,31,80,31,142,31,101,31,101,30,232,31,160,31,139,31,139,30,136,31,14,31,65,31,195,31,195,30,177,31,61,31,95,31,129,31,45,31,45,30,45,29,133,31,133,30,204,31,134,31,237,31,237,30,18,31,18,30,152,31,152,30,93,31,93,30,188,31,147,31,169,31,201,31,96,31,166,31,34,31,247,31,247,30,196,31,17,31,85,31,34,31,230,31,207,31,32,31,32,30,32,29,133,31,16,31,16,30,126,31,126,30,126,29,126,28,126,27,205,31,196,31,85,31,164,31,101,31,178,31,160,31,72,31,25,31,53,31,163,31,183,31,73,31,203,31,127,31,117,31,27,31,77,31,77,30,22,31,157,31,152,31,55,31,219,31,240,31,254,31,229,31,229,30,254,31,254,30,172,31,172,30,172,29,172,28,116,31,13,31,13,30,30,31,232,31,117,31,139,31,168,31,217,31,217,30,217,29,14,31,252,31,252,30,252,29,137,31,16,31,192,31,21,31,116,31,151,31,15,31,36,31,223,31,130,31,222,31,222,30,222,29,150,31,167,31,22,31,22,30,124,31,110,31,232,31,18,31,8,31,234,31,217,31,95,31,148,31,8,31,204,31,105,31,246,31,165,31,43,31,43,30,78,31,139,31,139,30,5,31,163,31,166,31,88,31,49,31,207,31,107,31,67,31,67,30,33,31,33,30,93,31,93,30,162,31,13,31,13,30,113,31,156,31,156,30,109,31,164,31,160,31,82,31,106,31,181,31,181,30,80,31,109,31,7,31,144,31,253,31,138,31,138,30,127,31,103,31,91,31,40,31,40,30,163,31,130,31,69,31,129,31,105,31,196,31,31,31,176,31,8,31,8,30,64,31,35,31,70,31,22,31,224,31,202,31,197,31,57,31,203,31,202,31,235,31,117,31,128,31,128,30,128,29,167,31,24,31,35,31,132,31,132,30,117,31,145,31,166,31,45,31,215,31,133,31,133,30,65,31,111,31,86,31,31,31,109,31,242,31,252,31,134,31,127,31,86,31,221,31,85,31,85,30,216,31,239,31,88,31,88,30,215,31,112,31,120,31,155,31,159,31,159,30,168,31,150,31,78,31,237,31,42,31,192,31,184,31,236,31,247,31,247,30,89,31,157,31,102,31,9,31,9,30,87,31,161,31,161,30,217,31,99,31,99,30,99,29,99,28,99,27,99,26,55,31,55,30,101,31,132,31,93,31,199,31,140,31,140,30,231,31,20,31,18,31,254,31,254,30,36,31,173,31,173,30,250,31,38,31,133,31,207,31,133,31,36,31,36,30,116,31,53,31,106,31,217,31,217,30,30,31,250,31,71,31,31,31,31,30,31,29,217,31,217,30,217,29,137,31,198,31,198,30,168,31,168,30,168,29,200,31,112,31,121,31,121,30,121,29,4,31,149,31,198,31,221,31,221,30,111,31,111,30,13,31,13,30,13,29,237,31,245,31,63,31,204,31,49,31,240,31,22,31,25,31,103,31,93,31,60,31,128,31,125,31,125,30,58,31,183,31,231,31,231,30,193,31,213,31,129,31,129,30,37,31,11,31,176,31,139,31,139,30,100,31,27,31,175,31,188,31,101,31,171,31,69,31,188,31,138,31,138,30,149,31,81,31,134,31,42,31,42,30,211,31,148,31,21,31,21,30,93,31,24,31,24,30,69,31,115,31,78,31,30,31,87,31,102,31,102,30,102,29,169,31,54,31,67,31,156,31,129,31,167,31,167,30,57,31,57,30,13,31,13,30,46,31,221,31,203,31,37,31,37,30,93,31,204,31,204,30,1,31,63,31,209,31,209,30,72,31,72,30,72,31,92,31,106,31,106,30,201,31,201,30,174,31,174,30,174,29,174,28,109,31,18,31,128,31,128,30,59,31,40,31,158,31,44,31,213,31,217,31,223,31,223,30,233,31,214,31,192,31,74,31,84,31,105,31,251,31,251,30,24,31,218,31,205,31,91,31,61,31,215,31,215,30,27,31,195,31,201,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
