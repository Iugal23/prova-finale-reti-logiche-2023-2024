-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_262 is
end project_tb_262;

architecture project_tb_arch_262 of project_tb_262 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 237;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,22,0,0,0,0,0,190,0,152,0,149,0,125,0,214,0,0,0,36,0,0,0,242,0,48,0,207,0,0,0,191,0,0,0,88,0,0,0,98,0,153,0,10,0,206,0,239,0,204,0,112,0,131,0,0,0,98,0,58,0,117,0,0,0,5,0,253,0,20,0,117,0,124,0,47,0,0,0,0,0,59,0,83,0,149,0,15,0,194,0,212,0,170,0,98,0,119,0,96,0,135,0,0,0,144,0,51,0,39,0,241,0,200,0,188,0,238,0,240,0,83,0,0,0,54,0,179,0,0,0,123,0,205,0,93,0,255,0,141,0,253,0,123,0,0,0,40,0,0,0,125,0,0,0,242,0,34,0,22,0,229,0,238,0,26,0,165,0,247,0,96,0,148,0,45,0,225,0,93,0,0,0,0,0,223,0,0,0,109,0,224,0,0,0,253,0,167,0,161,0,184,0,98,0,0,0,170,0,0,0,11,0,0,0,211,0,0,0,0,0,0,0,229,0,51,0,0,0,135,0,148,0,0,0,123,0,229,0,15,0,42,0,4,0,235,0,245,0,151,0,242,0,65,0,170,0,84,0,0,0,4,0,115,0,87,0,83,0,108,0,15,0,6,0,11,0,149,0,12,0,163,0,0,0,149,0,233,0,41,0,84,0,47,0,0,0,236,0,196,0,83,0,86,0,71,0,0,0,218,0,0,0,161,0,81,0,0,0,212,0,0,0,190,0,231,0,0,0,83,0,172,0,0,0,71,0,4,0,244,0,28,0,57,0,237,0,200,0,8,0,252,0,117,0,0,0,191,0,2,0,53,0,0,0,223,0,120,0,20,0,128,0,122,0,0,0,188,0,19,0,218,0,219,0,61,0,250,0,7,0,134,0,117,0,76,0,102,0,109,0,209,0,204,0,0,0,204,0,242,0,228,0,196,0,0,0,33,0,131,0,253,0,0,0,76,0,238,0,0,0,255,0,0,0,35,0,100,0,71,0,155,0,212,0,98,0,85,0,183,0,0,0,206,0,128,0,129,0,85,0,10,0,123,0,0,0,33,0,0,0,0,0);
signal scenario_full  : scenario_type := (128,31,22,31,22,30,22,29,190,31,152,31,149,31,125,31,214,31,214,30,36,31,36,30,242,31,48,31,207,31,207,30,191,31,191,30,88,31,88,30,98,31,153,31,10,31,206,31,239,31,204,31,112,31,131,31,131,30,98,31,58,31,117,31,117,30,5,31,253,31,20,31,117,31,124,31,47,31,47,30,47,29,59,31,83,31,149,31,15,31,194,31,212,31,170,31,98,31,119,31,96,31,135,31,135,30,144,31,51,31,39,31,241,31,200,31,188,31,238,31,240,31,83,31,83,30,54,31,179,31,179,30,123,31,205,31,93,31,255,31,141,31,253,31,123,31,123,30,40,31,40,30,125,31,125,30,242,31,34,31,22,31,229,31,238,31,26,31,165,31,247,31,96,31,148,31,45,31,225,31,93,31,93,30,93,29,223,31,223,30,109,31,224,31,224,30,253,31,167,31,161,31,184,31,98,31,98,30,170,31,170,30,11,31,11,30,211,31,211,30,211,29,211,28,229,31,51,31,51,30,135,31,148,31,148,30,123,31,229,31,15,31,42,31,4,31,235,31,245,31,151,31,242,31,65,31,170,31,84,31,84,30,4,31,115,31,87,31,83,31,108,31,15,31,6,31,11,31,149,31,12,31,163,31,163,30,149,31,233,31,41,31,84,31,47,31,47,30,236,31,196,31,83,31,86,31,71,31,71,30,218,31,218,30,161,31,81,31,81,30,212,31,212,30,190,31,231,31,231,30,83,31,172,31,172,30,71,31,4,31,244,31,28,31,57,31,237,31,200,31,8,31,252,31,117,31,117,30,191,31,2,31,53,31,53,30,223,31,120,31,20,31,128,31,122,31,122,30,188,31,19,31,218,31,219,31,61,31,250,31,7,31,134,31,117,31,76,31,102,31,109,31,209,31,204,31,204,30,204,31,242,31,228,31,196,31,196,30,33,31,131,31,253,31,253,30,76,31,238,31,238,30,255,31,255,30,35,31,100,31,71,31,155,31,212,31,98,31,85,31,183,31,183,30,206,31,128,31,129,31,85,31,10,31,123,31,123,30,33,31,33,30,33,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
