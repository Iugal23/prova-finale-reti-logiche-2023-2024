-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_83 is
end project_tb_83;

architecture project_tb_arch_83 of project_tb_83 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 493;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (79,0,236,0,137,0,220,0,147,0,134,0,240,0,206,0,2,0,0,0,189,0,233,0,189,0,63,0,135,0,217,0,0,0,153,0,174,0,96,0,91,0,41,0,73,0,32,0,1,0,131,0,239,0,121,0,136,0,39,0,19,0,180,0,158,0,50,0,253,0,48,0,84,0,248,0,0,0,71,0,0,0,184,0,184,0,87,0,178,0,40,0,0,0,63,0,114,0,122,0,234,0,113,0,94,0,249,0,242,0,82,0,185,0,23,0,0,0,74,0,181,0,122,0,155,0,119,0,122,0,66,0,223,0,166,0,154,0,142,0,108,0,0,0,58,0,17,0,26,0,202,0,108,0,121,0,107,0,0,0,82,0,210,0,22,0,255,0,240,0,140,0,25,0,244,0,207,0,216,0,161,0,125,0,32,0,152,0,180,0,114,0,210,0,250,0,134,0,97,0,131,0,237,0,171,0,144,0,181,0,30,0,45,0,248,0,71,0,203,0,135,0,188,0,0,0,60,0,249,0,249,0,19,0,71,0,18,0,0,0,0,0,11,0,0,0,69,0,76,0,94,0,83,0,179,0,234,0,0,0,82,0,15,0,246,0,0,0,207,0,230,0,191,0,134,0,0,0,67,0,232,0,247,0,170,0,65,0,0,0,7,0,62,0,49,0,0,0,40,0,183,0,140,0,98,0,212,0,166,0,182,0,65,0,164,0,118,0,0,0,86,0,86,0,156,0,63,0,17,0,84,0,113,0,0,0,192,0,191,0,70,0,102,0,249,0,163,0,66,0,46,0,0,0,238,0,110,0,174,0,71,0,244,0,80,0,0,0,0,0,30,0,49,0,146,0,189,0,80,0,231,0,75,0,0,0,79,0,146,0,92,0,62,0,0,0,104,0,116,0,9,0,220,0,245,0,49,0,6,0,71,0,129,0,0,0,28,0,101,0,224,0,0,0,0,0,0,0,0,0,79,0,56,0,9,0,60,0,101,0,27,0,213,0,194,0,67,0,162,0,0,0,253,0,24,0,234,0,63,0,171,0,47,0,12,0,120,0,178,0,40,0,26,0,0,0,55,0,133,0,198,0,0,0,2,0,207,0,12,0,230,0,220,0,0,0,0,0,245,0,240,0,0,0,225,0,0,0,163,0,208,0,187,0,75,0,74,0,0,0,36,0,139,0,186,0,229,0,0,0,132,0,0,0,179,0,0,0,0,0,0,0,12,0,192,0,121,0,169,0,0,0,125,0,89,0,248,0,193,0,0,0,172,0,207,0,150,0,139,0,176,0,206,0,31,0,9,0,158,0,0,0,139,0,21,0,192,0,128,0,92,0,27,0,110,0,39,0,40,0,65,0,53,0,0,0,0,0,241,0,0,0,107,0,0,0,183,0,0,0,135,0,98,0,160,0,191,0,157,0,204,0,68,0,124,0,71,0,98,0,10,0,101,0,216,0,67,0,0,0,195,0,234,0,200,0,0,0,0,0,119,0,162,0,0,0,123,0,216,0,0,0,200,0,86,0,0,0,156,0,0,0,0,0,62,0,26,0,0,0,57,0,168,0,191,0,0,0,117,0,12,0,85,0,19,0,153,0,0,0,159,0,0,0,116,0,67,0,25,0,139,0,201,0,136,0,0,0,243,0,205,0,21,0,182,0,131,0,79,0,0,0,0,0,251,0,126,0,0,0,207,0,230,0,121,0,19,0,0,0,0,0,0,0,189,0,168,0,165,0,14,0,0,0,130,0,191,0,0,0,198,0,0,0,250,0,161,0,189,0,4,0,0,0,197,0,212,0,117,0,220,0,53,0,0,0,0,0,166,0,169,0,96,0,226,0,183,0,182,0,159,0,25,0,0,0,72,0,149,0,179,0,0,0,0,0,99,0,204,0,53,0,79,0,255,0,0,0,234,0,110,0,21,0,0,0,161,0,27,0,214,0,124,0,144,0,21,0,57,0,251,0,212,0,245,0,237,0,10,0,41,0,83,0,202,0,125,0,27,0,162,0,1,0,10,0,0,0,79,0,216,0,0,0,49,0,92,0,143,0,136,0,0,0,0,0,13,0,254,0,154,0,92,0,174,0,38,0,235,0,86,0,53,0,0,0,105,0,9,0,0,0,11,0,33,0,0,0,187,0,87,0,63,0,78,0,234,0,46,0,0,0,116,0,140,0,173,0,110,0,227,0,148,0,109,0,0,0,169,0,4,0,179,0,238,0);
signal scenario_full  : scenario_type := (79,31,236,31,137,31,220,31,147,31,134,31,240,31,206,31,2,31,2,30,189,31,233,31,189,31,63,31,135,31,217,31,217,30,153,31,174,31,96,31,91,31,41,31,73,31,32,31,1,31,131,31,239,31,121,31,136,31,39,31,19,31,180,31,158,31,50,31,253,31,48,31,84,31,248,31,248,30,71,31,71,30,184,31,184,31,87,31,178,31,40,31,40,30,63,31,114,31,122,31,234,31,113,31,94,31,249,31,242,31,82,31,185,31,23,31,23,30,74,31,181,31,122,31,155,31,119,31,122,31,66,31,223,31,166,31,154,31,142,31,108,31,108,30,58,31,17,31,26,31,202,31,108,31,121,31,107,31,107,30,82,31,210,31,22,31,255,31,240,31,140,31,25,31,244,31,207,31,216,31,161,31,125,31,32,31,152,31,180,31,114,31,210,31,250,31,134,31,97,31,131,31,237,31,171,31,144,31,181,31,30,31,45,31,248,31,71,31,203,31,135,31,188,31,188,30,60,31,249,31,249,31,19,31,71,31,18,31,18,30,18,29,11,31,11,30,69,31,76,31,94,31,83,31,179,31,234,31,234,30,82,31,15,31,246,31,246,30,207,31,230,31,191,31,134,31,134,30,67,31,232,31,247,31,170,31,65,31,65,30,7,31,62,31,49,31,49,30,40,31,183,31,140,31,98,31,212,31,166,31,182,31,65,31,164,31,118,31,118,30,86,31,86,31,156,31,63,31,17,31,84,31,113,31,113,30,192,31,191,31,70,31,102,31,249,31,163,31,66,31,46,31,46,30,238,31,110,31,174,31,71,31,244,31,80,31,80,30,80,29,30,31,49,31,146,31,189,31,80,31,231,31,75,31,75,30,79,31,146,31,92,31,62,31,62,30,104,31,116,31,9,31,220,31,245,31,49,31,6,31,71,31,129,31,129,30,28,31,101,31,224,31,224,30,224,29,224,28,224,27,79,31,56,31,9,31,60,31,101,31,27,31,213,31,194,31,67,31,162,31,162,30,253,31,24,31,234,31,63,31,171,31,47,31,12,31,120,31,178,31,40,31,26,31,26,30,55,31,133,31,198,31,198,30,2,31,207,31,12,31,230,31,220,31,220,30,220,29,245,31,240,31,240,30,225,31,225,30,163,31,208,31,187,31,75,31,74,31,74,30,36,31,139,31,186,31,229,31,229,30,132,31,132,30,179,31,179,30,179,29,179,28,12,31,192,31,121,31,169,31,169,30,125,31,89,31,248,31,193,31,193,30,172,31,207,31,150,31,139,31,176,31,206,31,31,31,9,31,158,31,158,30,139,31,21,31,192,31,128,31,92,31,27,31,110,31,39,31,40,31,65,31,53,31,53,30,53,29,241,31,241,30,107,31,107,30,183,31,183,30,135,31,98,31,160,31,191,31,157,31,204,31,68,31,124,31,71,31,98,31,10,31,101,31,216,31,67,31,67,30,195,31,234,31,200,31,200,30,200,29,119,31,162,31,162,30,123,31,216,31,216,30,200,31,86,31,86,30,156,31,156,30,156,29,62,31,26,31,26,30,57,31,168,31,191,31,191,30,117,31,12,31,85,31,19,31,153,31,153,30,159,31,159,30,116,31,67,31,25,31,139,31,201,31,136,31,136,30,243,31,205,31,21,31,182,31,131,31,79,31,79,30,79,29,251,31,126,31,126,30,207,31,230,31,121,31,19,31,19,30,19,29,19,28,189,31,168,31,165,31,14,31,14,30,130,31,191,31,191,30,198,31,198,30,250,31,161,31,189,31,4,31,4,30,197,31,212,31,117,31,220,31,53,31,53,30,53,29,166,31,169,31,96,31,226,31,183,31,182,31,159,31,25,31,25,30,72,31,149,31,179,31,179,30,179,29,99,31,204,31,53,31,79,31,255,31,255,30,234,31,110,31,21,31,21,30,161,31,27,31,214,31,124,31,144,31,21,31,57,31,251,31,212,31,245,31,237,31,10,31,41,31,83,31,202,31,125,31,27,31,162,31,1,31,10,31,10,30,79,31,216,31,216,30,49,31,92,31,143,31,136,31,136,30,136,29,13,31,254,31,154,31,92,31,174,31,38,31,235,31,86,31,53,31,53,30,105,31,9,31,9,30,11,31,33,31,33,30,187,31,87,31,63,31,78,31,234,31,46,31,46,30,116,31,140,31,173,31,110,31,227,31,148,31,109,31,109,30,169,31,4,31,179,31,238,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
