-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_533 is
end project_tb_533;

architecture project_tb_arch_533 of project_tb_533 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 802;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (20,0,143,0,232,0,6,0,235,0,218,0,177,0,143,0,158,0,218,0,0,0,0,0,13,0,226,0,126,0,91,0,0,0,0,0,184,0,217,0,247,0,13,0,155,0,11,0,232,0,1,0,222,0,101,0,120,0,175,0,208,0,106,0,223,0,150,0,97,0,45,0,39,0,27,0,0,0,15,0,243,0,253,0,0,0,195,0,243,0,119,0,106,0,238,0,250,0,0,0,150,0,0,0,0,0,187,0,47,0,15,0,130,0,0,0,0,0,0,0,17,0,234,0,100,0,0,0,254,0,0,0,88,0,0,0,113,0,65,0,137,0,220,0,0,0,0,0,240,0,236,0,92,0,237,0,231,0,0,0,0,0,76,0,131,0,255,0,173,0,6,0,229,0,6,0,106,0,162,0,0,0,0,0,0,0,187,0,103,0,176,0,255,0,183,0,47,0,0,0,0,0,0,0,114,0,240,0,111,0,230,0,191,0,252,0,228,0,46,0,103,0,72,0,190,0,73,0,0,0,107,0,179,0,7,0,222,0,149,0,86,0,217,0,101,0,208,0,35,0,54,0,141,0,32,0,160,0,0,0,245,0,0,0,16,0,97,0,16,0,0,0,234,0,167,0,4,0,248,0,74,0,186,0,0,0,0,0,240,0,119,0,167,0,21,0,73,0,26,0,167,0,79,0,224,0,0,0,121,0,217,0,39,0,0,0,90,0,0,0,207,0,79,0,233,0,180,0,117,0,194,0,59,0,236,0,0,0,121,0,0,0,0,0,113,0,130,0,0,0,152,0,77,0,116,0,6,0,242,0,46,0,161,0,170,0,48,0,79,0,28,0,209,0,163,0,114,0,216,0,206,0,94,0,230,0,0,0,49,0,52,0,147,0,0,0,218,0,252,0,91,0,179,0,0,0,194,0,0,0,252,0,0,0,163,0,53,0,33,0,59,0,5,0,22,0,228,0,184,0,0,0,161,0,38,0,191,0,114,0,33,0,186,0,48,0,145,0,251,0,194,0,232,0,96,0,12,0,57,0,242,0,165,0,255,0,198,0,242,0,8,0,0,0,30,0,221,0,183,0,226,0,67,0,0,0,184,0,65,0,48,0,4,0,0,0,0,0,253,0,214,0,0,0,0,0,225,0,0,0,53,0,0,0,138,0,49,0,228,0,232,0,197,0,83,0,141,0,132,0,191,0,97,0,0,0,0,0,135,0,0,0,136,0,79,0,0,0,243,0,104,0,0,0,184,0,178,0,26,0,147,0,29,0,24,0,236,0,223,0,234,0,77,0,212,0,20,0,45,0,109,0,0,0,143,0,0,0,144,0,216,0,34,0,70,0,96,0,0,0,7,0,69,0,100,0,189,0,30,0,88,0,142,0,229,0,0,0,164,0,64,0,174,0,184,0,79,0,249,0,71,0,240,0,3,0,226,0,49,0,143,0,187,0,154,0,172,0,23,0,200,0,217,0,69,0,0,0,208,0,107,0,134,0,5,0,0,0,27,0,79,0,0,0,60,0,176,0,177,0,65,0,77,0,130,0,74,0,52,0,3,0,214,0,0,0,40,0,0,0,154,0,0,0,210,0,228,0,35,0,79,0,0,0,169,0,204,0,18,0,0,0,77,0,0,0,8,0,218,0,247,0,0,0,221,0,212,0,70,0,241,0,224,0,25,0,0,0,11,0,21,0,0,0,246,0,53,0,0,0,213,0,12,0,0,0,0,0,197,0,0,0,18,0,33,0,227,0,233,0,79,0,0,0,0,0,43,0,0,0,112,0,0,0,193,0,2,0,50,0,69,0,210,0,68,0,144,0,135,0,175,0,107,0,171,0,103,0,43,0,20,0,111,0,0,0,132,0,230,0,0,0,0,0,0,0,149,0,0,0,81,0,75,0,0,0,50,0,227,0,55,0,31,0,0,0,105,0,214,0,214,0,119,0,137,0,21,0,124,0,142,0,40,0,199,0,197,0,11,0,62,0,134,0,0,0,65,0,174,0,171,0,153,0,240,0,226,0,75,0,139,0,121,0,129,0,0,0,87,0,0,0,119,0,109,0,217,0,4,0,0,0,252,0,9,0,141,0,0,0,143,0,97,0,0,0,37,0,0,0,230,0,95,0,165,0,9,0,0,0,254,0,176,0,11,0,171,0,49,0,0,0,100,0,134,0,196,0,0,0,160,0,0,0,36,0,122,0,0,0,252,0,149,0,0,0,210,0,9,0,0,0,193,0,133,0,113,0,97,0,98,0,225,0,113,0,97,0,109,0,0,0,223,0,124,0,0,0,115,0,138,0,118,0,192,0,97,0,0,0,65,0,36,0,194,0,207,0,205,0,73,0,142,0,0,0,0,0,0,0,120,0,91,0,0,0,193,0,72,0,190,0,0,0,24,0,255,0,98,0,229,0,71,0,123,0,24,0,24,0,0,0,0,0,48,0,173,0,235,0,241,0,146,0,90,0,0,0,105,0,66,0,11,0,198,0,38,0,103,0,16,0,242,0,129,0,224,0,106,0,111,0,234,0,201,0,0,0,227,0,170,0,223,0,199,0,0,0,79,0,0,0,80,0,154,0,101,0,0,0,47,0,0,0,0,0,0,0,70,0,3,0,105,0,73,0,141,0,0,0,0,0,84,0,0,0,94,0,198,0,31,0,191,0,226,0,54,0,78,0,0,0,54,0,166,0,163,0,4,0,0,0,0,0,0,0,0,0,204,0,167,0,0,0,236,0,0,0,213,0,0,0,117,0,220,0,14,0,163,0,0,0,32,0,67,0,191,0,103,0,203,0,186,0,252,0,209,0,0,0,217,0,163,0,131,0,223,0,224,0,199,0,72,0,0,0,158,0,0,0,33,0,209,0,145,0,99,0,0,0,230,0,0,0,46,0,188,0,121,0,0,0,194,0,199,0,0,0,242,0,252,0,168,0,92,0,0,0,0,0,0,0,191,0,207,0,74,0,60,0,11,0,66,0,203,0,78,0,92,0,164,0,137,0,120,0,40,0,124,0,145,0,0,0,0,0,177,0,180,0,192,0,8,0,23,0,183,0,0,0,54,0,35,0,0,0,0,0,0,0,195,0,23,0,129,0,118,0,0,0,245,0,145,0,189,0,0,0,112,0,156,0,83,0,73,0,134,0,72,0,0,0,147,0,1,0,0,0,27,0,0,0,254,0,8,0,0,0,0,0,148,0,133,0,154,0,108,0,79,0,69,0,121,0,17,0,187,0,110,0,88,0,182,0,52,0,159,0,93,0,227,0,195,0,142,0,226,0,0,0,163,0,0,0,142,0,209,0,205,0,0,0,0,0,0,0,62,0,0,0,159,0,73,0,216,0,184,0,221,0,20,0,15,0,101,0,252,0,173,0,127,0,224,0,0,0,25,0,252,0,0,0,133,0,223,0,0,0,0,0,43,0,150,0,0,0,37,0,13,0,129,0,39,0,29,0,93,0,109,0,149,0,152,0,123,0,9,0,171,0,164,0,0,0,64,0,129,0,0,0,0,0,72,0,158,0,226,0,152,0,0,0,185,0,0,0,106,0,123,0,0,0,214,0,0,0,0,0,79,0,242,0,0,0,33,0,137,0,222,0,17,0,252,0);
signal scenario_full  : scenario_type := (20,31,143,31,232,31,6,31,235,31,218,31,177,31,143,31,158,31,218,31,218,30,218,29,13,31,226,31,126,31,91,31,91,30,91,29,184,31,217,31,247,31,13,31,155,31,11,31,232,31,1,31,222,31,101,31,120,31,175,31,208,31,106,31,223,31,150,31,97,31,45,31,39,31,27,31,27,30,15,31,243,31,253,31,253,30,195,31,243,31,119,31,106,31,238,31,250,31,250,30,150,31,150,30,150,29,187,31,47,31,15,31,130,31,130,30,130,29,130,28,17,31,234,31,100,31,100,30,254,31,254,30,88,31,88,30,113,31,65,31,137,31,220,31,220,30,220,29,240,31,236,31,92,31,237,31,231,31,231,30,231,29,76,31,131,31,255,31,173,31,6,31,229,31,6,31,106,31,162,31,162,30,162,29,162,28,187,31,103,31,176,31,255,31,183,31,47,31,47,30,47,29,47,28,114,31,240,31,111,31,230,31,191,31,252,31,228,31,46,31,103,31,72,31,190,31,73,31,73,30,107,31,179,31,7,31,222,31,149,31,86,31,217,31,101,31,208,31,35,31,54,31,141,31,32,31,160,31,160,30,245,31,245,30,16,31,97,31,16,31,16,30,234,31,167,31,4,31,248,31,74,31,186,31,186,30,186,29,240,31,119,31,167,31,21,31,73,31,26,31,167,31,79,31,224,31,224,30,121,31,217,31,39,31,39,30,90,31,90,30,207,31,79,31,233,31,180,31,117,31,194,31,59,31,236,31,236,30,121,31,121,30,121,29,113,31,130,31,130,30,152,31,77,31,116,31,6,31,242,31,46,31,161,31,170,31,48,31,79,31,28,31,209,31,163,31,114,31,216,31,206,31,94,31,230,31,230,30,49,31,52,31,147,31,147,30,218,31,252,31,91,31,179,31,179,30,194,31,194,30,252,31,252,30,163,31,53,31,33,31,59,31,5,31,22,31,228,31,184,31,184,30,161,31,38,31,191,31,114,31,33,31,186,31,48,31,145,31,251,31,194,31,232,31,96,31,12,31,57,31,242,31,165,31,255,31,198,31,242,31,8,31,8,30,30,31,221,31,183,31,226,31,67,31,67,30,184,31,65,31,48,31,4,31,4,30,4,29,253,31,214,31,214,30,214,29,225,31,225,30,53,31,53,30,138,31,49,31,228,31,232,31,197,31,83,31,141,31,132,31,191,31,97,31,97,30,97,29,135,31,135,30,136,31,79,31,79,30,243,31,104,31,104,30,184,31,178,31,26,31,147,31,29,31,24,31,236,31,223,31,234,31,77,31,212,31,20,31,45,31,109,31,109,30,143,31,143,30,144,31,216,31,34,31,70,31,96,31,96,30,7,31,69,31,100,31,189,31,30,31,88,31,142,31,229,31,229,30,164,31,64,31,174,31,184,31,79,31,249,31,71,31,240,31,3,31,226,31,49,31,143,31,187,31,154,31,172,31,23,31,200,31,217,31,69,31,69,30,208,31,107,31,134,31,5,31,5,30,27,31,79,31,79,30,60,31,176,31,177,31,65,31,77,31,130,31,74,31,52,31,3,31,214,31,214,30,40,31,40,30,154,31,154,30,210,31,228,31,35,31,79,31,79,30,169,31,204,31,18,31,18,30,77,31,77,30,8,31,218,31,247,31,247,30,221,31,212,31,70,31,241,31,224,31,25,31,25,30,11,31,21,31,21,30,246,31,53,31,53,30,213,31,12,31,12,30,12,29,197,31,197,30,18,31,33,31,227,31,233,31,79,31,79,30,79,29,43,31,43,30,112,31,112,30,193,31,2,31,50,31,69,31,210,31,68,31,144,31,135,31,175,31,107,31,171,31,103,31,43,31,20,31,111,31,111,30,132,31,230,31,230,30,230,29,230,28,149,31,149,30,81,31,75,31,75,30,50,31,227,31,55,31,31,31,31,30,105,31,214,31,214,31,119,31,137,31,21,31,124,31,142,31,40,31,199,31,197,31,11,31,62,31,134,31,134,30,65,31,174,31,171,31,153,31,240,31,226,31,75,31,139,31,121,31,129,31,129,30,87,31,87,30,119,31,109,31,217,31,4,31,4,30,252,31,9,31,141,31,141,30,143,31,97,31,97,30,37,31,37,30,230,31,95,31,165,31,9,31,9,30,254,31,176,31,11,31,171,31,49,31,49,30,100,31,134,31,196,31,196,30,160,31,160,30,36,31,122,31,122,30,252,31,149,31,149,30,210,31,9,31,9,30,193,31,133,31,113,31,97,31,98,31,225,31,113,31,97,31,109,31,109,30,223,31,124,31,124,30,115,31,138,31,118,31,192,31,97,31,97,30,65,31,36,31,194,31,207,31,205,31,73,31,142,31,142,30,142,29,142,28,120,31,91,31,91,30,193,31,72,31,190,31,190,30,24,31,255,31,98,31,229,31,71,31,123,31,24,31,24,31,24,30,24,29,48,31,173,31,235,31,241,31,146,31,90,31,90,30,105,31,66,31,11,31,198,31,38,31,103,31,16,31,242,31,129,31,224,31,106,31,111,31,234,31,201,31,201,30,227,31,170,31,223,31,199,31,199,30,79,31,79,30,80,31,154,31,101,31,101,30,47,31,47,30,47,29,47,28,70,31,3,31,105,31,73,31,141,31,141,30,141,29,84,31,84,30,94,31,198,31,31,31,191,31,226,31,54,31,78,31,78,30,54,31,166,31,163,31,4,31,4,30,4,29,4,28,4,27,204,31,167,31,167,30,236,31,236,30,213,31,213,30,117,31,220,31,14,31,163,31,163,30,32,31,67,31,191,31,103,31,203,31,186,31,252,31,209,31,209,30,217,31,163,31,131,31,223,31,224,31,199,31,72,31,72,30,158,31,158,30,33,31,209,31,145,31,99,31,99,30,230,31,230,30,46,31,188,31,121,31,121,30,194,31,199,31,199,30,242,31,252,31,168,31,92,31,92,30,92,29,92,28,191,31,207,31,74,31,60,31,11,31,66,31,203,31,78,31,92,31,164,31,137,31,120,31,40,31,124,31,145,31,145,30,145,29,177,31,180,31,192,31,8,31,23,31,183,31,183,30,54,31,35,31,35,30,35,29,35,28,195,31,23,31,129,31,118,31,118,30,245,31,145,31,189,31,189,30,112,31,156,31,83,31,73,31,134,31,72,31,72,30,147,31,1,31,1,30,27,31,27,30,254,31,8,31,8,30,8,29,148,31,133,31,154,31,108,31,79,31,69,31,121,31,17,31,187,31,110,31,88,31,182,31,52,31,159,31,93,31,227,31,195,31,142,31,226,31,226,30,163,31,163,30,142,31,209,31,205,31,205,30,205,29,205,28,62,31,62,30,159,31,73,31,216,31,184,31,221,31,20,31,15,31,101,31,252,31,173,31,127,31,224,31,224,30,25,31,252,31,252,30,133,31,223,31,223,30,223,29,43,31,150,31,150,30,37,31,13,31,129,31,39,31,29,31,93,31,109,31,149,31,152,31,123,31,9,31,171,31,164,31,164,30,64,31,129,31,129,30,129,29,72,31,158,31,226,31,152,31,152,30,185,31,185,30,106,31,123,31,123,30,214,31,214,30,214,29,79,31,242,31,242,30,33,31,137,31,222,31,17,31,252,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
