-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 272;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,89,0,150,0,43,0,225,0,124,0,0,0,65,0,0,0,225,0,168,0,244,0,172,0,193,0,144,0,139,0,190,0,57,0,0,0,238,0,197,0,102,0,2,0,173,0,242,0,19,0,109,0,190,0,160,0,26,0,0,0,188,0,252,0,174,0,211,0,81,0,49,0,0,0,238,0,32,0,72,0,249,0,195,0,0,0,149,0,29,0,216,0,99,0,241,0,23,0,0,0,10,0,54,0,0,0,243,0,82,0,215,0,43,0,150,0,190,0,224,0,214,0,42,0,11,0,182,0,198,0,69,0,78,0,0,0,225,0,46,0,145,0,0,0,43,0,0,0,0,0,16,0,0,0,117,0,70,0,0,0,70,0,0,0,0,0,160,0,116,0,0,0,13,0,241,0,0,0,98,0,76,0,70,0,236,0,203,0,11,0,195,0,214,0,162,0,253,0,134,0,82,0,236,0,247,0,92,0,187,0,173,0,0,0,250,0,158,0,207,0,230,0,121,0,203,0,130,0,0,0,193,0,146,0,0,0,202,0,61,0,131,0,209,0,178,0,31,0,0,0,197,0,88,0,0,0,99,0,74,0,174,0,0,0,18,0,0,0,191,0,218,0,102,0,67,0,135,0,160,0,88,0,124,0,229,0,51,0,158,0,0,0,240,0,190,0,0,0,43,0,30,0,122,0,86,0,249,0,145,0,23,0,0,0,153,0,138,0,165,0,33,0,61,0,147,0,57,0,0,0,153,0,36,0,42,0,181,0,97,0,7,0,91,0,157,0,197,0,201,0,95,0,0,0,121,0,0,0,0,0,44,0,1,0,3,0,53,0,0,0,188,0,215,0,245,0,172,0,147,0,224,0,102,0,248,0,3,0,97,0,87,0,26,0,66,0,239,0,216,0,0,0,240,0,233,0,235,0,183,0,198,0,33,0,0,0,0,0,167,0,236,0,105,0,0,0,0,0,178,0,206,0,98,0,128,0,148,0,63,0,172,0,189,0,67,0,0,0,172,0,148,0,21,0,213,0,245,0,148,0,20,0,116,0,120,0,127,0,228,0,62,0,0,0,92,0,206,0,97,0,234,0,101,0,90,0,143,0,220,0,207,0,85,0,51,0,0,0,188,0,205,0,0,0,139,0,114,0,178,0,225,0,178,0,126,0,0,0,167,0,230,0,0,0,0,0,2,0,67,0,243,0,182,0,65,0,100,0,0,0,0,0);
signal scenario_full  : scenario_type := (102,31,89,31,150,31,43,31,225,31,124,31,124,30,65,31,65,30,225,31,168,31,244,31,172,31,193,31,144,31,139,31,190,31,57,31,57,30,238,31,197,31,102,31,2,31,173,31,242,31,19,31,109,31,190,31,160,31,26,31,26,30,188,31,252,31,174,31,211,31,81,31,49,31,49,30,238,31,32,31,72,31,249,31,195,31,195,30,149,31,29,31,216,31,99,31,241,31,23,31,23,30,10,31,54,31,54,30,243,31,82,31,215,31,43,31,150,31,190,31,224,31,214,31,42,31,11,31,182,31,198,31,69,31,78,31,78,30,225,31,46,31,145,31,145,30,43,31,43,30,43,29,16,31,16,30,117,31,70,31,70,30,70,31,70,30,70,29,160,31,116,31,116,30,13,31,241,31,241,30,98,31,76,31,70,31,236,31,203,31,11,31,195,31,214,31,162,31,253,31,134,31,82,31,236,31,247,31,92,31,187,31,173,31,173,30,250,31,158,31,207,31,230,31,121,31,203,31,130,31,130,30,193,31,146,31,146,30,202,31,61,31,131,31,209,31,178,31,31,31,31,30,197,31,88,31,88,30,99,31,74,31,174,31,174,30,18,31,18,30,191,31,218,31,102,31,67,31,135,31,160,31,88,31,124,31,229,31,51,31,158,31,158,30,240,31,190,31,190,30,43,31,30,31,122,31,86,31,249,31,145,31,23,31,23,30,153,31,138,31,165,31,33,31,61,31,147,31,57,31,57,30,153,31,36,31,42,31,181,31,97,31,7,31,91,31,157,31,197,31,201,31,95,31,95,30,121,31,121,30,121,29,44,31,1,31,3,31,53,31,53,30,188,31,215,31,245,31,172,31,147,31,224,31,102,31,248,31,3,31,97,31,87,31,26,31,66,31,239,31,216,31,216,30,240,31,233,31,235,31,183,31,198,31,33,31,33,30,33,29,167,31,236,31,105,31,105,30,105,29,178,31,206,31,98,31,128,31,148,31,63,31,172,31,189,31,67,31,67,30,172,31,148,31,21,31,213,31,245,31,148,31,20,31,116,31,120,31,127,31,228,31,62,31,62,30,92,31,206,31,97,31,234,31,101,31,90,31,143,31,220,31,207,31,85,31,51,31,51,30,188,31,205,31,205,30,139,31,114,31,178,31,225,31,178,31,126,31,126,30,167,31,230,31,230,30,230,29,2,31,67,31,243,31,182,31,65,31,100,31,100,30,100,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
