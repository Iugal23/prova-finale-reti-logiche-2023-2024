-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_802 is
end project_tb_802;

architecture project_tb_arch_802 of project_tb_802 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 705;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,47,0,89,0,0,0,150,0,166,0,133,0,157,0,130,0,44,0,42,0,0,0,29,0,242,0,191,0,0,0,40,0,229,0,121,0,99,0,25,0,218,0,22,0,70,0,0,0,0,0,95,0,249,0,42,0,0,0,145,0,171,0,43,0,0,0,76,0,58,0,0,0,48,0,64,0,251,0,109,0,12,0,140,0,145,0,0,0,0,0,0,0,90,0,0,0,253,0,40,0,8,0,0,0,5,0,212,0,199,0,2,0,0,0,79,0,20,0,107,0,69,0,58,0,0,0,0,0,57,0,42,0,6,0,90,0,94,0,230,0,163,0,186,0,7,0,0,0,31,0,242,0,220,0,117,0,149,0,171,0,0,0,0,0,40,0,0,0,252,0,195,0,203,0,100,0,0,0,9,0,42,0,232,0,138,0,194,0,157,0,0,0,190,0,215,0,0,0,187,0,0,0,141,0,195,0,15,0,0,0,61,0,0,0,36,0,253,0,0,0,131,0,0,0,0,0,114,0,162,0,85,0,0,0,119,0,35,0,35,0,126,0,206,0,80,0,240,0,140,0,134,0,67,0,0,0,58,0,136,0,250,0,97,0,148,0,112,0,35,0,0,0,215,0,202,0,245,0,0,0,141,0,61,0,99,0,23,0,4,0,30,0,147,0,233,0,100,0,19,0,172,0,0,0,118,0,0,0,228,0,72,0,226,0,0,0,74,0,225,0,239,0,200,0,222,0,83,0,70,0,30,0,70,0,14,0,75,0,34,0,143,0,119,0,134,0,60,0,246,0,81,0,39,0,0,0,7,0,114,0,78,0,5,0,240,0,65,0,0,0,0,0,30,0,0,0,1,0,191,0,0,0,0,0,18,0,156,0,158,0,161,0,84,0,156,0,122,0,245,0,209,0,4,0,18,0,62,0,205,0,0,0,177,0,131,0,209,0,5,0,0,0,6,0,253,0,43,0,87,0,56,0,70,0,0,0,47,0,253,0,0,0,74,0,0,0,0,0,0,0,116,0,0,0,98,0,142,0,33,0,26,0,87,0,131,0,229,0,0,0,40,0,107,0,173,0,229,0,78,0,0,0,149,0,244,0,139,0,113,0,97,0,149,0,170,0,0,0,50,0,182,0,59,0,0,0,206,0,255,0,255,0,228,0,238,0,0,0,107,0,215,0,70,0,203,0,43,0,27,0,25,0,249,0,0,0,25,0,72,0,4,0,115,0,75,0,242,0,0,0,0,0,74,0,94,0,182,0,237,0,30,0,155,0,0,0,107,0,94,0,235,0,0,0,0,0,145,0,225,0,115,0,217,0,0,0,132,0,6,0,164,0,0,0,186,0,0,0,66,0,139,0,254,0,24,0,0,0,0,0,95,0,185,0,114,0,76,0,9,0,170,0,240,0,37,0,96,0,35,0,146,0,248,0,248,0,62,0,87,0,143,0,84,0,153,0,59,0,94,0,111,0,69,0,61,0,0,0,20,0,51,0,0,0,152,0,176,0,0,0,155,0,0,0,48,0,144,0,30,0,36,0,8,0,252,0,219,0,0,0,0,0,0,0,249,0,202,0,31,0,10,0,0,0,0,0,76,0,55,0,0,0,132,0,118,0,55,0,0,0,154,0,157,0,162,0,136,0,103,0,172,0,58,0,128,0,205,0,76,0,61,0,0,0,0,0,0,0,0,0,87,0,117,0,0,0,144,0,20,0,10,0,4,0,79,0,100,0,221,0,146,0,3,0,0,0,0,0,15,0,30,0,226,0,141,0,84,0,0,0,53,0,241,0,0,0,169,0,212,0,252,0,141,0,83,0,185,0,173,0,0,0,246,0,216,0,233,0,0,0,159,0,233,0,38,0,143,0,51,0,0,0,242,0,55,0,0,0,72,0,111,0,84,0,146,0,140,0,118,0,15,0,62,0,152,0,234,0,105,0,123,0,208,0,0,0,150,0,156,0,49,0,6,0,0,0,0,0,0,0,185,0,171,0,126,0,233,0,255,0,88,0,72,0,0,0,201,0,0,0,179,0,155,0,0,0,1,0,227,0,81,0,33,0,112,0,176,0,255,0,182,0,198,0,0,0,250,0,30,0,0,0,85,0,39,0,95,0,0,0,153,0,66,0,210,0,110,0,168,0,0,0,189,0,99,0,88,0,18,0,0,0,80,0,184,0,237,0,168,0,195,0,187,0,34,0,134,0,35,0,175,0,246,0,52,0,156,0,0,0,71,0,0,0,0,0,0,0,39,0,0,0,0,0,246,0,123,0,107,0,201,0,179,0,0,0,29,0,141,0,253,0,161,0,0,0,95,0,160,0,206,0,0,0,51,0,0,0,202,0,88,0,113,0,65,0,0,0,149,0,0,0,121,0,0,0,83,0,228,0,108,0,241,0,39,0,57,0,218,0,87,0,0,0,145,0,0,0,76,0,250,0,204,0,51,0,255,0,0,0,45,0,53,0,79,0,135,0,88,0,150,0,215,0,117,0,46,0,166,0,243,0,232,0,195,0,4,0,52,0,228,0,108,0,75,0,244,0,90,0,0,0,0,0,92,0,0,0,149,0,0,0,67,0,82,0,0,0,226,0,120,0,0,0,179,0,20,0,164,0,100,0,127,0,250,0,39,0,216,0,62,0,56,0,0,0,117,0,22,0,0,0,0,0,48,0,77,0,0,0,0,0,206,0,29,0,115,0,185,0,170,0,0,0,0,0,243,0,21,0,65,0,217,0,199,0,202,0,0,0,169,0,196,0,129,0,91,0,100,0,0,0,47,0,10,0,0,0,110,0,0,0,29,0,164,0,0,0,47,0,35,0,16,0,112,0,0,0,0,0,135,0,44,0,147,0,247,0,229,0,212,0,0,0,65,0,176,0,135,0,153,0,236,0,124,0,60,0,0,0,105,0,239,0,95,0,164,0,130,0,102,0,81,0,182,0,133,0,51,0,20,0,0,0,22,0,0,0,41,0,38,0,230,0,63,0,0,0,0,0,32,0,127,0,241,0,96,0,0,0,219,0,0,0,3,0,166,0,23,0,0,0,0,0,155,0,176,0,50,0,49,0,0,0,16,0,193,0,181,0,104,0,51,0,0,0,52,0,5,0,182,0,90,0,253,0,0,0,195,0,131,0,55,0,232,0,216,0,0,0,5,0,0,0,0,0,129,0);
signal scenario_full  : scenario_type := (0,0,47,31,89,31,89,30,150,31,166,31,133,31,157,31,130,31,44,31,42,31,42,30,29,31,242,31,191,31,191,30,40,31,229,31,121,31,99,31,25,31,218,31,22,31,70,31,70,30,70,29,95,31,249,31,42,31,42,30,145,31,171,31,43,31,43,30,76,31,58,31,58,30,48,31,64,31,251,31,109,31,12,31,140,31,145,31,145,30,145,29,145,28,90,31,90,30,253,31,40,31,8,31,8,30,5,31,212,31,199,31,2,31,2,30,79,31,20,31,107,31,69,31,58,31,58,30,58,29,57,31,42,31,6,31,90,31,94,31,230,31,163,31,186,31,7,31,7,30,31,31,242,31,220,31,117,31,149,31,171,31,171,30,171,29,40,31,40,30,252,31,195,31,203,31,100,31,100,30,9,31,42,31,232,31,138,31,194,31,157,31,157,30,190,31,215,31,215,30,187,31,187,30,141,31,195,31,15,31,15,30,61,31,61,30,36,31,253,31,253,30,131,31,131,30,131,29,114,31,162,31,85,31,85,30,119,31,35,31,35,31,126,31,206,31,80,31,240,31,140,31,134,31,67,31,67,30,58,31,136,31,250,31,97,31,148,31,112,31,35,31,35,30,215,31,202,31,245,31,245,30,141,31,61,31,99,31,23,31,4,31,30,31,147,31,233,31,100,31,19,31,172,31,172,30,118,31,118,30,228,31,72,31,226,31,226,30,74,31,225,31,239,31,200,31,222,31,83,31,70,31,30,31,70,31,14,31,75,31,34,31,143,31,119,31,134,31,60,31,246,31,81,31,39,31,39,30,7,31,114,31,78,31,5,31,240,31,65,31,65,30,65,29,30,31,30,30,1,31,191,31,191,30,191,29,18,31,156,31,158,31,161,31,84,31,156,31,122,31,245,31,209,31,4,31,18,31,62,31,205,31,205,30,177,31,131,31,209,31,5,31,5,30,6,31,253,31,43,31,87,31,56,31,70,31,70,30,47,31,253,31,253,30,74,31,74,30,74,29,74,28,116,31,116,30,98,31,142,31,33,31,26,31,87,31,131,31,229,31,229,30,40,31,107,31,173,31,229,31,78,31,78,30,149,31,244,31,139,31,113,31,97,31,149,31,170,31,170,30,50,31,182,31,59,31,59,30,206,31,255,31,255,31,228,31,238,31,238,30,107,31,215,31,70,31,203,31,43,31,27,31,25,31,249,31,249,30,25,31,72,31,4,31,115,31,75,31,242,31,242,30,242,29,74,31,94,31,182,31,237,31,30,31,155,31,155,30,107,31,94,31,235,31,235,30,235,29,145,31,225,31,115,31,217,31,217,30,132,31,6,31,164,31,164,30,186,31,186,30,66,31,139,31,254,31,24,31,24,30,24,29,95,31,185,31,114,31,76,31,9,31,170,31,240,31,37,31,96,31,35,31,146,31,248,31,248,31,62,31,87,31,143,31,84,31,153,31,59,31,94,31,111,31,69,31,61,31,61,30,20,31,51,31,51,30,152,31,176,31,176,30,155,31,155,30,48,31,144,31,30,31,36,31,8,31,252,31,219,31,219,30,219,29,219,28,249,31,202,31,31,31,10,31,10,30,10,29,76,31,55,31,55,30,132,31,118,31,55,31,55,30,154,31,157,31,162,31,136,31,103,31,172,31,58,31,128,31,205,31,76,31,61,31,61,30,61,29,61,28,61,27,87,31,117,31,117,30,144,31,20,31,10,31,4,31,79,31,100,31,221,31,146,31,3,31,3,30,3,29,15,31,30,31,226,31,141,31,84,31,84,30,53,31,241,31,241,30,169,31,212,31,252,31,141,31,83,31,185,31,173,31,173,30,246,31,216,31,233,31,233,30,159,31,233,31,38,31,143,31,51,31,51,30,242,31,55,31,55,30,72,31,111,31,84,31,146,31,140,31,118,31,15,31,62,31,152,31,234,31,105,31,123,31,208,31,208,30,150,31,156,31,49,31,6,31,6,30,6,29,6,28,185,31,171,31,126,31,233,31,255,31,88,31,72,31,72,30,201,31,201,30,179,31,155,31,155,30,1,31,227,31,81,31,33,31,112,31,176,31,255,31,182,31,198,31,198,30,250,31,30,31,30,30,85,31,39,31,95,31,95,30,153,31,66,31,210,31,110,31,168,31,168,30,189,31,99,31,88,31,18,31,18,30,80,31,184,31,237,31,168,31,195,31,187,31,34,31,134,31,35,31,175,31,246,31,52,31,156,31,156,30,71,31,71,30,71,29,71,28,39,31,39,30,39,29,246,31,123,31,107,31,201,31,179,31,179,30,29,31,141,31,253,31,161,31,161,30,95,31,160,31,206,31,206,30,51,31,51,30,202,31,88,31,113,31,65,31,65,30,149,31,149,30,121,31,121,30,83,31,228,31,108,31,241,31,39,31,57,31,218,31,87,31,87,30,145,31,145,30,76,31,250,31,204,31,51,31,255,31,255,30,45,31,53,31,79,31,135,31,88,31,150,31,215,31,117,31,46,31,166,31,243,31,232,31,195,31,4,31,52,31,228,31,108,31,75,31,244,31,90,31,90,30,90,29,92,31,92,30,149,31,149,30,67,31,82,31,82,30,226,31,120,31,120,30,179,31,20,31,164,31,100,31,127,31,250,31,39,31,216,31,62,31,56,31,56,30,117,31,22,31,22,30,22,29,48,31,77,31,77,30,77,29,206,31,29,31,115,31,185,31,170,31,170,30,170,29,243,31,21,31,65,31,217,31,199,31,202,31,202,30,169,31,196,31,129,31,91,31,100,31,100,30,47,31,10,31,10,30,110,31,110,30,29,31,164,31,164,30,47,31,35,31,16,31,112,31,112,30,112,29,135,31,44,31,147,31,247,31,229,31,212,31,212,30,65,31,176,31,135,31,153,31,236,31,124,31,60,31,60,30,105,31,239,31,95,31,164,31,130,31,102,31,81,31,182,31,133,31,51,31,20,31,20,30,22,31,22,30,41,31,38,31,230,31,63,31,63,30,63,29,32,31,127,31,241,31,96,31,96,30,219,31,219,30,3,31,166,31,23,31,23,30,23,29,155,31,176,31,50,31,49,31,49,30,16,31,193,31,181,31,104,31,51,31,51,30,52,31,5,31,182,31,90,31,253,31,253,30,195,31,131,31,55,31,232,31,216,31,216,30,5,31,5,30,5,29,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
