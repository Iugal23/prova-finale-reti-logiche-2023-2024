-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 959;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,205,0,4,0,106,0,158,0,248,0,218,0,20,0,140,0,252,0,188,0,153,0,0,0,152,0,16,0,147,0,97,0,4,0,23,0,14,0,0,0,129,0,12,0,0,0,0,0,0,0,162,0,0,0,192,0,116,0,1,0,152,0,227,0,0,0,0,0,30,0,54,0,216,0,123,0,17,0,0,0,109,0,176,0,59,0,0,0,220,0,159,0,249,0,232,0,5,0,0,0,0,0,233,0,110,0,226,0,0,0,231,0,0,0,250,0,96,0,122,0,206,0,6,0,160,0,250,0,184,0,0,0,66,0,0,0,156,0,73,0,125,0,174,0,0,0,202,0,140,0,0,0,0,0,210,0,23,0,0,0,3,0,132,0,0,0,0,0,150,0,194,0,0,0,167,0,132,0,0,0,203,0,196,0,39,0,246,0,61,0,206,0,190,0,144,0,72,0,0,0,189,0,29,0,80,0,0,0,39,0,0,0,158,0,86,0,228,0,211,0,251,0,95,0,238,0,0,0,0,0,250,0,177,0,0,0,185,0,0,0,0,0,216,0,191,0,5,0,123,0,167,0,81,0,70,0,192,0,127,0,156,0,106,0,110,0,0,0,212,0,0,0,142,0,176,0,194,0,156,0,16,0,212,0,72,0,57,0,196,0,50,0,206,0,74,0,242,0,0,0,119,0,0,0,0,0,0,0,0,0,0,0,133,0,153,0,212,0,223,0,155,0,196,0,172,0,170,0,182,0,227,0,225,0,154,0,0,0,0,0,44,0,132,0,124,0,60,0,200,0,0,0,0,0,59,0,0,0,226,0,66,0,63,0,0,0,51,0,0,0,170,0,0,0,0,0,242,0,116,0,236,0,162,0,0,0,246,0,67,0,48,0,89,0,0,0,46,0,190,0,35,0,76,0,112,0,139,0,65,0,232,0,0,0,0,0,198,0,139,0,245,0,99,0,157,0,0,0,221,0,53,0,0,0,255,0,115,0,38,0,197,0,122,0,80,0,149,0,100,0,26,0,7,0,0,0,189,0,198,0,151,0,122,0,42,0,0,0,116,0,249,0,51,0,87,0,237,0,199,0,0,0,0,0,44,0,112,0,32,0,237,0,222,0,67,0,203,0,0,0,0,0,0,0,227,0,210,0,94,0,151,0,36,0,85,0,147,0,197,0,251,0,99,0,251,0,36,0,30,0,131,0,0,0,145,0,0,0,43,0,235,0,189,0,246,0,20,0,0,0,0,0,0,0,26,0,0,0,50,0,62,0,28,0,114,0,0,0,181,0,0,0,0,0,0,0,231,0,0,0,0,0,175,0,74,0,110,0,0,0,242,0,166,0,116,0,0,0,128,0,0,0,0,0,98,0,16,0,0,0,153,0,161,0,221,0,25,0,0,0,58,0,99,0,18,0,168,0,87,0,245,0,0,0,5,0,133,0,197,0,76,0,0,0,73,0,0,0,161,0,75,0,129,0,64,0,31,0,228,0,79,0,53,0,0,0,0,0,5,0,234,0,213,0,62,0,87,0,108,0,240,0,211,0,0,0,18,0,84,0,36,0,0,0,42,0,52,0,196,0,11,0,0,0,63,0,186,0,139,0,234,0,210,0,0,0,83,0,0,0,209,0,0,0,184,0,0,0,178,0,67,0,178,0,0,0,198,0,0,0,237,0,0,0,0,0,24,0,206,0,133,0,193,0,55,0,153,0,188,0,178,0,92,0,184,0,0,0,25,0,0,0,21,0,196,0,0,0,234,0,162,0,0,0,141,0,0,0,215,0,18,0,91,0,0,0,68,0,81,0,182,0,240,0,228,0,190,0,0,0,117,0,10,0,0,0,0,0,229,0,0,0,13,0,80,0,148,0,143,0,135,0,226,0,212,0,128,0,5,0,64,0,62,0,168,0,5,0,72,0,236,0,96,0,0,0,0,0,120,0,178,0,47,0,20,0,249,0,1,0,80,0,0,0,214,0,29,0,65,0,253,0,255,0,0,0,123,0,151,0,0,0,139,0,12,0,0,0,175,0,47,0,32,0,53,0,0,0,7,0,86,0,0,0,194,0,8,0,119,0,198,0,157,0,227,0,185,0,163,0,28,0,94,0,0,0,147,0,46,0,0,0,145,0,244,0,66,0,121,0,244,0,40,0,0,0,142,0,135,0,179,0,179,0,90,0,105,0,249,0,17,0,41,0,95,0,0,0,143,0,230,0,121,0,4,0,114,0,73,0,253,0,0,0,97,0,156,0,88,0,78,0,211,0,0,0,67,0,0,0,15,0,70,0,0,0,122,0,176,0,37,0,171,0,160,0,187,0,235,0,165,0,142,0,117,0,211,0,166,0,102,0,157,0,165,0,139,0,172,0,198,0,142,0,90,0,24,0,0,0,0,0,74,0,17,0,38,0,69,0,0,0,4,0,170,0,132,0,252,0,104,0,0,0,251,0,55,0,0,0,212,0,0,0,134,0,237,0,58,0,23,0,71,0,187,0,0,0,0,0,248,0,242,0,51,0,0,0,118,0,202,0,99,0,139,0,0,0,35,0,69,0,97,0,206,0,141,0,53,0,137,0,233,0,40,0,246,0,0,0,128,0,213,0,44,0,31,0,107,0,61,0,130,0,13,0,34,0,9,0,66,0,243,0,0,0,54,0,29,0,0,0,159,0,190,0,130,0,153,0,0,0,129,0,75,0,0,0,12,0,45,0,124,0,251,0,0,0,63,0,0,0,168,0,235,0,173,0,0,0,0,0,0,0,0,0,104,0,184,0,225,0,188,0,216,0,0,0,213,0,157,0,72,0,244,0,0,0,143,0,40,0,74,0,205,0,235,0,170,0,163,0,0,0,0,0,0,0,54,0,62,0,0,0,198,0,0,0,222,0,53,0,125,0,40,0,3,0,172,0,0,0,83,0,13,0,97,0,86,0,216,0,235,0,58,0,0,0,16,0,23,0,57,0,14,0,48,0,127,0,188,0,187,0,142,0,0,0,215,0,118,0,160,0,113,0,17,0,110,0,17,0,0,0,214,0,0,0,0,0,223,0,0,0,153,0,0,0,86,0,0,0,192,0,47,0,54,0,193,0,227,0,183,0,210,0,0,0,248,0,94,0,189,0,0,0,42,0,0,0,53,0,247,0,186,0,0,0,97,0,71,0,198,0,0,0,105,0,0,0,86,0,0,0,35,0,96,0,30,0,182,0,156,0,6,0,0,0,202,0,191,0,226,0,152,0,205,0,0,0,0,0,243,0,216,0,0,0,14,0,123,0,154,0,0,0,0,0,165,0,51,0,134,0,135,0,202,0,97,0,15,0,0,0,0,0,61,0,245,0,8,0,177,0,37,0,5,0,191,0,21,0,0,0,92,0,89,0,54,0,10,0,59,0,61,0,58,0,149,0,0,0,134,0,41,0,221,0,0,0,74,0,0,0,93,0,237,0,165,0,212,0,219,0,124,0,85,0,53,0,0,0,0,0,166,0,5,0,192,0,188,0,194,0,64,0,60,0,165,0,85,0,12,0,222,0,0,0,246,0,67,0,53,0,165,0,124,0,114,0,0,0,163,0,0,0,220,0,92,0,110,0,110,0,194,0,245,0,0,0,46,0,159,0,102,0,0,0,224,0,0,0,81,0,7,0,11,0,206,0,95,0,109,0,72,0,113,0,0,0,183,0,68,0,53,0,7,0,78,0,87,0,23,0,192,0,0,0,35,0,245,0,0,0,113,0,223,0,159,0,237,0,0,0,0,0,165,0,228,0,135,0,225,0,0,0,130,0,0,0,0,0,0,0,6,0,218,0,91,0,0,0,46,0,253,0,217,0,51,0,0,0,240,0,16,0,0,0,0,0,132,0,8,0,37,0,127,0,63,0,197,0,62,0,201,0,0,0,184,0,115,0,24,0,214,0,7,0,174,0,0,0,0,0,210,0,209,0,205,0,243,0,126,0,113,0,178,0,83,0,215,0,80,0,223,0,141,0,248,0,210,0,83,0,185,0,0,0,199,0,132,0,142,0,130,0,186,0,141,0,9,0,0,0,7,0,144,0,222,0,15,0,185,0,255,0,143,0,117,0,25,0,141,0,215,0,61,0,13,0,16,0,169,0,94,0,209,0,247,0,124,0,96,0,0,0,200,0,141,0,165,0,101,0,228,0,15,0,172,0,0,0,0,0,91,0,44,0,215,0,194,0,0,0,204,0,248,0,111,0,0,0,228,0,11,0,0,0,0,0,190,0,231,0,20,0,0,0,241,0,161,0,132,0,0,0,0,0,227,0,236,0,69,0,155,0,180,0,59,0,168,0,64,0,250,0);
signal scenario_full  : scenario_type := (0,0,205,31,4,31,106,31,158,31,248,31,218,31,20,31,140,31,252,31,188,31,153,31,153,30,152,31,16,31,147,31,97,31,4,31,23,31,14,31,14,30,129,31,12,31,12,30,12,29,12,28,162,31,162,30,192,31,116,31,1,31,152,31,227,31,227,30,227,29,30,31,54,31,216,31,123,31,17,31,17,30,109,31,176,31,59,31,59,30,220,31,159,31,249,31,232,31,5,31,5,30,5,29,233,31,110,31,226,31,226,30,231,31,231,30,250,31,96,31,122,31,206,31,6,31,160,31,250,31,184,31,184,30,66,31,66,30,156,31,73,31,125,31,174,31,174,30,202,31,140,31,140,30,140,29,210,31,23,31,23,30,3,31,132,31,132,30,132,29,150,31,194,31,194,30,167,31,132,31,132,30,203,31,196,31,39,31,246,31,61,31,206,31,190,31,144,31,72,31,72,30,189,31,29,31,80,31,80,30,39,31,39,30,158,31,86,31,228,31,211,31,251,31,95,31,238,31,238,30,238,29,250,31,177,31,177,30,185,31,185,30,185,29,216,31,191,31,5,31,123,31,167,31,81,31,70,31,192,31,127,31,156,31,106,31,110,31,110,30,212,31,212,30,142,31,176,31,194,31,156,31,16,31,212,31,72,31,57,31,196,31,50,31,206,31,74,31,242,31,242,30,119,31,119,30,119,29,119,28,119,27,119,26,133,31,153,31,212,31,223,31,155,31,196,31,172,31,170,31,182,31,227,31,225,31,154,31,154,30,154,29,44,31,132,31,124,31,60,31,200,31,200,30,200,29,59,31,59,30,226,31,66,31,63,31,63,30,51,31,51,30,170,31,170,30,170,29,242,31,116,31,236,31,162,31,162,30,246,31,67,31,48,31,89,31,89,30,46,31,190,31,35,31,76,31,112,31,139,31,65,31,232,31,232,30,232,29,198,31,139,31,245,31,99,31,157,31,157,30,221,31,53,31,53,30,255,31,115,31,38,31,197,31,122,31,80,31,149,31,100,31,26,31,7,31,7,30,189,31,198,31,151,31,122,31,42,31,42,30,116,31,249,31,51,31,87,31,237,31,199,31,199,30,199,29,44,31,112,31,32,31,237,31,222,31,67,31,203,31,203,30,203,29,203,28,227,31,210,31,94,31,151,31,36,31,85,31,147,31,197,31,251,31,99,31,251,31,36,31,30,31,131,31,131,30,145,31,145,30,43,31,235,31,189,31,246,31,20,31,20,30,20,29,20,28,26,31,26,30,50,31,62,31,28,31,114,31,114,30,181,31,181,30,181,29,181,28,231,31,231,30,231,29,175,31,74,31,110,31,110,30,242,31,166,31,116,31,116,30,128,31,128,30,128,29,98,31,16,31,16,30,153,31,161,31,221,31,25,31,25,30,58,31,99,31,18,31,168,31,87,31,245,31,245,30,5,31,133,31,197,31,76,31,76,30,73,31,73,30,161,31,75,31,129,31,64,31,31,31,228,31,79,31,53,31,53,30,53,29,5,31,234,31,213,31,62,31,87,31,108,31,240,31,211,31,211,30,18,31,84,31,36,31,36,30,42,31,52,31,196,31,11,31,11,30,63,31,186,31,139,31,234,31,210,31,210,30,83,31,83,30,209,31,209,30,184,31,184,30,178,31,67,31,178,31,178,30,198,31,198,30,237,31,237,30,237,29,24,31,206,31,133,31,193,31,55,31,153,31,188,31,178,31,92,31,184,31,184,30,25,31,25,30,21,31,196,31,196,30,234,31,162,31,162,30,141,31,141,30,215,31,18,31,91,31,91,30,68,31,81,31,182,31,240,31,228,31,190,31,190,30,117,31,10,31,10,30,10,29,229,31,229,30,13,31,80,31,148,31,143,31,135,31,226,31,212,31,128,31,5,31,64,31,62,31,168,31,5,31,72,31,236,31,96,31,96,30,96,29,120,31,178,31,47,31,20,31,249,31,1,31,80,31,80,30,214,31,29,31,65,31,253,31,255,31,255,30,123,31,151,31,151,30,139,31,12,31,12,30,175,31,47,31,32,31,53,31,53,30,7,31,86,31,86,30,194,31,8,31,119,31,198,31,157,31,227,31,185,31,163,31,28,31,94,31,94,30,147,31,46,31,46,30,145,31,244,31,66,31,121,31,244,31,40,31,40,30,142,31,135,31,179,31,179,31,90,31,105,31,249,31,17,31,41,31,95,31,95,30,143,31,230,31,121,31,4,31,114,31,73,31,253,31,253,30,97,31,156,31,88,31,78,31,211,31,211,30,67,31,67,30,15,31,70,31,70,30,122,31,176,31,37,31,171,31,160,31,187,31,235,31,165,31,142,31,117,31,211,31,166,31,102,31,157,31,165,31,139,31,172,31,198,31,142,31,90,31,24,31,24,30,24,29,74,31,17,31,38,31,69,31,69,30,4,31,170,31,132,31,252,31,104,31,104,30,251,31,55,31,55,30,212,31,212,30,134,31,237,31,58,31,23,31,71,31,187,31,187,30,187,29,248,31,242,31,51,31,51,30,118,31,202,31,99,31,139,31,139,30,35,31,69,31,97,31,206,31,141,31,53,31,137,31,233,31,40,31,246,31,246,30,128,31,213,31,44,31,31,31,107,31,61,31,130,31,13,31,34,31,9,31,66,31,243,31,243,30,54,31,29,31,29,30,159,31,190,31,130,31,153,31,153,30,129,31,75,31,75,30,12,31,45,31,124,31,251,31,251,30,63,31,63,30,168,31,235,31,173,31,173,30,173,29,173,28,173,27,104,31,184,31,225,31,188,31,216,31,216,30,213,31,157,31,72,31,244,31,244,30,143,31,40,31,74,31,205,31,235,31,170,31,163,31,163,30,163,29,163,28,54,31,62,31,62,30,198,31,198,30,222,31,53,31,125,31,40,31,3,31,172,31,172,30,83,31,13,31,97,31,86,31,216,31,235,31,58,31,58,30,16,31,23,31,57,31,14,31,48,31,127,31,188,31,187,31,142,31,142,30,215,31,118,31,160,31,113,31,17,31,110,31,17,31,17,30,214,31,214,30,214,29,223,31,223,30,153,31,153,30,86,31,86,30,192,31,47,31,54,31,193,31,227,31,183,31,210,31,210,30,248,31,94,31,189,31,189,30,42,31,42,30,53,31,247,31,186,31,186,30,97,31,71,31,198,31,198,30,105,31,105,30,86,31,86,30,35,31,96,31,30,31,182,31,156,31,6,31,6,30,202,31,191,31,226,31,152,31,205,31,205,30,205,29,243,31,216,31,216,30,14,31,123,31,154,31,154,30,154,29,165,31,51,31,134,31,135,31,202,31,97,31,15,31,15,30,15,29,61,31,245,31,8,31,177,31,37,31,5,31,191,31,21,31,21,30,92,31,89,31,54,31,10,31,59,31,61,31,58,31,149,31,149,30,134,31,41,31,221,31,221,30,74,31,74,30,93,31,237,31,165,31,212,31,219,31,124,31,85,31,53,31,53,30,53,29,166,31,5,31,192,31,188,31,194,31,64,31,60,31,165,31,85,31,12,31,222,31,222,30,246,31,67,31,53,31,165,31,124,31,114,31,114,30,163,31,163,30,220,31,92,31,110,31,110,31,194,31,245,31,245,30,46,31,159,31,102,31,102,30,224,31,224,30,81,31,7,31,11,31,206,31,95,31,109,31,72,31,113,31,113,30,183,31,68,31,53,31,7,31,78,31,87,31,23,31,192,31,192,30,35,31,245,31,245,30,113,31,223,31,159,31,237,31,237,30,237,29,165,31,228,31,135,31,225,31,225,30,130,31,130,30,130,29,130,28,6,31,218,31,91,31,91,30,46,31,253,31,217,31,51,31,51,30,240,31,16,31,16,30,16,29,132,31,8,31,37,31,127,31,63,31,197,31,62,31,201,31,201,30,184,31,115,31,24,31,214,31,7,31,174,31,174,30,174,29,210,31,209,31,205,31,243,31,126,31,113,31,178,31,83,31,215,31,80,31,223,31,141,31,248,31,210,31,83,31,185,31,185,30,199,31,132,31,142,31,130,31,186,31,141,31,9,31,9,30,7,31,144,31,222,31,15,31,185,31,255,31,143,31,117,31,25,31,141,31,215,31,61,31,13,31,16,31,169,31,94,31,209,31,247,31,124,31,96,31,96,30,200,31,141,31,165,31,101,31,228,31,15,31,172,31,172,30,172,29,91,31,44,31,215,31,194,31,194,30,204,31,248,31,111,31,111,30,228,31,11,31,11,30,11,29,190,31,231,31,20,31,20,30,241,31,161,31,132,31,132,30,132,29,227,31,236,31,69,31,155,31,180,31,59,31,168,31,64,31,250,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
