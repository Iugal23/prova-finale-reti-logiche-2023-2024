-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_915 is
end project_tb_915;

architecture project_tb_arch_915 of project_tb_915 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 980;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,48,0,16,0,170,0,19,0,204,0,0,0,0,0,124,0,58,0,50,0,12,0,166,0,124,0,225,0,161,0,154,0,253,0,211,0,66,0,0,0,0,0,152,0,68,0,54,0,0,0,15,0,107,0,237,0,36,0,27,0,119,0,255,0,238,0,133,0,21,0,85,0,128,0,0,0,240,0,0,0,98,0,75,0,0,0,0,0,239,0,0,0,69,0,78,0,162,0,130,0,0,0,161,0,150,0,176,0,141,0,232,0,23,0,228,0,47,0,192,0,109,0,198,0,229,0,10,0,0,0,18,0,234,0,131,0,215,0,0,0,71,0,87,0,174,0,89,0,0,0,0,0,75,0,70,0,58,0,47,0,215,0,168,0,239,0,104,0,166,0,46,0,96,0,48,0,67,0,172,0,242,0,177,0,23,0,239,0,79,0,182,0,190,0,47,0,0,0,204,0,74,0,162,0,221,0,36,0,105,0,165,0,5,0,149,0,40,0,0,0,0,0,244,0,0,0,33,0,203,0,252,0,121,0,122,0,158,0,65,0,24,0,223,0,186,0,205,0,11,0,187,0,159,0,112,0,41,0,120,0,85,0,105,0,13,0,57,0,34,0,0,0,114,0,118,0,108,0,0,0,0,0,0,0,143,0,0,0,186,0,31,0,66,0,155,0,102,0,210,0,0,0,17,0,4,0,16,0,195,0,197,0,133,0,48,0,0,0,9,0,94,0,107,0,141,0,0,0,96,0,92,0,0,0,31,0,99,0,16,0,200,0,121,0,43,0,26,0,190,0,221,0,117,0,28,0,194,0,243,0,94,0,0,0,89,0,0,0,94,0,165,0,225,0,0,0,8,0,164,0,233,0,214,0,22,0,192,0,146,0,104,0,0,0,116,0,0,0,14,0,0,0,117,0,214,0,131,0,171,0,69,0,22,0,0,0,24,0,0,0,95,0,163,0,0,0,96,0,185,0,89,0,53,0,0,0,15,0,223,0,99,0,63,0,178,0,0,0,28,0,92,0,75,0,116,0,228,0,253,0,0,0,68,0,155,0,157,0,175,0,0,0,190,0,0,0,225,0,152,0,0,0,149,0,24,0,204,0,0,0,128,0,0,0,0,0,0,0,0,0,91,0,179,0,80,0,214,0,125,0,8,0,96,0,52,0,62,0,110,0,6,0,13,0,235,0,169,0,13,0,49,0,118,0,2,0,3,0,219,0,0,0,211,0,0,0,187,0,18,0,93,0,99,0,120,0,106,0,151,0,0,0,132,0,156,0,68,0,71,0,0,0,0,0,0,0,77,0,0,0,184,0,208,0,185,0,176,0,224,0,81,0,0,0,213,0,21,0,73,0,37,0,0,0,69,0,134,0,36,0,0,0,124,0,181,0,162,0,101,0,0,0,246,0,0,0,12,0,175,0,0,0,109,0,42,0,45,0,194,0,0,0,0,0,105,0,153,0,89,0,68,0,252,0,0,0,1,0,137,0,0,0,85,0,215,0,54,0,127,0,207,0,0,0,188,0,161,0,87,0,84,0,136,0,82,0,0,0,192,0,243,0,20,0,0,0,252,0,53,0,221,0,80,0,0,0,121,0,243,0,234,0,87,0,195,0,0,0,3,0,0,0,0,0,98,0,0,0,0,0,0,0,53,0,223,0,0,0,90,0,0,0,226,0,0,0,0,0,7,0,89,0,194,0,230,0,85,0,41,0,0,0,1,0,240,0,25,0,89,0,128,0,0,0,0,0,239,0,105,0,18,0,44,0,169,0,47,0,114,0,81,0,119,0,110,0,128,0,132,0,233,0,3,0,31,0,16,0,200,0,69,0,25,0,137,0,0,0,0,0,0,0,48,0,0,0,251,0,0,0,7,0,0,0,50,0,131,0,250,0,115,0,141,0,0,0,0,0,156,0,15,0,38,0,224,0,235,0,109,0,0,0,221,0,184,0,154,0,76,0,177,0,116,0,5,0,1,0,211,0,195,0,47,0,0,0,104,0,92,0,132,0,0,0,128,0,158,0,42,0,35,0,116,0,0,0,117,0,180,0,175,0,107,0,235,0,0,0,247,0,234,0,115,0,248,0,70,0,14,0,2,0,212,0,96,0,116,0,81,0,84,0,0,0,0,0,237,0,0,0,24,0,134,0,170,0,223,0,232,0,29,0,105,0,0,0,109,0,111,0,215,0,189,0,144,0,0,0,191,0,0,0,255,0,0,0,0,0,213,0,208,0,26,0,0,0,86,0,0,0,118,0,125,0,0,0,94,0,2,0,247,0,177,0,54,0,46,0,83,0,0,0,104,0,161,0,108,0,178,0,60,0,0,0,150,0,59,0,213,0,158,0,0,0,135,0,0,0,0,0,59,0,27,0,0,0,28,0,0,0,213,0,79,0,131,0,124,0,73,0,0,0,224,0,219,0,236,0,192,0,217,0,0,0,0,0,99,0,136,0,159,0,66,0,0,0,68,0,62,0,203,0,63,0,28,0,213,0,38,0,209,0,187,0,33,0,0,0,134,0,88,0,158,0,80,0,102,0,55,0,171,0,89,0,200,0,214,0,0,0,0,0,165,0,3,0,187,0,55,0,106,0,46,0,122,0,0,0,21,0,140,0,145,0,0,0,147,0,239,0,228,0,0,0,0,0,126,0,230,0,182,0,176,0,202,0,224,0,138,0,52,0,0,0,0,0,206,0,0,0,154,0,102,0,0,0,150,0,186,0,0,0,0,0,179,0,223,0,231,0,158,0,247,0,22,0,95,0,29,0,168,0,70,0,210,0,136,0,206,0,0,0,122,0,26,0,12,0,0,0,142,0,116,0,153,0,0,0,205,0,97,0,104,0,81,0,100,0,115,0,8,0,160,0,26,0,190,0,115,0,118,0,93,0,234,0,129,0,0,0,120,0,170,0,14,0,0,0,0,0,146,0,158,0,0,0,39,0,32,0,0,0,200,0,177,0,202,0,0,0,76,0,0,0,0,0,23,0,11,0,210,0,98,0,240,0,169,0,187,0,136,0,141,0,0,0,66,0,9,0,217,0,0,0,0,0,243,0,167,0,161,0,126,0,0,0,143,0,86,0,242,0,63,0,33,0,247,0,47,0,11,0,0,0,128,0,252,0,227,0,65,0,128,0,0,0,63,0,0,0,115,0,62,0,160,0,39,0,76,0,158,0,201,0,239,0,72,0,166,0,0,0,35,0,222,0,7,0,40,0,110,0,50,0,97,0,140,0,125,0,96,0,62,0,189,0,73,0,0,0,62,0,105,0,29,0,147,0,179,0,225,0,53,0,252,0,0,0,0,0,72,0,102,0,242,0,70,0,45,0,60,0,0,0,247,0,0,0,146,0,102,0,12,0,0,0,168,0,44,0,169,0,0,0,0,0,0,0,126,0,180,0,88,0,105,0,200,0,95,0,0,0,54,0,136,0,87,0,0,0,105,0,49,0,82,0,0,0,14,0,0,0,0,0,146,0,92,0,196,0,127,0,15,0,61,0,0,0,159,0,0,0,182,0,0,0,0,0,9,0,72,0,157,0,228,0,0,0,121,0,0,0,181,0,98,0,0,0,0,0,0,0,92,0,232,0,0,0,87,0,151,0,0,0,116,0,254,0,193,0,0,0,161,0,76,0,0,0,0,0,115,0,62,0,0,0,196,0,176,0,110,0,109,0,149,0,69,0,146,0,0,0,255,0,0,0,64,0,0,0,0,0,209,0,0,0,0,0,255,0,31,0,30,0,249,0,178,0,92,0,205,0,197,0,112,0,252,0,107,0,131,0,0,0,131,0,156,0,225,0,0,0,74,0,0,0,238,0,46,0,0,0,40,0,79,0,121,0,245,0,171,0,218,0,115,0,212,0,84,0,37,0,0,0,59,0,235,0,0,0,98,0,236,0,228,0,0,0,5,0,210,0,124,0,0,0,145,0,12,0,227,0,35,0,115,0,156,0,11,0,192,0,0,0,0,0,81,0,0,0,68,0,78,0,85,0,137,0,0,0,57,0,4,0,80,0,79,0,92,0,0,0,0,0,237,0,101,0,60,0,186,0,35,0,180,0,251,0,234,0,121,0,186,0,171,0,104,0,57,0,166,0,0,0,27,0,0,0,52,0,85,0,104,0,29,0,179,0,220,0,104,0,186,0,51,0,162,0,91,0,0,0,228,0,166,0,0,0,0,0,211,0,172,0,30,0,32,0,202,0,183,0,61,0,0,0,168,0,17,0,180,0,178,0,0,0,115,0,247,0,122,0,221,0,0,0,239,0,0,0,189,0,76,0,212,0,0,0,10,0,197,0,110,0,254,0,156,0,192,0,58,0,0,0,252,0,214,0,219,0,145,0,214,0,144,0,117,0,0,0,255,0,63,0,16,0,201,0,230,0,0,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,48,31,16,31,170,31,19,31,204,31,204,30,204,29,124,31,58,31,50,31,12,31,166,31,124,31,225,31,161,31,154,31,253,31,211,31,66,31,66,30,66,29,152,31,68,31,54,31,54,30,15,31,107,31,237,31,36,31,27,31,119,31,255,31,238,31,133,31,21,31,85,31,128,31,128,30,240,31,240,30,98,31,75,31,75,30,75,29,239,31,239,30,69,31,78,31,162,31,130,31,130,30,161,31,150,31,176,31,141,31,232,31,23,31,228,31,47,31,192,31,109,31,198,31,229,31,10,31,10,30,18,31,234,31,131,31,215,31,215,30,71,31,87,31,174,31,89,31,89,30,89,29,75,31,70,31,58,31,47,31,215,31,168,31,239,31,104,31,166,31,46,31,96,31,48,31,67,31,172,31,242,31,177,31,23,31,239,31,79,31,182,31,190,31,47,31,47,30,204,31,74,31,162,31,221,31,36,31,105,31,165,31,5,31,149,31,40,31,40,30,40,29,244,31,244,30,33,31,203,31,252,31,121,31,122,31,158,31,65,31,24,31,223,31,186,31,205,31,11,31,187,31,159,31,112,31,41,31,120,31,85,31,105,31,13,31,57,31,34,31,34,30,114,31,118,31,108,31,108,30,108,29,108,28,143,31,143,30,186,31,31,31,66,31,155,31,102,31,210,31,210,30,17,31,4,31,16,31,195,31,197,31,133,31,48,31,48,30,9,31,94,31,107,31,141,31,141,30,96,31,92,31,92,30,31,31,99,31,16,31,200,31,121,31,43,31,26,31,190,31,221,31,117,31,28,31,194,31,243,31,94,31,94,30,89,31,89,30,94,31,165,31,225,31,225,30,8,31,164,31,233,31,214,31,22,31,192,31,146,31,104,31,104,30,116,31,116,30,14,31,14,30,117,31,214,31,131,31,171,31,69,31,22,31,22,30,24,31,24,30,95,31,163,31,163,30,96,31,185,31,89,31,53,31,53,30,15,31,223,31,99,31,63,31,178,31,178,30,28,31,92,31,75,31,116,31,228,31,253,31,253,30,68,31,155,31,157,31,175,31,175,30,190,31,190,30,225,31,152,31,152,30,149,31,24,31,204,31,204,30,128,31,128,30,128,29,128,28,128,27,91,31,179,31,80,31,214,31,125,31,8,31,96,31,52,31,62,31,110,31,6,31,13,31,235,31,169,31,13,31,49,31,118,31,2,31,3,31,219,31,219,30,211,31,211,30,187,31,18,31,93,31,99,31,120,31,106,31,151,31,151,30,132,31,156,31,68,31,71,31,71,30,71,29,71,28,77,31,77,30,184,31,208,31,185,31,176,31,224,31,81,31,81,30,213,31,21,31,73,31,37,31,37,30,69,31,134,31,36,31,36,30,124,31,181,31,162,31,101,31,101,30,246,31,246,30,12,31,175,31,175,30,109,31,42,31,45,31,194,31,194,30,194,29,105,31,153,31,89,31,68,31,252,31,252,30,1,31,137,31,137,30,85,31,215,31,54,31,127,31,207,31,207,30,188,31,161,31,87,31,84,31,136,31,82,31,82,30,192,31,243,31,20,31,20,30,252,31,53,31,221,31,80,31,80,30,121,31,243,31,234,31,87,31,195,31,195,30,3,31,3,30,3,29,98,31,98,30,98,29,98,28,53,31,223,31,223,30,90,31,90,30,226,31,226,30,226,29,7,31,89,31,194,31,230,31,85,31,41,31,41,30,1,31,240,31,25,31,89,31,128,31,128,30,128,29,239,31,105,31,18,31,44,31,169,31,47,31,114,31,81,31,119,31,110,31,128,31,132,31,233,31,3,31,31,31,16,31,200,31,69,31,25,31,137,31,137,30,137,29,137,28,48,31,48,30,251,31,251,30,7,31,7,30,50,31,131,31,250,31,115,31,141,31,141,30,141,29,156,31,15,31,38,31,224,31,235,31,109,31,109,30,221,31,184,31,154,31,76,31,177,31,116,31,5,31,1,31,211,31,195,31,47,31,47,30,104,31,92,31,132,31,132,30,128,31,158,31,42,31,35,31,116,31,116,30,117,31,180,31,175,31,107,31,235,31,235,30,247,31,234,31,115,31,248,31,70,31,14,31,2,31,212,31,96,31,116,31,81,31,84,31,84,30,84,29,237,31,237,30,24,31,134,31,170,31,223,31,232,31,29,31,105,31,105,30,109,31,111,31,215,31,189,31,144,31,144,30,191,31,191,30,255,31,255,30,255,29,213,31,208,31,26,31,26,30,86,31,86,30,118,31,125,31,125,30,94,31,2,31,247,31,177,31,54,31,46,31,83,31,83,30,104,31,161,31,108,31,178,31,60,31,60,30,150,31,59,31,213,31,158,31,158,30,135,31,135,30,135,29,59,31,27,31,27,30,28,31,28,30,213,31,79,31,131,31,124,31,73,31,73,30,224,31,219,31,236,31,192,31,217,31,217,30,217,29,99,31,136,31,159,31,66,31,66,30,68,31,62,31,203,31,63,31,28,31,213,31,38,31,209,31,187,31,33,31,33,30,134,31,88,31,158,31,80,31,102,31,55,31,171,31,89,31,200,31,214,31,214,30,214,29,165,31,3,31,187,31,55,31,106,31,46,31,122,31,122,30,21,31,140,31,145,31,145,30,147,31,239,31,228,31,228,30,228,29,126,31,230,31,182,31,176,31,202,31,224,31,138,31,52,31,52,30,52,29,206,31,206,30,154,31,102,31,102,30,150,31,186,31,186,30,186,29,179,31,223,31,231,31,158,31,247,31,22,31,95,31,29,31,168,31,70,31,210,31,136,31,206,31,206,30,122,31,26,31,12,31,12,30,142,31,116,31,153,31,153,30,205,31,97,31,104,31,81,31,100,31,115,31,8,31,160,31,26,31,190,31,115,31,118,31,93,31,234,31,129,31,129,30,120,31,170,31,14,31,14,30,14,29,146,31,158,31,158,30,39,31,32,31,32,30,200,31,177,31,202,31,202,30,76,31,76,30,76,29,23,31,11,31,210,31,98,31,240,31,169,31,187,31,136,31,141,31,141,30,66,31,9,31,217,31,217,30,217,29,243,31,167,31,161,31,126,31,126,30,143,31,86,31,242,31,63,31,33,31,247,31,47,31,11,31,11,30,128,31,252,31,227,31,65,31,128,31,128,30,63,31,63,30,115,31,62,31,160,31,39,31,76,31,158,31,201,31,239,31,72,31,166,31,166,30,35,31,222,31,7,31,40,31,110,31,50,31,97,31,140,31,125,31,96,31,62,31,189,31,73,31,73,30,62,31,105,31,29,31,147,31,179,31,225,31,53,31,252,31,252,30,252,29,72,31,102,31,242,31,70,31,45,31,60,31,60,30,247,31,247,30,146,31,102,31,12,31,12,30,168,31,44,31,169,31,169,30,169,29,169,28,126,31,180,31,88,31,105,31,200,31,95,31,95,30,54,31,136,31,87,31,87,30,105,31,49,31,82,31,82,30,14,31,14,30,14,29,146,31,92,31,196,31,127,31,15,31,61,31,61,30,159,31,159,30,182,31,182,30,182,29,9,31,72,31,157,31,228,31,228,30,121,31,121,30,181,31,98,31,98,30,98,29,98,28,92,31,232,31,232,30,87,31,151,31,151,30,116,31,254,31,193,31,193,30,161,31,76,31,76,30,76,29,115,31,62,31,62,30,196,31,176,31,110,31,109,31,149,31,69,31,146,31,146,30,255,31,255,30,64,31,64,30,64,29,209,31,209,30,209,29,255,31,31,31,30,31,249,31,178,31,92,31,205,31,197,31,112,31,252,31,107,31,131,31,131,30,131,31,156,31,225,31,225,30,74,31,74,30,238,31,46,31,46,30,40,31,79,31,121,31,245,31,171,31,218,31,115,31,212,31,84,31,37,31,37,30,59,31,235,31,235,30,98,31,236,31,228,31,228,30,5,31,210,31,124,31,124,30,145,31,12,31,227,31,35,31,115,31,156,31,11,31,192,31,192,30,192,29,81,31,81,30,68,31,78,31,85,31,137,31,137,30,57,31,4,31,80,31,79,31,92,31,92,30,92,29,237,31,101,31,60,31,186,31,35,31,180,31,251,31,234,31,121,31,186,31,171,31,104,31,57,31,166,31,166,30,27,31,27,30,52,31,85,31,104,31,29,31,179,31,220,31,104,31,186,31,51,31,162,31,91,31,91,30,228,31,166,31,166,30,166,29,211,31,172,31,30,31,32,31,202,31,183,31,61,31,61,30,168,31,17,31,180,31,178,31,178,30,115,31,247,31,122,31,221,31,221,30,239,31,239,30,189,31,76,31,212,31,212,30,10,31,197,31,110,31,254,31,156,31,192,31,58,31,58,30,252,31,214,31,219,31,145,31,214,31,144,31,117,31,117,30,255,31,63,31,16,31,201,31,230,31,230,30,230,29,230,28,230,27);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
