-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 799;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (198,0,228,0,62,0,131,0,202,0,22,0,226,0,167,0,180,0,165,0,0,0,138,0,51,0,247,0,0,0,0,0,179,0,58,0,180,0,231,0,251,0,133,0,68,0,40,0,0,0,211,0,180,0,2,0,112,0,48,0,217,0,197,0,2,0,146,0,36,0,130,0,0,0,83,0,248,0,243,0,146,0,112,0,0,0,160,0,122,0,10,0,0,0,140,0,234,0,132,0,103,0,0,0,0,0,0,0,103,0,72,0,228,0,0,0,95,0,129,0,133,0,0,0,9,0,0,0,127,0,42,0,162,0,27,0,191,0,132,0,187,0,121,0,0,0,177,0,113,0,0,0,194,0,78,0,0,0,4,0,32,0,186,0,0,0,216,0,250,0,0,0,0,0,9,0,235,0,152,0,14,0,0,0,93,0,0,0,105,0,165,0,0,0,125,0,160,0,223,0,210,0,210,0,204,0,0,0,157,0,241,0,0,0,22,0,49,0,0,0,0,0,243,0,90,0,110,0,0,0,48,0,28,0,60,0,163,0,241,0,243,0,0,0,0,0,237,0,6,0,213,0,186,0,203,0,0,0,0,0,94,0,129,0,160,0,70,0,128,0,0,0,9,0,65,0,0,0,8,0,23,0,41,0,246,0,124,0,149,0,184,0,57,0,153,0,142,0,249,0,215,0,0,0,78,0,21,0,0,0,211,0,245,0,122,0,174,0,58,0,0,0,164,0,108,0,205,0,91,0,0,0,96,0,0,0,103,0,77,0,0,0,108,0,180,0,55,0,162,0,0,0,199,0,0,0,139,0,166,0,82,0,0,0,66,0,202,0,129,0,212,0,241,0,158,0,75,0,148,0,126,0,210,0,73,0,18,0,105,0,0,0,75,0,241,0,214,0,0,0,209,0,165,0,61,0,253,0,111,0,102,0,162,0,0,0,214,0,149,0,126,0,76,0,0,0,159,0,0,0,60,0,187,0,48,0,9,0,0,0,36,0,59,0,111,0,74,0,237,0,205,0,143,0,0,0,122,0,175,0,65,0,120,0,169,0,122,0,218,0,237,0,0,0,227,0,225,0,61,0,106,0,23,0,109,0,39,0,47,0,102,0,0,0,173,0,19,0,3,0,56,0,218,0,182,0,109,0,245,0,202,0,25,0,106,0,19,0,225,0,241,0,46,0,16,0,98,0,45,0,240,0,131,0,34,0,0,0,141,0,176,0,128,0,205,0,101,0,44,0,233,0,9,0,234,0,0,0,155,0,44,0,137,0,150,0,0,0,120,0,59,0,180,0,168,0,49,0,95,0,229,0,0,0,71,0,44,0,215,0,0,0,0,0,0,0,51,0,11,0,0,0,125,0,30,0,39,0,215,0,158,0,0,0,221,0,119,0,132,0,196,0,59,0,0,0,0,0,0,0,72,0,0,0,163,0,57,0,0,0,133,0,142,0,181,0,55,0,121,0,33,0,169,0,3,0,26,0,0,0,81,0,127,0,192,0,0,0,0,0,48,0,0,0,176,0,0,0,91,0,84,0,39,0,109,0,15,0,37,0,0,0,137,0,213,0,0,0,0,0,0,0,248,0,120,0,40,0,0,0,221,0,0,0,0,0,202,0,133,0,165,0,36,0,0,0,96,0,20,0,220,0,236,0,142,0,255,0,181,0,221,0,254,0,90,0,0,0,224,0,251,0,54,0,71,0,0,0,255,0,0,0,161,0,158,0,239,0,85,0,151,0,223,0,133,0,230,0,0,0,70,0,79,0,255,0,0,0,203,0,167,0,42,0,161,0,125,0,7,0,161,0,165,0,98,0,227,0,108,0,54,0,243,0,0,0,162,0,216,0,1,0,0,0,106,0,240,0,232,0,244,0,0,0,109,0,111,0,0,0,254,0,75,0,149,0,215,0,145,0,232,0,28,0,9,0,79,0,93,0,216,0,183,0,3,0,79,0,110,0,0,0,157,0,84,0,149,0,216,0,17,0,141,0,25,0,139,0,244,0,35,0,0,0,178,0,0,0,69,0,0,0,0,0,0,0,212,0,109,0,172,0,0,0,153,0,99,0,94,0,179,0,121,0,36,0,44,0,0,0,0,0,0,0,0,0,84,0,71,0,113,0,130,0,0,0,122,0,137,0,0,0,0,0,213,0,144,0,135,0,165,0,40,0,0,0,44,0,0,0,154,0,231,0,212,0,157,0,218,0,9,0,78,0,112,0,109,0,83,0,162,0,136,0,185,0,136,0,4,0,245,0,120,0,0,0,147,0,124,0,101,0,0,0,111,0,181,0,249,0,193,0,0,0,31,0,157,0,0,0,0,0,178,0,204,0,126,0,180,0,198,0,94,0,210,0,133,0,0,0,155,0,89,0,90,0,0,0,0,0,209,0,233,0,41,0,0,0,160,0,238,0,136,0,108,0,113,0,92,0,67,0,246,0,23,0,212,0,75,0,145,0,77,0,99,0,62,0,0,0,0,0,129,0,113,0,55,0,83,0,149,0,242,0,0,0,27,0,126,0,0,0,218,0,89,0,99,0,200,0,205,0,227,0,59,0,75,0,210,0,241,0,82,0,183,0,0,0,19,0,2,0,126,0,56,0,47,0,247,0,127,0,47,0,16,0,196,0,197,0,89,0,124,0,184,0,19,0,0,0,68,0,112,0,0,0,196,0,0,0,0,0,0,0,47,0,86,0,226,0,245,0,110,0,0,0,0,0,212,0,184,0,167,0,187,0,87,0,237,0,29,0,6,0,254,0,32,0,43,0,126,0,85,0,129,0,219,0,90,0,166,0,0,0,39,0,17,0,84,0,11,0,0,0,226,0,144,0,40,0,252,0,116,0,196,0,163,0,190,0,98,0,228,0,0,0,245,0,45,0,0,0,0,0,8,0,176,0,94,0,40,0,0,0,0,0,200,0,149,0,197,0,211,0,127,0,135,0,0,0,78,0,208,0,141,0,0,0,143,0,171,0,213,0,137,0,178,0,0,0,0,0,0,0,17,0,207,0,232,0,247,0,0,0,51,0,237,0,225,0,0,0,159,0,111,0,0,0,102,0,22,0,0,0,210,0,198,0,197,0,241,0,17,0,0,0,0,0,212,0,214,0,214,0,93,0,0,0,40,0,150,0,12,0,92,0,44,0,165,0,0,0,224,0,24,0,106,0,0,0,76,0,0,0,244,0,33,0,155,0,0,0,86,0,190,0,229,0,110,0,148,0,97,0,0,0,96,0,200,0,255,0,31,0,190,0,0,0,52,0,0,0,0,0,132,0,34,0,77,0,1,0,154,0,67,0,232,0,121,0,74,0,48,0,0,0,23,0,0,0,148,0,0,0,105,0,243,0,48,0,0,0,47,0,134,0,0,0,238,0,96,0,177,0,25,0,4,0,210,0,142,0,181,0,0,0,0,0,80,0,0,0,92,0,231,0,5,0,240,0,135,0,113,0,0,0,11,0,0,0,118,0,0,0,53,0,232,0,204,0,2,0,209,0,14,0,0,0,145,0,68,0,14,0,196,0,252,0,95,0,181,0,248,0,0,0,127,0,144,0,198,0,115,0,30,0,29,0,187,0,225,0,132,0,43,0,233,0);
signal scenario_full  : scenario_type := (198,31,228,31,62,31,131,31,202,31,22,31,226,31,167,31,180,31,165,31,165,30,138,31,51,31,247,31,247,30,247,29,179,31,58,31,180,31,231,31,251,31,133,31,68,31,40,31,40,30,211,31,180,31,2,31,112,31,48,31,217,31,197,31,2,31,146,31,36,31,130,31,130,30,83,31,248,31,243,31,146,31,112,31,112,30,160,31,122,31,10,31,10,30,140,31,234,31,132,31,103,31,103,30,103,29,103,28,103,31,72,31,228,31,228,30,95,31,129,31,133,31,133,30,9,31,9,30,127,31,42,31,162,31,27,31,191,31,132,31,187,31,121,31,121,30,177,31,113,31,113,30,194,31,78,31,78,30,4,31,32,31,186,31,186,30,216,31,250,31,250,30,250,29,9,31,235,31,152,31,14,31,14,30,93,31,93,30,105,31,165,31,165,30,125,31,160,31,223,31,210,31,210,31,204,31,204,30,157,31,241,31,241,30,22,31,49,31,49,30,49,29,243,31,90,31,110,31,110,30,48,31,28,31,60,31,163,31,241,31,243,31,243,30,243,29,237,31,6,31,213,31,186,31,203,31,203,30,203,29,94,31,129,31,160,31,70,31,128,31,128,30,9,31,65,31,65,30,8,31,23,31,41,31,246,31,124,31,149,31,184,31,57,31,153,31,142,31,249,31,215,31,215,30,78,31,21,31,21,30,211,31,245,31,122,31,174,31,58,31,58,30,164,31,108,31,205,31,91,31,91,30,96,31,96,30,103,31,77,31,77,30,108,31,180,31,55,31,162,31,162,30,199,31,199,30,139,31,166,31,82,31,82,30,66,31,202,31,129,31,212,31,241,31,158,31,75,31,148,31,126,31,210,31,73,31,18,31,105,31,105,30,75,31,241,31,214,31,214,30,209,31,165,31,61,31,253,31,111,31,102,31,162,31,162,30,214,31,149,31,126,31,76,31,76,30,159,31,159,30,60,31,187,31,48,31,9,31,9,30,36,31,59,31,111,31,74,31,237,31,205,31,143,31,143,30,122,31,175,31,65,31,120,31,169,31,122,31,218,31,237,31,237,30,227,31,225,31,61,31,106,31,23,31,109,31,39,31,47,31,102,31,102,30,173,31,19,31,3,31,56,31,218,31,182,31,109,31,245,31,202,31,25,31,106,31,19,31,225,31,241,31,46,31,16,31,98,31,45,31,240,31,131,31,34,31,34,30,141,31,176,31,128,31,205,31,101,31,44,31,233,31,9,31,234,31,234,30,155,31,44,31,137,31,150,31,150,30,120,31,59,31,180,31,168,31,49,31,95,31,229,31,229,30,71,31,44,31,215,31,215,30,215,29,215,28,51,31,11,31,11,30,125,31,30,31,39,31,215,31,158,31,158,30,221,31,119,31,132,31,196,31,59,31,59,30,59,29,59,28,72,31,72,30,163,31,57,31,57,30,133,31,142,31,181,31,55,31,121,31,33,31,169,31,3,31,26,31,26,30,81,31,127,31,192,31,192,30,192,29,48,31,48,30,176,31,176,30,91,31,84,31,39,31,109,31,15,31,37,31,37,30,137,31,213,31,213,30,213,29,213,28,248,31,120,31,40,31,40,30,221,31,221,30,221,29,202,31,133,31,165,31,36,31,36,30,96,31,20,31,220,31,236,31,142,31,255,31,181,31,221,31,254,31,90,31,90,30,224,31,251,31,54,31,71,31,71,30,255,31,255,30,161,31,158,31,239,31,85,31,151,31,223,31,133,31,230,31,230,30,70,31,79,31,255,31,255,30,203,31,167,31,42,31,161,31,125,31,7,31,161,31,165,31,98,31,227,31,108,31,54,31,243,31,243,30,162,31,216,31,1,31,1,30,106,31,240,31,232,31,244,31,244,30,109,31,111,31,111,30,254,31,75,31,149,31,215,31,145,31,232,31,28,31,9,31,79,31,93,31,216,31,183,31,3,31,79,31,110,31,110,30,157,31,84,31,149,31,216,31,17,31,141,31,25,31,139,31,244,31,35,31,35,30,178,31,178,30,69,31,69,30,69,29,69,28,212,31,109,31,172,31,172,30,153,31,99,31,94,31,179,31,121,31,36,31,44,31,44,30,44,29,44,28,44,27,84,31,71,31,113,31,130,31,130,30,122,31,137,31,137,30,137,29,213,31,144,31,135,31,165,31,40,31,40,30,44,31,44,30,154,31,231,31,212,31,157,31,218,31,9,31,78,31,112,31,109,31,83,31,162,31,136,31,185,31,136,31,4,31,245,31,120,31,120,30,147,31,124,31,101,31,101,30,111,31,181,31,249,31,193,31,193,30,31,31,157,31,157,30,157,29,178,31,204,31,126,31,180,31,198,31,94,31,210,31,133,31,133,30,155,31,89,31,90,31,90,30,90,29,209,31,233,31,41,31,41,30,160,31,238,31,136,31,108,31,113,31,92,31,67,31,246,31,23,31,212,31,75,31,145,31,77,31,99,31,62,31,62,30,62,29,129,31,113,31,55,31,83,31,149,31,242,31,242,30,27,31,126,31,126,30,218,31,89,31,99,31,200,31,205,31,227,31,59,31,75,31,210,31,241,31,82,31,183,31,183,30,19,31,2,31,126,31,56,31,47,31,247,31,127,31,47,31,16,31,196,31,197,31,89,31,124,31,184,31,19,31,19,30,68,31,112,31,112,30,196,31,196,30,196,29,196,28,47,31,86,31,226,31,245,31,110,31,110,30,110,29,212,31,184,31,167,31,187,31,87,31,237,31,29,31,6,31,254,31,32,31,43,31,126,31,85,31,129,31,219,31,90,31,166,31,166,30,39,31,17,31,84,31,11,31,11,30,226,31,144,31,40,31,252,31,116,31,196,31,163,31,190,31,98,31,228,31,228,30,245,31,45,31,45,30,45,29,8,31,176,31,94,31,40,31,40,30,40,29,200,31,149,31,197,31,211,31,127,31,135,31,135,30,78,31,208,31,141,31,141,30,143,31,171,31,213,31,137,31,178,31,178,30,178,29,178,28,17,31,207,31,232,31,247,31,247,30,51,31,237,31,225,31,225,30,159,31,111,31,111,30,102,31,22,31,22,30,210,31,198,31,197,31,241,31,17,31,17,30,17,29,212,31,214,31,214,31,93,31,93,30,40,31,150,31,12,31,92,31,44,31,165,31,165,30,224,31,24,31,106,31,106,30,76,31,76,30,244,31,33,31,155,31,155,30,86,31,190,31,229,31,110,31,148,31,97,31,97,30,96,31,200,31,255,31,31,31,190,31,190,30,52,31,52,30,52,29,132,31,34,31,77,31,1,31,154,31,67,31,232,31,121,31,74,31,48,31,48,30,23,31,23,30,148,31,148,30,105,31,243,31,48,31,48,30,47,31,134,31,134,30,238,31,96,31,177,31,25,31,4,31,210,31,142,31,181,31,181,30,181,29,80,31,80,30,92,31,231,31,5,31,240,31,135,31,113,31,113,30,11,31,11,30,118,31,118,30,53,31,232,31,204,31,2,31,209,31,14,31,14,30,145,31,68,31,14,31,196,31,252,31,95,31,181,31,248,31,248,30,127,31,144,31,198,31,115,31,30,31,29,31,187,31,225,31,132,31,43,31,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
