-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_519 is
end project_tb_519;

architecture project_tb_arch_519 of project_tb_519 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 992;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (38,0,113,0,84,0,180,0,184,0,0,0,113,0,50,0,10,0,44,0,148,0,113,0,82,0,0,0,0,0,160,0,0,0,169,0,0,0,183,0,146,0,60,0,48,0,99,0,0,0,17,0,137,0,128,0,114,0,16,0,0,0,134,0,230,0,40,0,200,0,224,0,0,0,10,0,0,0,207,0,151,0,6,0,198,0,0,0,6,0,188,0,199,0,72,0,0,0,183,0,135,0,0,0,137,0,108,0,182,0,0,0,156,0,130,0,3,0,58,0,83,0,175,0,0,0,8,0,222,0,0,0,0,0,197,0,176,0,251,0,173,0,186,0,137,0,165,0,53,0,0,0,201,0,0,0,225,0,202,0,174,0,102,0,222,0,85,0,203,0,197,0,0,0,0,0,85,0,0,0,0,0,145,0,129,0,152,0,117,0,224,0,222,0,9,0,244,0,104,0,216,0,227,0,7,0,87,0,199,0,25,0,207,0,0,0,50,0,0,0,105,0,0,0,52,0,219,0,39,0,6,0,21,0,0,0,191,0,36,0,214,0,103,0,0,0,179,0,160,0,241,0,96,0,0,0,0,0,173,0,59,0,74,0,133,0,30,0,100,0,106,0,58,0,0,0,195,0,0,0,171,0,0,0,172,0,0,0,33,0,79,0,217,0,0,0,0,0,16,0,65,0,24,0,0,0,33,0,6,0,51,0,239,0,238,0,142,0,0,0,220,0,0,0,12,0,110,0,210,0,26,0,16,0,26,0,107,0,101,0,246,0,185,0,140,0,128,0,5,0,163,0,0,0,213,0,94,0,255,0,5,0,122,0,237,0,200,0,86,0,25,0,252,0,40,0,59,0,138,0,68,0,126,0,238,0,67,0,180,0,10,0,171,0,69,0,139,0,17,0,0,0,56,0,0,0,20,0,0,0,13,0,0,0,141,0,20,0,159,0,0,0,0,0,39,0,0,0,243,0,0,0,129,0,0,0,211,0,106,0,143,0,37,0,197,0,170,0,160,0,2,0,127,0,1,0,233,0,0,0,169,0,97,0,119,0,233,0,0,0,166,0,0,0,97,0,10,0,33,0,23,0,0,0,86,0,68,0,12,0,172,0,0,0,127,0,0,0,103,0,160,0,178,0,129,0,25,0,174,0,227,0,167,0,240,0,0,0,210,0,60,0,154,0,152,0,0,0,127,0,0,0,201,0,17,0,0,0,112,0,64,0,80,0,39,0,220,0,0,0,129,0,250,0,111,0,21,0,63,0,138,0,0,0,246,0,162,0,14,0,23,0,79,0,0,0,195,0,143,0,186,0,66,0,66,0,7,0,19,0,49,0,79,0,108,0,200,0,44,0,93,0,144,0,128,0,0,0,39,0,182,0,193,0,15,0,138,0,2,0,0,0,184,0,34,0,0,0,116,0,168,0,0,0,166,0,86,0,198,0,0,0,92,0,0,0,240,0,194,0,0,0,181,0,98,0,196,0,117,0,22,0,253,0,153,0,101,0,0,0,0,0,17,0,92,0,178,0,171,0,115,0,0,0,217,0,141,0,0,0,179,0,28,0,49,0,0,0,105,0,0,0,253,0,93,0,49,0,160,0,219,0,134,0,121,0,177,0,0,0,193,0,0,0,212,0,210,0,233,0,59,0,0,0,115,0,125,0,133,0,194,0,247,0,0,0,234,0,102,0,0,0,206,0,191,0,173,0,35,0,191,0,137,0,0,0,98,0,81,0,40,0,200,0,5,0,35,0,253,0,131,0,0,0,0,0,0,0,236,0,48,0,178,0,167,0,168,0,156,0,144,0,8,0,215,0,54,0,35,0,162,0,151,0,167,0,159,0,0,0,0,0,184,0,182,0,146,0,0,0,89,0,0,0,169,0,141,0,68,0,0,0,84,0,0,0,247,0,84,0,173,0,248,0,224,0,0,0,152,0,0,0,0,0,210,0,212,0,46,0,155,0,85,0,196,0,186,0,0,0,0,0,75,0,14,0,0,0,62,0,251,0,207,0,0,0,97,0,0,0,196,0,0,0,0,0,17,0,0,0,150,0,73,0,104,0,0,0,210,0,13,0,176,0,38,0,0,0,0,0,150,0,242,0,72,0,242,0,4,0,148,0,189,0,151,0,55,0,12,0,196,0,180,0,194,0,0,0,10,0,45,0,97,0,0,0,84,0,0,0,255,0,0,0,115,0,237,0,234,0,210,0,152,0,5,0,68,0,42,0,249,0,178,0,237,0,189,0,103,0,0,0,227,0,141,0,0,0,176,0,0,0,6,0,223,0,0,0,144,0,183,0,13,0,145,0,57,0,233,0,102,0,0,0,0,0,68,0,73,0,5,0,0,0,0,0,179,0,0,0,0,0,162,0,42,0,93,0,212,0,247,0,177,0,173,0,178,0,41,0,19,0,88,0,99,0,170,0,238,0,183,0,0,0,114,0,248,0,0,0,229,0,0,0,0,0,0,0,0,0,144,0,75,0,0,0,48,0,158,0,75,0,182,0,252,0,0,0,0,0,23,0,92,0,211,0,33,0,0,0,250,0,189,0,224,0,159,0,114,0,221,0,0,0,85,0,151,0,52,0,102,0,41,0,155,0,14,0,221,0,40,0,118,0,0,0,79,0,83,0,13,0,98,0,144,0,166,0,127,0,122,0,96,0,0,0,180,0,196,0,0,0,173,0,131,0,114,0,63,0,153,0,133,0,206,0,196,0,192,0,0,0,248,0,0,0,212,0,17,0,217,0,195,0,51,0,0,0,39,0,0,0,190,0,0,0,110,0,102,0,227,0,223,0,192,0,181,0,0,0,13,0,0,0,29,0,83,0,254,0,0,0,227,0,252,0,9,0,202,0,79,0,103,0,189,0,158,0,8,0,0,0,0,0,222,0,213,0,0,0,222,0,157,0,0,0,248,0,171,0,0,0,146,0,32,0,77,0,153,0,100,0,59,0,181,0,0,0,62,0,39,0,112,0,0,0,53,0,113,0,246,0,212,0,249,0,0,0,150,0,0,0,155,0,0,0,228,0,227,0,12,0,197,0,127,0,0,0,0,0,171,0,12,0,40,0,150,0,85,0,217,0,0,0,217,0,0,0,12,0,0,0,222,0,110,0,0,0,0,0,104,0,140,0,119,0,0,0,9,0,207,0,129,0,164,0,21,0,203,0,0,0,146,0,0,0,0,0,65,0,0,0,64,0,170,0,0,0,213,0,0,0,142,0,123,0,0,0,0,0,244,0,123,0,160,0,150,0,13,0,0,0,0,0,151,0,176,0,192,0,127,0,233,0,163,0,26,0,151,0,87,0,230,0,238,0,210,0,0,0,206,0,197,0,215,0,226,0,0,0,122,0,0,0,246,0,16,0,23,0,0,0,176,0,65,0,0,0,192,0,44,0,50,0,30,0,11,0,234,0,0,0,13,0,138,0,208,0,205,0,0,0,83,0,93,0,204,0,238,0,177,0,0,0,229,0,254,0,164,0,242,0,5,0,229,0,209,0,81,0,228,0,210,0,3,0,122,0,0,0,103,0,121,0,43,0,0,0,9,0,159,0,135,0,237,0,186,0,200,0,51,0,96,0,11,0,240,0,224,0,42,0,215,0,0,0,128,0,172,0,160,0,133,0,0,0,208,0,30,0,94,0,0,0,0,0,85,0,93,0,251,0,80,0,0,0,96,0,95,0,0,0,0,0,7,0,133,0,141,0,0,0,106,0,175,0,210,0,47,0,151,0,189,0,255,0,63,0,136,0,0,0,106,0,37,0,25,0,138,0,252,0,50,0,173,0,225,0,0,0,174,0,115,0,63,0,243,0,87,0,166,0,110,0,156,0,116,0,147,0,0,0,245,0,44,0,191,0,111,0,198,0,210,0,202,0,111,0,173,0,170,0,13,0,80,0,0,0,200,0,0,0,184,0,27,0,0,0,0,0,53,0,128,0,28,0,191,0,3,0,0,0,225,0,218,0,0,0,74,0,0,0,10,0,39,0,11,0,185,0,155,0,240,0,38,0,82,0,80,0,19,0,0,0,0,0,109,0,19,0,229,0,104,0,0,0,114,0,126,0,0,0,40,0,0,0,30,0,213,0,123,0,170,0,189,0,0,0,0,0,0,0,92,0,1,0,150,0,147,0,9,0,32,0,65,0,34,0,205,0,57,0,0,0,203,0,32,0,7,0,236,0,172,0,0,0,216,0,189,0,0,0,81,0,203,0,201,0,164,0,129,0,42,0,82,0,0,0,97,0,74,0,78,0,189,0,243,0,178,0,156,0,113,0,215,0,70,0,176,0,79,0,20,0,94,0,0,0,191,0,190,0,62,0,31,0,180,0,0,0,0,0,37,0,127,0,237,0,135,0,142,0,255,0,88,0,174,0,205,0,182,0,211,0,0,0,140,0,138,0,245,0,207,0,201,0,15,0,21,0,89,0,198,0,255,0,0,0,0,0,0,0,44,0);
signal scenario_full  : scenario_type := (38,31,113,31,84,31,180,31,184,31,184,30,113,31,50,31,10,31,44,31,148,31,113,31,82,31,82,30,82,29,160,31,160,30,169,31,169,30,183,31,146,31,60,31,48,31,99,31,99,30,17,31,137,31,128,31,114,31,16,31,16,30,134,31,230,31,40,31,200,31,224,31,224,30,10,31,10,30,207,31,151,31,6,31,198,31,198,30,6,31,188,31,199,31,72,31,72,30,183,31,135,31,135,30,137,31,108,31,182,31,182,30,156,31,130,31,3,31,58,31,83,31,175,31,175,30,8,31,222,31,222,30,222,29,197,31,176,31,251,31,173,31,186,31,137,31,165,31,53,31,53,30,201,31,201,30,225,31,202,31,174,31,102,31,222,31,85,31,203,31,197,31,197,30,197,29,85,31,85,30,85,29,145,31,129,31,152,31,117,31,224,31,222,31,9,31,244,31,104,31,216,31,227,31,7,31,87,31,199,31,25,31,207,31,207,30,50,31,50,30,105,31,105,30,52,31,219,31,39,31,6,31,21,31,21,30,191,31,36,31,214,31,103,31,103,30,179,31,160,31,241,31,96,31,96,30,96,29,173,31,59,31,74,31,133,31,30,31,100,31,106,31,58,31,58,30,195,31,195,30,171,31,171,30,172,31,172,30,33,31,79,31,217,31,217,30,217,29,16,31,65,31,24,31,24,30,33,31,6,31,51,31,239,31,238,31,142,31,142,30,220,31,220,30,12,31,110,31,210,31,26,31,16,31,26,31,107,31,101,31,246,31,185,31,140,31,128,31,5,31,163,31,163,30,213,31,94,31,255,31,5,31,122,31,237,31,200,31,86,31,25,31,252,31,40,31,59,31,138,31,68,31,126,31,238,31,67,31,180,31,10,31,171,31,69,31,139,31,17,31,17,30,56,31,56,30,20,31,20,30,13,31,13,30,141,31,20,31,159,31,159,30,159,29,39,31,39,30,243,31,243,30,129,31,129,30,211,31,106,31,143,31,37,31,197,31,170,31,160,31,2,31,127,31,1,31,233,31,233,30,169,31,97,31,119,31,233,31,233,30,166,31,166,30,97,31,10,31,33,31,23,31,23,30,86,31,68,31,12,31,172,31,172,30,127,31,127,30,103,31,160,31,178,31,129,31,25,31,174,31,227,31,167,31,240,31,240,30,210,31,60,31,154,31,152,31,152,30,127,31,127,30,201,31,17,31,17,30,112,31,64,31,80,31,39,31,220,31,220,30,129,31,250,31,111,31,21,31,63,31,138,31,138,30,246,31,162,31,14,31,23,31,79,31,79,30,195,31,143,31,186,31,66,31,66,31,7,31,19,31,49,31,79,31,108,31,200,31,44,31,93,31,144,31,128,31,128,30,39,31,182,31,193,31,15,31,138,31,2,31,2,30,184,31,34,31,34,30,116,31,168,31,168,30,166,31,86,31,198,31,198,30,92,31,92,30,240,31,194,31,194,30,181,31,98,31,196,31,117,31,22,31,253,31,153,31,101,31,101,30,101,29,17,31,92,31,178,31,171,31,115,31,115,30,217,31,141,31,141,30,179,31,28,31,49,31,49,30,105,31,105,30,253,31,93,31,49,31,160,31,219,31,134,31,121,31,177,31,177,30,193,31,193,30,212,31,210,31,233,31,59,31,59,30,115,31,125,31,133,31,194,31,247,31,247,30,234,31,102,31,102,30,206,31,191,31,173,31,35,31,191,31,137,31,137,30,98,31,81,31,40,31,200,31,5,31,35,31,253,31,131,31,131,30,131,29,131,28,236,31,48,31,178,31,167,31,168,31,156,31,144,31,8,31,215,31,54,31,35,31,162,31,151,31,167,31,159,31,159,30,159,29,184,31,182,31,146,31,146,30,89,31,89,30,169,31,141,31,68,31,68,30,84,31,84,30,247,31,84,31,173,31,248,31,224,31,224,30,152,31,152,30,152,29,210,31,212,31,46,31,155,31,85,31,196,31,186,31,186,30,186,29,75,31,14,31,14,30,62,31,251,31,207,31,207,30,97,31,97,30,196,31,196,30,196,29,17,31,17,30,150,31,73,31,104,31,104,30,210,31,13,31,176,31,38,31,38,30,38,29,150,31,242,31,72,31,242,31,4,31,148,31,189,31,151,31,55,31,12,31,196,31,180,31,194,31,194,30,10,31,45,31,97,31,97,30,84,31,84,30,255,31,255,30,115,31,237,31,234,31,210,31,152,31,5,31,68,31,42,31,249,31,178,31,237,31,189,31,103,31,103,30,227,31,141,31,141,30,176,31,176,30,6,31,223,31,223,30,144,31,183,31,13,31,145,31,57,31,233,31,102,31,102,30,102,29,68,31,73,31,5,31,5,30,5,29,179,31,179,30,179,29,162,31,42,31,93,31,212,31,247,31,177,31,173,31,178,31,41,31,19,31,88,31,99,31,170,31,238,31,183,31,183,30,114,31,248,31,248,30,229,31,229,30,229,29,229,28,229,27,144,31,75,31,75,30,48,31,158,31,75,31,182,31,252,31,252,30,252,29,23,31,92,31,211,31,33,31,33,30,250,31,189,31,224,31,159,31,114,31,221,31,221,30,85,31,151,31,52,31,102,31,41,31,155,31,14,31,221,31,40,31,118,31,118,30,79,31,83,31,13,31,98,31,144,31,166,31,127,31,122,31,96,31,96,30,180,31,196,31,196,30,173,31,131,31,114,31,63,31,153,31,133,31,206,31,196,31,192,31,192,30,248,31,248,30,212,31,17,31,217,31,195,31,51,31,51,30,39,31,39,30,190,31,190,30,110,31,102,31,227,31,223,31,192,31,181,31,181,30,13,31,13,30,29,31,83,31,254,31,254,30,227,31,252,31,9,31,202,31,79,31,103,31,189,31,158,31,8,31,8,30,8,29,222,31,213,31,213,30,222,31,157,31,157,30,248,31,171,31,171,30,146,31,32,31,77,31,153,31,100,31,59,31,181,31,181,30,62,31,39,31,112,31,112,30,53,31,113,31,246,31,212,31,249,31,249,30,150,31,150,30,155,31,155,30,228,31,227,31,12,31,197,31,127,31,127,30,127,29,171,31,12,31,40,31,150,31,85,31,217,31,217,30,217,31,217,30,12,31,12,30,222,31,110,31,110,30,110,29,104,31,140,31,119,31,119,30,9,31,207,31,129,31,164,31,21,31,203,31,203,30,146,31,146,30,146,29,65,31,65,30,64,31,170,31,170,30,213,31,213,30,142,31,123,31,123,30,123,29,244,31,123,31,160,31,150,31,13,31,13,30,13,29,151,31,176,31,192,31,127,31,233,31,163,31,26,31,151,31,87,31,230,31,238,31,210,31,210,30,206,31,197,31,215,31,226,31,226,30,122,31,122,30,246,31,16,31,23,31,23,30,176,31,65,31,65,30,192,31,44,31,50,31,30,31,11,31,234,31,234,30,13,31,138,31,208,31,205,31,205,30,83,31,93,31,204,31,238,31,177,31,177,30,229,31,254,31,164,31,242,31,5,31,229,31,209,31,81,31,228,31,210,31,3,31,122,31,122,30,103,31,121,31,43,31,43,30,9,31,159,31,135,31,237,31,186,31,200,31,51,31,96,31,11,31,240,31,224,31,42,31,215,31,215,30,128,31,172,31,160,31,133,31,133,30,208,31,30,31,94,31,94,30,94,29,85,31,93,31,251,31,80,31,80,30,96,31,95,31,95,30,95,29,7,31,133,31,141,31,141,30,106,31,175,31,210,31,47,31,151,31,189,31,255,31,63,31,136,31,136,30,106,31,37,31,25,31,138,31,252,31,50,31,173,31,225,31,225,30,174,31,115,31,63,31,243,31,87,31,166,31,110,31,156,31,116,31,147,31,147,30,245,31,44,31,191,31,111,31,198,31,210,31,202,31,111,31,173,31,170,31,13,31,80,31,80,30,200,31,200,30,184,31,27,31,27,30,27,29,53,31,128,31,28,31,191,31,3,31,3,30,225,31,218,31,218,30,74,31,74,30,10,31,39,31,11,31,185,31,155,31,240,31,38,31,82,31,80,31,19,31,19,30,19,29,109,31,19,31,229,31,104,31,104,30,114,31,126,31,126,30,40,31,40,30,30,31,213,31,123,31,170,31,189,31,189,30,189,29,189,28,92,31,1,31,150,31,147,31,9,31,32,31,65,31,34,31,205,31,57,31,57,30,203,31,32,31,7,31,236,31,172,31,172,30,216,31,189,31,189,30,81,31,203,31,201,31,164,31,129,31,42,31,82,31,82,30,97,31,74,31,78,31,189,31,243,31,178,31,156,31,113,31,215,31,70,31,176,31,79,31,20,31,94,31,94,30,191,31,190,31,62,31,31,31,180,31,180,30,180,29,37,31,127,31,237,31,135,31,142,31,255,31,88,31,174,31,205,31,182,31,211,31,211,30,140,31,138,31,245,31,207,31,201,31,15,31,21,31,89,31,198,31,255,31,255,30,255,29,255,28,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
