-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_322 is
end project_tb_322;

architecture project_tb_arch_322 of project_tb_322 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 972;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,0,0,57,0,224,0,0,0,0,0,87,0,0,0,127,0,118,0,3,0,113,0,0,0,85,0,0,0,0,0,246,0,184,0,0,0,69,0,195,0,142,0,59,0,86,0,252,0,208,0,25,0,166,0,87,0,251,0,17,0,9,0,181,0,170,0,5,0,102,0,82,0,235,0,157,0,2,0,58,0,85,0,0,0,206,0,148,0,164,0,157,0,0,0,66,0,0,0,23,0,225,0,22,0,0,0,48,0,171,0,0,0,101,0,0,0,74,0,18,0,0,0,47,0,29,0,197,0,177,0,31,0,17,0,36,0,0,0,0,0,111,0,61,0,0,0,125,0,153,0,96,0,20,0,144,0,69,0,50,0,216,0,244,0,170,0,183,0,234,0,124,0,118,0,0,0,58,0,83,0,125,0,1,0,102,0,144,0,245,0,176,0,0,0,41,0,177,0,228,0,23,0,238,0,61,0,0,0,162,0,243,0,123,0,228,0,71,0,0,0,53,0,189,0,201,0,169,0,131,0,238,0,33,0,122,0,136,0,20,0,42,0,23,0,62,0,0,0,203,0,22,0,221,0,228,0,182,0,18,0,156,0,223,0,41,0,142,0,168,0,122,0,231,0,102,0,168,0,148,0,148,0,199,0,119,0,0,0,94,0,17,0,43,0,128,0,59,0,79,0,11,0,179,0,171,0,137,0,19,0,154,0,0,0,9,0,61,0,119,0,33,0,103,0,22,0,115,0,0,0,139,0,28,0,111,0,194,0,9,0,46,0,161,0,182,0,185,0,226,0,60,0,30,0,179,0,166,0,103,0,0,0,0,0,161,0,0,0,253,0,21,0,227,0,60,0,238,0,37,0,212,0,49,0,94,0,81,0,108,0,69,0,83,0,244,0,229,0,184,0,221,0,0,0,5,0,195,0,0,0,37,0,137,0,64,0,14,0,178,0,138,0,24,0,194,0,30,0,25,0,25,0,0,0,180,0,215,0,0,0,17,0,143,0,132,0,88,0,9,0,141,0,80,0,12,0,147,0,0,0,23,0,137,0,204,0,163,0,0,0,0,0,0,0,107,0,161,0,154,0,0,0,210,0,123,0,50,0,12,0,0,0,162,0,88,0,55,0,187,0,168,0,44,0,110,0,216,0,240,0,241,0,123,0,115,0,54,0,232,0,180,0,125,0,22,0,238,0,81,0,48,0,175,0,111,0,124,0,46,0,64,0,91,0,61,0,11,0,192,0,88,0,48,0,49,0,73,0,233,0,214,0,154,0,254,0,252,0,0,0,3,0,247,0,0,0,182,0,0,0,11,0,114,0,134,0,108,0,246,0,0,0,232,0,81,0,5,0,0,0,98,0,135,0,104,0,0,0,193,0,98,0,193,0,140,0,209,0,146,0,0,0,27,0,224,0,60,0,126,0,46,0,162,0,0,0,94,0,243,0,227,0,227,0,239,0,78,0,0,0,123,0,85,0,89,0,71,0,0,0,69,0,0,0,183,0,220,0,154,0,0,0,85,0,15,0,84,0,50,0,0,0,3,0,46,0,2,0,241,0,114,0,119,0,0,0,60,0,0,0,0,0,176,0,197,0,82,0,63,0,0,0,92,0,188,0,22,0,53,0,79,0,178,0,0,0,189,0,205,0,234,0,1,0,170,0,0,0,78,0,0,0,228,0,92,0,0,0,33,0,62,0,49,0,0,0,0,0,0,0,0,0,235,0,12,0,164,0,149,0,0,0,135,0,175,0,0,0,206,0,148,0,210,0,207,0,123,0,0,0,203,0,249,0,0,0,51,0,111,0,228,0,221,0,211,0,58,0,199,0,142,0,53,0,6,0,254,0,0,0,158,0,0,0,1,0,24,0,72,0,0,0,227,0,92,0,188,0,134,0,47,0,160,0,52,0,0,0,0,0,0,0,140,0,255,0,51,0,183,0,197,0,201,0,105,0,71,0,124,0,0,0,14,0,146,0,239,0,75,0,50,0,193,0,30,0,0,0,40,0,43,0,195,0,122,0,18,0,31,0,195,0,229,0,209,0,10,0,218,0,7,0,0,0,0,0,116,0,10,0,240,0,75,0,20,0,47,0,0,0,167,0,11,0,159,0,0,0,166,0,77,0,67,0,0,0,0,0,58,0,197,0,235,0,100,0,170,0,0,0,221,0,126,0,254,0,23,0,215,0,252,0,223,0,193,0,205,0,60,0,124,0,81,0,219,0,202,0,0,0,179,0,220,0,26,0,54,0,99,0,199,0,24,0,151,0,123,0,0,0,218,0,212,0,53,0,85,0,27,0,165,0,216,0,101,0,38,0,253,0,60,0,17,0,92,0,25,0,3,0,0,0,184,0,224,0,159,0,142,0,176,0,101,0,2,0,90,0,11,0,10,0,95,0,88,0,195,0,37,0,191,0,0,0,75,0,171,0,0,0,159,0,209,0,0,0,65,0,120,0,239,0,165,0,223,0,0,0,86,0,214,0,166,0,59,0,220,0,181,0,0,0,198,0,150,0,42,0,178,0,66,0,109,0,0,0,157,0,240,0,0,0,230,0,0,0,91,0,0,0,1,0,235,0,105,0,158,0,0,0,237,0,117,0,100,0,44,0,87,0,2,0,138,0,0,0,133,0,128,0,21,0,246,0,80,0,206,0,106,0,252,0,150,0,0,0,151,0,47,0,0,0,96,0,200,0,156,0,0,0,131,0,127,0,0,0,218,0,0,0,0,0,130,0,161,0,158,0,118,0,254,0,23,0,86,0,185,0,4,0,0,0,0,0,0,0,220,0,54,0,12,0,139,0,90,0,189,0,0,0,187,0,90,0,141,0,165,0,157,0,0,0,176,0,16,0,242,0,27,0,0,0,157,0,55,0,11,0,226,0,78,0,164,0,179,0,124,0,205,0,0,0,0,0,0,0,50,0,91,0,0,0,0,0,102,0,216,0,128,0,0,0,171,0,157,0,156,0,25,0,136,0,219,0,131,0,30,0,229,0,182,0,133,0,229,0,185,0,251,0,72,0,59,0,157,0,185,0,0,0,0,0,0,0,237,0,197,0,219,0,190,0,123,0,108,0,82,0,144,0,226,0,23,0,243,0,83,0,0,0,18,0,0,0,0,0,49,0,1,0,175,0,55,0,199,0,198,0,94,0,0,0,254,0,89,0,84,0,130,0,114,0,9,0,64,0,71,0,133,0,174,0,235,0,61,0,137,0,206,0,179,0,60,0,0,0,54,0,128,0,168,0,162,0,0,0,0,0,0,0,0,0,37,0,0,0,222,0,52,0,33,0,124,0,126,0,166,0,128,0,46,0,0,0,213,0,62,0,16,0,146,0,75,0,201,0,0,0,61,0,250,0,186,0,0,0,24,0,0,0,4,0,65,0,239,0,245,0,211,0,72,0,42,0,0,0,253,0,72,0,79,0,239,0,226,0,32,0,0,0,80,0,6,0,154,0,70,0,0,0,109,0,0,0,130,0,0,0,10,0,132,0,136,0,111,0,44,0,72,0,0,0,180,0,65,0,151,0,0,0,158,0,191,0,244,0,216,0,209,0,235,0,184,0,154,0,229,0,201,0,0,0,195,0,13,0,223,0,63,0,0,0,237,0,1,0,169,0,110,0,143,0,139,0,198,0,58,0,220,0,55,0,124,0,18,0,91,0,162,0,59,0,106,0,0,0,0,0,156,0,249,0,0,0,71,0,167,0,111,0,0,0,194,0,19,0,228,0,0,0,139,0,4,0,17,0,33,0,126,0,0,0,93,0,253,0,203,0,0,0,0,0,190,0,235,0,174,0,62,0,205,0,110,0,0,0,0,0,25,0,188,0,0,0,0,0,120,0,98,0,158,0,225,0,141,0,241,0,244,0,0,0,104,0,118,0,101,0,76,0,0,0,0,0,24,0,0,0,150,0,253,0,0,0,0,0,118,0,0,0,203,0,67,0,124,0,17,0,218,0,0,0,101,0,152,0,121,0,29,0,1,0,187,0,64,0,87,0,208,0,121,0,113,0,233,0,225,0,199,0,0,0,18,0,171,0,173,0,197,0,236,0,190,0,176,0,36,0,224,0,66,0,55,0,189,0,0,0,13,0,238,0,165,0,10,0,0,0,138,0,31,0,0,0,0,0,0,0,100,0,133,0,0,0,247,0,73,0,146,0,0,0,240,0,0,0,0,0,220,0,0,0,44,0,0,0,0,0,166,0,0,0,26,0,173,0,97,0,89,0,70,0,0,0,213,0,0,0,148,0,2,0,0,0,199,0,50,0,0,0,150,0,27,0,115,0,33,0,0,0,26,0,225,0,51,0,0,0,0,0,0,0,12,0,59,0,159,0,159,0,162,0,232,0,140,0,52,0,42,0,48,0);
signal scenario_full  : scenario_type := (169,31,169,30,57,31,224,31,224,30,224,29,87,31,87,30,127,31,118,31,3,31,113,31,113,30,85,31,85,30,85,29,246,31,184,31,184,30,69,31,195,31,142,31,59,31,86,31,252,31,208,31,25,31,166,31,87,31,251,31,17,31,9,31,181,31,170,31,5,31,102,31,82,31,235,31,157,31,2,31,58,31,85,31,85,30,206,31,148,31,164,31,157,31,157,30,66,31,66,30,23,31,225,31,22,31,22,30,48,31,171,31,171,30,101,31,101,30,74,31,18,31,18,30,47,31,29,31,197,31,177,31,31,31,17,31,36,31,36,30,36,29,111,31,61,31,61,30,125,31,153,31,96,31,20,31,144,31,69,31,50,31,216,31,244,31,170,31,183,31,234,31,124,31,118,31,118,30,58,31,83,31,125,31,1,31,102,31,144,31,245,31,176,31,176,30,41,31,177,31,228,31,23,31,238,31,61,31,61,30,162,31,243,31,123,31,228,31,71,31,71,30,53,31,189,31,201,31,169,31,131,31,238,31,33,31,122,31,136,31,20,31,42,31,23,31,62,31,62,30,203,31,22,31,221,31,228,31,182,31,18,31,156,31,223,31,41,31,142,31,168,31,122,31,231,31,102,31,168,31,148,31,148,31,199,31,119,31,119,30,94,31,17,31,43,31,128,31,59,31,79,31,11,31,179,31,171,31,137,31,19,31,154,31,154,30,9,31,61,31,119,31,33,31,103,31,22,31,115,31,115,30,139,31,28,31,111,31,194,31,9,31,46,31,161,31,182,31,185,31,226,31,60,31,30,31,179,31,166,31,103,31,103,30,103,29,161,31,161,30,253,31,21,31,227,31,60,31,238,31,37,31,212,31,49,31,94,31,81,31,108,31,69,31,83,31,244,31,229,31,184,31,221,31,221,30,5,31,195,31,195,30,37,31,137,31,64,31,14,31,178,31,138,31,24,31,194,31,30,31,25,31,25,31,25,30,180,31,215,31,215,30,17,31,143,31,132,31,88,31,9,31,141,31,80,31,12,31,147,31,147,30,23,31,137,31,204,31,163,31,163,30,163,29,163,28,107,31,161,31,154,31,154,30,210,31,123,31,50,31,12,31,12,30,162,31,88,31,55,31,187,31,168,31,44,31,110,31,216,31,240,31,241,31,123,31,115,31,54,31,232,31,180,31,125,31,22,31,238,31,81,31,48,31,175,31,111,31,124,31,46,31,64,31,91,31,61,31,11,31,192,31,88,31,48,31,49,31,73,31,233,31,214,31,154,31,254,31,252,31,252,30,3,31,247,31,247,30,182,31,182,30,11,31,114,31,134,31,108,31,246,31,246,30,232,31,81,31,5,31,5,30,98,31,135,31,104,31,104,30,193,31,98,31,193,31,140,31,209,31,146,31,146,30,27,31,224,31,60,31,126,31,46,31,162,31,162,30,94,31,243,31,227,31,227,31,239,31,78,31,78,30,123,31,85,31,89,31,71,31,71,30,69,31,69,30,183,31,220,31,154,31,154,30,85,31,15,31,84,31,50,31,50,30,3,31,46,31,2,31,241,31,114,31,119,31,119,30,60,31,60,30,60,29,176,31,197,31,82,31,63,31,63,30,92,31,188,31,22,31,53,31,79,31,178,31,178,30,189,31,205,31,234,31,1,31,170,31,170,30,78,31,78,30,228,31,92,31,92,30,33,31,62,31,49,31,49,30,49,29,49,28,49,27,235,31,12,31,164,31,149,31,149,30,135,31,175,31,175,30,206,31,148,31,210,31,207,31,123,31,123,30,203,31,249,31,249,30,51,31,111,31,228,31,221,31,211,31,58,31,199,31,142,31,53,31,6,31,254,31,254,30,158,31,158,30,1,31,24,31,72,31,72,30,227,31,92,31,188,31,134,31,47,31,160,31,52,31,52,30,52,29,52,28,140,31,255,31,51,31,183,31,197,31,201,31,105,31,71,31,124,31,124,30,14,31,146,31,239,31,75,31,50,31,193,31,30,31,30,30,40,31,43,31,195,31,122,31,18,31,31,31,195,31,229,31,209,31,10,31,218,31,7,31,7,30,7,29,116,31,10,31,240,31,75,31,20,31,47,31,47,30,167,31,11,31,159,31,159,30,166,31,77,31,67,31,67,30,67,29,58,31,197,31,235,31,100,31,170,31,170,30,221,31,126,31,254,31,23,31,215,31,252,31,223,31,193,31,205,31,60,31,124,31,81,31,219,31,202,31,202,30,179,31,220,31,26,31,54,31,99,31,199,31,24,31,151,31,123,31,123,30,218,31,212,31,53,31,85,31,27,31,165,31,216,31,101,31,38,31,253,31,60,31,17,31,92,31,25,31,3,31,3,30,184,31,224,31,159,31,142,31,176,31,101,31,2,31,90,31,11,31,10,31,95,31,88,31,195,31,37,31,191,31,191,30,75,31,171,31,171,30,159,31,209,31,209,30,65,31,120,31,239,31,165,31,223,31,223,30,86,31,214,31,166,31,59,31,220,31,181,31,181,30,198,31,150,31,42,31,178,31,66,31,109,31,109,30,157,31,240,31,240,30,230,31,230,30,91,31,91,30,1,31,235,31,105,31,158,31,158,30,237,31,117,31,100,31,44,31,87,31,2,31,138,31,138,30,133,31,128,31,21,31,246,31,80,31,206,31,106,31,252,31,150,31,150,30,151,31,47,31,47,30,96,31,200,31,156,31,156,30,131,31,127,31,127,30,218,31,218,30,218,29,130,31,161,31,158,31,118,31,254,31,23,31,86,31,185,31,4,31,4,30,4,29,4,28,220,31,54,31,12,31,139,31,90,31,189,31,189,30,187,31,90,31,141,31,165,31,157,31,157,30,176,31,16,31,242,31,27,31,27,30,157,31,55,31,11,31,226,31,78,31,164,31,179,31,124,31,205,31,205,30,205,29,205,28,50,31,91,31,91,30,91,29,102,31,216,31,128,31,128,30,171,31,157,31,156,31,25,31,136,31,219,31,131,31,30,31,229,31,182,31,133,31,229,31,185,31,251,31,72,31,59,31,157,31,185,31,185,30,185,29,185,28,237,31,197,31,219,31,190,31,123,31,108,31,82,31,144,31,226,31,23,31,243,31,83,31,83,30,18,31,18,30,18,29,49,31,1,31,175,31,55,31,199,31,198,31,94,31,94,30,254,31,89,31,84,31,130,31,114,31,9,31,64,31,71,31,133,31,174,31,235,31,61,31,137,31,206,31,179,31,60,31,60,30,54,31,128,31,168,31,162,31,162,30,162,29,162,28,162,27,37,31,37,30,222,31,52,31,33,31,124,31,126,31,166,31,128,31,46,31,46,30,213,31,62,31,16,31,146,31,75,31,201,31,201,30,61,31,250,31,186,31,186,30,24,31,24,30,4,31,65,31,239,31,245,31,211,31,72,31,42,31,42,30,253,31,72,31,79,31,239,31,226,31,32,31,32,30,80,31,6,31,154,31,70,31,70,30,109,31,109,30,130,31,130,30,10,31,132,31,136,31,111,31,44,31,72,31,72,30,180,31,65,31,151,31,151,30,158,31,191,31,244,31,216,31,209,31,235,31,184,31,154,31,229,31,201,31,201,30,195,31,13,31,223,31,63,31,63,30,237,31,1,31,169,31,110,31,143,31,139,31,198,31,58,31,220,31,55,31,124,31,18,31,91,31,162,31,59,31,106,31,106,30,106,29,156,31,249,31,249,30,71,31,167,31,111,31,111,30,194,31,19,31,228,31,228,30,139,31,4,31,17,31,33,31,126,31,126,30,93,31,253,31,203,31,203,30,203,29,190,31,235,31,174,31,62,31,205,31,110,31,110,30,110,29,25,31,188,31,188,30,188,29,120,31,98,31,158,31,225,31,141,31,241,31,244,31,244,30,104,31,118,31,101,31,76,31,76,30,76,29,24,31,24,30,150,31,253,31,253,30,253,29,118,31,118,30,203,31,67,31,124,31,17,31,218,31,218,30,101,31,152,31,121,31,29,31,1,31,187,31,64,31,87,31,208,31,121,31,113,31,233,31,225,31,199,31,199,30,18,31,171,31,173,31,197,31,236,31,190,31,176,31,36,31,224,31,66,31,55,31,189,31,189,30,13,31,238,31,165,31,10,31,10,30,138,31,31,31,31,30,31,29,31,28,100,31,133,31,133,30,247,31,73,31,146,31,146,30,240,31,240,30,240,29,220,31,220,30,44,31,44,30,44,29,166,31,166,30,26,31,173,31,97,31,89,31,70,31,70,30,213,31,213,30,148,31,2,31,2,30,199,31,50,31,50,30,150,31,27,31,115,31,33,31,33,30,26,31,225,31,51,31,51,30,51,29,51,28,12,31,59,31,159,31,159,31,162,31,232,31,140,31,52,31,42,31,48,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
