-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 751;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (194,0,0,0,244,0,235,0,0,0,47,0,131,0,77,0,7,0,109,0,0,0,144,0,81,0,171,0,82,0,38,0,220,0,248,0,12,0,176,0,0,0,14,0,0,0,8,0,171,0,225,0,199,0,240,0,104,0,245,0,112,0,168,0,1,0,7,0,178,0,65,0,0,0,20,0,125,0,201,0,0,0,0,0,0,0,231,0,218,0,168,0,62,0,118,0,164,0,82,0,173,0,58,0,0,0,45,0,216,0,74,0,226,0,0,0,186,0,37,0,0,0,114,0,131,0,81,0,0,0,124,0,182,0,216,0,193,0,109,0,221,0,0,0,184,0,143,0,94,0,38,0,0,0,58,0,95,0,193,0,0,0,237,0,35,0,0,0,36,0,161,0,162,0,93,0,56,0,21,0,230,0,100,0,121,0,69,0,120,0,178,0,63,0,78,0,0,0,83,0,113,0,233,0,191,0,160,0,0,0,251,0,0,0,105,0,159,0,0,0,0,0,159,0,183,0,104,0,0,0,132,0,255,0,67,0,0,0,62,0,64,0,234,0,0,0,152,0,5,0,75,0,0,0,0,0,19,0,0,0,0,0,239,0,0,0,216,0,142,0,48,0,0,0,8,0,0,0,111,0,25,0,26,0,0,0,231,0,18,0,11,0,226,0,19,0,118,0,69,0,0,0,163,0,234,0,32,0,117,0,0,0,57,0,175,0,181,0,0,0,44,0,155,0,158,0,41,0,222,0,251,0,0,0,252,0,88,0,237,0,0,0,6,0,165,0,12,0,134,0,173,0,239,0,0,0,0,0,0,0,189,0,45,0,142,0,239,0,255,0,13,0,48,0,219,0,63,0,0,0,178,0,228,0,7,0,0,0,66,0,0,0,245,0,71,0,203,0,0,0,122,0,133,0,0,0,21,0,226,0,226,0,0,0,4,0,0,0,251,0,160,0,0,0,25,0,77,0,54,0,1,0,190,0,0,0,231,0,187,0,44,0,89,0,0,0,104,0,190,0,9,0,0,0,83,0,0,0,0,0,202,0,151,0,0,0,85,0,183,0,136,0,197,0,0,0,0,0,33,0,18,0,140,0,0,0,15,0,4,0,93,0,0,0,215,0,9,0,81,0,0,0,159,0,122,0,175,0,180,0,0,0,146,0,225,0,0,0,216,0,173,0,62,0,253,0,79,0,0,0,0,0,0,0,147,0,70,0,122,0,0,0,221,0,0,0,168,0,147,0,0,0,119,0,216,0,0,0,0,0,130,0,185,0,205,0,87,0,232,0,183,0,0,0,43,0,0,0,234,0,210,0,8,0,0,0,190,0,0,0,149,0,34,0,144,0,107,0,0,0,38,0,173,0,2,0,0,0,57,0,0,0,207,0,101,0,49,0,6,0,0,0,196,0,15,0,241,0,219,0,134,0,0,0,54,0,0,0,0,0,79,0,199,0,0,0,143,0,227,0,15,0,0,0,181,0,253,0,141,0,102,0,73,0,0,0,54,0,9,0,0,0,0,0,0,0,67,0,205,0,138,0,116,0,114,0,0,0,0,0,34,0,0,0,0,0,47,0,229,0,13,0,52,0,235,0,70,0,217,0,167,0,208,0,32,0,205,0,54,0,197,0,34,0,0,0,0,0,146,0,113,0,22,0,148,0,44,0,0,0,0,0,171,0,188,0,83,0,0,0,28,0,0,0,0,0,76,0,0,0,72,0,58,0,69,0,95,0,221,0,18,0,227,0,34,0,140,0,144,0,97,0,39,0,147,0,8,0,57,0,83,0,210,0,238,0,4,0,138,0,0,0,144,0,0,0,224,0,79,0,0,0,0,0,0,0,217,0,47,0,118,0,188,0,72,0,81,0,143,0,0,0,92,0,115,0,231,0,192,0,239,0,0,0,87,0,86,0,45,0,70,0,218,0,0,0,87,0,89,0,0,0,0,0,203,0,60,0,10,0,5,0,55,0,0,0,225,0,239,0,135,0,15,0,138,0,185,0,184,0,12,0,189,0,25,0,170,0,153,0,125,0,114,0,25,0,72,0,185,0,175,0,111,0,154,0,149,0,47,0,166,0,161,0,88,0,93,0,4,0,0,0,0,0,190,0,43,0,15,0,34,0,3,0,57,0,62,0,189,0,16,0,36,0,138,0,6,0,23,0,157,0,0,0,202,0,6,0,213,0,223,0,81,0,0,0,0,0,247,0,162,0,127,0,201,0,55,0,164,0,27,0,131,0,172,0,44,0,32,0,197,0,0,0,206,0,188,0,80,0,188,0,0,0,0,0,61,0,138,0,0,0,236,0,140,0,27,0,34,0,166,0,69,0,164,0,6,0,163,0,77,0,0,0,188,0,97,0,0,0,233,0,230,0,239,0,0,0,2,0,164,0,146,0,244,0,119,0,181,0,230,0,31,0,81,0,131,0,40,0,169,0,0,0,186,0,148,0,0,0,0,0,68,0,234,0,63,0,188,0,224,0,129,0,124,0,123,0,147,0,80,0,170,0,204,0,0,0,50,0,103,0,27,0,131,0,0,0,252,0,0,0,102,0,0,0,203,0,0,0,117,0,188,0,0,0,214,0,232,0,74,0,0,0,0,0,124,0,81,0,43,0,135,0,13,0,0,0,33,0,164,0,120,0,211,0,129,0,46,0,205,0,26,0,0,0,74,0,126,0,23,0,13,0,0,0,217,0,153,0,80,0,128,0,37,0,109,0,159,0,59,0,38,0,0,0,143,0,0,0,15,0,135,0,96,0,93,0,239,0,140,0,172,0,160,0,106,0,52,0,80,0,69,0,118,0,0,0,11,0,121,0,31,0,10,0,243,0,48,0,82,0,83,0,0,0,24,0,2,0,224,0,15,0,207,0,106,0,234,0,254,0,4,0,78,0,132,0,15,0,107,0,23,0,0,0,87,0,0,0,0,0,150,0,77,0,22,0,54,0,0,0,166,0,131,0,134,0,110,0,0,0,0,0,0,0,250,0,115,0,59,0,90,0,248,0,0,0,0,0,215,0,239,0,203,0,74,0,240,0,29,0,246,0,179,0,0,0,107,0,190,0,162,0,161,0,0,0,219,0,1,0,15,0,155,0,0,0,87,0,104,0,0,0,0,0,105,0,242,0,203,0,226,0,234,0,74,0,214,0,94,0,68,0,0,0,202,0,151,0,8,0,238,0,0,0,234,0,97,0,108,0,185,0,159,0,180,0,157,0,165,0,115,0,0,0,148,0,0,0,80,0,42,0,146,0,42,0,152,0,183,0,255,0,184,0,0,0,0,0,196,0,0,0,76,0,17,0,0,0,216,0,0,0,0,0,206,0,36,0,220,0,173,0,75,0,131,0,153,0,0,0,145,0,223,0,250,0,179,0,0,0);
signal scenario_full  : scenario_type := (194,31,194,30,244,31,235,31,235,30,47,31,131,31,77,31,7,31,109,31,109,30,144,31,81,31,171,31,82,31,38,31,220,31,248,31,12,31,176,31,176,30,14,31,14,30,8,31,171,31,225,31,199,31,240,31,104,31,245,31,112,31,168,31,1,31,7,31,178,31,65,31,65,30,20,31,125,31,201,31,201,30,201,29,201,28,231,31,218,31,168,31,62,31,118,31,164,31,82,31,173,31,58,31,58,30,45,31,216,31,74,31,226,31,226,30,186,31,37,31,37,30,114,31,131,31,81,31,81,30,124,31,182,31,216,31,193,31,109,31,221,31,221,30,184,31,143,31,94,31,38,31,38,30,58,31,95,31,193,31,193,30,237,31,35,31,35,30,36,31,161,31,162,31,93,31,56,31,21,31,230,31,100,31,121,31,69,31,120,31,178,31,63,31,78,31,78,30,83,31,113,31,233,31,191,31,160,31,160,30,251,31,251,30,105,31,159,31,159,30,159,29,159,31,183,31,104,31,104,30,132,31,255,31,67,31,67,30,62,31,64,31,234,31,234,30,152,31,5,31,75,31,75,30,75,29,19,31,19,30,19,29,239,31,239,30,216,31,142,31,48,31,48,30,8,31,8,30,111,31,25,31,26,31,26,30,231,31,18,31,11,31,226,31,19,31,118,31,69,31,69,30,163,31,234,31,32,31,117,31,117,30,57,31,175,31,181,31,181,30,44,31,155,31,158,31,41,31,222,31,251,31,251,30,252,31,88,31,237,31,237,30,6,31,165,31,12,31,134,31,173,31,239,31,239,30,239,29,239,28,189,31,45,31,142,31,239,31,255,31,13,31,48,31,219,31,63,31,63,30,178,31,228,31,7,31,7,30,66,31,66,30,245,31,71,31,203,31,203,30,122,31,133,31,133,30,21,31,226,31,226,31,226,30,4,31,4,30,251,31,160,31,160,30,25,31,77,31,54,31,1,31,190,31,190,30,231,31,187,31,44,31,89,31,89,30,104,31,190,31,9,31,9,30,83,31,83,30,83,29,202,31,151,31,151,30,85,31,183,31,136,31,197,31,197,30,197,29,33,31,18,31,140,31,140,30,15,31,4,31,93,31,93,30,215,31,9,31,81,31,81,30,159,31,122,31,175,31,180,31,180,30,146,31,225,31,225,30,216,31,173,31,62,31,253,31,79,31,79,30,79,29,79,28,147,31,70,31,122,31,122,30,221,31,221,30,168,31,147,31,147,30,119,31,216,31,216,30,216,29,130,31,185,31,205,31,87,31,232,31,183,31,183,30,43,31,43,30,234,31,210,31,8,31,8,30,190,31,190,30,149,31,34,31,144,31,107,31,107,30,38,31,173,31,2,31,2,30,57,31,57,30,207,31,101,31,49,31,6,31,6,30,196,31,15,31,241,31,219,31,134,31,134,30,54,31,54,30,54,29,79,31,199,31,199,30,143,31,227,31,15,31,15,30,181,31,253,31,141,31,102,31,73,31,73,30,54,31,9,31,9,30,9,29,9,28,67,31,205,31,138,31,116,31,114,31,114,30,114,29,34,31,34,30,34,29,47,31,229,31,13,31,52,31,235,31,70,31,217,31,167,31,208,31,32,31,205,31,54,31,197,31,34,31,34,30,34,29,146,31,113,31,22,31,148,31,44,31,44,30,44,29,171,31,188,31,83,31,83,30,28,31,28,30,28,29,76,31,76,30,72,31,58,31,69,31,95,31,221,31,18,31,227,31,34,31,140,31,144,31,97,31,39,31,147,31,8,31,57,31,83,31,210,31,238,31,4,31,138,31,138,30,144,31,144,30,224,31,79,31,79,30,79,29,79,28,217,31,47,31,118,31,188,31,72,31,81,31,143,31,143,30,92,31,115,31,231,31,192,31,239,31,239,30,87,31,86,31,45,31,70,31,218,31,218,30,87,31,89,31,89,30,89,29,203,31,60,31,10,31,5,31,55,31,55,30,225,31,239,31,135,31,15,31,138,31,185,31,184,31,12,31,189,31,25,31,170,31,153,31,125,31,114,31,25,31,72,31,185,31,175,31,111,31,154,31,149,31,47,31,166,31,161,31,88,31,93,31,4,31,4,30,4,29,190,31,43,31,15,31,34,31,3,31,57,31,62,31,189,31,16,31,36,31,138,31,6,31,23,31,157,31,157,30,202,31,6,31,213,31,223,31,81,31,81,30,81,29,247,31,162,31,127,31,201,31,55,31,164,31,27,31,131,31,172,31,44,31,32,31,197,31,197,30,206,31,188,31,80,31,188,31,188,30,188,29,61,31,138,31,138,30,236,31,140,31,27,31,34,31,166,31,69,31,164,31,6,31,163,31,77,31,77,30,188,31,97,31,97,30,233,31,230,31,239,31,239,30,2,31,164,31,146,31,244,31,119,31,181,31,230,31,31,31,81,31,131,31,40,31,169,31,169,30,186,31,148,31,148,30,148,29,68,31,234,31,63,31,188,31,224,31,129,31,124,31,123,31,147,31,80,31,170,31,204,31,204,30,50,31,103,31,27,31,131,31,131,30,252,31,252,30,102,31,102,30,203,31,203,30,117,31,188,31,188,30,214,31,232,31,74,31,74,30,74,29,124,31,81,31,43,31,135,31,13,31,13,30,33,31,164,31,120,31,211,31,129,31,46,31,205,31,26,31,26,30,74,31,126,31,23,31,13,31,13,30,217,31,153,31,80,31,128,31,37,31,109,31,159,31,59,31,38,31,38,30,143,31,143,30,15,31,135,31,96,31,93,31,239,31,140,31,172,31,160,31,106,31,52,31,80,31,69,31,118,31,118,30,11,31,121,31,31,31,10,31,243,31,48,31,82,31,83,31,83,30,24,31,2,31,224,31,15,31,207,31,106,31,234,31,254,31,4,31,78,31,132,31,15,31,107,31,23,31,23,30,87,31,87,30,87,29,150,31,77,31,22,31,54,31,54,30,166,31,131,31,134,31,110,31,110,30,110,29,110,28,250,31,115,31,59,31,90,31,248,31,248,30,248,29,215,31,239,31,203,31,74,31,240,31,29,31,246,31,179,31,179,30,107,31,190,31,162,31,161,31,161,30,219,31,1,31,15,31,155,31,155,30,87,31,104,31,104,30,104,29,105,31,242,31,203,31,226,31,234,31,74,31,214,31,94,31,68,31,68,30,202,31,151,31,8,31,238,31,238,30,234,31,97,31,108,31,185,31,159,31,180,31,157,31,165,31,115,31,115,30,148,31,148,30,80,31,42,31,146,31,42,31,152,31,183,31,255,31,184,31,184,30,184,29,196,31,196,30,76,31,17,31,17,30,216,31,216,30,216,29,206,31,36,31,220,31,173,31,75,31,131,31,153,31,153,30,145,31,223,31,250,31,179,31,179,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
