-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_65 is
end project_tb_65;

architecture project_tb_arch_65 of project_tb_65 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 867;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,226,0,211,0,41,0,190,0,0,0,132,0,173,0,66,0,64,0,107,0,124,0,17,0,4,0,175,0,0,0,152,0,0,0,87,0,74,0,169,0,0,0,251,0,180,0,9,0,179,0,118,0,175,0,119,0,0,0,169,0,1,0,220,0,0,0,120,0,189,0,70,0,0,0,0,0,0,0,222,0,24,0,225,0,89,0,248,0,0,0,158,0,0,0,111,0,44,0,154,0,123,0,0,0,23,0,65,0,17,0,27,0,252,0,44,0,130,0,224,0,184,0,114,0,145,0,213,0,156,0,0,0,5,0,102,0,244,0,160,0,0,0,15,0,215,0,0,0,90,0,129,0,151,0,215,0,14,0,0,0,0,0,243,0,172,0,76,0,227,0,197,0,242,0,155,0,167,0,72,0,0,0,0,0,215,0,20,0,67,0,15,0,121,0,136,0,222,0,167,0,0,0,9,0,9,0,0,0,38,0,0,0,245,0,134,0,89,0,54,0,47,0,146,0,111,0,45,0,153,0,84,0,0,0,53,0,181,0,94,0,32,0,44,0,151,0,201,0,21,0,72,0,117,0,135,0,0,0,111,0,0,0,0,0,63,0,236,0,0,0,223,0,198,0,0,0,221,0,202,0,248,0,91,0,17,0,148,0,73,0,129,0,154,0,61,0,85,0,233,0,0,0,28,0,252,0,59,0,0,0,251,0,147,0,48,0,126,0,243,0,28,0,0,0,122,0,162,0,31,0,70,0,64,0,59,0,53,0,223,0,16,0,0,0,0,0,24,0,0,0,220,0,9,0,45,0,0,0,0,0,166,0,249,0,122,0,179,0,12,0,0,0,0,0,227,0,44,0,120,0,239,0,0,0,111,0,0,0,155,0,228,0,26,0,30,0,226,0,222,0,169,0,224,0,183,0,134,0,43,0,84,0,161,0,0,0,160,0,26,0,0,0,238,0,53,0,139,0,0,0,174,0,62,0,132,0,9,0,63,0,103,0,124,0,108,0,0,0,68,0,136,0,113,0,0,0,60,0,59,0,0,0,242,0,110,0,76,0,114,0,57,0,141,0,19,0,217,0,68,0,111,0,30,0,21,0,99,0,207,0,30,0,0,0,248,0,190,0,58,0,0,0,183,0,98,0,225,0,111,0,0,0,126,0,0,0,0,0,176,0,165,0,8,0,174,0,117,0,4,0,36,0,70,0,246,0,0,0,0,0,19,0,168,0,0,0,70,0,0,0,158,0,68,0,129,0,235,0,143,0,26,0,219,0,0,0,200,0,203,0,159,0,0,0,229,0,109,0,0,0,99,0,249,0,148,0,196,0,87,0,150,0,159,0,232,0,189,0,35,0,229,0,132,0,168,0,25,0,162,0,103,0,122,0,90,0,74,0,0,0,0,0,0,0,0,0,23,0,175,0,214,0,240,0,201,0,0,0,0,0,58,0,100,0,129,0,250,0,255,0,236,0,227,0,170,0,34,0,18,0,242,0,11,0,169,0,241,0,124,0,0,0,216,0,175,0,0,0,66,0,218,0,152,0,9,0,179,0,71,0,18,0,0,0,153,0,7,0,112,0,0,0,0,0,51,0,0,0,84,0,159,0,0,0,0,0,9,0,210,0,60,0,96,0,198,0,0,0,205,0,0,0,0,0,87,0,77,0,221,0,0,0,137,0,87,0,158,0,151,0,166,0,0,0,120,0,0,0,67,0,77,0,0,0,101,0,93,0,83,0,223,0,132,0,0,0,228,0,251,0,200,0,153,0,118,0,156,0,0,0,142,0,147,0,127,0,0,0,106,0,193,0,0,0,135,0,12,0,235,0,225,0,227,0,127,0,160,0,149,0,200,0,35,0,0,0,88,0,251,0,107,0,24,0,32,0,253,0,84,0,215,0,0,0,36,0,0,0,0,0,56,0,246,0,9,0,0,0,0,0,196,0,44,0,226,0,77,0,207,0,220,0,230,0,40,0,219,0,251,0,78,0,45,0,105,0,113,0,92,0,10,0,113,0,187,0,99,0,220,0,104,0,176,0,250,0,221,0,108,0,201,0,228,0,0,0,239,0,0,0,18,0,75,0,126,0,125,0,231,0,255,0,161,0,95,0,140,0,0,0,232,0,233,0,130,0,245,0,22,0,97,0,119,0,193,0,75,0,97,0,224,0,225,0,94,0,0,0,171,0,122,0,154,0,13,0,121,0,0,0,200,0,34,0,0,0,108,0,0,0,0,0,144,0,27,0,99,0,141,0,62,0,0,0,206,0,98,0,0,0,25,0,222,0,139,0,0,0,0,0,0,0,118,0,134,0,21,0,247,0,221,0,209,0,183,0,52,0,135,0,20,0,250,0,0,0,146,0,35,0,62,0,53,0,0,0,0,0,0,0,0,0,255,0,136,0,204,0,149,0,0,0,19,0,229,0,183,0,0,0,221,0,50,0,128,0,135,0,184,0,148,0,0,0,0,0,0,0,197,0,187,0,1,0,0,0,0,0,18,0,100,0,145,0,55,0,57,0,139,0,205,0,171,0,3,0,72,0,8,0,155,0,0,0,0,0,0,0,235,0,107,0,177,0,0,0,9,0,0,0,80,0,224,0,79,0,78,0,160,0,60,0,188,0,0,0,0,0,55,0,150,0,0,0,210,0,25,0,124,0,124,0,227,0,0,0,0,0,63,0,218,0,204,0,3,0,52,0,205,0,95,0,0,0,183,0,158,0,94,0,23,0,101,0,115,0,212,0,121,0,12,0,199,0,240,0,169,0,105,0,39,0,0,0,177,0,69,0,179,0,24,0,170,0,173,0,20,0,48,0,0,0,239,0,157,0,189,0,0,0,0,0,6,0,90,0,0,0,208,0,144,0,254,0,187,0,80,0,99,0,121,0,8,0,139,0,16,0,6,0,0,0,20,0,0,0,0,0,142,0,135,0,155,0,250,0,72,0,238,0,163,0,0,0,0,0,0,0,244,0,85,0,255,0,35,0,246,0,128,0,253,0,103,0,160,0,67,0,144,0,0,0,93,0,52,0,217,0,44,0,67,0,0,0,41,0,230,0,140,0,0,0,248,0,31,0,57,0,215,0,67,0,29,0,29,0,0,0,209,0,184,0,0,0,193,0,204,0,71,0,238,0,198,0,176,0,0,0,140,0,149,0,231,0,34,0,23,0,157,0,56,0,28,0,222,0,193,0,178,0,0,0,115,0,150,0,86,0,212,0,149,0,170,0,135,0,0,0,0,0,100,0,146,0,44,0,162,0,167,0,0,0,198,0,84,0,204,0,231,0,94,0,0,0,16,0,203,0,23,0,101,0,58,0,162,0,252,0,75,0,0,0,145,0,76,0,56,0,216,0,13,0,84,0,191,0,52,0,113,0,148,0,11,0,143,0,0,0,10,0,205,0,48,0,49,0,136,0,67,0,0,0,78,0,40,0,244,0,141,0,153,0,133,0,0,0,71,0,205,0,35,0,16,0,132,0,244,0,0,0,106,0,141,0,0,0,76,0,169,0,190,0,0,0,45,0,196,0,22,0,104,0,56,0,174,0,213,0,143,0,59,0,102,0,35,0,0,0,132,0,204,0,111,0,254,0,228,0,82,0,32,0,69,0,140,0,94,0,17,0,34,0,157,0,86,0,98,0,58,0,196,0,22,0,90,0,55,0,86,0,47,0,180,0,7,0,0,0,153,0,165,0,206,0,0,0,60,0,152,0,0,0,0,0,42,0,0,0,0,0,9,0,158,0,245,0,209,0,219,0,0,0,208,0,127,0,112,0,157,0,0,0,25,0,44,0,101,0,92,0,194,0,36,0,166,0,21,0,38,0,251,0,0,0,212,0,181,0,180,0,224,0,0,0,0,0,96,0,0,0,195,0,113,0,201,0,204,0,63,0);
signal scenario_full  : scenario_type := (0,0,0,0,226,31,211,31,41,31,190,31,190,30,132,31,173,31,66,31,64,31,107,31,124,31,17,31,4,31,175,31,175,30,152,31,152,30,87,31,74,31,169,31,169,30,251,31,180,31,9,31,179,31,118,31,175,31,119,31,119,30,169,31,1,31,220,31,220,30,120,31,189,31,70,31,70,30,70,29,70,28,222,31,24,31,225,31,89,31,248,31,248,30,158,31,158,30,111,31,44,31,154,31,123,31,123,30,23,31,65,31,17,31,27,31,252,31,44,31,130,31,224,31,184,31,114,31,145,31,213,31,156,31,156,30,5,31,102,31,244,31,160,31,160,30,15,31,215,31,215,30,90,31,129,31,151,31,215,31,14,31,14,30,14,29,243,31,172,31,76,31,227,31,197,31,242,31,155,31,167,31,72,31,72,30,72,29,215,31,20,31,67,31,15,31,121,31,136,31,222,31,167,31,167,30,9,31,9,31,9,30,38,31,38,30,245,31,134,31,89,31,54,31,47,31,146,31,111,31,45,31,153,31,84,31,84,30,53,31,181,31,94,31,32,31,44,31,151,31,201,31,21,31,72,31,117,31,135,31,135,30,111,31,111,30,111,29,63,31,236,31,236,30,223,31,198,31,198,30,221,31,202,31,248,31,91,31,17,31,148,31,73,31,129,31,154,31,61,31,85,31,233,31,233,30,28,31,252,31,59,31,59,30,251,31,147,31,48,31,126,31,243,31,28,31,28,30,122,31,162,31,31,31,70,31,64,31,59,31,53,31,223,31,16,31,16,30,16,29,24,31,24,30,220,31,9,31,45,31,45,30,45,29,166,31,249,31,122,31,179,31,12,31,12,30,12,29,227,31,44,31,120,31,239,31,239,30,111,31,111,30,155,31,228,31,26,31,30,31,226,31,222,31,169,31,224,31,183,31,134,31,43,31,84,31,161,31,161,30,160,31,26,31,26,30,238,31,53,31,139,31,139,30,174,31,62,31,132,31,9,31,63,31,103,31,124,31,108,31,108,30,68,31,136,31,113,31,113,30,60,31,59,31,59,30,242,31,110,31,76,31,114,31,57,31,141,31,19,31,217,31,68,31,111,31,30,31,21,31,99,31,207,31,30,31,30,30,248,31,190,31,58,31,58,30,183,31,98,31,225,31,111,31,111,30,126,31,126,30,126,29,176,31,165,31,8,31,174,31,117,31,4,31,36,31,70,31,246,31,246,30,246,29,19,31,168,31,168,30,70,31,70,30,158,31,68,31,129,31,235,31,143,31,26,31,219,31,219,30,200,31,203,31,159,31,159,30,229,31,109,31,109,30,99,31,249,31,148,31,196,31,87,31,150,31,159,31,232,31,189,31,35,31,229,31,132,31,168,31,25,31,162,31,103,31,122,31,90,31,74,31,74,30,74,29,74,28,74,27,23,31,175,31,214,31,240,31,201,31,201,30,201,29,58,31,100,31,129,31,250,31,255,31,236,31,227,31,170,31,34,31,18,31,242,31,11,31,169,31,241,31,124,31,124,30,216,31,175,31,175,30,66,31,218,31,152,31,9,31,179,31,71,31,18,31,18,30,153,31,7,31,112,31,112,30,112,29,51,31,51,30,84,31,159,31,159,30,159,29,9,31,210,31,60,31,96,31,198,31,198,30,205,31,205,30,205,29,87,31,77,31,221,31,221,30,137,31,87,31,158,31,151,31,166,31,166,30,120,31,120,30,67,31,77,31,77,30,101,31,93,31,83,31,223,31,132,31,132,30,228,31,251,31,200,31,153,31,118,31,156,31,156,30,142,31,147,31,127,31,127,30,106,31,193,31,193,30,135,31,12,31,235,31,225,31,227,31,127,31,160,31,149,31,200,31,35,31,35,30,88,31,251,31,107,31,24,31,32,31,253,31,84,31,215,31,215,30,36,31,36,30,36,29,56,31,246,31,9,31,9,30,9,29,196,31,44,31,226,31,77,31,207,31,220,31,230,31,40,31,219,31,251,31,78,31,45,31,105,31,113,31,92,31,10,31,113,31,187,31,99,31,220,31,104,31,176,31,250,31,221,31,108,31,201,31,228,31,228,30,239,31,239,30,18,31,75,31,126,31,125,31,231,31,255,31,161,31,95,31,140,31,140,30,232,31,233,31,130,31,245,31,22,31,97,31,119,31,193,31,75,31,97,31,224,31,225,31,94,31,94,30,171,31,122,31,154,31,13,31,121,31,121,30,200,31,34,31,34,30,108,31,108,30,108,29,144,31,27,31,99,31,141,31,62,31,62,30,206,31,98,31,98,30,25,31,222,31,139,31,139,30,139,29,139,28,118,31,134,31,21,31,247,31,221,31,209,31,183,31,52,31,135,31,20,31,250,31,250,30,146,31,35,31,62,31,53,31,53,30,53,29,53,28,53,27,255,31,136,31,204,31,149,31,149,30,19,31,229,31,183,31,183,30,221,31,50,31,128,31,135,31,184,31,148,31,148,30,148,29,148,28,197,31,187,31,1,31,1,30,1,29,18,31,100,31,145,31,55,31,57,31,139,31,205,31,171,31,3,31,72,31,8,31,155,31,155,30,155,29,155,28,235,31,107,31,177,31,177,30,9,31,9,30,80,31,224,31,79,31,78,31,160,31,60,31,188,31,188,30,188,29,55,31,150,31,150,30,210,31,25,31,124,31,124,31,227,31,227,30,227,29,63,31,218,31,204,31,3,31,52,31,205,31,95,31,95,30,183,31,158,31,94,31,23,31,101,31,115,31,212,31,121,31,12,31,199,31,240,31,169,31,105,31,39,31,39,30,177,31,69,31,179,31,24,31,170,31,173,31,20,31,48,31,48,30,239,31,157,31,189,31,189,30,189,29,6,31,90,31,90,30,208,31,144,31,254,31,187,31,80,31,99,31,121,31,8,31,139,31,16,31,6,31,6,30,20,31,20,30,20,29,142,31,135,31,155,31,250,31,72,31,238,31,163,31,163,30,163,29,163,28,244,31,85,31,255,31,35,31,246,31,128,31,253,31,103,31,160,31,67,31,144,31,144,30,93,31,52,31,217,31,44,31,67,31,67,30,41,31,230,31,140,31,140,30,248,31,31,31,57,31,215,31,67,31,29,31,29,31,29,30,209,31,184,31,184,30,193,31,204,31,71,31,238,31,198,31,176,31,176,30,140,31,149,31,231,31,34,31,23,31,157,31,56,31,28,31,222,31,193,31,178,31,178,30,115,31,150,31,86,31,212,31,149,31,170,31,135,31,135,30,135,29,100,31,146,31,44,31,162,31,167,31,167,30,198,31,84,31,204,31,231,31,94,31,94,30,16,31,203,31,23,31,101,31,58,31,162,31,252,31,75,31,75,30,145,31,76,31,56,31,216,31,13,31,84,31,191,31,52,31,113,31,148,31,11,31,143,31,143,30,10,31,205,31,48,31,49,31,136,31,67,31,67,30,78,31,40,31,244,31,141,31,153,31,133,31,133,30,71,31,205,31,35,31,16,31,132,31,244,31,244,30,106,31,141,31,141,30,76,31,169,31,190,31,190,30,45,31,196,31,22,31,104,31,56,31,174,31,213,31,143,31,59,31,102,31,35,31,35,30,132,31,204,31,111,31,254,31,228,31,82,31,32,31,69,31,140,31,94,31,17,31,34,31,157,31,86,31,98,31,58,31,196,31,22,31,90,31,55,31,86,31,47,31,180,31,7,31,7,30,153,31,165,31,206,31,206,30,60,31,152,31,152,30,152,29,42,31,42,30,42,29,9,31,158,31,245,31,209,31,219,31,219,30,208,31,127,31,112,31,157,31,157,30,25,31,44,31,101,31,92,31,194,31,36,31,166,31,21,31,38,31,251,31,251,30,212,31,181,31,180,31,224,31,224,30,224,29,96,31,96,30,195,31,113,31,201,31,204,31,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
