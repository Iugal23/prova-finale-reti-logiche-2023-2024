-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 611;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,95,0,0,0,186,0,0,0,54,0,60,0,55,0,0,0,111,0,153,0,73,0,0,0,204,0,79,0,178,0,206,0,199,0,92,0,0,0,26,0,0,0,0,0,116,0,233,0,42,0,84,0,86,0,173,0,160,0,184,0,220,0,145,0,0,0,30,0,38,0,0,0,31,0,88,0,158,0,0,0,0,0,145,0,178,0,57,0,209,0,0,0,64,0,86,0,189,0,249,0,204,0,111,0,4,0,37,0,3,0,56,0,141,0,0,0,152,0,157,0,174,0,0,0,0,0,0,0,126,0,153,0,150,0,0,0,0,0,187,0,205,0,4,0,238,0,241,0,253,0,0,0,249,0,60,0,83,0,104,0,232,0,29,0,35,0,171,0,0,0,184,0,0,0,17,0,231,0,212,0,190,0,248,0,244,0,242,0,186,0,209,0,155,0,0,0,0,0,224,0,0,0,50,0,0,0,149,0,216,0,0,0,167,0,167,0,53,0,162,0,208,0,8,0,0,0,86,0,69,0,0,0,165,0,36,0,222,0,42,0,0,0,137,0,0,0,159,0,108,0,94,0,75,0,222,0,0,0,210,0,211,0,104,0,111,0,238,0,80,0,181,0,62,0,233,0,234,0,126,0,0,0,218,0,49,0,108,0,47,0,44,0,42,0,214,0,192,0,211,0,0,0,196,0,45,0,43,0,120,0,19,0,77,0,147,0,122,0,114,0,251,0,0,0,133,0,103,0,234,0,46,0,0,0,188,0,48,0,0,0,207,0,151,0,0,0,43,0,249,0,97,0,127,0,61,0,0,0,0,0,0,0,127,0,164,0,100,0,129,0,139,0,177,0,16,0,70,0,233,0,34,0,38,0,52,0,56,0,127,0,0,0,67,0,146,0,226,0,192,0,1,0,27,0,201,0,166,0,81,0,0,0,30,0,77,0,6,0,194,0,169,0,194,0,122,0,222,0,167,0,163,0,0,0,228,0,0,0,50,0,45,0,0,0,193,0,4,0,121,0,0,0,195,0,0,0,0,0,0,0,149,0,84,0,181,0,0,0,62,0,77,0,232,0,142,0,49,0,0,0,71,0,181,0,213,0,0,0,17,0,53,0,6,0,207,0,242,0,18,0,202,0,240,0,53,0,91,0,67,0,0,0,162,0,0,0,222,0,0,0,240,0,29,0,193,0,0,0,225,0,0,0,52,0,139,0,113,0,122,0,222,0,143,0,0,0,118,0,127,0,226,0,0,0,219,0,85,0,136,0,105,0,0,0,143,0,0,0,250,0,31,0,0,0,223,0,77,0,239,0,162,0,177,0,177,0,0,0,205,0,175,0,20,0,28,0,21,0,0,0,159,0,106,0,219,0,0,0,207,0,254,0,32,0,178,0,131,0,78,0,121,0,80,0,0,0,0,0,167,0,0,0,240,0,0,0,208,0,13,0,86,0,0,0,185,0,211,0,0,0,19,0,113,0,155,0,30,0,126,0,217,0,160,0,0,0,191,0,63,0,147,0,12,0,0,0,246,0,26,0,0,0,188,0,203,0,1,0,138,0,27,0,13,0,35,0,197,0,0,0,128,0,58,0,0,0,0,0,59,0,15,0,13,0,115,0,0,0,147,0,135,0,0,0,45,0,248,0,0,0,30,0,25,0,246,0,36,0,114,0,0,0,81,0,193,0,0,0,188,0,12,0,137,0,216,0,28,0,53,0,232,0,0,0,0,0,49,0,157,0,122,0,23,0,22,0,0,0,21,0,100,0,0,0,0,0,134,0,153,0,179,0,0,0,13,0,2,0,198,0,22,0,109,0,0,0,161,0,104,0,9,0,35,0,0,0,0,0,25,0,0,0,0,0,72,0,64,0,0,0,200,0,0,0,10,0,160,0,242,0,205,0,0,0,253,0,24,0,183,0,197,0,33,0,245,0,160,0,0,0,94,0,62,0,176,0,177,0,200,0,170,0,240,0,0,0,0,0,137,0,134,0,12,0,0,0,145,0,0,0,127,0,46,0,0,0,160,0,0,0,243,0,125,0,219,0,0,0,37,0,133,0,0,0,152,0,0,0,0,0,238,0,0,0,0,0,168,0,149,0,143,0,88,0,191,0,216,0,161,0,118,0,75,0,0,0,37,0,178,0,104,0,127,0,6,0,200,0,0,0,0,0,0,0,161,0,56,0,65,0,52,0,211,0,0,0,232,0,240,0,14,0,31,0,193,0,234,0,99,0,76,0,119,0,60,0,164,0,105,0,173,0,234,0,207,0,0,0,253,0,101,0,0,0,83,0,142,0,176,0,5,0,66,0,144,0,217,0,113,0,180,0,71,0,75,0,2,0,59,0,244,0,50,0,33,0,71,0,0,0,0,0,0,0,0,0,12,0,91,0,212,0,0,0,82,0,90,0,141,0,0,0,176,0,129,0,0,0,102,0,9,0,0,0,156,0,181,0,0,0,39,0,254,0,251,0,78,0,226,0,39,0,126,0,220,0,172,0,213,0,225,0,98,0,0,0,51,0,250,0,37,0,120,0,153,0,102,0,0,0,39,0,0,0,38,0,226,0,209,0,150,0,106,0,0,0,0,0,115,0,163,0,0,0,70,0,240,0,134,0,6,0,84,0,87,0,208,0,179,0,93,0,21,0,55,0,10,0,227,0,155,0,0,0,15,0,166,0,108,0,218,0,144,0,148,0,20,0,35,0,0,0,122,0,197,0,22,0,29,0,216,0,122,0,227,0,43,0,215,0);
signal scenario_full  : scenario_type := (0,0,95,31,95,30,186,31,186,30,54,31,60,31,55,31,55,30,111,31,153,31,73,31,73,30,204,31,79,31,178,31,206,31,199,31,92,31,92,30,26,31,26,30,26,29,116,31,233,31,42,31,84,31,86,31,173,31,160,31,184,31,220,31,145,31,145,30,30,31,38,31,38,30,31,31,88,31,158,31,158,30,158,29,145,31,178,31,57,31,209,31,209,30,64,31,86,31,189,31,249,31,204,31,111,31,4,31,37,31,3,31,56,31,141,31,141,30,152,31,157,31,174,31,174,30,174,29,174,28,126,31,153,31,150,31,150,30,150,29,187,31,205,31,4,31,238,31,241,31,253,31,253,30,249,31,60,31,83,31,104,31,232,31,29,31,35,31,171,31,171,30,184,31,184,30,17,31,231,31,212,31,190,31,248,31,244,31,242,31,186,31,209,31,155,31,155,30,155,29,224,31,224,30,50,31,50,30,149,31,216,31,216,30,167,31,167,31,53,31,162,31,208,31,8,31,8,30,86,31,69,31,69,30,165,31,36,31,222,31,42,31,42,30,137,31,137,30,159,31,108,31,94,31,75,31,222,31,222,30,210,31,211,31,104,31,111,31,238,31,80,31,181,31,62,31,233,31,234,31,126,31,126,30,218,31,49,31,108,31,47,31,44,31,42,31,214,31,192,31,211,31,211,30,196,31,45,31,43,31,120,31,19,31,77,31,147,31,122,31,114,31,251,31,251,30,133,31,103,31,234,31,46,31,46,30,188,31,48,31,48,30,207,31,151,31,151,30,43,31,249,31,97,31,127,31,61,31,61,30,61,29,61,28,127,31,164,31,100,31,129,31,139,31,177,31,16,31,70,31,233,31,34,31,38,31,52,31,56,31,127,31,127,30,67,31,146,31,226,31,192,31,1,31,27,31,201,31,166,31,81,31,81,30,30,31,77,31,6,31,194,31,169,31,194,31,122,31,222,31,167,31,163,31,163,30,228,31,228,30,50,31,45,31,45,30,193,31,4,31,121,31,121,30,195,31,195,30,195,29,195,28,149,31,84,31,181,31,181,30,62,31,77,31,232,31,142,31,49,31,49,30,71,31,181,31,213,31,213,30,17,31,53,31,6,31,207,31,242,31,18,31,202,31,240,31,53,31,91,31,67,31,67,30,162,31,162,30,222,31,222,30,240,31,29,31,193,31,193,30,225,31,225,30,52,31,139,31,113,31,122,31,222,31,143,31,143,30,118,31,127,31,226,31,226,30,219,31,85,31,136,31,105,31,105,30,143,31,143,30,250,31,31,31,31,30,223,31,77,31,239,31,162,31,177,31,177,31,177,30,205,31,175,31,20,31,28,31,21,31,21,30,159,31,106,31,219,31,219,30,207,31,254,31,32,31,178,31,131,31,78,31,121,31,80,31,80,30,80,29,167,31,167,30,240,31,240,30,208,31,13,31,86,31,86,30,185,31,211,31,211,30,19,31,113,31,155,31,30,31,126,31,217,31,160,31,160,30,191,31,63,31,147,31,12,31,12,30,246,31,26,31,26,30,188,31,203,31,1,31,138,31,27,31,13,31,35,31,197,31,197,30,128,31,58,31,58,30,58,29,59,31,15,31,13,31,115,31,115,30,147,31,135,31,135,30,45,31,248,31,248,30,30,31,25,31,246,31,36,31,114,31,114,30,81,31,193,31,193,30,188,31,12,31,137,31,216,31,28,31,53,31,232,31,232,30,232,29,49,31,157,31,122,31,23,31,22,31,22,30,21,31,100,31,100,30,100,29,134,31,153,31,179,31,179,30,13,31,2,31,198,31,22,31,109,31,109,30,161,31,104,31,9,31,35,31,35,30,35,29,25,31,25,30,25,29,72,31,64,31,64,30,200,31,200,30,10,31,160,31,242,31,205,31,205,30,253,31,24,31,183,31,197,31,33,31,245,31,160,31,160,30,94,31,62,31,176,31,177,31,200,31,170,31,240,31,240,30,240,29,137,31,134,31,12,31,12,30,145,31,145,30,127,31,46,31,46,30,160,31,160,30,243,31,125,31,219,31,219,30,37,31,133,31,133,30,152,31,152,30,152,29,238,31,238,30,238,29,168,31,149,31,143,31,88,31,191,31,216,31,161,31,118,31,75,31,75,30,37,31,178,31,104,31,127,31,6,31,200,31,200,30,200,29,200,28,161,31,56,31,65,31,52,31,211,31,211,30,232,31,240,31,14,31,31,31,193,31,234,31,99,31,76,31,119,31,60,31,164,31,105,31,173,31,234,31,207,31,207,30,253,31,101,31,101,30,83,31,142,31,176,31,5,31,66,31,144,31,217,31,113,31,180,31,71,31,75,31,2,31,59,31,244,31,50,31,33,31,71,31,71,30,71,29,71,28,71,27,12,31,91,31,212,31,212,30,82,31,90,31,141,31,141,30,176,31,129,31,129,30,102,31,9,31,9,30,156,31,181,31,181,30,39,31,254,31,251,31,78,31,226,31,39,31,126,31,220,31,172,31,213,31,225,31,98,31,98,30,51,31,250,31,37,31,120,31,153,31,102,31,102,30,39,31,39,30,38,31,226,31,209,31,150,31,106,31,106,30,106,29,115,31,163,31,163,30,70,31,240,31,134,31,6,31,84,31,87,31,208,31,179,31,93,31,21,31,55,31,10,31,227,31,155,31,155,30,15,31,166,31,108,31,218,31,144,31,148,31,20,31,35,31,35,30,122,31,197,31,22,31,29,31,216,31,122,31,227,31,43,31,215,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
