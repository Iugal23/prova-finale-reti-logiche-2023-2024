-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 981;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,0,0,35,0,62,0,129,0,141,0,71,0,153,0,60,0,32,0,224,0,0,0,235,0,0,0,215,0,132,0,0,0,154,0,117,0,0,0,0,0,207,0,102,0,9,0,14,0,136,0,224,0,135,0,0,0,0,0,21,0,0,0,102,0,0,0,85,0,109,0,173,0,136,0,125,0,91,0,0,0,126,0,183,0,4,0,92,0,114,0,0,0,112,0,239,0,74,0,0,0,46,0,82,0,0,0,39,0,0,0,111,0,119,0,107,0,198,0,30,0,219,0,106,0,204,0,0,0,5,0,231,0,155,0,179,0,126,0,8,0,253,0,195,0,90,0,97,0,255,0,89,0,64,0,0,0,0,0,226,0,148,0,182,0,67,0,250,0,118,0,148,0,164,0,174,0,10,0,112,0,229,0,148,0,0,0,9,0,226,0,220,0,0,0,167,0,243,0,58,0,117,0,119,0,94,0,64,0,220,0,169,0,0,0,45,0,103,0,140,0,208,0,0,0,98,0,95,0,227,0,218,0,81,0,44,0,212,0,111,0,0,0,82,0,98,0,46,0,0,0,58,0,30,0,82,0,200,0,119,0,204,0,19,0,64,0,171,0,205,0,231,0,155,0,24,0,221,0,171,0,160,0,0,0,235,0,133,0,70,0,0,0,89,0,0,0,30,0,126,0,132,0,89,0,207,0,138,0,25,0,0,0,149,0,0,0,0,0,8,0,0,0,206,0,67,0,141,0,0,0,0,0,75,0,0,0,196,0,247,0,6,0,143,0,0,0,132,0,34,0,0,0,183,0,214,0,139,0,224,0,0,0,172,0,180,0,167,0,170,0,60,0,147,0,0,0,189,0,0,0,4,0,0,0,60,0,176,0,29,0,0,0,0,0,77,0,68,0,58,0,74,0,151,0,0,0,0,0,0,0,0,0,0,0,199,0,0,0,0,0,54,0,232,0,77,0,254,0,191,0,234,0,240,0,4,0,190,0,48,0,0,0,0,0,146,0,61,0,38,0,49,0,109,0,239,0,165,0,242,0,200,0,30,0,59,0,0,0,243,0,102,0,111,0,213,0,57,0,8,0,247,0,0,0,79,0,10,0,179,0,194,0,133,0,181,0,202,0,158,0,0,0,0,0,130,0,4,0,142,0,250,0,141,0,116,0,53,0,0,0,105,0,0,0,249,0,202,0,0,0,136,0,236,0,95,0,210,0,85,0,157,0,0,0,96,0,0,0,182,0,22,0,203,0,0,0,218,0,0,0,170,0,19,0,147,0,0,0,0,0,0,0,219,0,0,0,137,0,197,0,13,0,244,0,255,0,81,0,171,0,41,0,243,0,0,0,11,0,0,0,198,0,33,0,188,0,43,0,40,0,12,0,110,0,31,0,189,0,30,0,90,0,67,0,142,0,151,0,152,0,174,0,7,0,71,0,41,0,124,0,248,0,126,0,81,0,0,0,170,0,217,0,127,0,0,0,65,0,0,0,150,0,0,0,0,0,146,0,236,0,246,0,58,0,0,0,71,0,9,0,235,0,93,0,254,0,0,0,18,0,114,0,247,0,0,0,0,0,0,0,62,0,90,0,0,0,0,0,20,0,127,0,243,0,0,0,0,0,122,0,76,0,7,0,28,0,7,0,0,0,60,0,109,0,162,0,197,0,133,0,59,0,67,0,197,0,21,0,67,0,46,0,22,0,186,0,0,0,152,0,71,0,29,0,0,0,0,0,102,0,120,0,150,0,101,0,93,0,0,0,204,0,41,0,79,0,71,0,97,0,19,0,220,0,0,0,188,0,40,0,151,0,80,0,188,0,0,0,85,0,0,0,37,0,87,0,250,0,93,0,147,0,33,0,66,0,110,0,124,0,0,0,0,0,81,0,26,0,127,0,43,0,35,0,0,0,130,0,0,0,44,0,12,0,0,0,0,0,224,0,117,0,49,0,0,0,142,0,68,0,149,0,39,0,215,0,0,0,13,0,13,0,123,0,206,0,79,0,0,0,59,0,0,0,0,0,168,0,255,0,91,0,77,0,0,0,76,0,127,0,0,0,243,0,173,0,0,0,85,0,182,0,155,0,45,0,0,0,0,0,129,0,0,0,0,0,0,0,147,0,0,0,234,0,226,0,0,0,142,0,183,0,50,0,43,0,119,0,95,0,0,0,211,0,0,0,75,0,0,0,87,0,0,0,0,0,43,0,148,0,154,0,31,0,103,0,0,0,0,0,31,0,65,0,244,0,173,0,106,0,50,0,232,0,0,0,152,0,154,0,0,0,78,0,188,0,169,0,0,0,0,0,149,0,224,0,0,0,84,0,141,0,0,0,0,0,36,0,196,0,0,0,6,0,178,0,206,0,105,0,96,0,77,0,18,0,0,0,117,0,36,0,207,0,251,0,127,0,205,0,111,0,192,0,55,0,10,0,132,0,96,0,162,0,0,0,0,0,220,0,0,0,0,0,152,0,36,0,48,0,88,0,183,0,33,0,171,0,0,0,235,0,0,0,0,0,0,0,121,0,91,0,185,0,35,0,245,0,140,0,31,0,0,0,0,0,102,0,238,0,113,0,46,0,0,0,200,0,0,0,0,0,0,0,0,0,82,0,0,0,100,0,0,0,138,0,190,0,0,0,157,0,41,0,0,0,0,0,209,0,73,0,220,0,144,0,0,0,197,0,144,0,0,0,167,0,178,0,35,0,0,0,205,0,0,0,0,0,226,0,75,0,29,0,17,0,138,0,151,0,37,0,198,0,140,0,135,0,181,0,197,0,74,0,119,0,0,0,87,0,131,0,240,0,165,0,25,0,47,0,208,0,140,0,0,0,193,0,180,0,141,0,36,0,0,0,223,0,21,0,117,0,7,0,53,0,81,0,14,0,208,0,168,0,204,0,83,0,40,0,16,0,238,0,0,0,36,0,39,0,109,0,232,0,12,0,43,0,190,0,132,0,236,0,41,0,17,0,0,0,175,0,111,0,12,0,17,0,184,0,41,0,208,0,2,0,0,0,113,0,25,0,64,0,19,0,0,0,168,0,116,0,4,0,53,0,236,0,12,0,0,0,0,0,0,0,107,0,0,0,115,0,38,0,196,0,81,0,114,0,207,0,37,0,0,0,0,0,0,0,246,0,196,0,124,0,181,0,0,0,171,0,102,0,0,0,128,0,122,0,147,0,30,0,0,0,0,0,44,0,28,0,183,0,64,0,36,0,188,0,124,0,0,0,216,0,108,0,109,0,0,0,203,0,68,0,241,0,5,0,0,0,135,0,236,0,37,0,216,0,119,0,136,0,163,0,108,0,170,0,243,0,132,0,37,0,28,0,0,0,25,0,226,0,99,0,161,0,217,0,212,0,33,0,14,0,193,0,161,0,228,0,0,0,65,0,207,0,86,0,51,0,162,0,0,0,208,0,91,0,75,0,96,0,168,0,76,0,0,0,0,0,0,0,0,0,142,0,146,0,0,0,0,0,170,0,246,0,138,0,123,0,0,0,71,0,0,0,0,0,212,0,13,0,129,0,26,0,75,0,45,0,0,0,84,0,152,0,72,0,172,0,0,0,0,0,0,0,192,0,0,0,215,0,192,0,0,0,100,0,214,0,77,0,0,0,0,0,251,0,0,0,54,0,58,0,189,0,189,0,0,0,0,0,243,0,174,0,72,0,28,0,168,0,0,0,28,0,107,0,57,0,74,0,152,0,128,0,44,0,0,0,0,0,60,0,143,0,194,0,64,0,60,0,174,0,112,0,223,0,36,0,145,0,17,0,209,0,89,0,64,0,0,0,22,0,0,0,18,0,0,0,15,0,87,0,145,0,161,0,146,0,246,0,23,0,0,0,0,0,23,0,63,0,145,0,223,0,172,0,135,0,155,0,68,0,183,0,246,0,246,0,67,0,0,0,0,0,68,0,58,0,165,0,0,0,92,0,0,0,247,0,243,0,249,0,169,0,0,0,58,0,57,0,35,0,0,0,182,0,252,0,193,0,57,0,0,0,171,0,0,0,85,0,21,0,131,0,55,0,0,0,77,0,246,0,236,0,58,0,210,0,142,0,105,0,230,0,0,0,0,0,220,0,99,0,129,0,70,0,181,0,0,0,0,0,254,0,218,0,240,0,52,0,0,0,0,0,0,0,0,0,0,0,146,0,14,0,165,0,167,0,48,0,118,0,0,0,43,0,0,0,184,0,76,0,137,0,254,0,45,0,194,0,65,0,0,0,94,0,250,0,0,0,0,0,76,0,155,0,51,0,159,0,2,0,170,0,255,0,119,0,182,0,57,0,99,0,137,0,110,0,9,0,44,0,119,0,172,0,88,0,0,0,27,0,23,0,245,0,141,0,191,0,0,0,156,0,119,0,15,0,184,0,211,0,100,0,169,0,24,0,251,0,135,0,203,0,101,0);
signal scenario_full  : scenario_type := (219,31,219,30,35,31,62,31,129,31,141,31,71,31,153,31,60,31,32,31,224,31,224,30,235,31,235,30,215,31,132,31,132,30,154,31,117,31,117,30,117,29,207,31,102,31,9,31,14,31,136,31,224,31,135,31,135,30,135,29,21,31,21,30,102,31,102,30,85,31,109,31,173,31,136,31,125,31,91,31,91,30,126,31,183,31,4,31,92,31,114,31,114,30,112,31,239,31,74,31,74,30,46,31,82,31,82,30,39,31,39,30,111,31,119,31,107,31,198,31,30,31,219,31,106,31,204,31,204,30,5,31,231,31,155,31,179,31,126,31,8,31,253,31,195,31,90,31,97,31,255,31,89,31,64,31,64,30,64,29,226,31,148,31,182,31,67,31,250,31,118,31,148,31,164,31,174,31,10,31,112,31,229,31,148,31,148,30,9,31,226,31,220,31,220,30,167,31,243,31,58,31,117,31,119,31,94,31,64,31,220,31,169,31,169,30,45,31,103,31,140,31,208,31,208,30,98,31,95,31,227,31,218,31,81,31,44,31,212,31,111,31,111,30,82,31,98,31,46,31,46,30,58,31,30,31,82,31,200,31,119,31,204,31,19,31,64,31,171,31,205,31,231,31,155,31,24,31,221,31,171,31,160,31,160,30,235,31,133,31,70,31,70,30,89,31,89,30,30,31,126,31,132,31,89,31,207,31,138,31,25,31,25,30,149,31,149,30,149,29,8,31,8,30,206,31,67,31,141,31,141,30,141,29,75,31,75,30,196,31,247,31,6,31,143,31,143,30,132,31,34,31,34,30,183,31,214,31,139,31,224,31,224,30,172,31,180,31,167,31,170,31,60,31,147,31,147,30,189,31,189,30,4,31,4,30,60,31,176,31,29,31,29,30,29,29,77,31,68,31,58,31,74,31,151,31,151,30,151,29,151,28,151,27,151,26,199,31,199,30,199,29,54,31,232,31,77,31,254,31,191,31,234,31,240,31,4,31,190,31,48,31,48,30,48,29,146,31,61,31,38,31,49,31,109,31,239,31,165,31,242,31,200,31,30,31,59,31,59,30,243,31,102,31,111,31,213,31,57,31,8,31,247,31,247,30,79,31,10,31,179,31,194,31,133,31,181,31,202,31,158,31,158,30,158,29,130,31,4,31,142,31,250,31,141,31,116,31,53,31,53,30,105,31,105,30,249,31,202,31,202,30,136,31,236,31,95,31,210,31,85,31,157,31,157,30,96,31,96,30,182,31,22,31,203,31,203,30,218,31,218,30,170,31,19,31,147,31,147,30,147,29,147,28,219,31,219,30,137,31,197,31,13,31,244,31,255,31,81,31,171,31,41,31,243,31,243,30,11,31,11,30,198,31,33,31,188,31,43,31,40,31,12,31,110,31,31,31,189,31,30,31,90,31,67,31,142,31,151,31,152,31,174,31,7,31,71,31,41,31,124,31,248,31,126,31,81,31,81,30,170,31,217,31,127,31,127,30,65,31,65,30,150,31,150,30,150,29,146,31,236,31,246,31,58,31,58,30,71,31,9,31,235,31,93,31,254,31,254,30,18,31,114,31,247,31,247,30,247,29,247,28,62,31,90,31,90,30,90,29,20,31,127,31,243,31,243,30,243,29,122,31,76,31,7,31,28,31,7,31,7,30,60,31,109,31,162,31,197,31,133,31,59,31,67,31,197,31,21,31,67,31,46,31,22,31,186,31,186,30,152,31,71,31,29,31,29,30,29,29,102,31,120,31,150,31,101,31,93,31,93,30,204,31,41,31,79,31,71,31,97,31,19,31,220,31,220,30,188,31,40,31,151,31,80,31,188,31,188,30,85,31,85,30,37,31,87,31,250,31,93,31,147,31,33,31,66,31,110,31,124,31,124,30,124,29,81,31,26,31,127,31,43,31,35,31,35,30,130,31,130,30,44,31,12,31,12,30,12,29,224,31,117,31,49,31,49,30,142,31,68,31,149,31,39,31,215,31,215,30,13,31,13,31,123,31,206,31,79,31,79,30,59,31,59,30,59,29,168,31,255,31,91,31,77,31,77,30,76,31,127,31,127,30,243,31,173,31,173,30,85,31,182,31,155,31,45,31,45,30,45,29,129,31,129,30,129,29,129,28,147,31,147,30,234,31,226,31,226,30,142,31,183,31,50,31,43,31,119,31,95,31,95,30,211,31,211,30,75,31,75,30,87,31,87,30,87,29,43,31,148,31,154,31,31,31,103,31,103,30,103,29,31,31,65,31,244,31,173,31,106,31,50,31,232,31,232,30,152,31,154,31,154,30,78,31,188,31,169,31,169,30,169,29,149,31,224,31,224,30,84,31,141,31,141,30,141,29,36,31,196,31,196,30,6,31,178,31,206,31,105,31,96,31,77,31,18,31,18,30,117,31,36,31,207,31,251,31,127,31,205,31,111,31,192,31,55,31,10,31,132,31,96,31,162,31,162,30,162,29,220,31,220,30,220,29,152,31,36,31,48,31,88,31,183,31,33,31,171,31,171,30,235,31,235,30,235,29,235,28,121,31,91,31,185,31,35,31,245,31,140,31,31,31,31,30,31,29,102,31,238,31,113,31,46,31,46,30,200,31,200,30,200,29,200,28,200,27,82,31,82,30,100,31,100,30,138,31,190,31,190,30,157,31,41,31,41,30,41,29,209,31,73,31,220,31,144,31,144,30,197,31,144,31,144,30,167,31,178,31,35,31,35,30,205,31,205,30,205,29,226,31,75,31,29,31,17,31,138,31,151,31,37,31,198,31,140,31,135,31,181,31,197,31,74,31,119,31,119,30,87,31,131,31,240,31,165,31,25,31,47,31,208,31,140,31,140,30,193,31,180,31,141,31,36,31,36,30,223,31,21,31,117,31,7,31,53,31,81,31,14,31,208,31,168,31,204,31,83,31,40,31,16,31,238,31,238,30,36,31,39,31,109,31,232,31,12,31,43,31,190,31,132,31,236,31,41,31,17,31,17,30,175,31,111,31,12,31,17,31,184,31,41,31,208,31,2,31,2,30,113,31,25,31,64,31,19,31,19,30,168,31,116,31,4,31,53,31,236,31,12,31,12,30,12,29,12,28,107,31,107,30,115,31,38,31,196,31,81,31,114,31,207,31,37,31,37,30,37,29,37,28,246,31,196,31,124,31,181,31,181,30,171,31,102,31,102,30,128,31,122,31,147,31,30,31,30,30,30,29,44,31,28,31,183,31,64,31,36,31,188,31,124,31,124,30,216,31,108,31,109,31,109,30,203,31,68,31,241,31,5,31,5,30,135,31,236,31,37,31,216,31,119,31,136,31,163,31,108,31,170,31,243,31,132,31,37,31,28,31,28,30,25,31,226,31,99,31,161,31,217,31,212,31,33,31,14,31,193,31,161,31,228,31,228,30,65,31,207,31,86,31,51,31,162,31,162,30,208,31,91,31,75,31,96,31,168,31,76,31,76,30,76,29,76,28,76,27,142,31,146,31,146,30,146,29,170,31,246,31,138,31,123,31,123,30,71,31,71,30,71,29,212,31,13,31,129,31,26,31,75,31,45,31,45,30,84,31,152,31,72,31,172,31,172,30,172,29,172,28,192,31,192,30,215,31,192,31,192,30,100,31,214,31,77,31,77,30,77,29,251,31,251,30,54,31,58,31,189,31,189,31,189,30,189,29,243,31,174,31,72,31,28,31,168,31,168,30,28,31,107,31,57,31,74,31,152,31,128,31,44,31,44,30,44,29,60,31,143,31,194,31,64,31,60,31,174,31,112,31,223,31,36,31,145,31,17,31,209,31,89,31,64,31,64,30,22,31,22,30,18,31,18,30,15,31,87,31,145,31,161,31,146,31,246,31,23,31,23,30,23,29,23,31,63,31,145,31,223,31,172,31,135,31,155,31,68,31,183,31,246,31,246,31,67,31,67,30,67,29,68,31,58,31,165,31,165,30,92,31,92,30,247,31,243,31,249,31,169,31,169,30,58,31,57,31,35,31,35,30,182,31,252,31,193,31,57,31,57,30,171,31,171,30,85,31,21,31,131,31,55,31,55,30,77,31,246,31,236,31,58,31,210,31,142,31,105,31,230,31,230,30,230,29,220,31,99,31,129,31,70,31,181,31,181,30,181,29,254,31,218,31,240,31,52,31,52,30,52,29,52,28,52,27,52,26,146,31,14,31,165,31,167,31,48,31,118,31,118,30,43,31,43,30,184,31,76,31,137,31,254,31,45,31,194,31,65,31,65,30,94,31,250,31,250,30,250,29,76,31,155,31,51,31,159,31,2,31,170,31,255,31,119,31,182,31,57,31,99,31,137,31,110,31,9,31,44,31,119,31,172,31,88,31,88,30,27,31,23,31,245,31,141,31,191,31,191,30,156,31,119,31,15,31,184,31,211,31,100,31,169,31,24,31,251,31,135,31,203,31,101,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
