-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_607 is
end project_tb_607;

architecture project_tb_arch_607 of project_tb_607 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 637;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (174,0,0,0,127,0,135,0,179,0,0,0,95,0,132,0,4,0,174,0,52,0,122,0,0,0,44,0,0,0,194,0,199,0,129,0,228,0,0,0,79,0,172,0,193,0,0,0,86,0,91,0,166,0,233,0,0,0,218,0,101,0,0,0,87,0,217,0,0,0,101,0,0,0,248,0,158,0,121,0,160,0,0,0,223,0,139,0,50,0,20,0,53,0,115,0,241,0,107,0,0,0,0,0,230,0,153,0,0,0,4,0,120,0,176,0,15,0,0,0,41,0,147,0,0,0,214,0,250,0,32,0,64,0,0,0,68,0,19,0,73,0,0,0,190,0,35,0,128,0,141,0,103,0,28,0,162,0,93,0,10,0,159,0,25,0,68,0,109,0,222,0,78,0,16,0,59,0,0,0,0,0,39,0,0,0,65,0,193,0,193,0,84,0,37,0,153,0,76,0,214,0,0,0,50,0,0,0,0,0,176,0,82,0,175,0,4,0,13,0,239,0,42,0,86,0,213,0,103,0,0,0,0,0,170,0,133,0,224,0,0,0,0,0,235,0,0,0,3,0,118,0,73,0,185,0,192,0,25,0,226,0,237,0,27,0,190,0,50,0,0,0,149,0,155,0,155,0,69,0,130,0,52,0,211,0,15,0,164,0,96,0,204,0,35,0,49,0,174,0,32,0,167,0,89,0,222,0,211,0,232,0,190,0,63,0,189,0,69,0,220,0,54,0,167,0,198,0,254,0,117,0,147,0,0,0,23,0,149,0,130,0,180,0,39,0,196,0,174,0,1,0,114,0,188,0,0,0,162,0,0,0,75,0,174,0,0,0,215,0,115,0,191,0,0,0,159,0,114,0,232,0,247,0,0,0,0,0,182,0,201,0,163,0,196,0,46,0,0,0,165,0,146,0,157,0,48,0,119,0,198,0,0,0,52,0,99,0,126,0,38,0,255,0,59,0,55,0,72,0,234,0,115,0,255,0,21,0,73,0,225,0,157,0,93,0,39,0,227,0,78,0,199,0,253,0,209,0,0,0,51,0,0,0,124,0,77,0,123,0,0,0,76,0,150,0,0,0,194,0,60,0,110,0,0,0,147,0,0,0,70,0,0,0,44,0,182,0,175,0,197,0,228,0,214,0,69,0,206,0,42,0,204,0,209,0,116,0,190,0,25,0,161,0,67,0,0,0,155,0,209,0,0,0,224,0,65,0,0,0,217,0,206,0,13,0,112,0,155,0,87,0,0,0,0,0,20,0,0,0,120,0,210,0,251,0,173,0,168,0,4,0,0,0,0,0,122,0,0,0,190,0,37,0,113,0,251,0,0,0,41,0,0,0,117,0,12,0,0,0,95,0,0,0,69,0,0,0,0,0,126,0,125,0,182,0,184,0,8,0,0,0,230,0,4,0,64,0,237,0,246,0,0,0,133,0,224,0,23,0,136,0,211,0,0,0,141,0,30,0,211,0,196,0,175,0,225,0,195,0,0,0,95,0,99,0,138,0,31,0,0,0,212,0,89,0,147,0,3,0,128,0,0,0,0,0,0,0,134,0,124,0,116,0,27,0,11,0,251,0,0,0,117,0,253,0,17,0,158,0,18,0,68,0,0,0,162,0,22,0,111,0,173,0,207,0,118,0,189,0,168,0,27,0,88,0,35,0,148,0,0,0,36,0,62,0,136,0,235,0,143,0,238,0,0,0,120,0,0,0,238,0,0,0,54,0,133,0,177,0,0,0,77,0,149,0,95,0,167,0,188,0,7,0,245,0,61,0,186,0,145,0,57,0,175,0,21,0,169,0,166,0,236,0,71,0,96,0,246,0,109,0,116,0,0,0,138,0,136,0,0,0,78,0,124,0,193,0,9,0,199,0,0,0,58,0,68,0,25,0,194,0,175,0,250,0,202,0,129,0,91,0,173,0,79,0,35,0,191,0,116,0,83,0,0,0,44,0,113,0,191,0,22,0,106,0,157,0,82,0,0,0,0,0,92,0,0,0,170,0,118,0,45,0,196,0,254,0,0,0,0,0,215,0,38,0,110,0,0,0,248,0,38,0,136,0,146,0,0,0,113,0,65,0,0,0,188,0,0,0,248,0,21,0,168,0,214,0,91,0,114,0,48,0,0,0,99,0,0,0,226,0,0,0,148,0,0,0,76,0,155,0,61,0,157,0,254,0,252,0,73,0,91,0,124,0,108,0,25,0,8,0,115,0,0,0,0,0,157,0,167,0,195,0,130,0,145,0,193,0,180,0,0,0,200,0,98,0,42,0,0,0,176,0,219,0,26,0,5,0,127,0,96,0,75,0,72,0,188,0,129,0,134,0,12,0,107,0,0,0,0,0,112,0,125,0,208,0,45,0,14,0,248,0,8,0,236,0,228,0,0,0,0,0,0,0,0,0,146,0,143,0,177,0,24,0,203,0,0,0,0,0,99,0,66,0,81,0,41,0,0,0,18,0,207,0,235,0,40,0,0,0,31,0,0,0,110,0,167,0,156,0,174,0,9,0,0,0,56,0,183,0,34,0,97,0,156,0,95,0,0,0,115,0,40,0,251,0,0,0,129,0,127,0,9,0,208,0,178,0,0,0,250,0,240,0,139,0,228,0,92,0,70,0,175,0,124,0,170,0,194,0,128,0,79,0,232,0,242,0,190,0,102,0,100,0,22,0,148,0,201,0,0,0,223,0,25,0,0,0,249,0,0,0,209,0,104,0,0,0,0,0,90,0,62,0,15,0,236,0,48,0,247,0,171,0,16,0,0,0,211,0,24,0,138,0,209,0,252,0,203,0,58,0,149,0,85,0,48,0,177,0,66,0,0,0,0,0,20,0,129,0,179,0,217,0,84,0,123,0,122,0,56,0);
signal scenario_full  : scenario_type := (174,31,174,30,127,31,135,31,179,31,179,30,95,31,132,31,4,31,174,31,52,31,122,31,122,30,44,31,44,30,194,31,199,31,129,31,228,31,228,30,79,31,172,31,193,31,193,30,86,31,91,31,166,31,233,31,233,30,218,31,101,31,101,30,87,31,217,31,217,30,101,31,101,30,248,31,158,31,121,31,160,31,160,30,223,31,139,31,50,31,20,31,53,31,115,31,241,31,107,31,107,30,107,29,230,31,153,31,153,30,4,31,120,31,176,31,15,31,15,30,41,31,147,31,147,30,214,31,250,31,32,31,64,31,64,30,68,31,19,31,73,31,73,30,190,31,35,31,128,31,141,31,103,31,28,31,162,31,93,31,10,31,159,31,25,31,68,31,109,31,222,31,78,31,16,31,59,31,59,30,59,29,39,31,39,30,65,31,193,31,193,31,84,31,37,31,153,31,76,31,214,31,214,30,50,31,50,30,50,29,176,31,82,31,175,31,4,31,13,31,239,31,42,31,86,31,213,31,103,31,103,30,103,29,170,31,133,31,224,31,224,30,224,29,235,31,235,30,3,31,118,31,73,31,185,31,192,31,25,31,226,31,237,31,27,31,190,31,50,31,50,30,149,31,155,31,155,31,69,31,130,31,52,31,211,31,15,31,164,31,96,31,204,31,35,31,49,31,174,31,32,31,167,31,89,31,222,31,211,31,232,31,190,31,63,31,189,31,69,31,220,31,54,31,167,31,198,31,254,31,117,31,147,31,147,30,23,31,149,31,130,31,180,31,39,31,196,31,174,31,1,31,114,31,188,31,188,30,162,31,162,30,75,31,174,31,174,30,215,31,115,31,191,31,191,30,159,31,114,31,232,31,247,31,247,30,247,29,182,31,201,31,163,31,196,31,46,31,46,30,165,31,146,31,157,31,48,31,119,31,198,31,198,30,52,31,99,31,126,31,38,31,255,31,59,31,55,31,72,31,234,31,115,31,255,31,21,31,73,31,225,31,157,31,93,31,39,31,227,31,78,31,199,31,253,31,209,31,209,30,51,31,51,30,124,31,77,31,123,31,123,30,76,31,150,31,150,30,194,31,60,31,110,31,110,30,147,31,147,30,70,31,70,30,44,31,182,31,175,31,197,31,228,31,214,31,69,31,206,31,42,31,204,31,209,31,116,31,190,31,25,31,161,31,67,31,67,30,155,31,209,31,209,30,224,31,65,31,65,30,217,31,206,31,13,31,112,31,155,31,87,31,87,30,87,29,20,31,20,30,120,31,210,31,251,31,173,31,168,31,4,31,4,30,4,29,122,31,122,30,190,31,37,31,113,31,251,31,251,30,41,31,41,30,117,31,12,31,12,30,95,31,95,30,69,31,69,30,69,29,126,31,125,31,182,31,184,31,8,31,8,30,230,31,4,31,64,31,237,31,246,31,246,30,133,31,224,31,23,31,136,31,211,31,211,30,141,31,30,31,211,31,196,31,175,31,225,31,195,31,195,30,95,31,99,31,138,31,31,31,31,30,212,31,89,31,147,31,3,31,128,31,128,30,128,29,128,28,134,31,124,31,116,31,27,31,11,31,251,31,251,30,117,31,253,31,17,31,158,31,18,31,68,31,68,30,162,31,22,31,111,31,173,31,207,31,118,31,189,31,168,31,27,31,88,31,35,31,148,31,148,30,36,31,62,31,136,31,235,31,143,31,238,31,238,30,120,31,120,30,238,31,238,30,54,31,133,31,177,31,177,30,77,31,149,31,95,31,167,31,188,31,7,31,245,31,61,31,186,31,145,31,57,31,175,31,21,31,169,31,166,31,236,31,71,31,96,31,246,31,109,31,116,31,116,30,138,31,136,31,136,30,78,31,124,31,193,31,9,31,199,31,199,30,58,31,68,31,25,31,194,31,175,31,250,31,202,31,129,31,91,31,173,31,79,31,35,31,191,31,116,31,83,31,83,30,44,31,113,31,191,31,22,31,106,31,157,31,82,31,82,30,82,29,92,31,92,30,170,31,118,31,45,31,196,31,254,31,254,30,254,29,215,31,38,31,110,31,110,30,248,31,38,31,136,31,146,31,146,30,113,31,65,31,65,30,188,31,188,30,248,31,21,31,168,31,214,31,91,31,114,31,48,31,48,30,99,31,99,30,226,31,226,30,148,31,148,30,76,31,155,31,61,31,157,31,254,31,252,31,73,31,91,31,124,31,108,31,25,31,8,31,115,31,115,30,115,29,157,31,167,31,195,31,130,31,145,31,193,31,180,31,180,30,200,31,98,31,42,31,42,30,176,31,219,31,26,31,5,31,127,31,96,31,75,31,72,31,188,31,129,31,134,31,12,31,107,31,107,30,107,29,112,31,125,31,208,31,45,31,14,31,248,31,8,31,236,31,228,31,228,30,228,29,228,28,228,27,146,31,143,31,177,31,24,31,203,31,203,30,203,29,99,31,66,31,81,31,41,31,41,30,18,31,207,31,235,31,40,31,40,30,31,31,31,30,110,31,167,31,156,31,174,31,9,31,9,30,56,31,183,31,34,31,97,31,156,31,95,31,95,30,115,31,40,31,251,31,251,30,129,31,127,31,9,31,208,31,178,31,178,30,250,31,240,31,139,31,228,31,92,31,70,31,175,31,124,31,170,31,194,31,128,31,79,31,232,31,242,31,190,31,102,31,100,31,22,31,148,31,201,31,201,30,223,31,25,31,25,30,249,31,249,30,209,31,104,31,104,30,104,29,90,31,62,31,15,31,236,31,48,31,247,31,171,31,16,31,16,30,211,31,24,31,138,31,209,31,252,31,203,31,58,31,149,31,85,31,48,31,177,31,66,31,66,30,66,29,20,31,129,31,179,31,217,31,84,31,123,31,122,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
