-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 885;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,129,0,249,0,120,0,19,0,70,0,176,0,241,0,176,0,252,0,87,0,0,0,144,0,42,0,145,0,57,0,61,0,201,0,43,0,220,0,238,0,159,0,43,0,143,0,0,0,229,0,116,0,0,0,182,0,120,0,26,0,182,0,0,0,101,0,109,0,148,0,181,0,34,0,0,0,38,0,133,0,226,0,163,0,0,0,184,0,87,0,249,0,58,0,144,0,0,0,0,0,0,0,0,0,145,0,218,0,0,0,48,0,84,0,0,0,0,0,102,0,144,0,0,0,120,0,244,0,0,0,3,0,120,0,77,0,77,0,191,0,138,0,0,0,81,0,0,0,196,0,0,0,0,0,108,0,0,0,0,0,0,0,0,0,81,0,0,0,7,0,0,0,45,0,225,0,70,0,218,0,0,0,159,0,106,0,0,0,46,0,220,0,103,0,118,0,105,0,15,0,233,0,55,0,140,0,162,0,34,0,0,0,0,0,0,0,148,0,123,0,61,0,115,0,99,0,197,0,183,0,0,0,104,0,8,0,0,0,20,0,196,0,0,0,119,0,3,0,127,0,0,0,20,0,0,0,243,0,0,0,132,0,220,0,228,0,14,0,186,0,83,0,178,0,140,0,0,0,193,0,137,0,8,0,21,0,157,0,180,0,243,0,16,0,0,0,160,0,0,0,97,0,166,0,0,0,0,0,254,0,166,0,0,0,56,0,72,0,23,0,83,0,29,0,136,0,109,0,144,0,116,0,195,0,111,0,229,0,8,0,90,0,44,0,121,0,205,0,0,0,75,0,0,0,153,0,0,0,78,0,92,0,231,0,81,0,66,0,180,0,38,0,92,0,208,0,74,0,102,0,96,0,195,0,0,0,238,0,0,0,15,0,188,0,0,0,116,0,21,0,241,0,114,0,0,0,95,0,0,0,0,0,5,0,61,0,148,0,0,0,160,0,91,0,88,0,155,0,175,0,37,0,0,0,85,0,14,0,100,0,0,0,12,0,10,0,75,0,112,0,17,0,67,0,124,0,32,0,134,0,8,0,111,0,77,0,0,0,62,0,170,0,125,0,0,0,125,0,161,0,196,0,57,0,116,0,110,0,4,0,0,0,128,0,108,0,125,0,113,0,221,0,57,0,166,0,253,0,0,0,19,0,75,0,2,0,36,0,231,0,0,0,76,0,242,0,169,0,205,0,255,0,77,0,206,0,98,0,0,0,201,0,165,0,147,0,188,0,60,0,0,0,229,0,0,0,8,0,116,0,22,0,99,0,243,0,216,0,0,0,131,0,243,0,242,0,245,0,197,0,32,0,34,0,22,0,235,0,235,0,0,0,149,0,161,0,247,0,1,0,50,0,171,0,0,0,0,0,149,0,239,0,0,0,21,0,169,0,0,0,229,0,129,0,0,0,0,0,105,0,97,0,0,0,154,0,189,0,136,0,94,0,156,0,0,0,202,0,0,0,181,0,0,0,0,0,219,0,21,0,39,0,9,0,96,0,16,0,74,0,122,0,120,0,0,0,39,0,235,0,132,0,119,0,141,0,203,0,228,0,173,0,231,0,44,0,0,0,0,0,253,0,0,0,207,0,230,0,0,0,145,0,250,0,0,0,150,0,176,0,220,0,0,0,112,0,145,0,72,0,157,0,150,0,218,0,52,0,158,0,108,0,54,0,0,0,98,0,0,0,103,0,179,0,231,0,117,0,227,0,34,0,150,0,41,0,144,0,144,0,0,0,151,0,5,0,0,0,92,0,163,0,161,0,204,0,45,0,236,0,106,0,0,0,81,0,243,0,12,0,190,0,231,0,62,0,0,0,174,0,226,0,15,0,138,0,218,0,236,0,26,0,179,0,162,0,168,0,26,0,71,0,0,0,191,0,0,0,33,0,123,0,117,0,88,0,249,0,0,0,0,0,0,0,86,0,13,0,218,0,0,0,233,0,94,0,77,0,63,0,64,0,0,0,215,0,249,0,21,0,98,0,182,0,0,0,0,0,0,0,156,0,160,0,84,0,0,0,160,0,228,0,0,0,0,0,12,0,0,0,251,0,185,0,0,0,46,0,82,0,0,0,235,0,152,0,122,0,0,0,179,0,19,0,232,0,0,0,72,0,151,0,48,0,142,0,64,0,88,0,116,0,194,0,130,0,199,0,104,0,115,0,142,0,19,0,223,0,50,0,56,0,0,0,169,0,183,0,0,0,0,0,80,0,21,0,117,0,105,0,122,0,0,0,123,0,61,0,105,0,214,0,87,0,196,0,45,0,67,0,97,0,0,0,180,0,214,0,96,0,205,0,97,0,248,0,136,0,130,0,162,0,204,0,115,0,0,0,121,0,0,0,239,0,0,0,11,0,202,0,246,0,0,0,153,0,56,0,113,0,229,0,189,0,109,0,121,0,0,0,163,0,0,0,0,0,164,0,212,0,101,0,64,0,83,0,73,0,170,0,113,0,122,0,83,0,96,0,148,0,0,0,209,0,146,0,126,0,195,0,155,0,167,0,167,0,204,0,0,0,179,0,207,0,60,0,187,0,0,0,188,0,210,0,42,0,72,0,85,0,133,0,0,0,94,0,135,0,98,0,120,0,141,0,233,0,246,0,0,0,0,0,0,0,21,0,0,0,96,0,61,0,41,0,0,0,186,0,207,0,230,0,118,0,71,0,47,0,236,0,94,0,93,0,157,0,199,0,194,0,225,0,125,0,0,0,82,0,0,0,5,0,165,0,90,0,0,0,229,0,112,0,88,0,135,0,255,0,173,0,2,0,83,0,174,0,92,0,0,0,217,0,132,0,37,0,246,0,106,0,165,0,210,0,76,0,42,0,57,0,124,0,144,0,128,0,51,0,112,0,184,0,220,0,188,0,114,0,16,0,0,0,0,0,55,0,250,0,172,0,0,0,152,0,0,0,60,0,92,0,233,0,48,0,138,0,182,0,228,0,237,0,52,0,146,0,83,0,0,0,169,0,122,0,210,0,42,0,48,0,175,0,121,0,39,0,233,0,124,0,163,0,150,0,83,0,0,0,0,0,4,0,231,0,0,0,145,0,0,0,195,0,0,0,0,0,64,0,5,0,0,0,184,0,0,0,36,0,200,0,0,0,171,0,240,0,0,0,200,0,112,0,61,0,250,0,227,0,175,0,0,0,0,0,69,0,152,0,42,0,51,0,89,0,0,0,0,0,0,0,146,0,19,0,191,0,119,0,139,0,194,0,83,0,94,0,53,0,163,0,248,0,214,0,0,0,142,0,30,0,3,0,40,0,223,0,202,0,0,0,36,0,106,0,60,0,37,0,46,0,57,0,236,0,0,0,246,0,0,0,211,0,75,0,92,0,222,0,68,0,110,0,158,0,0,0,108,0,17,0,193,0,247,0,80,0,234,0,171,0,243,0,0,0,126,0,120,0,17,0,57,0,98,0,48,0,198,0,95,0,173,0,173,0,109,0,206,0,0,0,121,0,0,0,86,0,92,0,159,0,0,0,196,0,137,0,34,0,164,0,15,0,238,0,124,0,0,0,41,0,48,0,219,0,133,0,105,0,166,0,171,0,180,0,54,0,20,0,60,0,196,0,168,0,161,0,225,0,239,0,185,0,109,0,109,0,0,0,70,0,194,0,56,0,10,0,90,0,103,0,99,0,147,0,88,0,119,0,160,0,0,0,0,0,34,0,118,0,216,0,78,0,166,0,0,0,56,0,0,0,0,0,0,0,59,0,112,0,0,0,0,0,61,0,100,0,130,0,0,0,149,0,132,0,223,0,64,0,133,0,44,0,0,0,137,0,226,0,100,0,57,0,95,0,0,0,247,0,183,0,243,0,91,0,124,0,73,0,0,0,189,0,0,0,160,0,212,0,211,0,183,0,5,0,0,0,189,0,28,0,138,0,69,0,246,0,24,0,21,0,0,0,28,0,13,0,219,0,187,0,29,0,6,0,227,0,0,0,65,0,18,0,117,0,51,0,0,0);
signal scenario_full  : scenario_type := (0,0,129,31,249,31,120,31,19,31,70,31,176,31,241,31,176,31,252,31,87,31,87,30,144,31,42,31,145,31,57,31,61,31,201,31,43,31,220,31,238,31,159,31,43,31,143,31,143,30,229,31,116,31,116,30,182,31,120,31,26,31,182,31,182,30,101,31,109,31,148,31,181,31,34,31,34,30,38,31,133,31,226,31,163,31,163,30,184,31,87,31,249,31,58,31,144,31,144,30,144,29,144,28,144,27,145,31,218,31,218,30,48,31,84,31,84,30,84,29,102,31,144,31,144,30,120,31,244,31,244,30,3,31,120,31,77,31,77,31,191,31,138,31,138,30,81,31,81,30,196,31,196,30,196,29,108,31,108,30,108,29,108,28,108,27,81,31,81,30,7,31,7,30,45,31,225,31,70,31,218,31,218,30,159,31,106,31,106,30,46,31,220,31,103,31,118,31,105,31,15,31,233,31,55,31,140,31,162,31,34,31,34,30,34,29,34,28,148,31,123,31,61,31,115,31,99,31,197,31,183,31,183,30,104,31,8,31,8,30,20,31,196,31,196,30,119,31,3,31,127,31,127,30,20,31,20,30,243,31,243,30,132,31,220,31,228,31,14,31,186,31,83,31,178,31,140,31,140,30,193,31,137,31,8,31,21,31,157,31,180,31,243,31,16,31,16,30,160,31,160,30,97,31,166,31,166,30,166,29,254,31,166,31,166,30,56,31,72,31,23,31,83,31,29,31,136,31,109,31,144,31,116,31,195,31,111,31,229,31,8,31,90,31,44,31,121,31,205,31,205,30,75,31,75,30,153,31,153,30,78,31,92,31,231,31,81,31,66,31,180,31,38,31,92,31,208,31,74,31,102,31,96,31,195,31,195,30,238,31,238,30,15,31,188,31,188,30,116,31,21,31,241,31,114,31,114,30,95,31,95,30,95,29,5,31,61,31,148,31,148,30,160,31,91,31,88,31,155,31,175,31,37,31,37,30,85,31,14,31,100,31,100,30,12,31,10,31,75,31,112,31,17,31,67,31,124,31,32,31,134,31,8,31,111,31,77,31,77,30,62,31,170,31,125,31,125,30,125,31,161,31,196,31,57,31,116,31,110,31,4,31,4,30,128,31,108,31,125,31,113,31,221,31,57,31,166,31,253,31,253,30,19,31,75,31,2,31,36,31,231,31,231,30,76,31,242,31,169,31,205,31,255,31,77,31,206,31,98,31,98,30,201,31,165,31,147,31,188,31,60,31,60,30,229,31,229,30,8,31,116,31,22,31,99,31,243,31,216,31,216,30,131,31,243,31,242,31,245,31,197,31,32,31,34,31,22,31,235,31,235,31,235,30,149,31,161,31,247,31,1,31,50,31,171,31,171,30,171,29,149,31,239,31,239,30,21,31,169,31,169,30,229,31,129,31,129,30,129,29,105,31,97,31,97,30,154,31,189,31,136,31,94,31,156,31,156,30,202,31,202,30,181,31,181,30,181,29,219,31,21,31,39,31,9,31,96,31,16,31,74,31,122,31,120,31,120,30,39,31,235,31,132,31,119,31,141,31,203,31,228,31,173,31,231,31,44,31,44,30,44,29,253,31,253,30,207,31,230,31,230,30,145,31,250,31,250,30,150,31,176,31,220,31,220,30,112,31,145,31,72,31,157,31,150,31,218,31,52,31,158,31,108,31,54,31,54,30,98,31,98,30,103,31,179,31,231,31,117,31,227,31,34,31,150,31,41,31,144,31,144,31,144,30,151,31,5,31,5,30,92,31,163,31,161,31,204,31,45,31,236,31,106,31,106,30,81,31,243,31,12,31,190,31,231,31,62,31,62,30,174,31,226,31,15,31,138,31,218,31,236,31,26,31,179,31,162,31,168,31,26,31,71,31,71,30,191,31,191,30,33,31,123,31,117,31,88,31,249,31,249,30,249,29,249,28,86,31,13,31,218,31,218,30,233,31,94,31,77,31,63,31,64,31,64,30,215,31,249,31,21,31,98,31,182,31,182,30,182,29,182,28,156,31,160,31,84,31,84,30,160,31,228,31,228,30,228,29,12,31,12,30,251,31,185,31,185,30,46,31,82,31,82,30,235,31,152,31,122,31,122,30,179,31,19,31,232,31,232,30,72,31,151,31,48,31,142,31,64,31,88,31,116,31,194,31,130,31,199,31,104,31,115,31,142,31,19,31,223,31,50,31,56,31,56,30,169,31,183,31,183,30,183,29,80,31,21,31,117,31,105,31,122,31,122,30,123,31,61,31,105,31,214,31,87,31,196,31,45,31,67,31,97,31,97,30,180,31,214,31,96,31,205,31,97,31,248,31,136,31,130,31,162,31,204,31,115,31,115,30,121,31,121,30,239,31,239,30,11,31,202,31,246,31,246,30,153,31,56,31,113,31,229,31,189,31,109,31,121,31,121,30,163,31,163,30,163,29,164,31,212,31,101,31,64,31,83,31,73,31,170,31,113,31,122,31,83,31,96,31,148,31,148,30,209,31,146,31,126,31,195,31,155,31,167,31,167,31,204,31,204,30,179,31,207,31,60,31,187,31,187,30,188,31,210,31,42,31,72,31,85,31,133,31,133,30,94,31,135,31,98,31,120,31,141,31,233,31,246,31,246,30,246,29,246,28,21,31,21,30,96,31,61,31,41,31,41,30,186,31,207,31,230,31,118,31,71,31,47,31,236,31,94,31,93,31,157,31,199,31,194,31,225,31,125,31,125,30,82,31,82,30,5,31,165,31,90,31,90,30,229,31,112,31,88,31,135,31,255,31,173,31,2,31,83,31,174,31,92,31,92,30,217,31,132,31,37,31,246,31,106,31,165,31,210,31,76,31,42,31,57,31,124,31,144,31,128,31,51,31,112,31,184,31,220,31,188,31,114,31,16,31,16,30,16,29,55,31,250,31,172,31,172,30,152,31,152,30,60,31,92,31,233,31,48,31,138,31,182,31,228,31,237,31,52,31,146,31,83,31,83,30,169,31,122,31,210,31,42,31,48,31,175,31,121,31,39,31,233,31,124,31,163,31,150,31,83,31,83,30,83,29,4,31,231,31,231,30,145,31,145,30,195,31,195,30,195,29,64,31,5,31,5,30,184,31,184,30,36,31,200,31,200,30,171,31,240,31,240,30,200,31,112,31,61,31,250,31,227,31,175,31,175,30,175,29,69,31,152,31,42,31,51,31,89,31,89,30,89,29,89,28,146,31,19,31,191,31,119,31,139,31,194,31,83,31,94,31,53,31,163,31,248,31,214,31,214,30,142,31,30,31,3,31,40,31,223,31,202,31,202,30,36,31,106,31,60,31,37,31,46,31,57,31,236,31,236,30,246,31,246,30,211,31,75,31,92,31,222,31,68,31,110,31,158,31,158,30,108,31,17,31,193,31,247,31,80,31,234,31,171,31,243,31,243,30,126,31,120,31,17,31,57,31,98,31,48,31,198,31,95,31,173,31,173,31,109,31,206,31,206,30,121,31,121,30,86,31,92,31,159,31,159,30,196,31,137,31,34,31,164,31,15,31,238,31,124,31,124,30,41,31,48,31,219,31,133,31,105,31,166,31,171,31,180,31,54,31,20,31,60,31,196,31,168,31,161,31,225,31,239,31,185,31,109,31,109,31,109,30,70,31,194,31,56,31,10,31,90,31,103,31,99,31,147,31,88,31,119,31,160,31,160,30,160,29,34,31,118,31,216,31,78,31,166,31,166,30,56,31,56,30,56,29,56,28,59,31,112,31,112,30,112,29,61,31,100,31,130,31,130,30,149,31,132,31,223,31,64,31,133,31,44,31,44,30,137,31,226,31,100,31,57,31,95,31,95,30,247,31,183,31,243,31,91,31,124,31,73,31,73,30,189,31,189,30,160,31,212,31,211,31,183,31,5,31,5,30,189,31,28,31,138,31,69,31,246,31,24,31,21,31,21,30,28,31,13,31,219,31,187,31,29,31,6,31,227,31,227,30,65,31,18,31,117,31,51,31,51,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
