-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_136 is
end project_tb_136;

architecture project_tb_arch_136 of project_tb_136 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 763;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,19,0,169,0,124,0,0,0,212,0,0,0,2,0,144,0,17,0,191,0,35,0,0,0,24,0,33,0,31,0,0,0,230,0,7,0,0,0,161,0,8,0,137,0,17,0,195,0,0,0,131,0,185,0,0,0,82,0,140,0,173,0,20,0,252,0,166,0,91,0,118,0,63,0,108,0,92,0,81,0,109,0,229,0,28,0,198,0,186,0,233,0,220,0,27,0,139,0,139,0,254,0,74,0,36,0,55,0,0,0,87,0,32,0,128,0,194,0,0,0,198,0,36,0,0,0,93,0,161,0,3,0,0,0,110,0,0,0,123,0,0,0,66,0,170,0,119,0,0,0,143,0,69,0,231,0,0,0,146,0,209,0,186,0,166,0,92,0,0,0,137,0,0,0,0,0,150,0,228,0,208,0,230,0,147,0,242,0,223,0,17,0,177,0,194,0,206,0,31,0,181,0,157,0,103,0,81,0,174,0,0,0,9,0,17,0,153,0,113,0,60,0,241,0,0,0,0,0,34,0,241,0,178,0,0,0,0,0,243,0,242,0,79,0,0,0,0,0,230,0,0,0,252,0,54,0,32,0,0,0,155,0,0,0,61,0,0,0,17,0,118,0,211,0,191,0,75,0,0,0,0,0,63,0,0,0,0,0,0,0,119,0,0,0,19,0,47,0,136,0,91,0,0,0,126,0,0,0,183,0,2,0,163,0,160,0,175,0,239,0,187,0,0,0,43,0,186,0,30,0,49,0,0,0,0,0,14,0,198,0,174,0,116,0,0,0,129,0,0,0,0,0,111,0,0,0,110,0,172,0,0,0,202,0,0,0,88,0,176,0,116,0,0,0,99,0,241,0,0,0,0,0,0,0,74,0,95,0,223,0,218,0,123,0,0,0,14,0,136,0,71,0,197,0,0,0,55,0,131,0,245,0,135,0,92,0,22,0,154,0,0,0,238,0,160,0,31,0,196,0,147,0,138,0,64,0,0,0,0,0,225,0,197,0,101,0,193,0,220,0,93,0,127,0,215,0,172,0,246,0,6,0,38,0,56,0,35,0,150,0,152,0,53,0,0,0,0,0,0,0,205,0,219,0,212,0,173,0,61,0,215,0,141,0,198,0,46,0,184,0,161,0,109,0,0,0,62,0,23,0,0,0,0,0,1,0,0,0,201,0,121,0,165,0,186,0,234,0,80,0,253,0,177,0,100,0,1,0,68,0,36,0,195,0,197,0,110,0,37,0,116,0,116,0,65,0,192,0,100,0,0,0,45,0,0,0,80,0,149,0,195,0,0,0,181,0,126,0,7,0,172,0,252,0,26,0,32,0,204,0,89,0,174,0,0,0,184,0,0,0,65,0,181,0,72,0,242,0,72,0,0,0,250,0,17,0,19,0,164,0,250,0,28,0,4,0,193,0,208,0,176,0,75,0,38,0,21,0,3,0,28,0,177,0,108,0,244,0,196,0,51,0,184,0,124,0,198,0,184,0,0,0,37,0,147,0,141,0,80,0,223,0,227,0,188,0,156,0,154,0,66,0,184,0,125,0,6,0,84,0,0,0,113,0,250,0,95,0,46,0,116,0,255,0,61,0,53,0,150,0,188,0,223,0,37,0,238,0,205,0,9,0,232,0,83,0,202,0,0,0,0,0,27,0,86,0,135,0,196,0,113,0,165,0,0,0,23,0,0,0,113,0,0,0,107,0,0,0,0,0,0,0,126,0,191,0,156,0,157,0,0,0,0,0,9,0,222,0,176,0,66,0,220,0,237,0,0,0,0,0,239,0,123,0,0,0,0,0,81,0,112,0,69,0,0,0,38,0,161,0,75,0,55,0,98,0,0,0,69,0,5,0,37,0,0,0,85,0,136,0,58,0,132,0,182,0,35,0,0,0,220,0,0,0,0,0,140,0,63,0,226,0,147,0,0,0,140,0,91,0,163,0,0,0,100,0,60,0,0,0,119,0,189,0,131,0,165,0,0,0,0,0,0,0,0,0,37,0,254,0,222,0,120,0,0,0,214,0,184,0,200,0,120,0,0,0,0,0,53,0,160,0,0,0,16,0,55,0,0,0,104,0,0,0,163,0,122,0,0,0,159,0,199,0,169,0,194,0,0,0,18,0,0,0,211,0,123,0,109,0,125,0,118,0,102,0,0,0,40,0,29,0,139,0,0,0,60,0,161,0,0,0,197,0,134,0,242,0,35,0,129,0,75,0,73,0,236,0,229,0,143,0,9,0,0,0,173,0,30,0,46,0,7,0,204,0,0,0,0,0,127,0,178,0,240,0,18,0,251,0,71,0,131,0,0,0,57,0,225,0,0,0,66,0,27,0,251,0,171,0,249,0,0,0,0,0,188,0,207,0,73,0,128,0,253,0,0,0,49,0,107,0,132,0,231,0,207,0,40,0,59,0,213,0,121,0,179,0,238,0,0,0,0,0,88,0,103,0,13,0,86,0,185,0,198,0,0,0,105,0,200,0,22,0,115,0,125,0,0,0,25,0,183,0,179,0,0,0,0,0,148,0,101,0,0,0,98,0,100,0,0,0,51,0,0,0,0,0,233,0,11,0,0,0,80,0,241,0,0,0,241,0,211,0,156,0,0,0,147,0,156,0,0,0,188,0,244,0,0,0,92,0,135,0,141,0,141,0,244,0,164,0,0,0,60,0,135,0,249,0,41,0,212,0,169,0,218,0,232,0,243,0,204,0,0,0,115,0,176,0,144,0,222,0,23,0,0,0,21,0,188,0,47,0,35,0,0,0,7,0,36,0,37,0,231,0,70,0,40,0,136,0,0,0,195,0,50,0,13,0,174,0,190,0,0,0,94,0,103,0,100,0,51,0,130,0,184,0,36,0,1,0,149,0,0,0,180,0,0,0,160,0,241,0,29,0,164,0,0,0,45,0,178,0,232,0,0,0,138,0,181,0,99,0,105,0,90,0,177,0,187,0,49,0,166,0,145,0,77,0,18,0,153,0,78,0,20,0,232,0,170,0,59,0,128,0,0,0,160,0,230,0,171,0,152,0,0,0,0,0,22,0,204,0,239,0,0,0,86,0,236,0,236,0,0,0,100,0,162,0,192,0,109,0,0,0,0,0,0,0,58,0,0,0,94,0,12,0,133,0,240,0,233,0,148,0,45,0,0,0,249,0,57,0,118,0,137,0,245,0,133,0,0,0,12,0,0,0,196,0,16,0,111,0,191,0,195,0,0,0,249,0,12,0,183,0,0,0,252,0,169,0,173,0,1,0,155,0,240,0,52,0,90,0,75,0,220,0,191,0,80,0,188,0,229,0,0,0,52,0,80,0,40,0,37,0,0,0,65,0,102,0,68,0,187,0,112,0,68,0,244,0,131,0,34,0,36,0,0,0,25,0,0,0,0,0,0,0,222,0,0,0,168,0,0,0,67,0,172,0,116,0,45,0);
signal scenario_full  : scenario_type := (0,0,19,31,169,31,124,31,124,30,212,31,212,30,2,31,144,31,17,31,191,31,35,31,35,30,24,31,33,31,31,31,31,30,230,31,7,31,7,30,161,31,8,31,137,31,17,31,195,31,195,30,131,31,185,31,185,30,82,31,140,31,173,31,20,31,252,31,166,31,91,31,118,31,63,31,108,31,92,31,81,31,109,31,229,31,28,31,198,31,186,31,233,31,220,31,27,31,139,31,139,31,254,31,74,31,36,31,55,31,55,30,87,31,32,31,128,31,194,31,194,30,198,31,36,31,36,30,93,31,161,31,3,31,3,30,110,31,110,30,123,31,123,30,66,31,170,31,119,31,119,30,143,31,69,31,231,31,231,30,146,31,209,31,186,31,166,31,92,31,92,30,137,31,137,30,137,29,150,31,228,31,208,31,230,31,147,31,242,31,223,31,17,31,177,31,194,31,206,31,31,31,181,31,157,31,103,31,81,31,174,31,174,30,9,31,17,31,153,31,113,31,60,31,241,31,241,30,241,29,34,31,241,31,178,31,178,30,178,29,243,31,242,31,79,31,79,30,79,29,230,31,230,30,252,31,54,31,32,31,32,30,155,31,155,30,61,31,61,30,17,31,118,31,211,31,191,31,75,31,75,30,75,29,63,31,63,30,63,29,63,28,119,31,119,30,19,31,47,31,136,31,91,31,91,30,126,31,126,30,183,31,2,31,163,31,160,31,175,31,239,31,187,31,187,30,43,31,186,31,30,31,49,31,49,30,49,29,14,31,198,31,174,31,116,31,116,30,129,31,129,30,129,29,111,31,111,30,110,31,172,31,172,30,202,31,202,30,88,31,176,31,116,31,116,30,99,31,241,31,241,30,241,29,241,28,74,31,95,31,223,31,218,31,123,31,123,30,14,31,136,31,71,31,197,31,197,30,55,31,131,31,245,31,135,31,92,31,22,31,154,31,154,30,238,31,160,31,31,31,196,31,147,31,138,31,64,31,64,30,64,29,225,31,197,31,101,31,193,31,220,31,93,31,127,31,215,31,172,31,246,31,6,31,38,31,56,31,35,31,150,31,152,31,53,31,53,30,53,29,53,28,205,31,219,31,212,31,173,31,61,31,215,31,141,31,198,31,46,31,184,31,161,31,109,31,109,30,62,31,23,31,23,30,23,29,1,31,1,30,201,31,121,31,165,31,186,31,234,31,80,31,253,31,177,31,100,31,1,31,68,31,36,31,195,31,197,31,110,31,37,31,116,31,116,31,65,31,192,31,100,31,100,30,45,31,45,30,80,31,149,31,195,31,195,30,181,31,126,31,7,31,172,31,252,31,26,31,32,31,204,31,89,31,174,31,174,30,184,31,184,30,65,31,181,31,72,31,242,31,72,31,72,30,250,31,17,31,19,31,164,31,250,31,28,31,4,31,193,31,208,31,176,31,75,31,38,31,21,31,3,31,28,31,177,31,108,31,244,31,196,31,51,31,184,31,124,31,198,31,184,31,184,30,37,31,147,31,141,31,80,31,223,31,227,31,188,31,156,31,154,31,66,31,184,31,125,31,6,31,84,31,84,30,113,31,250,31,95,31,46,31,116,31,255,31,61,31,53,31,150,31,188,31,223,31,37,31,238,31,205,31,9,31,232,31,83,31,202,31,202,30,202,29,27,31,86,31,135,31,196,31,113,31,165,31,165,30,23,31,23,30,113,31,113,30,107,31,107,30,107,29,107,28,126,31,191,31,156,31,157,31,157,30,157,29,9,31,222,31,176,31,66,31,220,31,237,31,237,30,237,29,239,31,123,31,123,30,123,29,81,31,112,31,69,31,69,30,38,31,161,31,75,31,55,31,98,31,98,30,69,31,5,31,37,31,37,30,85,31,136,31,58,31,132,31,182,31,35,31,35,30,220,31,220,30,220,29,140,31,63,31,226,31,147,31,147,30,140,31,91,31,163,31,163,30,100,31,60,31,60,30,119,31,189,31,131,31,165,31,165,30,165,29,165,28,165,27,37,31,254,31,222,31,120,31,120,30,214,31,184,31,200,31,120,31,120,30,120,29,53,31,160,31,160,30,16,31,55,31,55,30,104,31,104,30,163,31,122,31,122,30,159,31,199,31,169,31,194,31,194,30,18,31,18,30,211,31,123,31,109,31,125,31,118,31,102,31,102,30,40,31,29,31,139,31,139,30,60,31,161,31,161,30,197,31,134,31,242,31,35,31,129,31,75,31,73,31,236,31,229,31,143,31,9,31,9,30,173,31,30,31,46,31,7,31,204,31,204,30,204,29,127,31,178,31,240,31,18,31,251,31,71,31,131,31,131,30,57,31,225,31,225,30,66,31,27,31,251,31,171,31,249,31,249,30,249,29,188,31,207,31,73,31,128,31,253,31,253,30,49,31,107,31,132,31,231,31,207,31,40,31,59,31,213,31,121,31,179,31,238,31,238,30,238,29,88,31,103,31,13,31,86,31,185,31,198,31,198,30,105,31,200,31,22,31,115,31,125,31,125,30,25,31,183,31,179,31,179,30,179,29,148,31,101,31,101,30,98,31,100,31,100,30,51,31,51,30,51,29,233,31,11,31,11,30,80,31,241,31,241,30,241,31,211,31,156,31,156,30,147,31,156,31,156,30,188,31,244,31,244,30,92,31,135,31,141,31,141,31,244,31,164,31,164,30,60,31,135,31,249,31,41,31,212,31,169,31,218,31,232,31,243,31,204,31,204,30,115,31,176,31,144,31,222,31,23,31,23,30,21,31,188,31,47,31,35,31,35,30,7,31,36,31,37,31,231,31,70,31,40,31,136,31,136,30,195,31,50,31,13,31,174,31,190,31,190,30,94,31,103,31,100,31,51,31,130,31,184,31,36,31,1,31,149,31,149,30,180,31,180,30,160,31,241,31,29,31,164,31,164,30,45,31,178,31,232,31,232,30,138,31,181,31,99,31,105,31,90,31,177,31,187,31,49,31,166,31,145,31,77,31,18,31,153,31,78,31,20,31,232,31,170,31,59,31,128,31,128,30,160,31,230,31,171,31,152,31,152,30,152,29,22,31,204,31,239,31,239,30,86,31,236,31,236,31,236,30,100,31,162,31,192,31,109,31,109,30,109,29,109,28,58,31,58,30,94,31,12,31,133,31,240,31,233,31,148,31,45,31,45,30,249,31,57,31,118,31,137,31,245,31,133,31,133,30,12,31,12,30,196,31,16,31,111,31,191,31,195,31,195,30,249,31,12,31,183,31,183,30,252,31,169,31,173,31,1,31,155,31,240,31,52,31,90,31,75,31,220,31,191,31,80,31,188,31,229,31,229,30,52,31,80,31,40,31,37,31,37,30,65,31,102,31,68,31,187,31,112,31,68,31,244,31,131,31,34,31,36,31,36,30,25,31,25,30,25,29,25,28,222,31,222,30,168,31,168,30,67,31,172,31,116,31,45,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
