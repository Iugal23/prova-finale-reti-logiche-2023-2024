-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_974 is
end project_tb_974;

architecture project_tb_arch_974 of project_tb_974 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 845;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (244,0,0,0,0,0,71,0,131,0,86,0,18,0,137,0,207,0,151,0,5,0,172,0,0,0,25,0,64,0,0,0,0,0,0,0,236,0,0,0,56,0,0,0,127,0,244,0,223,0,0,0,181,0,54,0,17,0,145,0,93,0,177,0,246,0,159,0,230,0,0,0,198,0,101,0,187,0,42,0,127,0,0,0,0,0,0,0,27,0,0,0,168,0,58,0,144,0,116,0,253,0,44,0,61,0,47,0,2,0,239,0,0,0,40,0,227,0,0,0,30,0,91,0,253,0,202,0,105,0,0,0,106,0,0,0,34,0,114,0,0,0,0,0,149,0,97,0,125,0,138,0,215,0,174,0,26,0,131,0,57,0,25,0,115,0,170,0,183,0,0,0,100,0,112,0,0,0,162,0,68,0,14,0,69,0,225,0,195,0,0,0,248,0,48,0,254,0,0,0,0,0,175,0,151,0,113,0,212,0,85,0,135,0,105,0,0,0,188,0,143,0,137,0,175,0,0,0,43,0,204,0,186,0,79,0,94,0,187,0,27,0,253,0,181,0,56,0,248,0,190,0,187,0,242,0,159,0,244,0,205,0,0,0,110,0,174,0,125,0,145,0,64,0,0,0,0,0,201,0,153,0,147,0,119,0,162,0,126,0,0,0,236,0,195,0,0,0,195,0,168,0,0,0,0,0,11,0,0,0,97,0,201,0,244,0,0,0,110,0,139,0,7,0,26,0,130,0,117,0,109,0,222,0,18,0,0,0,48,0,117,0,0,0,169,0,238,0,29,0,66,0,0,0,81,0,166,0,74,0,15,0,56,0,0,0,124,0,0,0,135,0,57,0,59,0,56,0,128,0,91,0,12,0,15,0,235,0,222,0,125,0,0,0,0,0,194,0,2,0,29,0,0,0,227,0,0,0,0,0,224,0,215,0,120,0,0,0,123,0,104,0,202,0,194,0,17,0,47,0,82,0,87,0,105,0,115,0,0,0,47,0,197,0,179,0,216,0,216,0,77,0,179,0,96,0,88,0,6,0,11,0,81,0,25,0,217,0,38,0,0,0,90,0,49,0,226,0,166,0,253,0,120,0,0,0,0,0,0,0,0,0,0,0,169,0,135,0,90,0,0,0,254,0,19,0,96,0,129,0,111,0,0,0,1,0,81,0,250,0,47,0,166,0,62,0,204,0,5,0,33,0,155,0,228,0,242,0,164,0,18,0,203,0,161,0,105,0,0,0,107,0,0,0,0,0,120,0,37,0,0,0,43,0,0,0,120,0,0,0,239,0,0,0,154,0,249,0,63,0,129,0,233,0,184,0,0,0,39,0,0,0,75,0,240,0,151,0,233,0,0,0,36,0,133,0,204,0,31,0,106,0,193,0,26,0,0,0,8,0,153,0,0,0,0,0,95,0,96,0,13,0,253,0,254,0,177,0,208,0,255,0,0,0,152,0,146,0,252,0,107,0,211,0,131,0,144,0,164,0,0,0,96,0,44,0,61,0,0,0,3,0,32,0,142,0,0,0,20,0,15,0,0,0,0,0,0,0,53,0,95,0,162,0,157,0,18,0,41,0,151,0,230,0,167,0,9,0,0,0,35,0,0,0,199,0,55,0,17,0,0,0,62,0,91,0,0,0,34,0,0,0,88,0,27,0,65,0,0,0,94,0,0,0,187,0,79,0,0,0,86,0,89,0,91,0,31,0,71,0,130,0,235,0,0,0,81,0,109,0,204,0,251,0,0,0,247,0,116,0,0,0,0,0,162,0,121,0,0,0,0,0,143,0,177,0,58,0,245,0,122,0,0,0,237,0,20,0,0,0,0,0,91,0,0,0,0,0,0,0,0,0,82,0,174,0,109,0,13,0,124,0,0,0,254,0,137,0,225,0,38,0,24,0,99,0,230,0,220,0,213,0,10,0,37,0,12,0,81,0,190,0,15,0,60,0,132,0,233,0,0,0,11,0,135,0,56,0,163,0,209,0,98,0,225,0,122,0,13,0,39,0,45,0,98,0,0,0,33,0,106,0,210,0,63,0,145,0,0,0,19,0,0,0,171,0,126,0,115,0,25,0,105,0,153,0,99,0,249,0,248,0,87,0,7,0,235,0,240,0,11,0,128,0,35,0,32,0,104,0,249,0,0,0,45,0,147,0,239,0,208,0,0,0,110,0,247,0,200,0,70,0,159,0,51,0,234,0,227,0,238,0,105,0,215,0,18,0,42,0,248,0,63,0,11,0,152,0,76,0,69,0,56,0,173,0,111,0,150,0,251,0,0,0,132,0,7,0,239,0,132,0,34,0,47,0,137,0,0,0,0,0,42,0,178,0,26,0,66,0,0,0,137,0,196,0,46,0,27,0,200,0,0,0,255,0,0,0,200,0,98,0,88,0,174,0,142,0,68,0,105,0,189,0,124,0,244,0,214,0,169,0,96,0,61,0,96,0,143,0,0,0,99,0,83,0,239,0,254,0,145,0,248,0,14,0,1,0,150,0,190,0,63,0,10,0,134,0,62,0,127,0,159,0,54,0,0,0,227,0,96,0,65,0,175,0,205,0,214,0,44,0,21,0,170,0,38,0,128,0,0,0,0,0,210,0,212,0,100,0,216,0,32,0,34,0,111,0,174,0,0,0,194,0,226,0,92,0,0,0,120,0,196,0,142,0,129,0,216,0,0,0,195,0,41,0,0,0,208,0,156,0,150,0,199,0,0,0,152,0,0,0,11,0,117,0,19,0,0,0,221,0,0,0,42,0,234,0,159,0,242,0,135,0,129,0,0,0,149,0,203,0,184,0,0,0,94,0,40,0,101,0,100,0,214,0,138,0,159,0,89,0,167,0,47,0,139,0,253,0,0,0,8,0,134,0,127,0,203,0,98,0,0,0,18,0,7,0,155,0,49,0,94,0,242,0,220,0,0,0,0,0,238,0,173,0,72,0,230,0,252,0,56,0,0,0,137,0,195,0,121,0,31,0,0,0,0,0,138,0,21,0,0,0,148,0,214,0,196,0,144,0,138,0,171,0,83,0,148,0,0,0,0,0,106,0,0,0,217,0,0,0,184,0,130,0,37,0,94,0,238,0,135,0,201,0,104,0,0,0,179,0,0,0,101,0,93,0,154,0,246,0,102,0,155,0,193,0,46,0,0,0,99,0,157,0,0,0,0,0,0,0,60,0,196,0,30,0,86,0,165,0,225,0,15,0,210,0,0,0,20,0,68,0,255,0,42,0,196,0,121,0,35,0,148,0,68,0,0,0,71,0,224,0,84,0,164,0,111,0,173,0,62,0,0,0,123,0,203,0,235,0,185,0,233,0,32,0,57,0,171,0,189,0,129,0,193,0,151,0,56,0,219,0,103,0,249,0,209,0,140,0,245,0,127,0,119,0,211,0,104,0,0,0,0,0,89,0,81,0,131,0,32,0,24,0,0,0,14,0,165,0,146,0,144,0,0,0,135,0,0,0,81,0,0,0,0,0,48,0,112,0,236,0,232,0,150,0,95,0,134,0,44,0,152,0,114,0,0,0,0,0,75,0,143,0,206,0,92,0,140,0,226,0,159,0,221,0,150,0,242,0,0,0,69,0,196,0,0,0,179,0,193,0,0,0,0,0,153,0,131,0,0,0,220,0,47,0,4,0,123,0,0,0,0,0,115,0,121,0,0,0,60,0,254,0,182,0,84,0,164,0,160,0,152,0,228,0,12,0,31,0,189,0,72,0,196,0,116,0,64,0,65,0,220,0,168,0,40,0,238,0,0,0,0,0,9,0,0,0,60,0,0,0,126,0,61,0,188,0);
signal scenario_full  : scenario_type := (244,31,244,30,244,29,71,31,131,31,86,31,18,31,137,31,207,31,151,31,5,31,172,31,172,30,25,31,64,31,64,30,64,29,64,28,236,31,236,30,56,31,56,30,127,31,244,31,223,31,223,30,181,31,54,31,17,31,145,31,93,31,177,31,246,31,159,31,230,31,230,30,198,31,101,31,187,31,42,31,127,31,127,30,127,29,127,28,27,31,27,30,168,31,58,31,144,31,116,31,253,31,44,31,61,31,47,31,2,31,239,31,239,30,40,31,227,31,227,30,30,31,91,31,253,31,202,31,105,31,105,30,106,31,106,30,34,31,114,31,114,30,114,29,149,31,97,31,125,31,138,31,215,31,174,31,26,31,131,31,57,31,25,31,115,31,170,31,183,31,183,30,100,31,112,31,112,30,162,31,68,31,14,31,69,31,225,31,195,31,195,30,248,31,48,31,254,31,254,30,254,29,175,31,151,31,113,31,212,31,85,31,135,31,105,31,105,30,188,31,143,31,137,31,175,31,175,30,43,31,204,31,186,31,79,31,94,31,187,31,27,31,253,31,181,31,56,31,248,31,190,31,187,31,242,31,159,31,244,31,205,31,205,30,110,31,174,31,125,31,145,31,64,31,64,30,64,29,201,31,153,31,147,31,119,31,162,31,126,31,126,30,236,31,195,31,195,30,195,31,168,31,168,30,168,29,11,31,11,30,97,31,201,31,244,31,244,30,110,31,139,31,7,31,26,31,130,31,117,31,109,31,222,31,18,31,18,30,48,31,117,31,117,30,169,31,238,31,29,31,66,31,66,30,81,31,166,31,74,31,15,31,56,31,56,30,124,31,124,30,135,31,57,31,59,31,56,31,128,31,91,31,12,31,15,31,235,31,222,31,125,31,125,30,125,29,194,31,2,31,29,31,29,30,227,31,227,30,227,29,224,31,215,31,120,31,120,30,123,31,104,31,202,31,194,31,17,31,47,31,82,31,87,31,105,31,115,31,115,30,47,31,197,31,179,31,216,31,216,31,77,31,179,31,96,31,88,31,6,31,11,31,81,31,25,31,217,31,38,31,38,30,90,31,49,31,226,31,166,31,253,31,120,31,120,30,120,29,120,28,120,27,120,26,169,31,135,31,90,31,90,30,254,31,19,31,96,31,129,31,111,31,111,30,1,31,81,31,250,31,47,31,166,31,62,31,204,31,5,31,33,31,155,31,228,31,242,31,164,31,18,31,203,31,161,31,105,31,105,30,107,31,107,30,107,29,120,31,37,31,37,30,43,31,43,30,120,31,120,30,239,31,239,30,154,31,249,31,63,31,129,31,233,31,184,31,184,30,39,31,39,30,75,31,240,31,151,31,233,31,233,30,36,31,133,31,204,31,31,31,106,31,193,31,26,31,26,30,8,31,153,31,153,30,153,29,95,31,96,31,13,31,253,31,254,31,177,31,208,31,255,31,255,30,152,31,146,31,252,31,107,31,211,31,131,31,144,31,164,31,164,30,96,31,44,31,61,31,61,30,3,31,32,31,142,31,142,30,20,31,15,31,15,30,15,29,15,28,53,31,95,31,162,31,157,31,18,31,41,31,151,31,230,31,167,31,9,31,9,30,35,31,35,30,199,31,55,31,17,31,17,30,62,31,91,31,91,30,34,31,34,30,88,31,27,31,65,31,65,30,94,31,94,30,187,31,79,31,79,30,86,31,89,31,91,31,31,31,71,31,130,31,235,31,235,30,81,31,109,31,204,31,251,31,251,30,247,31,116,31,116,30,116,29,162,31,121,31,121,30,121,29,143,31,177,31,58,31,245,31,122,31,122,30,237,31,20,31,20,30,20,29,91,31,91,30,91,29,91,28,91,27,82,31,174,31,109,31,13,31,124,31,124,30,254,31,137,31,225,31,38,31,24,31,99,31,230,31,220,31,213,31,10,31,37,31,12,31,81,31,190,31,15,31,60,31,132,31,233,31,233,30,11,31,135,31,56,31,163,31,209,31,98,31,225,31,122,31,13,31,39,31,45,31,98,31,98,30,33,31,106,31,210,31,63,31,145,31,145,30,19,31,19,30,171,31,126,31,115,31,25,31,105,31,153,31,99,31,249,31,248,31,87,31,7,31,235,31,240,31,11,31,128,31,35,31,32,31,104,31,249,31,249,30,45,31,147,31,239,31,208,31,208,30,110,31,247,31,200,31,70,31,159,31,51,31,234,31,227,31,238,31,105,31,215,31,18,31,42,31,248,31,63,31,11,31,152,31,76,31,69,31,56,31,173,31,111,31,150,31,251,31,251,30,132,31,7,31,239,31,132,31,34,31,47,31,137,31,137,30,137,29,42,31,178,31,26,31,66,31,66,30,137,31,196,31,46,31,27,31,200,31,200,30,255,31,255,30,200,31,98,31,88,31,174,31,142,31,68,31,105,31,189,31,124,31,244,31,214,31,169,31,96,31,61,31,96,31,143,31,143,30,99,31,83,31,239,31,254,31,145,31,248,31,14,31,1,31,150,31,190,31,63,31,10,31,134,31,62,31,127,31,159,31,54,31,54,30,227,31,96,31,65,31,175,31,205,31,214,31,44,31,21,31,170,31,38,31,128,31,128,30,128,29,210,31,212,31,100,31,216,31,32,31,34,31,111,31,174,31,174,30,194,31,226,31,92,31,92,30,120,31,196,31,142,31,129,31,216,31,216,30,195,31,41,31,41,30,208,31,156,31,150,31,199,31,199,30,152,31,152,30,11,31,117,31,19,31,19,30,221,31,221,30,42,31,234,31,159,31,242,31,135,31,129,31,129,30,149,31,203,31,184,31,184,30,94,31,40,31,101,31,100,31,214,31,138,31,159,31,89,31,167,31,47,31,139,31,253,31,253,30,8,31,134,31,127,31,203,31,98,31,98,30,18,31,7,31,155,31,49,31,94,31,242,31,220,31,220,30,220,29,238,31,173,31,72,31,230,31,252,31,56,31,56,30,137,31,195,31,121,31,31,31,31,30,31,29,138,31,21,31,21,30,148,31,214,31,196,31,144,31,138,31,171,31,83,31,148,31,148,30,148,29,106,31,106,30,217,31,217,30,184,31,130,31,37,31,94,31,238,31,135,31,201,31,104,31,104,30,179,31,179,30,101,31,93,31,154,31,246,31,102,31,155,31,193,31,46,31,46,30,99,31,157,31,157,30,157,29,157,28,60,31,196,31,30,31,86,31,165,31,225,31,15,31,210,31,210,30,20,31,68,31,255,31,42,31,196,31,121,31,35,31,148,31,68,31,68,30,71,31,224,31,84,31,164,31,111,31,173,31,62,31,62,30,123,31,203,31,235,31,185,31,233,31,32,31,57,31,171,31,189,31,129,31,193,31,151,31,56,31,219,31,103,31,249,31,209,31,140,31,245,31,127,31,119,31,211,31,104,31,104,30,104,29,89,31,81,31,131,31,32,31,24,31,24,30,14,31,165,31,146,31,144,31,144,30,135,31,135,30,81,31,81,30,81,29,48,31,112,31,236,31,232,31,150,31,95,31,134,31,44,31,152,31,114,31,114,30,114,29,75,31,143,31,206,31,92,31,140,31,226,31,159,31,221,31,150,31,242,31,242,30,69,31,196,31,196,30,179,31,193,31,193,30,193,29,153,31,131,31,131,30,220,31,47,31,4,31,123,31,123,30,123,29,115,31,121,31,121,30,60,31,254,31,182,31,84,31,164,31,160,31,152,31,228,31,12,31,31,31,189,31,72,31,196,31,116,31,64,31,65,31,220,31,168,31,40,31,238,31,238,30,238,29,9,31,9,30,60,31,60,30,126,31,61,31,188,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
