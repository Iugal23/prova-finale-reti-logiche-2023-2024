-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_654 is
end project_tb_654;

architecture project_tb_arch_654 of project_tb_654 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 755;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,59,0,232,0,106,0,126,0,165,0,180,0,58,0,255,0,54,0,216,0,0,0,221,0,153,0,99,0,179,0,115,0,154,0,50,0,0,0,0,0,244,0,65,0,0,0,62,0,190,0,52,0,98,0,168,0,198,0,215,0,76,0,59,0,191,0,55,0,118,0,56,0,0,0,212,0,27,0,146,0,219,0,216,0,0,0,80,0,183,0,254,0,181,0,0,0,118,0,101,0,128,0,205,0,39,0,55,0,111,0,222,0,174,0,42,0,122,0,5,0,188,0,184,0,14,0,9,0,0,0,120,0,41,0,38,0,0,0,159,0,170,0,0,0,56,0,185,0,0,0,69,0,227,0,254,0,0,0,68,0,3,0,211,0,42,0,1,0,60,0,33,0,55,0,82,0,61,0,0,0,0,0,0,0,136,0,122,0,0,0,0,0,132,0,103,0,0,0,5,0,187,0,65,0,113,0,159,0,153,0,0,0,192,0,51,0,118,0,40,0,191,0,0,0,218,0,0,0,44,0,175,0,154,0,111,0,80,0,151,0,218,0,213,0,238,0,141,0,9,0,114,0,52,0,87,0,0,0,221,0,23,0,0,0,4,0,0,0,15,0,204,0,0,0,183,0,0,0,0,0,186,0,48,0,0,0,0,0,132,0,0,0,180,0,193,0,83,0,0,0,69,0,111,0,0,0,189,0,111,0,246,0,146,0,0,0,216,0,229,0,208,0,0,0,119,0,0,0,55,0,93,0,40,0,133,0,0,0,18,0,0,0,191,0,0,0,97,0,163,0,122,0,125,0,106,0,192,0,17,0,80,0,0,0,123,0,223,0,87,0,158,0,90,0,89,0,180,0,157,0,34,0,101,0,23,0,146,0,109,0,0,0,171,0,82,0,0,0,32,0,46,0,241,0,89,0,161,0,0,0,199,0,2,0,0,0,209,0,101,0,40,0,84,0,139,0,120,0,134,0,249,0,142,0,55,0,0,0,98,0,113,0,249,0,70,0,0,0,0,0,255,0,47,0,142,0,209,0,176,0,228,0,0,0,0,0,128,0,195,0,115,0,59,0,125,0,198,0,96,0,14,0,146,0,115,0,44,0,8,0,38,0,0,0,66,0,72,0,254,0,0,0,92,0,208,0,33,0,125,0,38,0,30,0,225,0,185,0,158,0,174,0,244,0,0,0,3,0,167,0,0,0,82,0,19,0,7,0,95,0,0,0,52,0,179,0,199,0,21,0,31,0,199,0,162,0,215,0,229,0,163,0,247,0,154,0,0,0,238,0,32,0,216,0,246,0,30,0,9,0,33,0,9,0,97,0,236,0,132,0,0,0,0,0,96,0,231,0,120,0,249,0,73,0,153,0,100,0,233,0,37,0,0,0,160,0,193,0,70,0,112,0,95,0,83,0,49,0,235,0,121,0,215,0,179,0,129,0,217,0,198,0,0,0,250,0,35,0,0,0,148,0,18,0,138,0,50,0,1,0,138,0,136,0,48,0,242,0,143,0,170,0,84,0,150,0,0,0,16,0,0,0,97,0,140,0,16,0,14,0,248,0,37,0,0,0,243,0,191,0,0,0,65,0,207,0,0,0,17,0,0,0,213,0,116,0,6,0,0,0,92,0,184,0,124,0,249,0,200,0,34,0,249,0,0,0,26,0,0,0,14,0,156,0,146,0,223,0,209,0,215,0,77,0,0,0,82,0,217,0,84,0,33,0,0,0,1,0,3,0,0,0,170,0,113,0,248,0,233,0,238,0,238,0,250,0,166,0,142,0,6,0,14,0,127,0,76,0,0,0,0,0,0,0,0,0,177,0,0,0,0,0,145,0,34,0,123,0,130,0,213,0,229,0,0,0,199,0,122,0,107,0,135,0,159,0,195,0,107,0,56,0,239,0,0,0,224,0,0,0,140,0,18,0,0,0,151,0,205,0,102,0,54,0,135,0,90,0,14,0,27,0,186,0,81,0,138,0,4,0,38,0,124,0,4,0,5,0,92,0,0,0,0,0,0,0,0,0,183,0,113,0,10,0,0,0,218,0,55,0,0,0,42,0,245,0,62,0,0,0,214,0,35,0,109,0,154,0,97,0,114,0,30,0,149,0,105,0,105,0,97,0,245,0,0,0,135,0,212,0,0,0,22,0,0,0,121,0,39,0,141,0,84,0,0,0,193,0,0,0,174,0,139,0,162,0,158,0,34,0,91,0,0,0,132,0,129,0,1,0,9,0,225,0,19,0,244,0,0,0,111,0,169,0,29,0,0,0,210,0,115,0,105,0,85,0,185,0,0,0,178,0,185,0,169,0,103,0,14,0,32,0,130,0,16,0,227,0,45,0,221,0,103,0,172,0,118,0,188,0,54,0,208,0,19,0,232,0,128,0,102,0,0,0,0,0,72,0,230,0,0,0,252,0,217,0,105,0,0,0,0,0,0,0,187,0,0,0,0,0,245,0,253,0,0,0,11,0,30,0,0,0,241,0,58,0,159,0,143,0,128,0,52,0,175,0,0,0,189,0,0,0,28,0,224,0,0,0,224,0,5,0,118,0,241,0,0,0,63,0,73,0,147,0,196,0,203,0,177,0,238,0,111,0,40,0,122,0,0,0,52,0,159,0,42,0,0,0,0,0,226,0,47,0,157,0,99,0,120,0,226,0,118,0,146,0,0,0,24,0,31,0,230,0,239,0,202,0,114,0,128,0,26,0,87,0,59,0,13,0,38,0,0,0,61,0,246,0,158,0,103,0,42,0,0,0,0,0,254,0,173,0,0,0,7,0,100,0,162,0,222,0,209,0,153,0,188,0,0,0,215,0,56,0,194,0,54,0,0,0,0,0,129,0,0,0,196,0,0,0,129,0,0,0,0,0,0,0,0,0,0,0,238,0,195,0,226,0,0,0,0,0,135,0,0,0,62,0,14,0,11,0,0,0,0,0,215,0,236,0,67,0,33,0,160,0,0,0,248,0,118,0,22,0,18,0,132,0,0,0,189,0,0,0,237,0,4,0,106,0,63,0,0,0,144,0,133,0,66,0,0,0,218,0,160,0,22,0,186,0,254,0,72,0,68,0,0,0,96,0,202,0,239,0,219,0,11,0,30,0,0,0,171,0,0,0,0,0,82,0,145,0,184,0,0,0,88,0,15,0,99,0,92,0,226,0,0,0,56,0,171,0,3,0,139,0,1,0,82,0,89,0,4,0,109,0,14,0,208,0,0,0,98,0,0,0,32,0,84,0,142,0,0,0,194,0,0,0,0,0,149,0,194,0,28,0,177,0,55,0,163,0,51,0,134,0,43,0,226,0,190,0,137,0,113,0,248,0,216,0,135,0,136,0,166,0,0,0,0,0,0,0,158,0,0,0,15,0,224,0,189,0,74,0,95,0,164,0);
signal scenario_full  : scenario_type := (0,0,59,31,232,31,106,31,126,31,165,31,180,31,58,31,255,31,54,31,216,31,216,30,221,31,153,31,99,31,179,31,115,31,154,31,50,31,50,30,50,29,244,31,65,31,65,30,62,31,190,31,52,31,98,31,168,31,198,31,215,31,76,31,59,31,191,31,55,31,118,31,56,31,56,30,212,31,27,31,146,31,219,31,216,31,216,30,80,31,183,31,254,31,181,31,181,30,118,31,101,31,128,31,205,31,39,31,55,31,111,31,222,31,174,31,42,31,122,31,5,31,188,31,184,31,14,31,9,31,9,30,120,31,41,31,38,31,38,30,159,31,170,31,170,30,56,31,185,31,185,30,69,31,227,31,254,31,254,30,68,31,3,31,211,31,42,31,1,31,60,31,33,31,55,31,82,31,61,31,61,30,61,29,61,28,136,31,122,31,122,30,122,29,132,31,103,31,103,30,5,31,187,31,65,31,113,31,159,31,153,31,153,30,192,31,51,31,118,31,40,31,191,31,191,30,218,31,218,30,44,31,175,31,154,31,111,31,80,31,151,31,218,31,213,31,238,31,141,31,9,31,114,31,52,31,87,31,87,30,221,31,23,31,23,30,4,31,4,30,15,31,204,31,204,30,183,31,183,30,183,29,186,31,48,31,48,30,48,29,132,31,132,30,180,31,193,31,83,31,83,30,69,31,111,31,111,30,189,31,111,31,246,31,146,31,146,30,216,31,229,31,208,31,208,30,119,31,119,30,55,31,93,31,40,31,133,31,133,30,18,31,18,30,191,31,191,30,97,31,163,31,122,31,125,31,106,31,192,31,17,31,80,31,80,30,123,31,223,31,87,31,158,31,90,31,89,31,180,31,157,31,34,31,101,31,23,31,146,31,109,31,109,30,171,31,82,31,82,30,32,31,46,31,241,31,89,31,161,31,161,30,199,31,2,31,2,30,209,31,101,31,40,31,84,31,139,31,120,31,134,31,249,31,142,31,55,31,55,30,98,31,113,31,249,31,70,31,70,30,70,29,255,31,47,31,142,31,209,31,176,31,228,31,228,30,228,29,128,31,195,31,115,31,59,31,125,31,198,31,96,31,14,31,146,31,115,31,44,31,8,31,38,31,38,30,66,31,72,31,254,31,254,30,92,31,208,31,33,31,125,31,38,31,30,31,225,31,185,31,158,31,174,31,244,31,244,30,3,31,167,31,167,30,82,31,19,31,7,31,95,31,95,30,52,31,179,31,199,31,21,31,31,31,199,31,162,31,215,31,229,31,163,31,247,31,154,31,154,30,238,31,32,31,216,31,246,31,30,31,9,31,33,31,9,31,97,31,236,31,132,31,132,30,132,29,96,31,231,31,120,31,249,31,73,31,153,31,100,31,233,31,37,31,37,30,160,31,193,31,70,31,112,31,95,31,83,31,49,31,235,31,121,31,215,31,179,31,129,31,217,31,198,31,198,30,250,31,35,31,35,30,148,31,18,31,138,31,50,31,1,31,138,31,136,31,48,31,242,31,143,31,170,31,84,31,150,31,150,30,16,31,16,30,97,31,140,31,16,31,14,31,248,31,37,31,37,30,243,31,191,31,191,30,65,31,207,31,207,30,17,31,17,30,213,31,116,31,6,31,6,30,92,31,184,31,124,31,249,31,200,31,34,31,249,31,249,30,26,31,26,30,14,31,156,31,146,31,223,31,209,31,215,31,77,31,77,30,82,31,217,31,84,31,33,31,33,30,1,31,3,31,3,30,170,31,113,31,248,31,233,31,238,31,238,31,250,31,166,31,142,31,6,31,14,31,127,31,76,31,76,30,76,29,76,28,76,27,177,31,177,30,177,29,145,31,34,31,123,31,130,31,213,31,229,31,229,30,199,31,122,31,107,31,135,31,159,31,195,31,107,31,56,31,239,31,239,30,224,31,224,30,140,31,18,31,18,30,151,31,205,31,102,31,54,31,135,31,90,31,14,31,27,31,186,31,81,31,138,31,4,31,38,31,124,31,4,31,5,31,92,31,92,30,92,29,92,28,92,27,183,31,113,31,10,31,10,30,218,31,55,31,55,30,42,31,245,31,62,31,62,30,214,31,35,31,109,31,154,31,97,31,114,31,30,31,149,31,105,31,105,31,97,31,245,31,245,30,135,31,212,31,212,30,22,31,22,30,121,31,39,31,141,31,84,31,84,30,193,31,193,30,174,31,139,31,162,31,158,31,34,31,91,31,91,30,132,31,129,31,1,31,9,31,225,31,19,31,244,31,244,30,111,31,169,31,29,31,29,30,210,31,115,31,105,31,85,31,185,31,185,30,178,31,185,31,169,31,103,31,14,31,32,31,130,31,16,31,227,31,45,31,221,31,103,31,172,31,118,31,188,31,54,31,208,31,19,31,232,31,128,31,102,31,102,30,102,29,72,31,230,31,230,30,252,31,217,31,105,31,105,30,105,29,105,28,187,31,187,30,187,29,245,31,253,31,253,30,11,31,30,31,30,30,241,31,58,31,159,31,143,31,128,31,52,31,175,31,175,30,189,31,189,30,28,31,224,31,224,30,224,31,5,31,118,31,241,31,241,30,63,31,73,31,147,31,196,31,203,31,177,31,238,31,111,31,40,31,122,31,122,30,52,31,159,31,42,31,42,30,42,29,226,31,47,31,157,31,99,31,120,31,226,31,118,31,146,31,146,30,24,31,31,31,230,31,239,31,202,31,114,31,128,31,26,31,87,31,59,31,13,31,38,31,38,30,61,31,246,31,158,31,103,31,42,31,42,30,42,29,254,31,173,31,173,30,7,31,100,31,162,31,222,31,209,31,153,31,188,31,188,30,215,31,56,31,194,31,54,31,54,30,54,29,129,31,129,30,196,31,196,30,129,31,129,30,129,29,129,28,129,27,129,26,238,31,195,31,226,31,226,30,226,29,135,31,135,30,62,31,14,31,11,31,11,30,11,29,215,31,236,31,67,31,33,31,160,31,160,30,248,31,118,31,22,31,18,31,132,31,132,30,189,31,189,30,237,31,4,31,106,31,63,31,63,30,144,31,133,31,66,31,66,30,218,31,160,31,22,31,186,31,254,31,72,31,68,31,68,30,96,31,202,31,239,31,219,31,11,31,30,31,30,30,171,31,171,30,171,29,82,31,145,31,184,31,184,30,88,31,15,31,99,31,92,31,226,31,226,30,56,31,171,31,3,31,139,31,1,31,82,31,89,31,4,31,109,31,14,31,208,31,208,30,98,31,98,30,32,31,84,31,142,31,142,30,194,31,194,30,194,29,149,31,194,31,28,31,177,31,55,31,163,31,51,31,134,31,43,31,226,31,190,31,137,31,113,31,248,31,216,31,135,31,136,31,166,31,166,30,166,29,166,28,158,31,158,30,15,31,224,31,189,31,74,31,95,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
