-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 795;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (230,0,216,0,0,0,137,0,14,0,123,0,229,0,184,0,0,0,19,0,0,0,81,0,16,0,21,0,172,0,81,0,6,0,117,0,0,0,146,0,54,0,0,0,152,0,82,0,0,0,7,0,10,0,89,0,173,0,66,0,0,0,17,0,221,0,152,0,171,0,188,0,186,0,108,0,124,0,134,0,139,0,0,0,37,0,0,0,62,0,130,0,21,0,111,0,250,0,206,0,16,0,23,0,0,0,217,0,134,0,182,0,192,0,50,0,79,0,192,0,103,0,0,0,157,0,0,0,191,0,112,0,26,0,191,0,119,0,213,0,0,0,71,0,40,0,183,0,203,0,0,0,245,0,135,0,26,0,0,0,0,0,0,0,0,0,254,0,133,0,91,0,0,0,106,0,133,0,0,0,155,0,81,0,234,0,0,0,170,0,172,0,127,0,185,0,14,0,31,0,146,0,0,0,16,0,49,0,73,0,237,0,248,0,200,0,75,0,120,0,32,0,101,0,42,0,137,0,0,0,216,0,227,0,85,0,0,0,35,0,187,0,0,0,44,0,0,0,222,0,101,0,33,0,189,0,152,0,0,0,80,0,0,0,201,0,166,0,39,0,250,0,0,0,120,0,74,0,118,0,21,0,78,0,0,0,151,0,0,0,0,0,103,0,62,0,0,0,0,0,0,0,204,0,204,0,0,0,0,0,154,0,0,0,71,0,109,0,64,0,90,0,54,0,118,0,5,0,217,0,74,0,0,0,140,0,0,0,125,0,176,0,94,0,102,0,204,0,239,0,32,0,135,0,164,0,140,0,126,0,71,0,83,0,51,0,16,0,253,0,32,0,252,0,62,0,0,0,0,0,0,0,16,0,227,0,228,0,215,0,121,0,35,0,251,0,164,0,196,0,97,0,30,0,0,0,159,0,119,0,112,0,216,0,157,0,189,0,163,0,0,0,248,0,111,0,0,0,206,0,111,0,41,0,222,0,216,0,0,0,5,0,21,0,222,0,26,0,0,0,37,0,234,0,215,0,226,0,0,0,0,0,65,0,216,0,58,0,212,0,0,0,170,0,108,0,101,0,114,0,0,0,0,0,97,0,21,0,0,0,200,0,251,0,114,0,1,0,83,0,135,0,178,0,0,0,222,0,0,0,73,0,192,0,102,0,244,0,180,0,161,0,0,0,37,0,154,0,121,0,0,0,0,0,164,0,83,0,0,0,0,0,0,0,154,0,0,0,197,0,17,0,0,0,235,0,108,0,0,0,96,0,169,0,144,0,201,0,66,0,19,0,122,0,10,0,228,0,0,0,149,0,249,0,125,0,156,0,73,0,114,0,0,0,102,0,106,0,0,0,149,0,235,0,0,0,0,0,0,0,68,0,20,0,0,0,98,0,87,0,0,0,80,0,229,0,154,0,240,0,31,0,86,0,106,0,168,0,51,0,0,0,82,0,151,0,17,0,2,0,126,0,241,0,0,0,225,0,21,0,0,0,172,0,28,0,212,0,0,0,186,0,56,0,0,0,36,0,151,0,237,0,209,0,0,0,4,0,123,0,0,0,33,0,226,0,238,0,7,0,180,0,70,0,27,0,0,0,254,0,40,0,189,0,93,0,0,0,49,0,21,0,30,0,61,0,169,0,47,0,0,0,65,0,244,0,151,0,0,0,124,0,0,0,206,0,33,0,47,0,42,0,228,0,251,0,0,0,0,0,21,0,124,0,205,0,33,0,250,0,75,0,137,0,64,0,197,0,0,0,61,0,171,0,7,0,225,0,70,0,0,0,37,0,52,0,45,0,218,0,154,0,11,0,42,0,240,0,134,0,142,0,27,0,44,0,56,0,130,0,51,0,0,0,25,0,69,0,190,0,66,0,239,0,207,0,183,0,179,0,244,0,87,0,121,0,202,0,236,0,122,0,251,0,59,0,9,0,135,0,0,0,0,0,159,0,178,0,207,0,109,0,249,0,0,0,214,0,244,0,28,0,156,0,149,0,45,0,39,0,0,0,0,0,0,0,39,0,203,0,217,0,2,0,0,0,128,0,192,0,193,0,157,0,178,0,197,0,204,0,0,0,25,0,12,0,0,0,206,0,164,0,84,0,54,0,116,0,144,0,63,0,248,0,7,0,216,0,76,0,0,0,84,0,246,0,142,0,240,0,0,0,152,0,88,0,0,0,252,0,0,0,222,0,159,0,93,0,223,0,78,0,216,0,18,0,53,0,67,0,64,0,214,0,241,0,116,0,244,0,203,0,56,0,171,0,17,0,127,0,174,0,255,0,31,0,110,0,62,0,188,0,244,0,231,0,17,0,37,0,9,0,106,0,128,0,153,0,82,0,238,0,225,0,0,0,205,0,74,0,10,0,137,0,191,0,76,0,0,0,0,0,74,0,125,0,34,0,66,0,0,0,200,0,0,0,0,0,0,0,131,0,113,0,93,0,170,0,239,0,171,0,172,0,169,0,51,0,96,0,195,0,253,0,147,0,77,0,26,0,0,0,194,0,0,0,143,0,0,0,195,0,168,0,0,0,121,0,221,0,0,0,174,0,0,0,116,0,46,0,20,0,147,0,251,0,214,0,0,0,0,0,0,0,66,0,141,0,118,0,72,0,179,0,150,0,126,0,217,0,0,0,84,0,23,0,158,0,43,0,206,0,0,0,0,0,13,0,164,0,166,0,152,0,0,0,93,0,0,0,146,0,0,0,104,0,120,0,97,0,0,0,33,0,197,0,0,0,0,0,0,0,127,0,53,0,254,0,7,0,244,0,0,0,253,0,14,0,89,0,0,0,0,0,142,0,250,0,245,0,103,0,119,0,26,0,75,0,159,0,196,0,157,0,217,0,218,0,180,0,165,0,71,0,82,0,248,0,49,0,0,0,0,0,0,0,0,0,118,0,23,0,219,0,110,0,0,0,127,0,213,0,0,0,0,0,0,0,19,0,108,0,0,0,102,0,41,0,0,0,230,0,209,0,26,0,172,0,0,0,66,0,61,0,73,0,215,0,248,0,118,0,0,0,69,0,0,0,36,0,0,0,127,0,210,0,179,0,193,0,142,0,214,0,0,0,47,0,0,0,83,0,110,0,127,0,38,0,127,0,0,0,60,0,186,0,117,0,47,0,151,0,1,0,67,0,215,0,19,0,201,0,0,0,146,0,25,0,215,0,59,0,0,0,61,0,14,0,124,0,15,0,245,0,245,0,188,0,241,0,255,0,22,0,93,0,0,0,84,0,172,0,0,0,56,0,87,0,156,0,87,0,76,0,228,0,0,0,227,0,0,0,16,0,0,0,116,0,220,0,45,0,209,0,76,0,45,0,127,0,76,0,43,0,123,0,185,0,200,0,240,0,50,0,0,0,113,0,0,0,193,0,196,0,9,0,146,0,97,0,12,0,0,0,10,0,156,0,0,0,224,0,113,0,19,0,184,0,197,0,0,0,171,0,189,0,0,0,31,0,0,0,66,0,0,0,106,0,0,0,68,0,209,0,113,0,63,0,119,0,185,0,41,0,198,0,112,0,137,0,119,0,192,0,239,0,69,0,0,0,114,0,109,0,10,0,11,0,76,0);
signal scenario_full  : scenario_type := (230,31,216,31,216,30,137,31,14,31,123,31,229,31,184,31,184,30,19,31,19,30,81,31,16,31,21,31,172,31,81,31,6,31,117,31,117,30,146,31,54,31,54,30,152,31,82,31,82,30,7,31,10,31,89,31,173,31,66,31,66,30,17,31,221,31,152,31,171,31,188,31,186,31,108,31,124,31,134,31,139,31,139,30,37,31,37,30,62,31,130,31,21,31,111,31,250,31,206,31,16,31,23,31,23,30,217,31,134,31,182,31,192,31,50,31,79,31,192,31,103,31,103,30,157,31,157,30,191,31,112,31,26,31,191,31,119,31,213,31,213,30,71,31,40,31,183,31,203,31,203,30,245,31,135,31,26,31,26,30,26,29,26,28,26,27,254,31,133,31,91,31,91,30,106,31,133,31,133,30,155,31,81,31,234,31,234,30,170,31,172,31,127,31,185,31,14,31,31,31,146,31,146,30,16,31,49,31,73,31,237,31,248,31,200,31,75,31,120,31,32,31,101,31,42,31,137,31,137,30,216,31,227,31,85,31,85,30,35,31,187,31,187,30,44,31,44,30,222,31,101,31,33,31,189,31,152,31,152,30,80,31,80,30,201,31,166,31,39,31,250,31,250,30,120,31,74,31,118,31,21,31,78,31,78,30,151,31,151,30,151,29,103,31,62,31,62,30,62,29,62,28,204,31,204,31,204,30,204,29,154,31,154,30,71,31,109,31,64,31,90,31,54,31,118,31,5,31,217,31,74,31,74,30,140,31,140,30,125,31,176,31,94,31,102,31,204,31,239,31,32,31,135,31,164,31,140,31,126,31,71,31,83,31,51,31,16,31,253,31,32,31,252,31,62,31,62,30,62,29,62,28,16,31,227,31,228,31,215,31,121,31,35,31,251,31,164,31,196,31,97,31,30,31,30,30,159,31,119,31,112,31,216,31,157,31,189,31,163,31,163,30,248,31,111,31,111,30,206,31,111,31,41,31,222,31,216,31,216,30,5,31,21,31,222,31,26,31,26,30,37,31,234,31,215,31,226,31,226,30,226,29,65,31,216,31,58,31,212,31,212,30,170,31,108,31,101,31,114,31,114,30,114,29,97,31,21,31,21,30,200,31,251,31,114,31,1,31,83,31,135,31,178,31,178,30,222,31,222,30,73,31,192,31,102,31,244,31,180,31,161,31,161,30,37,31,154,31,121,31,121,30,121,29,164,31,83,31,83,30,83,29,83,28,154,31,154,30,197,31,17,31,17,30,235,31,108,31,108,30,96,31,169,31,144,31,201,31,66,31,19,31,122,31,10,31,228,31,228,30,149,31,249,31,125,31,156,31,73,31,114,31,114,30,102,31,106,31,106,30,149,31,235,31,235,30,235,29,235,28,68,31,20,31,20,30,98,31,87,31,87,30,80,31,229,31,154,31,240,31,31,31,86,31,106,31,168,31,51,31,51,30,82,31,151,31,17,31,2,31,126,31,241,31,241,30,225,31,21,31,21,30,172,31,28,31,212,31,212,30,186,31,56,31,56,30,36,31,151,31,237,31,209,31,209,30,4,31,123,31,123,30,33,31,226,31,238,31,7,31,180,31,70,31,27,31,27,30,254,31,40,31,189,31,93,31,93,30,49,31,21,31,30,31,61,31,169,31,47,31,47,30,65,31,244,31,151,31,151,30,124,31,124,30,206,31,33,31,47,31,42,31,228,31,251,31,251,30,251,29,21,31,124,31,205,31,33,31,250,31,75,31,137,31,64,31,197,31,197,30,61,31,171,31,7,31,225,31,70,31,70,30,37,31,52,31,45,31,218,31,154,31,11,31,42,31,240,31,134,31,142,31,27,31,44,31,56,31,130,31,51,31,51,30,25,31,69,31,190,31,66,31,239,31,207,31,183,31,179,31,244,31,87,31,121,31,202,31,236,31,122,31,251,31,59,31,9,31,135,31,135,30,135,29,159,31,178,31,207,31,109,31,249,31,249,30,214,31,244,31,28,31,156,31,149,31,45,31,39,31,39,30,39,29,39,28,39,31,203,31,217,31,2,31,2,30,128,31,192,31,193,31,157,31,178,31,197,31,204,31,204,30,25,31,12,31,12,30,206,31,164,31,84,31,54,31,116,31,144,31,63,31,248,31,7,31,216,31,76,31,76,30,84,31,246,31,142,31,240,31,240,30,152,31,88,31,88,30,252,31,252,30,222,31,159,31,93,31,223,31,78,31,216,31,18,31,53,31,67,31,64,31,214,31,241,31,116,31,244,31,203,31,56,31,171,31,17,31,127,31,174,31,255,31,31,31,110,31,62,31,188,31,244,31,231,31,17,31,37,31,9,31,106,31,128,31,153,31,82,31,238,31,225,31,225,30,205,31,74,31,10,31,137,31,191,31,76,31,76,30,76,29,74,31,125,31,34,31,66,31,66,30,200,31,200,30,200,29,200,28,131,31,113,31,93,31,170,31,239,31,171,31,172,31,169,31,51,31,96,31,195,31,253,31,147,31,77,31,26,31,26,30,194,31,194,30,143,31,143,30,195,31,168,31,168,30,121,31,221,31,221,30,174,31,174,30,116,31,46,31,20,31,147,31,251,31,214,31,214,30,214,29,214,28,66,31,141,31,118,31,72,31,179,31,150,31,126,31,217,31,217,30,84,31,23,31,158,31,43,31,206,31,206,30,206,29,13,31,164,31,166,31,152,31,152,30,93,31,93,30,146,31,146,30,104,31,120,31,97,31,97,30,33,31,197,31,197,30,197,29,197,28,127,31,53,31,254,31,7,31,244,31,244,30,253,31,14,31,89,31,89,30,89,29,142,31,250,31,245,31,103,31,119,31,26,31,75,31,159,31,196,31,157,31,217,31,218,31,180,31,165,31,71,31,82,31,248,31,49,31,49,30,49,29,49,28,49,27,118,31,23,31,219,31,110,31,110,30,127,31,213,31,213,30,213,29,213,28,19,31,108,31,108,30,102,31,41,31,41,30,230,31,209,31,26,31,172,31,172,30,66,31,61,31,73,31,215,31,248,31,118,31,118,30,69,31,69,30,36,31,36,30,127,31,210,31,179,31,193,31,142,31,214,31,214,30,47,31,47,30,83,31,110,31,127,31,38,31,127,31,127,30,60,31,186,31,117,31,47,31,151,31,1,31,67,31,215,31,19,31,201,31,201,30,146,31,25,31,215,31,59,31,59,30,61,31,14,31,124,31,15,31,245,31,245,31,188,31,241,31,255,31,22,31,93,31,93,30,84,31,172,31,172,30,56,31,87,31,156,31,87,31,76,31,228,31,228,30,227,31,227,30,16,31,16,30,116,31,220,31,45,31,209,31,76,31,45,31,127,31,76,31,43,31,123,31,185,31,200,31,240,31,50,31,50,30,113,31,113,30,193,31,196,31,9,31,146,31,97,31,12,31,12,30,10,31,156,31,156,30,224,31,113,31,19,31,184,31,197,31,197,30,171,31,189,31,189,30,31,31,31,30,66,31,66,30,106,31,106,30,68,31,209,31,113,31,63,31,119,31,185,31,41,31,198,31,112,31,137,31,119,31,192,31,239,31,69,31,69,30,114,31,109,31,10,31,11,31,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
