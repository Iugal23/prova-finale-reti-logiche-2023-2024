-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_436 is
end project_tb_436;

architecture project_tb_arch_436 of project_tb_436 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 659;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (8,0,224,0,71,0,29,0,146,0,164,0,241,0,100,0,0,0,35,0,158,0,235,0,208,0,85,0,102,0,0,0,226,0,0,0,165,0,222,0,208,0,139,0,0,0,42,0,0,0,57,0,0,0,204,0,206,0,236,0,122,0,0,0,103,0,95,0,178,0,224,0,182,0,48,0,104,0,79,0,0,0,0,0,177,0,82,0,190,0,14,0,23,0,127,0,13,0,69,0,14,0,214,0,221,0,19,0,174,0,210,0,10,0,238,0,213,0,0,0,208,0,19,0,0,0,252,0,0,0,154,0,140,0,141,0,130,0,221,0,45,0,151,0,0,0,201,0,0,0,197,0,184,0,102,0,178,0,123,0,0,0,50,0,229,0,190,0,6,0,168,0,98,0,0,0,3,0,0,0,59,0,118,0,16,0,210,0,0,0,0,0,215,0,14,0,0,0,0,0,132,0,192,0,0,0,163,0,62,0,89,0,88,0,0,0,187,0,0,0,72,0,99,0,118,0,1,0,94,0,0,0,58,0,0,0,0,0,241,0,61,0,251,0,0,0,0,0,227,0,0,0,0,0,201,0,0,0,0,0,177,0,225,0,58,0,15,0,113,0,53,0,197,0,0,0,235,0,203,0,231,0,124,0,104,0,71,0,253,0,152,0,98,0,119,0,172,0,183,0,222,0,181,0,0,0,0,0,0,0,163,0,0,0,0,0,0,0,117,0,76,0,141,0,252,0,145,0,67,0,121,0,0,0,60,0,113,0,147,0,192,0,12,0,125,0,241,0,93,0,83,0,98,0,113,0,0,0,0,0,101,0,16,0,81,0,0,0,0,0,91,0,253,0,36,0,144,0,237,0,83,0,159,0,0,0,0,0,92,0,90,0,202,0,227,0,208,0,189,0,0,0,54,0,180,0,213,0,251,0,159,0,0,0,19,0,142,0,191,0,246,0,15,0,80,0,114,0,68,0,0,0,25,0,18,0,172,0,72,0,0,0,99,0,81,0,152,0,177,0,219,0,78,0,17,0,218,0,224,0,197,0,50,0,94,0,68,0,0,0,0,0,37,0,229,0,0,0,147,0,241,0,0,0,90,0,118,0,27,0,29,0,148,0,0,0,121,0,0,0,142,0,57,0,115,0,157,0,241,0,230,0,199,0,91,0,166,0,104,0,127,0,86,0,144,0,228,0,0,0,23,0,210,0,88,0,198,0,40,0,189,0,0,0,32,0,119,0,77,0,137,0,159,0,142,0,84,0,135,0,99,0,0,0,14,0,0,0,0,0,107,0,163,0,238,0,125,0,224,0,76,0,21,0,90,0,99,0,88,0,229,0,10,0,166,0,0,0,215,0,21,0,224,0,133,0,53,0,48,0,0,0,243,0,198,0,70,0,0,0,101,0,194,0,226,0,46,0,86,0,158,0,118,0,59,0,241,0,0,0,63,0,0,0,0,0,138,0,184,0,129,0,239,0,166,0,225,0,75,0,0,0,93,0,0,0,215,0,225,0,113,0,70,0,244,0,179,0,201,0,9,0,187,0,180,0,176,0,77,0,158,0,0,0,166,0,245,0,46,0,181,0,184,0,246,0,0,0,101,0,183,0,0,0,210,0,209,0,0,0,243,0,21,0,36,0,33,0,234,0,22,0,0,0,162,0,227,0,119,0,166,0,30,0,238,0,24,0,0,0,75,0,196,0,110,0,0,0,0,0,125,0,116,0,73,0,0,0,83,0,24,0,234,0,147,0,41,0,0,0,19,0,0,0,24,0,106,0,41,0,91,0,0,0,242,0,138,0,165,0,179,0,28,0,148,0,225,0,136,0,0,0,0,0,83,0,228,0,35,0,0,0,0,0,114,0,208,0,21,0,26,0,0,0,233,0,66,0,0,0,194,0,59,0,5,0,58,0,83,0,48,0,108,0,141,0,227,0,101,0,219,0,45,0,199,0,173,0,100,0,187,0,120,0,139,0,214,0,58,0,0,0,67,0,171,0,248,0,55,0,175,0,253,0,188,0,8,0,173,0,170,0,0,0,110,0,64,0,32,0,188,0,195,0,0,0,224,0,133,0,243,0,76,0,0,0,18,0,0,0,187,0,154,0,215,0,67,0,22,0,255,0,235,0,0,0,0,0,124,0,0,0,63,0,0,0,68,0,31,0,127,0,0,0,218,0,171,0,0,0,72,0,0,0,45,0,72,0,144,0,98,0,5,0,185,0,0,0,63,0,221,0,151,0,79,0,174,0,35,0,240,0,175,0,154,0,96,0,45,0,125,0,88,0,250,0,2,0,0,0,164,0,119,0,226,0,160,0,0,0,18,0,255,0,44,0,0,0,121,0,184,0,56,0,7,0,158,0,11,0,107,0,56,0,33,0,185,0,71,0,210,0,188,0,0,0,33,0,160,0,128,0,8,0,213,0,0,0,116,0,124,0,0,0,56,0,164,0,24,0,115,0,0,0,199,0,136,0,215,0,213,0,207,0,204,0,255,0,139,0,98,0,63,0,28,0,59,0,150,0,179,0,131,0,254,0,58,0,125,0,148,0,220,0,203,0,44,0,24,0,142,0,0,0,65,0,121,0,174,0,155,0,0,0,141,0,40,0,191,0,0,0,243,0,33,0,23,0,0,0,137,0,28,0,17,0,238,0,191,0,175,0,0,0,235,0,125,0,85,0,0,0,83,0,255,0,0,0,208,0,0,0,96,0,162,0,145,0,0,0,124,0,0,0,240,0,165,0,0,0,219,0,7,0,0,0,120,0,0,0,0,0,85,0,222,0,255,0,163,0,201,0,0,0,127,0,20,0,11,0,52,0,60,0,59,0,171,0,223,0,0,0,0,0,113,0,212,0,25,0,235,0,143,0,71,0,12,0,213,0,110,0,224,0,0,0,39,0,9,0,29,0,10,0,156,0,130,0,162,0,0,0,116,0,104,0,234,0,179,0,0,0,0,0,168,0,51,0);
signal scenario_full  : scenario_type := (8,31,224,31,71,31,29,31,146,31,164,31,241,31,100,31,100,30,35,31,158,31,235,31,208,31,85,31,102,31,102,30,226,31,226,30,165,31,222,31,208,31,139,31,139,30,42,31,42,30,57,31,57,30,204,31,206,31,236,31,122,31,122,30,103,31,95,31,178,31,224,31,182,31,48,31,104,31,79,31,79,30,79,29,177,31,82,31,190,31,14,31,23,31,127,31,13,31,69,31,14,31,214,31,221,31,19,31,174,31,210,31,10,31,238,31,213,31,213,30,208,31,19,31,19,30,252,31,252,30,154,31,140,31,141,31,130,31,221,31,45,31,151,31,151,30,201,31,201,30,197,31,184,31,102,31,178,31,123,31,123,30,50,31,229,31,190,31,6,31,168,31,98,31,98,30,3,31,3,30,59,31,118,31,16,31,210,31,210,30,210,29,215,31,14,31,14,30,14,29,132,31,192,31,192,30,163,31,62,31,89,31,88,31,88,30,187,31,187,30,72,31,99,31,118,31,1,31,94,31,94,30,58,31,58,30,58,29,241,31,61,31,251,31,251,30,251,29,227,31,227,30,227,29,201,31,201,30,201,29,177,31,225,31,58,31,15,31,113,31,53,31,197,31,197,30,235,31,203,31,231,31,124,31,104,31,71,31,253,31,152,31,98,31,119,31,172,31,183,31,222,31,181,31,181,30,181,29,181,28,163,31,163,30,163,29,163,28,117,31,76,31,141,31,252,31,145,31,67,31,121,31,121,30,60,31,113,31,147,31,192,31,12,31,125,31,241,31,93,31,83,31,98,31,113,31,113,30,113,29,101,31,16,31,81,31,81,30,81,29,91,31,253,31,36,31,144,31,237,31,83,31,159,31,159,30,159,29,92,31,90,31,202,31,227,31,208,31,189,31,189,30,54,31,180,31,213,31,251,31,159,31,159,30,19,31,142,31,191,31,246,31,15,31,80,31,114,31,68,31,68,30,25,31,18,31,172,31,72,31,72,30,99,31,81,31,152,31,177,31,219,31,78,31,17,31,218,31,224,31,197,31,50,31,94,31,68,31,68,30,68,29,37,31,229,31,229,30,147,31,241,31,241,30,90,31,118,31,27,31,29,31,148,31,148,30,121,31,121,30,142,31,57,31,115,31,157,31,241,31,230,31,199,31,91,31,166,31,104,31,127,31,86,31,144,31,228,31,228,30,23,31,210,31,88,31,198,31,40,31,189,31,189,30,32,31,119,31,77,31,137,31,159,31,142,31,84,31,135,31,99,31,99,30,14,31,14,30,14,29,107,31,163,31,238,31,125,31,224,31,76,31,21,31,90,31,99,31,88,31,229,31,10,31,166,31,166,30,215,31,21,31,224,31,133,31,53,31,48,31,48,30,243,31,198,31,70,31,70,30,101,31,194,31,226,31,46,31,86,31,158,31,118,31,59,31,241,31,241,30,63,31,63,30,63,29,138,31,184,31,129,31,239,31,166,31,225,31,75,31,75,30,93,31,93,30,215,31,225,31,113,31,70,31,244,31,179,31,201,31,9,31,187,31,180,31,176,31,77,31,158,31,158,30,166,31,245,31,46,31,181,31,184,31,246,31,246,30,101,31,183,31,183,30,210,31,209,31,209,30,243,31,21,31,36,31,33,31,234,31,22,31,22,30,162,31,227,31,119,31,166,31,30,31,238,31,24,31,24,30,75,31,196,31,110,31,110,30,110,29,125,31,116,31,73,31,73,30,83,31,24,31,234,31,147,31,41,31,41,30,19,31,19,30,24,31,106,31,41,31,91,31,91,30,242,31,138,31,165,31,179,31,28,31,148,31,225,31,136,31,136,30,136,29,83,31,228,31,35,31,35,30,35,29,114,31,208,31,21,31,26,31,26,30,233,31,66,31,66,30,194,31,59,31,5,31,58,31,83,31,48,31,108,31,141,31,227,31,101,31,219,31,45,31,199,31,173,31,100,31,187,31,120,31,139,31,214,31,58,31,58,30,67,31,171,31,248,31,55,31,175,31,253,31,188,31,8,31,173,31,170,31,170,30,110,31,64,31,32,31,188,31,195,31,195,30,224,31,133,31,243,31,76,31,76,30,18,31,18,30,187,31,154,31,215,31,67,31,22,31,255,31,235,31,235,30,235,29,124,31,124,30,63,31,63,30,68,31,31,31,127,31,127,30,218,31,171,31,171,30,72,31,72,30,45,31,72,31,144,31,98,31,5,31,185,31,185,30,63,31,221,31,151,31,79,31,174,31,35,31,240,31,175,31,154,31,96,31,45,31,125,31,88,31,250,31,2,31,2,30,164,31,119,31,226,31,160,31,160,30,18,31,255,31,44,31,44,30,121,31,184,31,56,31,7,31,158,31,11,31,107,31,56,31,33,31,185,31,71,31,210,31,188,31,188,30,33,31,160,31,128,31,8,31,213,31,213,30,116,31,124,31,124,30,56,31,164,31,24,31,115,31,115,30,199,31,136,31,215,31,213,31,207,31,204,31,255,31,139,31,98,31,63,31,28,31,59,31,150,31,179,31,131,31,254,31,58,31,125,31,148,31,220,31,203,31,44,31,24,31,142,31,142,30,65,31,121,31,174,31,155,31,155,30,141,31,40,31,191,31,191,30,243,31,33,31,23,31,23,30,137,31,28,31,17,31,238,31,191,31,175,31,175,30,235,31,125,31,85,31,85,30,83,31,255,31,255,30,208,31,208,30,96,31,162,31,145,31,145,30,124,31,124,30,240,31,165,31,165,30,219,31,7,31,7,30,120,31,120,30,120,29,85,31,222,31,255,31,163,31,201,31,201,30,127,31,20,31,11,31,52,31,60,31,59,31,171,31,223,31,223,30,223,29,113,31,212,31,25,31,235,31,143,31,71,31,12,31,213,31,110,31,224,31,224,30,39,31,9,31,29,31,10,31,156,31,130,31,162,31,162,30,116,31,104,31,234,31,179,31,179,30,179,29,168,31,51,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
