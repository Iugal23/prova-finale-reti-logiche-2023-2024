-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_643 is
end project_tb_643;

architecture project_tb_arch_643 of project_tb_643 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,11,0,163,0,32,0,85,0,43,0,0,0,0,0,43,0,101,0,207,0,0,0,39,0,199,0,124,0,125,0,11,0,46,0,0,0,100,0,181,0,141,0,46,0,0,0,113,0,235,0,9,0,209,0,0,0,164,0,157,0,0,0,78,0,238,0,175,0,71,0,158,0,122,0,133,0,3,0,60,0,200,0,0,0,97,0,0,0,164,0,67,0,0,0,11,0,182,0,105,0,52,0,221,0,26,0,106,0,9,0,171,0,9,0,53,0,33,0,192,0,134,0,173,0,166,0,109,0,224,0,53,0,121,0,21,0,105,0,224,0,181,0,159,0,163,0,83,0,69,0,155,0,0,0,215,0,162,0,242,0,0,0,0,0,51,0,0,0,0,0,224,0,0,0,135,0,0,0,117,0,101,0,191,0,0,0,247,0,90,0,147,0,143,0,219,0,98,0,180,0,217,0,0,0,147,0,182,0,10,0,0,0,160,0,0,0,235,0,209,0,167,0,159,0,232,0,155,0,77,0,0,0,0,0,166,0,0,0,231,0,0,0,178,0,241,0,16,0,0,0,161,0,174,0,0,0,0,0,201,0,231,0,243,0,237,0,0,0,184,0,247,0,100,0,110,0,233,0,125,0,82,0,226,0,216,0,79,0,202,0,118,0,130,0,32,0,15,0,175,0,190,0,139,0,126,0,80,0,152,0,0,0,181,0,130,0,94,0,85,0,0,0,116,0,0,0,202,0,0,0,12,0,239,0,207,0,0,0,97,0,0,0,0,0,0,0,0,0,112,0,22,0,0,0,156,0,12,0,186,0,203,0,0,0,38,0,68,0,0,0,0,0,218,0,119,0,0,0,27,0,0,0,16,0,149,0,244,0,64,0,199,0,239,0,17,0,2,0,148,0,86,0,95,0,47,0,96,0,120,0,0,0,67,0,0,0,80,0,232,0,180,0,225,0,218,0,44,0,127,0,0,0,217,0,145,0,200,0,188,0,200,0,83,0,117,0,13,0,189,0,5,0,242,0,0,0,0,0,192,0,208,0,6,0,29,0,0,0,0,0,160,0,50,0,167,0,225,0,142,0,211,0,228,0,0,0,191,0,26,0,121,0,0,0,15,0,44,0,0,0,0,0,60,0,33,0,49,0,151,0,0,0,0,0,188,0,76,0,185,0,166,0,23,0,215,0,47,0,119,0,229,0,0,0,55,0,0,0,93,0,160,0,225,0,1,0,248,0,211,0,103,0,233,0,153,0,144,0,180,0,204,0,121,0,59,0,199,0,1,0,154,0,127,0,241,0,159,0,48,0,43,0,181,0,234,0,20,0,188,0,185,0,185,0,18,0,46,0,154,0,90,0,0,0,50,0,0,0,183,0,132,0,187,0,152,0,114,0,12,0,1,0,173,0,0,0,142,0,81,0,0,0,181,0,152,0,208,0,91,0,0,0,128,0,24,0,140,0,0,0,170,0,39,0,0,0,0,0,22,0,69,0,205,0,0,0,80,0,0,0,0,0,0,0,169,0,67,0,192,0,156,0,124,0,0,0,187,0,0,0,139,0,9,0,0,0,222,0,199,0,101,0,202,0,119,0,108,0,100,0,0,0,0,0,187,0,98,0,81,0,52,0,0,0,101,0,167,0,166,0,0,0,185,0,172,0,118,0,150,0,70,0,0,0,123,0,240,0,43,0,207,0,45,0,111,0,0,0,169,0,41,0,131,0,0,0,61,0,22,0,62,0,0,0,233,0,40,0,221,0,6,0,0,0,166,0,45,0,250,0,0,0,21,0,206,0,69,0,247,0,242,0,0,0,154,0,176,0,223,0,180,0,0,0,198,0,134,0,72,0,78,0,3,0,0,0,224,0,3,0,204,0,112,0,244,0,24,0,65,0,0,0,0,0,38,0,7,0,229,0,203,0,137,0,19,0,0,0,77,0,94,0,49,0,145,0,24,0,202,0,106,0,0,0,100,0,61,0,38,0,3,0,101,0,20,0,205,0,14,0,39,0,27,0,114,0,117,0,127,0,102,0,97,0,113,0,101,0,240,0,117,0,0,0,248,0,124,0,0,0,131,0,71,0,98,0,47,0,252,0,0,0,167,0,241,0,28,0,142,0,0,0,186,0,81,0,226,0,88,0,204,0,207,0,0,0,119,0,213,0,218,0,241,0,84,0,105,0,41,0,3,0,35,0,226,0,144,0,73,0,84,0,87,0,195,0,0,0,0,0,104,0,190,0,240,0,105,0,245,0,20,0,31,0,65,0,0,0,239,0,136,0,0,0,0,0,236,0,0,0,122,0,150,0,10,0,53,0,0,0,0,0,17,0,111,0,182,0,107,0,3,0,184,0,189,0,204,0,192,0,0,0,255,0,101,0,195,0,71,0,0,0,202,0,0,0,221,0,244,0,0,0,196,0,28,0,25,0,135,0,42,0,0,0,135,0,0,0,0,0,213,0,247,0,67,0,0,0,0,0,0,0,158,0,137,0,37,0,222,0,111,0,102,0,100,0,43,0,216,0,12,0,15,0,122,0,7,0,71,0,0,0,159,0,0,0,0,0,138,0,100,0,23,0,0,0,185,0,205,0,62,0,17,0,205,0,115,0,223,0,125,0,150,0,112,0,66,0,40,0,218,0,70,0,93,0,229,0,241,0,220,0,189,0,142,0,21,0,48,0,0,0,0,0,96,0,0,0,252,0,217,0,142,0,200,0,0,0,255,0,169,0,0,0,85,0,136,0,219,0,74,0,134,0,0,0,0,0,54,0,100,0,99,0,0,0,163,0,45,0,149,0,134,0,141,0,42,0,96,0,137,0,199,0,181,0,255,0,241,0,252,0,105,0,30,0,0,0,81,0,206,0,72,0,12,0,185,0,147,0,71,0,61,0,0,0,81,0,208,0,0,0,183,0,150,0,246,0,44,0,160,0,45,0,51,0,170,0,59,0,13,0,0,0,249,0,128,0,27,0,3,0,26,0,91,0,71,0,27,0,144,0,116,0,160,0,152,0,0,0,242,0,234,0,0,0,43,0,157,0,224,0,9,0,182,0,40,0,23,0,109,0,157,0,151,0,214,0,131,0,59,0,38,0,0,0,220,0,246,0,145,0,55,0,169,0,204,0,149,0,251,0,235,0,225,0,214,0,251,0,0,0,203,0,0,0,77,0,228,0,183,0,0,0,85,0,142,0,0,0,147,0,0,0,0,0,207,0,51,0,10,0,99,0,151,0,0,0,0,0,114,0,188,0,123,0,204,0,0,0,33,0,0,0,118,0,154,0,64,0,240,0,122,0,122,0,0,0,24,0,11,0,213,0,0,0,86,0,123,0,81,0,143,0,87,0,0,0,89,0,0,0,133,0,0,0,187,0,39,0,117,0,68,0,199,0,219,0,154,0,223,0,3,0,121,0,101,0,203,0,253,0,219,0,110,0,19,0,122,0,245,0,221,0,108,0,0,0,181,0,16,0,0,0,1,0,115,0,0,0,244,0,73,0,70,0,39,0,154,0,165,0,204,0,144,0,0,0,245,0,94,0,225,0,196,0,131,0,206,0,241,0,237,0,231,0,163,0,134,0,170,0,86,0,89,0,0,0,3,0,112,0,58,0,11,0,136,0,22,0,119,0,201,0,202,0,201,0,105,0,0,0,212,0,0,0,52,0,41,0,0,0,55,0,3,0,0,0,158,0,141,0,0,0,171,0,0,0,165,0,56,0,85,0,75,0,87,0,32,0,74,0,218,0,85,0,69,0,181,0,218,0,103,0,0,0,80,0,0,0,89,0,248,0,172,0,252,0,138,0,0,0,139,0,121,0,59,0,164,0,126,0,89,0,38,0,74,0,187,0,133,0);
signal scenario_full  : scenario_type := (245,31,11,31,163,31,32,31,85,31,43,31,43,30,43,29,43,31,101,31,207,31,207,30,39,31,199,31,124,31,125,31,11,31,46,31,46,30,100,31,181,31,141,31,46,31,46,30,113,31,235,31,9,31,209,31,209,30,164,31,157,31,157,30,78,31,238,31,175,31,71,31,158,31,122,31,133,31,3,31,60,31,200,31,200,30,97,31,97,30,164,31,67,31,67,30,11,31,182,31,105,31,52,31,221,31,26,31,106,31,9,31,171,31,9,31,53,31,33,31,192,31,134,31,173,31,166,31,109,31,224,31,53,31,121,31,21,31,105,31,224,31,181,31,159,31,163,31,83,31,69,31,155,31,155,30,215,31,162,31,242,31,242,30,242,29,51,31,51,30,51,29,224,31,224,30,135,31,135,30,117,31,101,31,191,31,191,30,247,31,90,31,147,31,143,31,219,31,98,31,180,31,217,31,217,30,147,31,182,31,10,31,10,30,160,31,160,30,235,31,209,31,167,31,159,31,232,31,155,31,77,31,77,30,77,29,166,31,166,30,231,31,231,30,178,31,241,31,16,31,16,30,161,31,174,31,174,30,174,29,201,31,231,31,243,31,237,31,237,30,184,31,247,31,100,31,110,31,233,31,125,31,82,31,226,31,216,31,79,31,202,31,118,31,130,31,32,31,15,31,175,31,190,31,139,31,126,31,80,31,152,31,152,30,181,31,130,31,94,31,85,31,85,30,116,31,116,30,202,31,202,30,12,31,239,31,207,31,207,30,97,31,97,30,97,29,97,28,97,27,112,31,22,31,22,30,156,31,12,31,186,31,203,31,203,30,38,31,68,31,68,30,68,29,218,31,119,31,119,30,27,31,27,30,16,31,149,31,244,31,64,31,199,31,239,31,17,31,2,31,148,31,86,31,95,31,47,31,96,31,120,31,120,30,67,31,67,30,80,31,232,31,180,31,225,31,218,31,44,31,127,31,127,30,217,31,145,31,200,31,188,31,200,31,83,31,117,31,13,31,189,31,5,31,242,31,242,30,242,29,192,31,208,31,6,31,29,31,29,30,29,29,160,31,50,31,167,31,225,31,142,31,211,31,228,31,228,30,191,31,26,31,121,31,121,30,15,31,44,31,44,30,44,29,60,31,33,31,49,31,151,31,151,30,151,29,188,31,76,31,185,31,166,31,23,31,215,31,47,31,119,31,229,31,229,30,55,31,55,30,93,31,160,31,225,31,1,31,248,31,211,31,103,31,233,31,153,31,144,31,180,31,204,31,121,31,59,31,199,31,1,31,154,31,127,31,241,31,159,31,48,31,43,31,181,31,234,31,20,31,188,31,185,31,185,31,18,31,46,31,154,31,90,31,90,30,50,31,50,30,183,31,132,31,187,31,152,31,114,31,12,31,1,31,173,31,173,30,142,31,81,31,81,30,181,31,152,31,208,31,91,31,91,30,128,31,24,31,140,31,140,30,170,31,39,31,39,30,39,29,22,31,69,31,205,31,205,30,80,31,80,30,80,29,80,28,169,31,67,31,192,31,156,31,124,31,124,30,187,31,187,30,139,31,9,31,9,30,222,31,199,31,101,31,202,31,119,31,108,31,100,31,100,30,100,29,187,31,98,31,81,31,52,31,52,30,101,31,167,31,166,31,166,30,185,31,172,31,118,31,150,31,70,31,70,30,123,31,240,31,43,31,207,31,45,31,111,31,111,30,169,31,41,31,131,31,131,30,61,31,22,31,62,31,62,30,233,31,40,31,221,31,6,31,6,30,166,31,45,31,250,31,250,30,21,31,206,31,69,31,247,31,242,31,242,30,154,31,176,31,223,31,180,31,180,30,198,31,134,31,72,31,78,31,3,31,3,30,224,31,3,31,204,31,112,31,244,31,24,31,65,31,65,30,65,29,38,31,7,31,229,31,203,31,137,31,19,31,19,30,77,31,94,31,49,31,145,31,24,31,202,31,106,31,106,30,100,31,61,31,38,31,3,31,101,31,20,31,205,31,14,31,39,31,27,31,114,31,117,31,127,31,102,31,97,31,113,31,101,31,240,31,117,31,117,30,248,31,124,31,124,30,131,31,71,31,98,31,47,31,252,31,252,30,167,31,241,31,28,31,142,31,142,30,186,31,81,31,226,31,88,31,204,31,207,31,207,30,119,31,213,31,218,31,241,31,84,31,105,31,41,31,3,31,35,31,226,31,144,31,73,31,84,31,87,31,195,31,195,30,195,29,104,31,190,31,240,31,105,31,245,31,20,31,31,31,65,31,65,30,239,31,136,31,136,30,136,29,236,31,236,30,122,31,150,31,10,31,53,31,53,30,53,29,17,31,111,31,182,31,107,31,3,31,184,31,189,31,204,31,192,31,192,30,255,31,101,31,195,31,71,31,71,30,202,31,202,30,221,31,244,31,244,30,196,31,28,31,25,31,135,31,42,31,42,30,135,31,135,30,135,29,213,31,247,31,67,31,67,30,67,29,67,28,158,31,137,31,37,31,222,31,111,31,102,31,100,31,43,31,216,31,12,31,15,31,122,31,7,31,71,31,71,30,159,31,159,30,159,29,138,31,100,31,23,31,23,30,185,31,205,31,62,31,17,31,205,31,115,31,223,31,125,31,150,31,112,31,66,31,40,31,218,31,70,31,93,31,229,31,241,31,220,31,189,31,142,31,21,31,48,31,48,30,48,29,96,31,96,30,252,31,217,31,142,31,200,31,200,30,255,31,169,31,169,30,85,31,136,31,219,31,74,31,134,31,134,30,134,29,54,31,100,31,99,31,99,30,163,31,45,31,149,31,134,31,141,31,42,31,96,31,137,31,199,31,181,31,255,31,241,31,252,31,105,31,30,31,30,30,81,31,206,31,72,31,12,31,185,31,147,31,71,31,61,31,61,30,81,31,208,31,208,30,183,31,150,31,246,31,44,31,160,31,45,31,51,31,170,31,59,31,13,31,13,30,249,31,128,31,27,31,3,31,26,31,91,31,71,31,27,31,144,31,116,31,160,31,152,31,152,30,242,31,234,31,234,30,43,31,157,31,224,31,9,31,182,31,40,31,23,31,109,31,157,31,151,31,214,31,131,31,59,31,38,31,38,30,220,31,246,31,145,31,55,31,169,31,204,31,149,31,251,31,235,31,225,31,214,31,251,31,251,30,203,31,203,30,77,31,228,31,183,31,183,30,85,31,142,31,142,30,147,31,147,30,147,29,207,31,51,31,10,31,99,31,151,31,151,30,151,29,114,31,188,31,123,31,204,31,204,30,33,31,33,30,118,31,154,31,64,31,240,31,122,31,122,31,122,30,24,31,11,31,213,31,213,30,86,31,123,31,81,31,143,31,87,31,87,30,89,31,89,30,133,31,133,30,187,31,39,31,117,31,68,31,199,31,219,31,154,31,223,31,3,31,121,31,101,31,203,31,253,31,219,31,110,31,19,31,122,31,245,31,221,31,108,31,108,30,181,31,16,31,16,30,1,31,115,31,115,30,244,31,73,31,70,31,39,31,154,31,165,31,204,31,144,31,144,30,245,31,94,31,225,31,196,31,131,31,206,31,241,31,237,31,231,31,163,31,134,31,170,31,86,31,89,31,89,30,3,31,112,31,58,31,11,31,136,31,22,31,119,31,201,31,202,31,201,31,105,31,105,30,212,31,212,30,52,31,41,31,41,30,55,31,3,31,3,30,158,31,141,31,141,30,171,31,171,30,165,31,56,31,85,31,75,31,87,31,32,31,74,31,218,31,85,31,69,31,181,31,218,31,103,31,103,30,80,31,80,30,89,31,248,31,172,31,252,31,138,31,138,30,139,31,121,31,59,31,164,31,126,31,89,31,38,31,74,31,187,31,133,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
