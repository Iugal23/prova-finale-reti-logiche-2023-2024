-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_306 is
end project_tb_306;

architecture project_tb_arch_306 of project_tb_306 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 987;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (203,0,202,0,56,0,189,0,95,0,0,0,41,0,221,0,225,0,128,0,0,0,0,0,167,0,177,0,234,0,75,0,146,0,0,0,50,0,0,0,139,0,0,0,0,0,185,0,28,0,90,0,24,0,0,0,229,0,155,0,181,0,82,0,188,0,135,0,224,0,78,0,14,0,168,0,172,0,105,0,0,0,240,0,168,0,0,0,248,0,111,0,191,0,0,0,164,0,88,0,247,0,74,0,56,0,21,0,19,0,0,0,187,0,89,0,0,0,128,0,98,0,116,0,192,0,0,0,109,0,0,0,233,0,0,0,30,0,245,0,251,0,47,0,0,0,35,0,221,0,128,0,200,0,124,0,0,0,0,0,0,0,139,0,1,0,98,0,163,0,131,0,224,0,0,0,0,0,162,0,164,0,51,0,0,0,114,0,159,0,28,0,212,0,121,0,192,0,230,0,0,0,131,0,29,0,73,0,44,0,191,0,63,0,62,0,71,0,160,0,0,0,32,0,0,0,0,0,173,0,211,0,1,0,0,0,38,0,0,0,183,0,251,0,155,0,65,0,0,0,227,0,0,0,0,0,0,0,235,0,171,0,54,0,3,0,0,0,213,0,20,0,27,0,151,0,193,0,83,0,0,0,77,0,254,0,237,0,226,0,178,0,0,0,128,0,246,0,131,0,248,0,35,0,0,0,169,0,97,0,16,0,165,0,0,0,81,0,171,0,123,0,103,0,237,0,222,0,66,0,131,0,37,0,253,0,246,0,168,0,215,0,242,0,0,0,80,0,0,0,0,0,236,0,57,0,64,0,186,0,122,0,0,0,240,0,110,0,228,0,136,0,0,0,0,0,230,0,93,0,145,0,3,0,137,0,0,0,68,0,63,0,16,0,1,0,182,0,133,0,239,0,198,0,202,0,218,0,145,0,0,0,122,0,138,0,0,0,0,0,52,0,0,0,175,0,0,0,249,0,176,0,113,0,0,0,0,0,39,0,132,0,87,0,41,0,43,0,66,0,166,0,187,0,84,0,146,0,215,0,181,0,136,0,0,0,0,0,62,0,124,0,14,0,63,0,217,0,106,0,50,0,2,0,189,0,248,0,59,0,28,0,4,0,67,0,123,0,135,0,0,0,42,0,0,0,163,0,213,0,121,0,139,0,152,0,0,0,58,0,175,0,163,0,0,0,239,0,98,0,219,0,94,0,0,0,6,0,207,0,76,0,0,0,247,0,5,0,11,0,226,0,166,0,77,0,0,0,32,0,44,0,1,0,17,0,195,0,225,0,95,0,214,0,107,0,53,0,122,0,43,0,165,0,49,0,64,0,37,0,85,0,241,0,42,0,77,0,140,0,115,0,15,0,93,0,0,0,165,0,251,0,136,0,0,0,230,0,187,0,0,0,178,0,11,0,145,0,86,0,16,0,80,0,60,0,0,0,145,0,203,0,136,0,0,0,147,0,0,0,169,0,0,0,10,0,0,0,0,0,16,0,96,0,103,0,0,0,38,0,159,0,57,0,21,0,0,0,184,0,59,0,207,0,0,0,229,0,23,0,117,0,0,0,0,0,223,0,41,0,170,0,185,0,89,0,251,0,222,0,0,0,139,0,118,0,180,0,147,0,27,0,0,0,105,0,101,0,170,0,244,0,250,0,0,0,116,0,83,0,160,0,131,0,247,0,142,0,171,0,28,0,90,0,20,0,39,0,0,0,54,0,14,0,62,0,72,0,186,0,156,0,16,0,211,0,0,0,6,0,132,0,5,0,124,0,136,0,96,0,57,0,225,0,94,0,234,0,156,0,216,0,23,0,255,0,116,0,84,0,0,0,25,0,126,0,42,0,32,0,139,0,8,0,0,0,131,0,120,0,143,0,0,0,32,0,33,0,182,0,134,0,15,0,65,0,93,0,0,0,237,0,225,0,192,0,174,0,0,0,198,0,30,0,21,0,0,0,0,0,0,0,0,0,0,0,178,0,160,0,0,0,112,0,62,0,89,0,251,0,201,0,165,0,244,0,228,0,72,0,87,0,218,0,0,0,124,0,198,0,0,0,175,0,35,0,231,0,48,0,46,0,224,0,113,0,102,0,101,0,163,0,92,0,195,0,60,0,191,0,47,0,59,0,212,0,190,0,0,0,140,0,0,0,11,0,77,0,185,0,0,0,42,0,195,0,68,0,124,0,141,0,0,0,99,0,84,0,10,0,219,0,103,0,161,0,16,0,94,0,113,0,8,0,112,0,227,0,211,0,51,0,0,0,90,0,210,0,0,0,0,0,81,0,12,0,189,0,23,0,232,0,141,0,104,0,0,0,0,0,0,0,0,0,0,0,0,0,78,0,109,0,107,0,0,0,181,0,43,0,96,0,0,0,211,0,189,0,57,0,0,0,104,0,184,0,237,0,83,0,0,0,132,0,0,0,110,0,207,0,238,0,183,0,100,0,68,0,94,0,211,0,228,0,124,0,253,0,53,0,0,0,77,0,143,0,0,0,84,0,215,0,23,0,176,0,64,0,75,0,130,0,5,0,215,0,186,0,136,0,0,0,124,0,149,0,30,0,203,0,222,0,8,0,224,0,79,0,0,0,14,0,9,0,69,0,14,0,236,0,104,0,168,0,0,0,180,0,171,0,247,0,0,0,111,0,167,0,34,0,251,0,234,0,119,0,0,0,173,0,195,0,134,0,0,0,0,0,211,0,169,0,116,0,69,0,43,0,0,0,28,0,0,0,30,0,79,0,245,0,249,0,0,0,0,0,211,0,0,0,0,0,0,0,28,0,59,0,204,0,0,0,80,0,73,0,185,0,0,0,234,0,137,0,0,0,0,0,0,0,205,0,47,0,169,0,251,0,0,0,196,0,90,0,126,0,103,0,61,0,0,0,100,0,48,0,203,0,0,0,144,0,93,0,0,0,0,0,90,0,89,0,157,0,119,0,83,0,0,0,215,0,142,0,155,0,5,0,97,0,203,0,0,0,0,0,81,0,117,0,106,0,108,0,0,0,161,0,0,0,159,0,186,0,116,0,161,0,87,0,116,0,244,0,12,0,236,0,159,0,0,0,125,0,0,0,14,0,245,0,63,0,0,0,154,0,0,0,201,0,218,0,214,0,0,0,130,0,0,0,0,0,0,0,61,0,0,0,220,0,68,0,192,0,14,0,58,0,239,0,26,0,210,0,0,0,0,0,0,0,136,0,63,0,62,0,0,0,174,0,40,0,152,0,0,0,208,0,69,0,255,0,215,0,26,0,13,0,112,0,0,0,168,0,96,0,239,0,225,0,0,0,67,0,200,0,94,0,0,0,70,0,252,0,46,0,0,0,227,0,116,0,14,0,157,0,173,0,70,0,180,0,0,0,0,0,24,0,220,0,0,0,232,0,42,0,147,0,116,0,115,0,200,0,69,0,0,0,178,0,194,0,219,0,255,0,0,0,220,0,0,0,125,0,174,0,57,0,202,0,37,0,65,0,209,0,180,0,255,0,0,0,0,0,116,0,0,0,13,0,21,0,239,0,0,0,63,0,0,0,0,0,95,0,0,0,72,0,225,0,52,0,70,0,85,0,0,0,168,0,40,0,0,0,251,0,76,0,16,0,185,0,253,0,249,0,255,0,133,0,85,0,130,0,25,0,79,0,136,0,56,0,19,0,118,0,0,0,34,0,85,0,113,0,26,0,14,0,66,0,32,0,130,0,187,0,0,0,109,0,176,0,0,0,185,0,177,0,100,0,215,0,171,0,139,0,0,0,237,0,99,0,155,0,172,0,41,0,228,0,0,0,71,0,49,0,137,0,153,0,30,0,37,0,117,0,217,0,252,0,139,0,58,0,0,0,238,0,184,0,50,0,116,0,39,0,224,0,147,0,114,0,160,0,70,0,72,0,15,0,0,0,0,0,253,0,171,0,9,0,113,0,0,0,250,0,0,0,164,0,0,0,12,0,152,0,72,0,170,0,82,0,43,0,0,0,239,0,53,0,96,0,0,0,242,0,161,0,231,0,0,0,0,0,0,0,92,0,0,0,129,0,102,0,131,0,206,0,222,0,142,0,202,0,0,0,230,0,201,0,205,0,0,0,0,0,58,0,210,0,224,0,50,0,226,0,233,0,214,0,118,0,0,0,49,0,191,0,0,0,0,0,230,0,204,0,44,0,90,0,150,0,0,0,150,0,3,0,0,0,52,0,155,0,176,0,61,0,99,0,75,0,208,0,35,0,0,0,204,0,247,0,241,0,11,0,88,0,201,0,112,0,201,0,131,0,135,0,187,0,134,0,82,0,102,0,55,0,162,0,0,0,24,0,218,0,54,0,112,0,0,0,231,0,249,0,68,0,76,0,27,0,70,0,93,0,149,0,0,0,156,0,233,0,0,0,151,0,228,0,3,0,254,0,71,0,91,0,6,0,242,0,0,0,108,0,151,0,1,0,202,0,0,0);
signal scenario_full  : scenario_type := (203,31,202,31,56,31,189,31,95,31,95,30,41,31,221,31,225,31,128,31,128,30,128,29,167,31,177,31,234,31,75,31,146,31,146,30,50,31,50,30,139,31,139,30,139,29,185,31,28,31,90,31,24,31,24,30,229,31,155,31,181,31,82,31,188,31,135,31,224,31,78,31,14,31,168,31,172,31,105,31,105,30,240,31,168,31,168,30,248,31,111,31,191,31,191,30,164,31,88,31,247,31,74,31,56,31,21,31,19,31,19,30,187,31,89,31,89,30,128,31,98,31,116,31,192,31,192,30,109,31,109,30,233,31,233,30,30,31,245,31,251,31,47,31,47,30,35,31,221,31,128,31,200,31,124,31,124,30,124,29,124,28,139,31,1,31,98,31,163,31,131,31,224,31,224,30,224,29,162,31,164,31,51,31,51,30,114,31,159,31,28,31,212,31,121,31,192,31,230,31,230,30,131,31,29,31,73,31,44,31,191,31,63,31,62,31,71,31,160,31,160,30,32,31,32,30,32,29,173,31,211,31,1,31,1,30,38,31,38,30,183,31,251,31,155,31,65,31,65,30,227,31,227,30,227,29,227,28,235,31,171,31,54,31,3,31,3,30,213,31,20,31,27,31,151,31,193,31,83,31,83,30,77,31,254,31,237,31,226,31,178,31,178,30,128,31,246,31,131,31,248,31,35,31,35,30,169,31,97,31,16,31,165,31,165,30,81,31,171,31,123,31,103,31,237,31,222,31,66,31,131,31,37,31,253,31,246,31,168,31,215,31,242,31,242,30,80,31,80,30,80,29,236,31,57,31,64,31,186,31,122,31,122,30,240,31,110,31,228,31,136,31,136,30,136,29,230,31,93,31,145,31,3,31,137,31,137,30,68,31,63,31,16,31,1,31,182,31,133,31,239,31,198,31,202,31,218,31,145,31,145,30,122,31,138,31,138,30,138,29,52,31,52,30,175,31,175,30,249,31,176,31,113,31,113,30,113,29,39,31,132,31,87,31,41,31,43,31,66,31,166,31,187,31,84,31,146,31,215,31,181,31,136,31,136,30,136,29,62,31,124,31,14,31,63,31,217,31,106,31,50,31,2,31,189,31,248,31,59,31,28,31,4,31,67,31,123,31,135,31,135,30,42,31,42,30,163,31,213,31,121,31,139,31,152,31,152,30,58,31,175,31,163,31,163,30,239,31,98,31,219,31,94,31,94,30,6,31,207,31,76,31,76,30,247,31,5,31,11,31,226,31,166,31,77,31,77,30,32,31,44,31,1,31,17,31,195,31,225,31,95,31,214,31,107,31,53,31,122,31,43,31,165,31,49,31,64,31,37,31,85,31,241,31,42,31,77,31,140,31,115,31,15,31,93,31,93,30,165,31,251,31,136,31,136,30,230,31,187,31,187,30,178,31,11,31,145,31,86,31,16,31,80,31,60,31,60,30,145,31,203,31,136,31,136,30,147,31,147,30,169,31,169,30,10,31,10,30,10,29,16,31,96,31,103,31,103,30,38,31,159,31,57,31,21,31,21,30,184,31,59,31,207,31,207,30,229,31,23,31,117,31,117,30,117,29,223,31,41,31,170,31,185,31,89,31,251,31,222,31,222,30,139,31,118,31,180,31,147,31,27,31,27,30,105,31,101,31,170,31,244,31,250,31,250,30,116,31,83,31,160,31,131,31,247,31,142,31,171,31,28,31,90,31,20,31,39,31,39,30,54,31,14,31,62,31,72,31,186,31,156,31,16,31,211,31,211,30,6,31,132,31,5,31,124,31,136,31,96,31,57,31,225,31,94,31,234,31,156,31,216,31,23,31,255,31,116,31,84,31,84,30,25,31,126,31,42,31,32,31,139,31,8,31,8,30,131,31,120,31,143,31,143,30,32,31,33,31,182,31,134,31,15,31,65,31,93,31,93,30,237,31,225,31,192,31,174,31,174,30,198,31,30,31,21,31,21,30,21,29,21,28,21,27,21,26,178,31,160,31,160,30,112,31,62,31,89,31,251,31,201,31,165,31,244,31,228,31,72,31,87,31,218,31,218,30,124,31,198,31,198,30,175,31,35,31,231,31,48,31,46,31,224,31,113,31,102,31,101,31,163,31,92,31,195,31,60,31,191,31,47,31,59,31,212,31,190,31,190,30,140,31,140,30,11,31,77,31,185,31,185,30,42,31,195,31,68,31,124,31,141,31,141,30,99,31,84,31,10,31,219,31,103,31,161,31,16,31,94,31,113,31,8,31,112,31,227,31,211,31,51,31,51,30,90,31,210,31,210,30,210,29,81,31,12,31,189,31,23,31,232,31,141,31,104,31,104,30,104,29,104,28,104,27,104,26,104,25,78,31,109,31,107,31,107,30,181,31,43,31,96,31,96,30,211,31,189,31,57,31,57,30,104,31,184,31,237,31,83,31,83,30,132,31,132,30,110,31,207,31,238,31,183,31,100,31,68,31,94,31,211,31,228,31,124,31,253,31,53,31,53,30,77,31,143,31,143,30,84,31,215,31,23,31,176,31,64,31,75,31,130,31,5,31,215,31,186,31,136,31,136,30,124,31,149,31,30,31,203,31,222,31,8,31,224,31,79,31,79,30,14,31,9,31,69,31,14,31,236,31,104,31,168,31,168,30,180,31,171,31,247,31,247,30,111,31,167,31,34,31,251,31,234,31,119,31,119,30,173,31,195,31,134,31,134,30,134,29,211,31,169,31,116,31,69,31,43,31,43,30,28,31,28,30,30,31,79,31,245,31,249,31,249,30,249,29,211,31,211,30,211,29,211,28,28,31,59,31,204,31,204,30,80,31,73,31,185,31,185,30,234,31,137,31,137,30,137,29,137,28,205,31,47,31,169,31,251,31,251,30,196,31,90,31,126,31,103,31,61,31,61,30,100,31,48,31,203,31,203,30,144,31,93,31,93,30,93,29,90,31,89,31,157,31,119,31,83,31,83,30,215,31,142,31,155,31,5,31,97,31,203,31,203,30,203,29,81,31,117,31,106,31,108,31,108,30,161,31,161,30,159,31,186,31,116,31,161,31,87,31,116,31,244,31,12,31,236,31,159,31,159,30,125,31,125,30,14,31,245,31,63,31,63,30,154,31,154,30,201,31,218,31,214,31,214,30,130,31,130,30,130,29,130,28,61,31,61,30,220,31,68,31,192,31,14,31,58,31,239,31,26,31,210,31,210,30,210,29,210,28,136,31,63,31,62,31,62,30,174,31,40,31,152,31,152,30,208,31,69,31,255,31,215,31,26,31,13,31,112,31,112,30,168,31,96,31,239,31,225,31,225,30,67,31,200,31,94,31,94,30,70,31,252,31,46,31,46,30,227,31,116,31,14,31,157,31,173,31,70,31,180,31,180,30,180,29,24,31,220,31,220,30,232,31,42,31,147,31,116,31,115,31,200,31,69,31,69,30,178,31,194,31,219,31,255,31,255,30,220,31,220,30,125,31,174,31,57,31,202,31,37,31,65,31,209,31,180,31,255,31,255,30,255,29,116,31,116,30,13,31,21,31,239,31,239,30,63,31,63,30,63,29,95,31,95,30,72,31,225,31,52,31,70,31,85,31,85,30,168,31,40,31,40,30,251,31,76,31,16,31,185,31,253,31,249,31,255,31,133,31,85,31,130,31,25,31,79,31,136,31,56,31,19,31,118,31,118,30,34,31,85,31,113,31,26,31,14,31,66,31,32,31,130,31,187,31,187,30,109,31,176,31,176,30,185,31,177,31,100,31,215,31,171,31,139,31,139,30,237,31,99,31,155,31,172,31,41,31,228,31,228,30,71,31,49,31,137,31,153,31,30,31,37,31,117,31,217,31,252,31,139,31,58,31,58,30,238,31,184,31,50,31,116,31,39,31,224,31,147,31,114,31,160,31,70,31,72,31,15,31,15,30,15,29,253,31,171,31,9,31,113,31,113,30,250,31,250,30,164,31,164,30,12,31,152,31,72,31,170,31,82,31,43,31,43,30,239,31,53,31,96,31,96,30,242,31,161,31,231,31,231,30,231,29,231,28,92,31,92,30,129,31,102,31,131,31,206,31,222,31,142,31,202,31,202,30,230,31,201,31,205,31,205,30,205,29,58,31,210,31,224,31,50,31,226,31,233,31,214,31,118,31,118,30,49,31,191,31,191,30,191,29,230,31,204,31,44,31,90,31,150,31,150,30,150,31,3,31,3,30,52,31,155,31,176,31,61,31,99,31,75,31,208,31,35,31,35,30,204,31,247,31,241,31,11,31,88,31,201,31,112,31,201,31,131,31,135,31,187,31,134,31,82,31,102,31,55,31,162,31,162,30,24,31,218,31,54,31,112,31,112,30,231,31,249,31,68,31,76,31,27,31,70,31,93,31,149,31,149,30,156,31,233,31,233,30,151,31,228,31,3,31,254,31,71,31,91,31,6,31,242,31,242,30,108,31,151,31,1,31,202,31,202,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
