-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 287;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (143,0,10,0,121,0,132,0,0,0,97,0,161,0,105,0,245,0,229,0,236,0,18,0,5,0,0,0,50,0,14,0,23,0,0,0,78,0,119,0,223,0,161,0,233,0,10,0,102,0,107,0,0,0,254,0,25,0,62,0,61,0,237,0,113,0,232,0,168,0,239,0,0,0,176,0,56,0,72,0,41,0,57,0,232,0,205,0,0,0,128,0,0,0,31,0,162,0,137,0,48,0,208,0,239,0,93,0,177,0,199,0,0,0,0,0,200,0,0,0,70,0,17,0,246,0,78,0,0,0,57,0,114,0,0,0,0,0,109,0,58,0,238,0,0,0,230,0,63,0,226,0,0,0,46,0,214,0,111,0,249,0,0,0,10,0,153,0,17,0,137,0,19,0,1,0,0,0,200,0,0,0,0,0,0,0,108,0,186,0,64,0,0,0,0,0,31,0,55,0,205,0,165,0,145,0,115,0,181,0,57,0,0,0,126,0,0,0,221,0,237,0,241,0,0,0,158,0,1,0,108,0,43,0,14,0,156,0,139,0,183,0,0,0,17,0,0,0,246,0,18,0,172,0,148,0,132,0,253,0,171,0,211,0,0,0,207,0,142,0,138,0,222,0,204,0,0,0,170,0,216,0,212,0,38,0,99,0,168,0,53,0,178,0,43,0,115,0,204,0,253,0,63,0,255,0,115,0,196,0,0,0,14,0,156,0,0,0,132,0,185,0,0,0,0,0,13,0,67,0,155,0,5,0,251,0,114,0,0,0,243,0,1,0,0,0,96,0,228,0,58,0,109,0,1,0,0,0,86,0,178,0,113,0,248,0,43,0,94,0,238,0,0,0,0,0,216,0,0,0,226,0,231,0,0,0,195,0,191,0,189,0,46,0,216,0,136,0,55,0,8,0,251,0,223,0,229,0,187,0,113,0,0,0,39,0,0,0,0,0,139,0,143,0,13,0,202,0,0,0,157,0,190,0,90,0,132,0,0,0,230,0,204,0,150,0,226,0,0,0,49,0,101,0,198,0,32,0,69,0,208,0,63,0,254,0,136,0,67,0,223,0,0,0,76,0,138,0,0,0,223,0,211,0,0,0,255,0,151,0,0,0,215,0,87,0,144,0,0,0,0,0,137,0,0,0,46,0,251,0,84,0,221,0,234,0,215,0,160,0,15,0,252,0,245,0,176,0,227,0,16,0,150,0,168,0,23,0,25,0,136,0,53,0,45,0,87,0,227,0,0,0,75,0,149,0,157,0,99,0,92,0,225,0,0,0,135,0,0,0,229,0,58,0);
signal scenario_full  : scenario_type := (143,31,10,31,121,31,132,31,132,30,97,31,161,31,105,31,245,31,229,31,236,31,18,31,5,31,5,30,50,31,14,31,23,31,23,30,78,31,119,31,223,31,161,31,233,31,10,31,102,31,107,31,107,30,254,31,25,31,62,31,61,31,237,31,113,31,232,31,168,31,239,31,239,30,176,31,56,31,72,31,41,31,57,31,232,31,205,31,205,30,128,31,128,30,31,31,162,31,137,31,48,31,208,31,239,31,93,31,177,31,199,31,199,30,199,29,200,31,200,30,70,31,17,31,246,31,78,31,78,30,57,31,114,31,114,30,114,29,109,31,58,31,238,31,238,30,230,31,63,31,226,31,226,30,46,31,214,31,111,31,249,31,249,30,10,31,153,31,17,31,137,31,19,31,1,31,1,30,200,31,200,30,200,29,200,28,108,31,186,31,64,31,64,30,64,29,31,31,55,31,205,31,165,31,145,31,115,31,181,31,57,31,57,30,126,31,126,30,221,31,237,31,241,31,241,30,158,31,1,31,108,31,43,31,14,31,156,31,139,31,183,31,183,30,17,31,17,30,246,31,18,31,172,31,148,31,132,31,253,31,171,31,211,31,211,30,207,31,142,31,138,31,222,31,204,31,204,30,170,31,216,31,212,31,38,31,99,31,168,31,53,31,178,31,43,31,115,31,204,31,253,31,63,31,255,31,115,31,196,31,196,30,14,31,156,31,156,30,132,31,185,31,185,30,185,29,13,31,67,31,155,31,5,31,251,31,114,31,114,30,243,31,1,31,1,30,96,31,228,31,58,31,109,31,1,31,1,30,86,31,178,31,113,31,248,31,43,31,94,31,238,31,238,30,238,29,216,31,216,30,226,31,231,31,231,30,195,31,191,31,189,31,46,31,216,31,136,31,55,31,8,31,251,31,223,31,229,31,187,31,113,31,113,30,39,31,39,30,39,29,139,31,143,31,13,31,202,31,202,30,157,31,190,31,90,31,132,31,132,30,230,31,204,31,150,31,226,31,226,30,49,31,101,31,198,31,32,31,69,31,208,31,63,31,254,31,136,31,67,31,223,31,223,30,76,31,138,31,138,30,223,31,211,31,211,30,255,31,151,31,151,30,215,31,87,31,144,31,144,30,144,29,137,31,137,30,46,31,251,31,84,31,221,31,234,31,215,31,160,31,15,31,252,31,245,31,176,31,227,31,16,31,150,31,168,31,23,31,25,31,136,31,53,31,45,31,87,31,227,31,227,30,75,31,149,31,157,31,99,31,92,31,225,31,225,30,135,31,135,30,229,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
