-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_465 is
end project_tb_465;

architecture project_tb_arch_465 of project_tb_465 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 156;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (11,0,157,0,0,0,251,0,112,0,0,0,23,0,155,0,121,0,204,0,40,0,0,0,130,0,140,0,15,0,213,0,57,0,81,0,206,0,0,0,180,0,0,0,85,0,22,0,0,0,70,0,0,0,229,0,144,0,0,0,51,0,93,0,241,0,211,0,252,0,4,0,35,0,36,0,3,0,105,0,0,0,45,0,31,0,247,0,211,0,229,0,162,0,208,0,152,0,205,0,120,0,0,0,83,0,15,0,40,0,234,0,190,0,69,0,240,0,125,0,7,0,0,0,163,0,39,0,0,0,209,0,48,0,0,0,0,0,178,0,0,0,184,0,101,0,6,0,224,0,179,0,0,0,0,0,0,0,164,0,70,0,72,0,0,0,3,0,221,0,82,0,240,0,136,0,247,0,163,0,231,0,247,0,7,0,56,0,2,0,0,0,64,0,247,0,0,0,213,0,0,0,67,0,101,0,203,0,61,0,0,0,16,0,142,0,251,0,0,0,117,0,7,0,210,0,210,0,14,0,84,0,100,0,0,0,99,0,0,0,33,0,223,0,89,0,17,0,52,0,169,0,212,0,0,0,103,0,105,0,145,0,20,0,73,0,88,0,0,0,0,0,231,0,4,0,60,0,243,0,9,0,145,0,114,0,158,0,205,0,38,0,47,0,0,0,0,0,91,0,198,0,157,0,156,0,0,0,236,0,219,0);
signal scenario_full  : scenario_type := (11,31,157,31,157,30,251,31,112,31,112,30,23,31,155,31,121,31,204,31,40,31,40,30,130,31,140,31,15,31,213,31,57,31,81,31,206,31,206,30,180,31,180,30,85,31,22,31,22,30,70,31,70,30,229,31,144,31,144,30,51,31,93,31,241,31,211,31,252,31,4,31,35,31,36,31,3,31,105,31,105,30,45,31,31,31,247,31,211,31,229,31,162,31,208,31,152,31,205,31,120,31,120,30,83,31,15,31,40,31,234,31,190,31,69,31,240,31,125,31,7,31,7,30,163,31,39,31,39,30,209,31,48,31,48,30,48,29,178,31,178,30,184,31,101,31,6,31,224,31,179,31,179,30,179,29,179,28,164,31,70,31,72,31,72,30,3,31,221,31,82,31,240,31,136,31,247,31,163,31,231,31,247,31,7,31,56,31,2,31,2,30,64,31,247,31,247,30,213,31,213,30,67,31,101,31,203,31,61,31,61,30,16,31,142,31,251,31,251,30,117,31,7,31,210,31,210,31,14,31,84,31,100,31,100,30,99,31,99,30,33,31,223,31,89,31,17,31,52,31,169,31,212,31,212,30,103,31,105,31,145,31,20,31,73,31,88,31,88,30,88,29,231,31,4,31,60,31,243,31,9,31,145,31,114,31,158,31,205,31,38,31,47,31,47,30,47,29,91,31,198,31,157,31,156,31,156,30,236,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
