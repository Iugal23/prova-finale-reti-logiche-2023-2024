-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_742 is
end project_tb_742;

architecture project_tb_arch_742 of project_tb_742 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 826;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,0,0,0,0,0,0,0,0,0,0,63,0,50,0,135,0,217,0,70,0,128,0,21,0,195,0,11,0,147,0,249,0,180,0,55,0,13,0,175,0,145,0,26,0,185,0,148,0,125,0,0,0,205,0,174,0,216,0,5,0,181,0,170,0,35,0,209,0,107,0,194,0,0,0,118,0,196,0,82,0,150,0,227,0,0,0,135,0,211,0,72,0,217,0,143,0,138,0,136,0,250,0,166,0,43,0,145,0,84,0,146,0,0,0,248,0,92,0,123,0,224,0,96,0,39,0,133,0,140,0,0,0,0,0,61,0,0,0,27,0,19,0,13,0,89,0,91,0,147,0,0,0,192,0,0,0,0,0,47,0,30,0,0,0,17,0,17,0,10,0,179,0,236,0,69,0,10,0,3,0,93,0,189,0,59,0,112,0,220,0,52,0,46,0,150,0,0,0,250,0,2,0,96,0,32,0,89,0,181,0,182,0,186,0,0,0,57,0,164,0,129,0,178,0,219,0,189,0,70,0,94,0,0,0,94,0,172,0,253,0,0,0,60,0,0,0,166,0,22,0,0,0,26,0,29,0,75,0,0,0,73,0,206,0,0,0,129,0,20,0,227,0,226,0,0,0,0,0,205,0,65,0,173,0,144,0,0,0,120,0,69,0,181,0,90,0,93,0,250,0,106,0,7,0,7,0,9,0,130,0,81,0,0,0,242,0,239,0,157,0,246,0,148,0,102,0,137,0,155,0,52,0,216,0,1,0,207,0,34,0,0,0,205,0,38,0,166,0,63,0,179,0,62,0,24,0,236,0,205,0,122,0,0,0,0,0,50,0,149,0,120,0,76,0,42,0,221,0,35,0,225,0,212,0,113,0,0,0,0,0,217,0,182,0,196,0,196,0,102,0,196,0,157,0,54,0,223,0,84,0,0,0,0,0,102,0,226,0,0,0,47,0,201,0,48,0,49,0,151,0,148,0,14,0,0,0,252,0,239,0,74,0,0,0,61,0,32,0,0,0,224,0,0,0,0,0,0,0,114,0,1,0,0,0,185,0,167,0,146,0,197,0,0,0,32,0,0,0,0,0,222,0,119,0,163,0,162,0,89,0,64,0,251,0,0,0,147,0,14,0,143,0,143,0,84,0,226,0,59,0,46,0,103,0,96,0,34,0,0,0,75,0,159,0,151,0,15,0,248,0,0,0,0,0,200,0,0,0,0,0,204,0,72,0,156,0,141,0,0,0,252,0,0,0,63,0,0,0,0,0,244,0,201,0,116,0,98,0,0,0,206,0,72,0,228,0,68,0,69,0,119,0,34,0,147,0,0,0,113,0,81,0,48,0,0,0,254,0,127,0,228,0,187,0,138,0,32,0,29,0,0,0,246,0,222,0,0,0,0,0,234,0,120,0,32,0,212,0,167,0,33,0,0,0,170,0,235,0,170,0,236,0,27,0,144,0,134,0,69,0,243,0,140,0,219,0,147,0,0,0,94,0,210,0,65,0,12,0,230,0,43,0,51,0,202,0,0,0,0,0,53,0,0,0,20,0,212,0,186,0,118,0,157,0,12,0,219,0,20,0,0,0,0,0,221,0,138,0,15,0,0,0,0,0,229,0,129,0,156,0,75,0,56,0,0,0,0,0,0,0,108,0,98,0,128,0,33,0,23,0,0,0,0,0,215,0,207,0,90,0,178,0,141,0,195,0,0,0,95,0,169,0,19,0,205,0,210,0,79,0,204,0,142,0,0,0,60,0,117,0,48,0,64,0,124,0,37,0,0,0,216,0,169,0,61,0,201,0,66,0,0,0,75,0,163,0,133,0,0,0,80,0,204,0,79,0,27,0,54,0,46,0,96,0,67,0,190,0,4,0,174,0,215,0,51,0,105,0,98,0,0,0,183,0,50,0,31,0,83,0,165,0,49,0,0,0,90,0,0,0,217,0,0,0,80,0,92,0,68,0,9,0,105,0,167,0,14,0,220,0,0,0,0,0,178,0,50,0,10,0,38,0,0,0,221,0,210,0,50,0,226,0,0,0,210,0,27,0,0,0,221,0,0,0,0,0,251,0,66,0,107,0,147,0,69,0,90,0,0,0,0,0,24,0,124,0,49,0,177,0,135,0,91,0,89,0,223,0,224,0,0,0,126,0,148,0,214,0,70,0,15,0,127,0,212,0,62,0,21,0,173,0,36,0,185,0,0,0,123,0,70,0,0,0,63,0,187,0,67,0,0,0,34,0,44,0,25,0,141,0,0,0,144,0,79,0,0,0,17,0,111,0,221,0,82,0,83,0,46,0,181,0,200,0,101,0,84,0,194,0,150,0,101,0,158,0,221,0,178,0,0,0,39,0,212,0,205,0,153,0,5,0,71,0,218,0,0,0,45,0,69,0,206,0,29,0,135,0,113,0,181,0,66,0,0,0,0,0,3,0,87,0,225,0,141,0,38,0,113,0,248,0,55,0,196,0,209,0,0,0,0,0,133,0,235,0,0,0,110,0,0,0,201,0,154,0,206,0,34,0,47,0,243,0,93,0,112,0,12,0,22,0,34,0,232,0,242,0,140,0,190,0,32,0,197,0,142,0,0,0,0,0,232,0,250,0,94,0,0,0,72,0,141,0,161,0,0,0,16,0,155,0,0,0,202,0,167,0,121,0,248,0,203,0,154,0,227,0,254,0,180,0,0,0,35,0,90,0,240,0,156,0,232,0,72,0,39,0,42,0,0,0,109,0,0,0,234,0,80,0,200,0,0,0,0,0,0,0,11,0,235,0,234,0,117,0,47,0,217,0,99,0,250,0,111,0,244,0,0,0,108,0,0,0,11,0,0,0,54,0,226,0,0,0,83,0,0,0,0,0,206,0,128,0,70,0,158,0,212,0,51,0,194,0,215,0,152,0,210,0,52,0,182,0,98,0,38,0,0,0,0,0,115,0,47,0,30,0,61,0,135,0,187,0,0,0,34,0,6,0,86,0,145,0,114,0,187,0,43,0,51,0,52,0,47,0,0,0,47,0,207,0,0,0,0,0,250,0,134,0,55,0,66,0,50,0,182,0,135,0,0,0,0,0,239,0,223,0,119,0,189,0,147,0,186,0,0,0,0,0,58,0,198,0,227,0,165,0,31,0,0,0,40,0,0,0,180,0,27,0,0,0,114,0,166,0,169,0,204,0,42,0,180,0,235,0,60,0,44,0,242,0,97,0,199,0,0,0,0,0,183,0,0,0,224,0,154,0,8,0,184,0,242,0,129,0,201,0,242,0,150,0,21,0,105,0,0,0,229,0,81,0,64,0,0,0,111,0,0,0,0,0,0,0,68,0,123,0,218,0,156,0,205,0,83,0,243,0,249,0,0,0,250,0,153,0,96,0,72,0,190,0,84,0,69,0,111,0,213,0,48,0,0,0,229,0,103,0,14,0,0,0,148,0,160,0,79,0,0,0,13,0,44,0,215,0,203,0,120,0,137,0,0,0,40,0,151,0,142,0,149,0,12,0,0,0,0,0,4,0,59,0,85,0,74,0,64,0,189,0,224,0,198,0,75,0,136,0,21,0,0,0,0,0,0,0,8,0,229,0,137,0,200,0,17,0,39,0,124,0,147,0,72,0,152,0,0,0,9,0,216,0,236,0,97,0,50,0,0,0,29,0,102,0,166,0,98,0,59,0,209,0,71,0,23,0,228,0,54,0,74,0,152,0,4,0,206,0,14,0);
signal scenario_full  : scenario_type := (169,31,169,30,169,29,169,28,169,27,169,26,63,31,50,31,135,31,217,31,70,31,128,31,21,31,195,31,11,31,147,31,249,31,180,31,55,31,13,31,175,31,145,31,26,31,185,31,148,31,125,31,125,30,205,31,174,31,216,31,5,31,181,31,170,31,35,31,209,31,107,31,194,31,194,30,118,31,196,31,82,31,150,31,227,31,227,30,135,31,211,31,72,31,217,31,143,31,138,31,136,31,250,31,166,31,43,31,145,31,84,31,146,31,146,30,248,31,92,31,123,31,224,31,96,31,39,31,133,31,140,31,140,30,140,29,61,31,61,30,27,31,19,31,13,31,89,31,91,31,147,31,147,30,192,31,192,30,192,29,47,31,30,31,30,30,17,31,17,31,10,31,179,31,236,31,69,31,10,31,3,31,93,31,189,31,59,31,112,31,220,31,52,31,46,31,150,31,150,30,250,31,2,31,96,31,32,31,89,31,181,31,182,31,186,31,186,30,57,31,164,31,129,31,178,31,219,31,189,31,70,31,94,31,94,30,94,31,172,31,253,31,253,30,60,31,60,30,166,31,22,31,22,30,26,31,29,31,75,31,75,30,73,31,206,31,206,30,129,31,20,31,227,31,226,31,226,30,226,29,205,31,65,31,173,31,144,31,144,30,120,31,69,31,181,31,90,31,93,31,250,31,106,31,7,31,7,31,9,31,130,31,81,31,81,30,242,31,239,31,157,31,246,31,148,31,102,31,137,31,155,31,52,31,216,31,1,31,207,31,34,31,34,30,205,31,38,31,166,31,63,31,179,31,62,31,24,31,236,31,205,31,122,31,122,30,122,29,50,31,149,31,120,31,76,31,42,31,221,31,35,31,225,31,212,31,113,31,113,30,113,29,217,31,182,31,196,31,196,31,102,31,196,31,157,31,54,31,223,31,84,31,84,30,84,29,102,31,226,31,226,30,47,31,201,31,48,31,49,31,151,31,148,31,14,31,14,30,252,31,239,31,74,31,74,30,61,31,32,31,32,30,224,31,224,30,224,29,224,28,114,31,1,31,1,30,185,31,167,31,146,31,197,31,197,30,32,31,32,30,32,29,222,31,119,31,163,31,162,31,89,31,64,31,251,31,251,30,147,31,14,31,143,31,143,31,84,31,226,31,59,31,46,31,103,31,96,31,34,31,34,30,75,31,159,31,151,31,15,31,248,31,248,30,248,29,200,31,200,30,200,29,204,31,72,31,156,31,141,31,141,30,252,31,252,30,63,31,63,30,63,29,244,31,201,31,116,31,98,31,98,30,206,31,72,31,228,31,68,31,69,31,119,31,34,31,147,31,147,30,113,31,81,31,48,31,48,30,254,31,127,31,228,31,187,31,138,31,32,31,29,31,29,30,246,31,222,31,222,30,222,29,234,31,120,31,32,31,212,31,167,31,33,31,33,30,170,31,235,31,170,31,236,31,27,31,144,31,134,31,69,31,243,31,140,31,219,31,147,31,147,30,94,31,210,31,65,31,12,31,230,31,43,31,51,31,202,31,202,30,202,29,53,31,53,30,20,31,212,31,186,31,118,31,157,31,12,31,219,31,20,31,20,30,20,29,221,31,138,31,15,31,15,30,15,29,229,31,129,31,156,31,75,31,56,31,56,30,56,29,56,28,108,31,98,31,128,31,33,31,23,31,23,30,23,29,215,31,207,31,90,31,178,31,141,31,195,31,195,30,95,31,169,31,19,31,205,31,210,31,79,31,204,31,142,31,142,30,60,31,117,31,48,31,64,31,124,31,37,31,37,30,216,31,169,31,61,31,201,31,66,31,66,30,75,31,163,31,133,31,133,30,80,31,204,31,79,31,27,31,54,31,46,31,96,31,67,31,190,31,4,31,174,31,215,31,51,31,105,31,98,31,98,30,183,31,50,31,31,31,83,31,165,31,49,31,49,30,90,31,90,30,217,31,217,30,80,31,92,31,68,31,9,31,105,31,167,31,14,31,220,31,220,30,220,29,178,31,50,31,10,31,38,31,38,30,221,31,210,31,50,31,226,31,226,30,210,31,27,31,27,30,221,31,221,30,221,29,251,31,66,31,107,31,147,31,69,31,90,31,90,30,90,29,24,31,124,31,49,31,177,31,135,31,91,31,89,31,223,31,224,31,224,30,126,31,148,31,214,31,70,31,15,31,127,31,212,31,62,31,21,31,173,31,36,31,185,31,185,30,123,31,70,31,70,30,63,31,187,31,67,31,67,30,34,31,44,31,25,31,141,31,141,30,144,31,79,31,79,30,17,31,111,31,221,31,82,31,83,31,46,31,181,31,200,31,101,31,84,31,194,31,150,31,101,31,158,31,221,31,178,31,178,30,39,31,212,31,205,31,153,31,5,31,71,31,218,31,218,30,45,31,69,31,206,31,29,31,135,31,113,31,181,31,66,31,66,30,66,29,3,31,87,31,225,31,141,31,38,31,113,31,248,31,55,31,196,31,209,31,209,30,209,29,133,31,235,31,235,30,110,31,110,30,201,31,154,31,206,31,34,31,47,31,243,31,93,31,112,31,12,31,22,31,34,31,232,31,242,31,140,31,190,31,32,31,197,31,142,31,142,30,142,29,232,31,250,31,94,31,94,30,72,31,141,31,161,31,161,30,16,31,155,31,155,30,202,31,167,31,121,31,248,31,203,31,154,31,227,31,254,31,180,31,180,30,35,31,90,31,240,31,156,31,232,31,72,31,39,31,42,31,42,30,109,31,109,30,234,31,80,31,200,31,200,30,200,29,200,28,11,31,235,31,234,31,117,31,47,31,217,31,99,31,250,31,111,31,244,31,244,30,108,31,108,30,11,31,11,30,54,31,226,31,226,30,83,31,83,30,83,29,206,31,128,31,70,31,158,31,212,31,51,31,194,31,215,31,152,31,210,31,52,31,182,31,98,31,38,31,38,30,38,29,115,31,47,31,30,31,61,31,135,31,187,31,187,30,34,31,6,31,86,31,145,31,114,31,187,31,43,31,51,31,52,31,47,31,47,30,47,31,207,31,207,30,207,29,250,31,134,31,55,31,66,31,50,31,182,31,135,31,135,30,135,29,239,31,223,31,119,31,189,31,147,31,186,31,186,30,186,29,58,31,198,31,227,31,165,31,31,31,31,30,40,31,40,30,180,31,27,31,27,30,114,31,166,31,169,31,204,31,42,31,180,31,235,31,60,31,44,31,242,31,97,31,199,31,199,30,199,29,183,31,183,30,224,31,154,31,8,31,184,31,242,31,129,31,201,31,242,31,150,31,21,31,105,31,105,30,229,31,81,31,64,31,64,30,111,31,111,30,111,29,111,28,68,31,123,31,218,31,156,31,205,31,83,31,243,31,249,31,249,30,250,31,153,31,96,31,72,31,190,31,84,31,69,31,111,31,213,31,48,31,48,30,229,31,103,31,14,31,14,30,148,31,160,31,79,31,79,30,13,31,44,31,215,31,203,31,120,31,137,31,137,30,40,31,151,31,142,31,149,31,12,31,12,30,12,29,4,31,59,31,85,31,74,31,64,31,189,31,224,31,198,31,75,31,136,31,21,31,21,30,21,29,21,28,8,31,229,31,137,31,200,31,17,31,39,31,124,31,147,31,72,31,152,31,152,30,9,31,216,31,236,31,97,31,50,31,50,30,29,31,102,31,166,31,98,31,59,31,209,31,71,31,23,31,228,31,54,31,74,31,152,31,4,31,206,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
