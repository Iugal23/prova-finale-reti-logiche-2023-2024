-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_801 is
end project_tb_801;

architecture project_tb_arch_801 of project_tb_801 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 918;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,0,0,0,0,212,0,189,0,220,0,160,0,253,0,104,0,71,0,0,0,0,0,0,0,228,0,186,0,117,0,0,0,156,0,0,0,233,0,251,0,137,0,37,0,244,0,22,0,0,0,0,0,0,0,94,0,226,0,0,0,255,0,154,0,195,0,0,0,29,0,71,0,223,0,160,0,172,0,230,0,11,0,114,0,107,0,245,0,0,0,211,0,0,0,49,0,0,0,75,0,40,0,56,0,195,0,27,0,116,0,56,0,129,0,0,0,190,0,173,0,54,0,160,0,92,0,188,0,125,0,255,0,70,0,104,0,238,0,0,0,195,0,91,0,0,0,124,0,201,0,81,0,208,0,69,0,61,0,222,0,0,0,177,0,79,0,0,0,29,0,24,0,1,0,203,0,171,0,18,0,0,0,203,0,233,0,0,0,148,0,0,0,0,0,0,0,125,0,239,0,224,0,213,0,72,0,180,0,253,0,218,0,0,0,0,0,184,0,189,0,0,0,224,0,111,0,153,0,0,0,32,0,107,0,189,0,123,0,62,0,198,0,249,0,179,0,45,0,106,0,141,0,44,0,124,0,0,0,71,0,226,0,224,0,83,0,46,0,0,0,0,0,112,0,206,0,0,0,0,0,0,0,183,0,176,0,220,0,124,0,0,0,212,0,0,0,91,0,0,0,36,0,113,0,78,0,22,0,156,0,17,0,0,0,252,0,212,0,0,0,117,0,0,0,0,0,104,0,170,0,16,0,60,0,17,0,155,0,0,0,206,0,0,0,231,0,0,0,162,0,226,0,82,0,0,0,40,0,161,0,52,0,31,0,215,0,38,0,9,0,62,0,0,0,151,0,0,0,4,0,46,0,127,0,160,0,82,0,159,0,0,0,70,0,222,0,223,0,37,0,0,0,0,0,169,0,174,0,63,0,0,0,0,0,61,0,210,0,249,0,1,0,211,0,0,0,28,0,70,0,170,0,72,0,0,0,0,0,248,0,151,0,9,0,219,0,61,0,0,0,219,0,0,0,0,0,157,0,0,0,183,0,95,0,68,0,223,0,240,0,168,0,0,0,158,0,168,0,0,0,216,0,0,0,54,0,0,0,101,0,0,0,93,0,198,0,0,0,0,0,207,0,0,0,119,0,169,0,211,0,70,0,0,0,147,0,66,0,0,0,85,0,126,0,122,0,0,0,207,0,0,0,191,0,219,0,59,0,39,0,245,0,77,0,149,0,137,0,0,0,55,0,108,0,245,0,193,0,0,0,0,0,171,0,61,0,240,0,106,0,52,0,230,0,86,0,21,0,9,0,9,0,30,0,0,0,10,0,0,0,189,0,96,0,25,0,19,0,25,0,97,0,220,0,240,0,255,0,32,0,49,0,104,0,21,0,0,0,0,0,118,0,119,0,150,0,0,0,142,0,63,0,212,0,0,0,0,0,16,0,28,0,159,0,111,0,0,0,0,0,102,0,35,0,104,0,95,0,189,0,123,0,94,0,0,0,97,0,75,0,18,0,168,0,252,0,169,0,244,0,95,0,183,0,65,0,0,0,0,0,0,0,113,0,0,0,148,0,38,0,78,0,151,0,114,0,136,0,81,0,37,0,91,0,87,0,0,0,212,0,24,0,7,0,26,0,5,0,49,0,40,0,0,0,0,0,220,0,247,0,136,0,154,0,0,0,135,0,0,0,174,0,132,0,163,0,0,0,44,0,231,0,0,0,0,0,47,0,0,0,48,0,0,0,150,0,33,0,222,0,175,0,162,0,79,0,56,0,46,0,221,0,229,0,188,0,37,0,164,0,0,0,116,0,77,0,228,0,0,0,251,0,5,0,0,0,216,0,125,0,0,0,158,0,235,0,109,0,158,0,100,0,43,0,163,0,0,0,71,0,32,0,196,0,122,0,114,0,162,0,196,0,123,0,0,0,0,0,182,0,4,0,72,0,50,0,0,0,230,0,0,0,135,0,0,0,101,0,132,0,87,0,178,0,0,0,225,0,137,0,121,0,175,0,209,0,0,0,187,0,0,0,39,0,0,0,192,0,233,0,37,0,197,0,0,0,135,0,12,0,144,0,185,0,250,0,193,0,154,0,112,0,23,0,23,0,0,0,24,0,128,0,239,0,0,0,202,0,0,0,143,0,178,0,86,0,145,0,51,0,233,0,76,0,79,0,0,0,78,0,44,0,0,0,195,0,149,0,153,0,0,0,191,0,0,0,80,0,117,0,175,0,0,0,247,0,0,0,31,0,228,0,235,0,54,0,17,0,0,0,197,0,158,0,75,0,9,0,181,0,0,0,129,0,158,0,107,0,0,0,2,0,38,0,141,0,184,0,18,0,211,0,104,0,0,0,3,0,182,0,48,0,28,0,36,0,28,0,7,0,213,0,0,0,112,0,233,0,22,0,0,0,214,0,0,0,224,0,243,0,81,0,165,0,0,0,41,0,87,0,167,0,136,0,130,0,0,0,116,0,0,0,177,0,162,0,44,0,19,0,214,0,60,0,152,0,0,0,82,0,73,0,117,0,214,0,161,0,194,0,0,0,120,0,64,0,0,0,244,0,0,0,36,0,0,0,66,0,26,0,246,0,65,0,0,0,137,0,56,0,126,0,29,0,48,0,14,0,129,0,0,0,188,0,140,0,226,0,78,0,0,0,139,0,0,0,0,0,197,0,131,0,24,0,146,0,181,0,0,0,74,0,214,0,161,0,27,0,249,0,102,0,0,0,78,0,151,0,0,0,64,0,172,0,219,0,49,0,30,0,91,0,193,0,180,0,34,0,237,0,124,0,0,0,80,0,189,0,223,0,14,0,40,0,252,0,0,0,0,0,0,0,45,0,122,0,221,0,19,0,108,0,6,0,85,0,38,0,159,0,245,0,169,0,11,0,209,0,165,0,0,0,46,0,198,0,198,0,0,0,82,0,136,0,230,0,214,0,31,0,72,0,12,0,9,0,1,0,1,0,157,0,63,0,30,0,0,0,132,0,196,0,10,0,143,0,0,0,153,0,184,0,181,0,40,0,30,0,151,0,227,0,113,0,205,0,162,0,154,0,158,0,0,0,127,0,0,0,22,0,17,0,90,0,128,0,0,0,165,0,198,0,172,0,217,0,0,0,238,0,185,0,249,0,20,0,119,0,140,0,59,0,241,0,239,0,92,0,234,0,229,0,185,0,147,0,176,0,100,0,125,0,90,0,0,0,5,0,67,0,81,0,47,0,0,0,0,0,0,0,54,0,52,0,131,0,126,0,0,0,0,0,77,0,252,0,101,0,133,0,156,0,28,0,0,0,83,0,0,0,211,0,136,0,0,0,189,0,169,0,217,0,18,0,0,0,152,0,142,0,0,0,159,0,114,0,0,0,0,0,196,0,31,0,73,0,239,0,201,0,0,0,75,0,59,0,66,0,69,0,56,0,255,0,154,0,104,0,239,0,0,0,1,0,175,0,86,0,236,0,38,0,0,0,162,0,213,0,0,0,0,0,245,0,20,0,99,0,203,0,99,0,0,0,171,0,0,0,43,0,99,0,255,0,0,0,86,0,4,0,127,0,15,0,121,0,32,0,105,0,47,0,57,0,212,0,199,0,0,0,0,0,158,0,218,0,36,0,246,0,225,0,79,0,0,0,231,0,47,0,162,0,171,0,105,0,12,0,112,0,0,0,75,0,71,0,54,0,90,0,139,0,179,0,205,0,148,0,192,0,216,0,0,0,174,0,0,0,237,0,237,0,0,0,0,0,0,0,86,0,225,0,192,0,11,0,226,0,56,0,0,0,188,0,4,0,141,0,0,0,212,0,0,0,1,0,174,0,0,0,223,0,192,0,132,0,95,0,56,0,143,0,201,0,175,0,82,0,66,0,120,0,68,0,49,0,0,0,165,0,146,0,197,0,0,0,163,0,34,0,0,0,210,0,101,0,201,0,111,0,0,0,0,0,0,0,197,0,244,0,2,0,156,0,88,0,0,0,0,0,39,0,0,0,200,0,34,0,148,0,0,0,0,0,150,0,240,0,0,0,36,0,0,0,194,0,174,0,190,0,143,0,221,0,159,0,129,0,117,0,0,0,90,0,102,0,217,0,58,0,0,0,155,0,0,0,176,0,147,0,44,0,123,0);
signal scenario_full  : scenario_type := (93,31,93,30,93,29,212,31,189,31,220,31,160,31,253,31,104,31,71,31,71,30,71,29,71,28,228,31,186,31,117,31,117,30,156,31,156,30,233,31,251,31,137,31,37,31,244,31,22,31,22,30,22,29,22,28,94,31,226,31,226,30,255,31,154,31,195,31,195,30,29,31,71,31,223,31,160,31,172,31,230,31,11,31,114,31,107,31,245,31,245,30,211,31,211,30,49,31,49,30,75,31,40,31,56,31,195,31,27,31,116,31,56,31,129,31,129,30,190,31,173,31,54,31,160,31,92,31,188,31,125,31,255,31,70,31,104,31,238,31,238,30,195,31,91,31,91,30,124,31,201,31,81,31,208,31,69,31,61,31,222,31,222,30,177,31,79,31,79,30,29,31,24,31,1,31,203,31,171,31,18,31,18,30,203,31,233,31,233,30,148,31,148,30,148,29,148,28,125,31,239,31,224,31,213,31,72,31,180,31,253,31,218,31,218,30,218,29,184,31,189,31,189,30,224,31,111,31,153,31,153,30,32,31,107,31,189,31,123,31,62,31,198,31,249,31,179,31,45,31,106,31,141,31,44,31,124,31,124,30,71,31,226,31,224,31,83,31,46,31,46,30,46,29,112,31,206,31,206,30,206,29,206,28,183,31,176,31,220,31,124,31,124,30,212,31,212,30,91,31,91,30,36,31,113,31,78,31,22,31,156,31,17,31,17,30,252,31,212,31,212,30,117,31,117,30,117,29,104,31,170,31,16,31,60,31,17,31,155,31,155,30,206,31,206,30,231,31,231,30,162,31,226,31,82,31,82,30,40,31,161,31,52,31,31,31,215,31,38,31,9,31,62,31,62,30,151,31,151,30,4,31,46,31,127,31,160,31,82,31,159,31,159,30,70,31,222,31,223,31,37,31,37,30,37,29,169,31,174,31,63,31,63,30,63,29,61,31,210,31,249,31,1,31,211,31,211,30,28,31,70,31,170,31,72,31,72,30,72,29,248,31,151,31,9,31,219,31,61,31,61,30,219,31,219,30,219,29,157,31,157,30,183,31,95,31,68,31,223,31,240,31,168,31,168,30,158,31,168,31,168,30,216,31,216,30,54,31,54,30,101,31,101,30,93,31,198,31,198,30,198,29,207,31,207,30,119,31,169,31,211,31,70,31,70,30,147,31,66,31,66,30,85,31,126,31,122,31,122,30,207,31,207,30,191,31,219,31,59,31,39,31,245,31,77,31,149,31,137,31,137,30,55,31,108,31,245,31,193,31,193,30,193,29,171,31,61,31,240,31,106,31,52,31,230,31,86,31,21,31,9,31,9,31,30,31,30,30,10,31,10,30,189,31,96,31,25,31,19,31,25,31,97,31,220,31,240,31,255,31,32,31,49,31,104,31,21,31,21,30,21,29,118,31,119,31,150,31,150,30,142,31,63,31,212,31,212,30,212,29,16,31,28,31,159,31,111,31,111,30,111,29,102,31,35,31,104,31,95,31,189,31,123,31,94,31,94,30,97,31,75,31,18,31,168,31,252,31,169,31,244,31,95,31,183,31,65,31,65,30,65,29,65,28,113,31,113,30,148,31,38,31,78,31,151,31,114,31,136,31,81,31,37,31,91,31,87,31,87,30,212,31,24,31,7,31,26,31,5,31,49,31,40,31,40,30,40,29,220,31,247,31,136,31,154,31,154,30,135,31,135,30,174,31,132,31,163,31,163,30,44,31,231,31,231,30,231,29,47,31,47,30,48,31,48,30,150,31,33,31,222,31,175,31,162,31,79,31,56,31,46,31,221,31,229,31,188,31,37,31,164,31,164,30,116,31,77,31,228,31,228,30,251,31,5,31,5,30,216,31,125,31,125,30,158,31,235,31,109,31,158,31,100,31,43,31,163,31,163,30,71,31,32,31,196,31,122,31,114,31,162,31,196,31,123,31,123,30,123,29,182,31,4,31,72,31,50,31,50,30,230,31,230,30,135,31,135,30,101,31,132,31,87,31,178,31,178,30,225,31,137,31,121,31,175,31,209,31,209,30,187,31,187,30,39,31,39,30,192,31,233,31,37,31,197,31,197,30,135,31,12,31,144,31,185,31,250,31,193,31,154,31,112,31,23,31,23,31,23,30,24,31,128,31,239,31,239,30,202,31,202,30,143,31,178,31,86,31,145,31,51,31,233,31,76,31,79,31,79,30,78,31,44,31,44,30,195,31,149,31,153,31,153,30,191,31,191,30,80,31,117,31,175,31,175,30,247,31,247,30,31,31,228,31,235,31,54,31,17,31,17,30,197,31,158,31,75,31,9,31,181,31,181,30,129,31,158,31,107,31,107,30,2,31,38,31,141,31,184,31,18,31,211,31,104,31,104,30,3,31,182,31,48,31,28,31,36,31,28,31,7,31,213,31,213,30,112,31,233,31,22,31,22,30,214,31,214,30,224,31,243,31,81,31,165,31,165,30,41,31,87,31,167,31,136,31,130,31,130,30,116,31,116,30,177,31,162,31,44,31,19,31,214,31,60,31,152,31,152,30,82,31,73,31,117,31,214,31,161,31,194,31,194,30,120,31,64,31,64,30,244,31,244,30,36,31,36,30,66,31,26,31,246,31,65,31,65,30,137,31,56,31,126,31,29,31,48,31,14,31,129,31,129,30,188,31,140,31,226,31,78,31,78,30,139,31,139,30,139,29,197,31,131,31,24,31,146,31,181,31,181,30,74,31,214,31,161,31,27,31,249,31,102,31,102,30,78,31,151,31,151,30,64,31,172,31,219,31,49,31,30,31,91,31,193,31,180,31,34,31,237,31,124,31,124,30,80,31,189,31,223,31,14,31,40,31,252,31,252,30,252,29,252,28,45,31,122,31,221,31,19,31,108,31,6,31,85,31,38,31,159,31,245,31,169,31,11,31,209,31,165,31,165,30,46,31,198,31,198,31,198,30,82,31,136,31,230,31,214,31,31,31,72,31,12,31,9,31,1,31,1,31,157,31,63,31,30,31,30,30,132,31,196,31,10,31,143,31,143,30,153,31,184,31,181,31,40,31,30,31,151,31,227,31,113,31,205,31,162,31,154,31,158,31,158,30,127,31,127,30,22,31,17,31,90,31,128,31,128,30,165,31,198,31,172,31,217,31,217,30,238,31,185,31,249,31,20,31,119,31,140,31,59,31,241,31,239,31,92,31,234,31,229,31,185,31,147,31,176,31,100,31,125,31,90,31,90,30,5,31,67,31,81,31,47,31,47,30,47,29,47,28,54,31,52,31,131,31,126,31,126,30,126,29,77,31,252,31,101,31,133,31,156,31,28,31,28,30,83,31,83,30,211,31,136,31,136,30,189,31,169,31,217,31,18,31,18,30,152,31,142,31,142,30,159,31,114,31,114,30,114,29,196,31,31,31,73,31,239,31,201,31,201,30,75,31,59,31,66,31,69,31,56,31,255,31,154,31,104,31,239,31,239,30,1,31,175,31,86,31,236,31,38,31,38,30,162,31,213,31,213,30,213,29,245,31,20,31,99,31,203,31,99,31,99,30,171,31,171,30,43,31,99,31,255,31,255,30,86,31,4,31,127,31,15,31,121,31,32,31,105,31,47,31,57,31,212,31,199,31,199,30,199,29,158,31,218,31,36,31,246,31,225,31,79,31,79,30,231,31,47,31,162,31,171,31,105,31,12,31,112,31,112,30,75,31,71,31,54,31,90,31,139,31,179,31,205,31,148,31,192,31,216,31,216,30,174,31,174,30,237,31,237,31,237,30,237,29,237,28,86,31,225,31,192,31,11,31,226,31,56,31,56,30,188,31,4,31,141,31,141,30,212,31,212,30,1,31,174,31,174,30,223,31,192,31,132,31,95,31,56,31,143,31,201,31,175,31,82,31,66,31,120,31,68,31,49,31,49,30,165,31,146,31,197,31,197,30,163,31,34,31,34,30,210,31,101,31,201,31,111,31,111,30,111,29,111,28,197,31,244,31,2,31,156,31,88,31,88,30,88,29,39,31,39,30,200,31,34,31,148,31,148,30,148,29,150,31,240,31,240,30,36,31,36,30,194,31,174,31,190,31,143,31,221,31,159,31,129,31,117,31,117,30,90,31,102,31,217,31,58,31,58,30,155,31,155,30,176,31,147,31,44,31,123,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
