-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 369;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,47,0,86,0,118,0,0,0,39,0,0,0,133,0,0,0,0,0,183,0,102,0,66,0,112,0,99,0,163,0,170,0,159,0,0,0,115,0,0,0,179,0,80,0,155,0,34,0,122,0,214,0,51,0,239,0,0,0,191,0,41,0,41,0,125,0,47,0,197,0,0,0,0,0,131,0,89,0,249,0,65,0,209,0,0,0,235,0,148,0,0,0,19,0,10,0,113,0,0,0,200,0,134,0,134,0,194,0,174,0,90,0,88,0,108,0,208,0,152,0,17,0,174,0,40,0,17,0,143,0,188,0,113,0,111,0,129,0,0,0,17,0,188,0,45,0,97,0,33,0,23,0,71,0,27,0,157,0,0,0,0,0,167,0,145,0,115,0,129,0,0,0,153,0,249,0,0,0,245,0,5,0,81,0,189,0,182,0,156,0,177,0,0,0,190,0,208,0,154,0,226,0,94,0,50,0,111,0,169,0,194,0,91,0,0,0,57,0,190,0,0,0,0,0,50,0,0,0,0,0,0,0,28,0,4,0,171,0,148,0,40,0,21,0,188,0,0,0,61,0,120,0,162,0,0,0,139,0,51,0,0,0,185,0,159,0,114,0,202,0,33,0,0,0,213,0,228,0,120,0,5,0,163,0,138,0,201,0,0,0,167,0,0,0,113,0,80,0,211,0,18,0,50,0,157,0,159,0,136,0,213,0,218,0,227,0,157,0,0,0,0,0,163,0,0,0,115,0,243,0,91,0,40,0,24,0,90,0,220,0,206,0,0,0,37,0,174,0,186,0,0,0,72,0,139,0,39,0,168,0,201,0,107,0,201,0,16,0,0,0,58,0,245,0,165,0,115,0,84,0,0,0,149,0,206,0,0,0,64,0,0,0,158,0,135,0,0,0,114,0,8,0,36,0,221,0,0,0,131,0,23,0,114,0,192,0,132,0,22,0,30,0,221,0,62,0,127,0,0,0,192,0,9,0,246,0,0,0,87,0,164,0,2,0,252,0,87,0,66,0,202,0,111,0,139,0,155,0,248,0,81,0,0,0,148,0,157,0,0,0,211,0,197,0,168,0,136,0,25,0,82,0,0,0,0,0,0,0,5,0,164,0,220,0,130,0,158,0,0,0,0,0,123,0,31,0,36,0,142,0,0,0,28,0,185,0,246,0,0,0,61,0,112,0,0,0,189,0,0,0,145,0,233,0,74,0,154,0,119,0,52,0,68,0,154,0,235,0,152,0,171,0,176,0,178,0,46,0,241,0,138,0,88,0,0,0,190,0,246,0,96,0,112,0,100,0,14,0,207,0,40,0,220,0,173,0,224,0,0,0,242,0,157,0,216,0,191,0,255,0,5,0,85,0,121,0,102,0,35,0,34,0,54,0,244,0,0,0,16,0,199,0,29,0,0,0,0,0,0,0,0,0,58,0,31,0,234,0,198,0,192,0,140,0,107,0,189,0,131,0,61,0,189,0,56,0,178,0,167,0,205,0,0,0,101,0,0,0,9,0,0,0,247,0,246,0,162,0,0,0,186,0,187,0,0,0,0,0,68,0,0,0,25,0,0,0,251,0,0,0,125,0,0,0,34,0,240,0,214,0,75,0,9,0,100,0,197,0,66,0,116,0,69,0,184,0,200,0,60,0,196,0,0,0,69,0);
signal scenario_full  : scenario_type := (139,31,47,31,86,31,118,31,118,30,39,31,39,30,133,31,133,30,133,29,183,31,102,31,66,31,112,31,99,31,163,31,170,31,159,31,159,30,115,31,115,30,179,31,80,31,155,31,34,31,122,31,214,31,51,31,239,31,239,30,191,31,41,31,41,31,125,31,47,31,197,31,197,30,197,29,131,31,89,31,249,31,65,31,209,31,209,30,235,31,148,31,148,30,19,31,10,31,113,31,113,30,200,31,134,31,134,31,194,31,174,31,90,31,88,31,108,31,208,31,152,31,17,31,174,31,40,31,17,31,143,31,188,31,113,31,111,31,129,31,129,30,17,31,188,31,45,31,97,31,33,31,23,31,71,31,27,31,157,31,157,30,157,29,167,31,145,31,115,31,129,31,129,30,153,31,249,31,249,30,245,31,5,31,81,31,189,31,182,31,156,31,177,31,177,30,190,31,208,31,154,31,226,31,94,31,50,31,111,31,169,31,194,31,91,31,91,30,57,31,190,31,190,30,190,29,50,31,50,30,50,29,50,28,28,31,4,31,171,31,148,31,40,31,21,31,188,31,188,30,61,31,120,31,162,31,162,30,139,31,51,31,51,30,185,31,159,31,114,31,202,31,33,31,33,30,213,31,228,31,120,31,5,31,163,31,138,31,201,31,201,30,167,31,167,30,113,31,80,31,211,31,18,31,50,31,157,31,159,31,136,31,213,31,218,31,227,31,157,31,157,30,157,29,163,31,163,30,115,31,243,31,91,31,40,31,24,31,90,31,220,31,206,31,206,30,37,31,174,31,186,31,186,30,72,31,139,31,39,31,168,31,201,31,107,31,201,31,16,31,16,30,58,31,245,31,165,31,115,31,84,31,84,30,149,31,206,31,206,30,64,31,64,30,158,31,135,31,135,30,114,31,8,31,36,31,221,31,221,30,131,31,23,31,114,31,192,31,132,31,22,31,30,31,221,31,62,31,127,31,127,30,192,31,9,31,246,31,246,30,87,31,164,31,2,31,252,31,87,31,66,31,202,31,111,31,139,31,155,31,248,31,81,31,81,30,148,31,157,31,157,30,211,31,197,31,168,31,136,31,25,31,82,31,82,30,82,29,82,28,5,31,164,31,220,31,130,31,158,31,158,30,158,29,123,31,31,31,36,31,142,31,142,30,28,31,185,31,246,31,246,30,61,31,112,31,112,30,189,31,189,30,145,31,233,31,74,31,154,31,119,31,52,31,68,31,154,31,235,31,152,31,171,31,176,31,178,31,46,31,241,31,138,31,88,31,88,30,190,31,246,31,96,31,112,31,100,31,14,31,207,31,40,31,220,31,173,31,224,31,224,30,242,31,157,31,216,31,191,31,255,31,5,31,85,31,121,31,102,31,35,31,34,31,54,31,244,31,244,30,16,31,199,31,29,31,29,30,29,29,29,28,29,27,58,31,31,31,234,31,198,31,192,31,140,31,107,31,189,31,131,31,61,31,189,31,56,31,178,31,167,31,205,31,205,30,101,31,101,30,9,31,9,30,247,31,246,31,162,31,162,30,186,31,187,31,187,30,187,29,68,31,68,30,25,31,25,30,251,31,251,30,125,31,125,30,34,31,240,31,214,31,75,31,9,31,100,31,197,31,66,31,116,31,69,31,184,31,200,31,60,31,196,31,196,30,69,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
