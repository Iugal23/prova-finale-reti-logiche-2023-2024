-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 452;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,60,0,194,0,218,0,62,0,0,0,0,0,48,0,105,0,96,0,168,0,0,0,0,0,138,0,67,0,168,0,95,0,0,0,111,0,230,0,0,0,131,0,6,0,0,0,115,0,154,0,175,0,193,0,30,0,122,0,134,0,224,0,103,0,123,0,231,0,17,0,53,0,58,0,0,0,0,0,177,0,93,0,0,0,0,0,69,0,4,0,217,0,15,0,91,0,0,0,241,0,0,0,60,0,2,0,196,0,234,0,251,0,206,0,0,0,108,0,124,0,45,0,0,0,72,0,99,0,164,0,102,0,244,0,218,0,123,0,28,0,167,0,51,0,77,0,0,0,27,0,20,0,233,0,0,0,42,0,0,0,189,0,207,0,0,0,17,0,252,0,142,0,195,0,24,0,0,0,0,0,117,0,0,0,93,0,208,0,8,0,113,0,203,0,61,0,87,0,119,0,103,0,121,0,95,0,71,0,178,0,0,0,216,0,0,0,214,0,74,0,0,0,13,0,247,0,3,0,227,0,39,0,0,0,155,0,55,0,0,0,0,0,237,0,153,0,63,0,215,0,0,0,152,0,180,0,0,0,0,0,58,0,143,0,126,0,254,0,236,0,0,0,67,0,0,0,103,0,240,0,159,0,2,0,4,0,208,0,212,0,190,0,214,0,37,0,125,0,0,0,158,0,154,0,0,0,93,0,10,0,118,0,0,0,249,0,49,0,0,0,36,0,31,0,0,0,226,0,181,0,27,0,124,0,0,0,218,0,56,0,86,0,69,0,68,0,100,0,109,0,0,0,190,0,230,0,113,0,252,0,204,0,0,0,42,0,69,0,9,0,0,0,124,0,160,0,19,0,181,0,210,0,248,0,42,0,202,0,253,0,221,0,113,0,60,0,61,0,193,0,24,0,0,0,107,0,242,0,164,0,116,0,191,0,158,0,0,0,41,0,15,0,71,0,126,0,0,0,102,0,194,0,72,0,197,0,0,0,117,0,60,0,0,0,0,0,0,0,175,0,0,0,58,0,166,0,143,0,96,0,171,0,0,0,215,0,173,0,132,0,12,0,226,0,72,0,178,0,41,0,100,0,227,0,0,0,240,0,60,0,49,0,44,0,109,0,0,0,64,0,93,0,226,0,240,0,0,0,71,0,23,0,130,0,0,0,29,0,5,0,0,0,0,0,0,0,76,0,146,0,2,0,148,0,0,0,23,0,49,0,101,0,154,0,25,0,182,0,0,0,19,0,69,0,174,0,206,0,172,0,205,0,0,0,244,0,103,0,181,0,0,0,128,0,0,0,0,0,173,0,2,0,211,0,0,0,159,0,171,0,193,0,185,0,176,0,0,0,164,0,0,0,111,0,241,0,0,0,0,0,73,0,180,0,53,0,141,0,145,0,32,0,38,0,134,0,93,0,0,0,249,0,0,0,0,0,253,0,0,0,0,0,183,0,107,0,239,0,236,0,31,0,170,0,0,0,69,0,143,0,43,0,0,0,226,0,0,0,11,0,206,0,60,0,20,0,114,0,0,0,224,0,149,0,57,0,24,0,152,0,0,0,0,0,253,0,21,0,74,0,77,0,0,0,56,0,219,0,174,0,0,0,35,0,32,0,200,0,231,0,76,0,80,0,199,0,145,0,0,0,190,0,221,0,185,0,8,0,162,0,163,0,122,0,85,0,195,0,205,0,172,0,33,0,216,0,250,0,250,0,14,0,19,0,213,0,88,0,203,0,25,0,215,0,89,0,154,0,26,0,0,0,134,0,0,0,0,0,150,0,8,0,23,0,3,0,72,0,98,0,28,0,200,0,5,0,0,0,0,0,0,0,136,0,86,0,139,0,53,0,223,0,228,0,0,0,163,0,17,0,0,0,137,0,244,0,2,0,0,0,0,0,157,0,106,0,0,0,0,0,96,0,167,0,149,0,10,0,0,0,187,0,33,0,0,0,253,0,220,0,12,0,0,0,65,0,166,0,152,0,109,0,75,0,110,0,0,0,175,0,244,0,179,0,182,0,211,0,0,0,141,0);
signal scenario_full  : scenario_type := (245,31,60,31,194,31,218,31,62,31,62,30,62,29,48,31,105,31,96,31,168,31,168,30,168,29,138,31,67,31,168,31,95,31,95,30,111,31,230,31,230,30,131,31,6,31,6,30,115,31,154,31,175,31,193,31,30,31,122,31,134,31,224,31,103,31,123,31,231,31,17,31,53,31,58,31,58,30,58,29,177,31,93,31,93,30,93,29,69,31,4,31,217,31,15,31,91,31,91,30,241,31,241,30,60,31,2,31,196,31,234,31,251,31,206,31,206,30,108,31,124,31,45,31,45,30,72,31,99,31,164,31,102,31,244,31,218,31,123,31,28,31,167,31,51,31,77,31,77,30,27,31,20,31,233,31,233,30,42,31,42,30,189,31,207,31,207,30,17,31,252,31,142,31,195,31,24,31,24,30,24,29,117,31,117,30,93,31,208,31,8,31,113,31,203,31,61,31,87,31,119,31,103,31,121,31,95,31,71,31,178,31,178,30,216,31,216,30,214,31,74,31,74,30,13,31,247,31,3,31,227,31,39,31,39,30,155,31,55,31,55,30,55,29,237,31,153,31,63,31,215,31,215,30,152,31,180,31,180,30,180,29,58,31,143,31,126,31,254,31,236,31,236,30,67,31,67,30,103,31,240,31,159,31,2,31,4,31,208,31,212,31,190,31,214,31,37,31,125,31,125,30,158,31,154,31,154,30,93,31,10,31,118,31,118,30,249,31,49,31,49,30,36,31,31,31,31,30,226,31,181,31,27,31,124,31,124,30,218,31,56,31,86,31,69,31,68,31,100,31,109,31,109,30,190,31,230,31,113,31,252,31,204,31,204,30,42,31,69,31,9,31,9,30,124,31,160,31,19,31,181,31,210,31,248,31,42,31,202,31,253,31,221,31,113,31,60,31,61,31,193,31,24,31,24,30,107,31,242,31,164,31,116,31,191,31,158,31,158,30,41,31,15,31,71,31,126,31,126,30,102,31,194,31,72,31,197,31,197,30,117,31,60,31,60,30,60,29,60,28,175,31,175,30,58,31,166,31,143,31,96,31,171,31,171,30,215,31,173,31,132,31,12,31,226,31,72,31,178,31,41,31,100,31,227,31,227,30,240,31,60,31,49,31,44,31,109,31,109,30,64,31,93,31,226,31,240,31,240,30,71,31,23,31,130,31,130,30,29,31,5,31,5,30,5,29,5,28,76,31,146,31,2,31,148,31,148,30,23,31,49,31,101,31,154,31,25,31,182,31,182,30,19,31,69,31,174,31,206,31,172,31,205,31,205,30,244,31,103,31,181,31,181,30,128,31,128,30,128,29,173,31,2,31,211,31,211,30,159,31,171,31,193,31,185,31,176,31,176,30,164,31,164,30,111,31,241,31,241,30,241,29,73,31,180,31,53,31,141,31,145,31,32,31,38,31,134,31,93,31,93,30,249,31,249,30,249,29,253,31,253,30,253,29,183,31,107,31,239,31,236,31,31,31,170,31,170,30,69,31,143,31,43,31,43,30,226,31,226,30,11,31,206,31,60,31,20,31,114,31,114,30,224,31,149,31,57,31,24,31,152,31,152,30,152,29,253,31,21,31,74,31,77,31,77,30,56,31,219,31,174,31,174,30,35,31,32,31,200,31,231,31,76,31,80,31,199,31,145,31,145,30,190,31,221,31,185,31,8,31,162,31,163,31,122,31,85,31,195,31,205,31,172,31,33,31,216,31,250,31,250,31,14,31,19,31,213,31,88,31,203,31,25,31,215,31,89,31,154,31,26,31,26,30,134,31,134,30,134,29,150,31,8,31,23,31,3,31,72,31,98,31,28,31,200,31,5,31,5,30,5,29,5,28,136,31,86,31,139,31,53,31,223,31,228,31,228,30,163,31,17,31,17,30,137,31,244,31,2,31,2,30,2,29,157,31,106,31,106,30,106,29,96,31,167,31,149,31,10,31,10,30,187,31,33,31,33,30,253,31,220,31,12,31,12,30,65,31,166,31,152,31,109,31,75,31,110,31,110,30,175,31,244,31,179,31,182,31,211,31,211,30,141,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
