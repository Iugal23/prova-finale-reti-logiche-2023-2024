-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 726;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,185,0,174,0,0,0,92,0,109,0,241,0,85,0,48,0,38,0,141,0,213,0,42,0,150,0,196,0,254,0,160,0,252,0,0,0,190,0,108,0,56,0,0,0,21,0,185,0,137,0,87,0,0,0,46,0,179,0,138,0,131,0,122,0,236,0,147,0,0,0,78,0,249,0,42,0,33,0,216,0,225,0,226,0,98,0,247,0,0,0,71,0,98,0,198,0,49,0,186,0,79,0,0,0,112,0,67,0,81,0,4,0,156,0,47,0,237,0,88,0,0,0,0,0,94,0,161,0,82,0,163,0,170,0,0,0,0,0,117,0,175,0,254,0,63,0,58,0,209,0,254,0,0,0,0,0,131,0,76,0,72,0,104,0,242,0,72,0,191,0,115,0,225,0,155,0,0,0,0,0,70,0,117,0,69,0,164,0,87,0,136,0,9,0,0,0,129,0,9,0,0,0,122,0,0,0,0,0,0,0,0,0,17,0,138,0,76,0,135,0,123,0,0,0,225,0,0,0,179,0,50,0,146,0,193,0,188,0,78,0,179,0,158,0,52,0,0,0,83,0,162,0,59,0,184,0,23,0,155,0,118,0,193,0,148,0,122,0,0,0,14,0,6,0,38,0,11,0,194,0,151,0,0,0,106,0,0,0,229,0,47,0,0,0,122,0,29,0,172,0,241,0,195,0,137,0,31,0,0,0,229,0,41,0,243,0,165,0,71,0,45,0,122,0,68,0,125,0,5,0,125,0,0,0,0,0,232,0,6,0,154,0,0,0,0,0,5,0,242,0,0,0,29,0,0,0,104,0,188,0,0,0,243,0,43,0,24,0,0,0,2,0,11,0,184,0,110,0,0,0,94,0,8,0,7,0,117,0,77,0,62,0,31,0,204,0,129,0,66,0,88,0,133,0,0,0,82,0,0,0,0,0,48,0,97,0,0,0,124,0,215,0,0,0,136,0,232,0,0,0,0,0,137,0,217,0,1,0,99,0,231,0,218,0,222,0,53,0,137,0,180,0,25,0,54,0,250,0,147,0,181,0,178,0,76,0,0,0,231,0,12,0,240,0,0,0,0,0,252,0,245,0,7,0,168,0,24,0,0,0,32,0,25,0,204,0,53,0,134,0,216,0,40,0,141,0,239,0,0,0,74,0,123,0,87,0,215,0,149,0,160,0,49,0,8,0,0,0,224,0,105,0,0,0,15,0,0,0,0,0,102,0,164,0,113,0,149,0,60,0,36,0,12,0,0,0,157,0,149,0,130,0,249,0,57,0,216,0,183,0,0,0,81,0,29,0,0,0,50,0,138,0,191,0,0,0,16,0,210,0,0,0,129,0,165,0,0,0,0,0,134,0,0,0,241,0,108,0,76,0,78,0,191,0,194,0,209,0,32,0,0,0,0,0,0,0,125,0,229,0,158,0,25,0,105,0,86,0,247,0,0,0,119,0,81,0,228,0,125,0,190,0,171,0,228,0,0,0,11,0,112,0,77,0,93,0,124,0,0,0,10,0,180,0,61,0,218,0,191,0,176,0,0,0,0,0,73,0,39,0,191,0,0,0,45,0,38,0,0,0,0,0,204,0,253,0,37,0,234,0,132,0,81,0,117,0,0,0,103,0,183,0,148,0,0,0,133,0,0,0,0,0,241,0,144,0,44,0,126,0,66,0,20,0,0,0,0,0,240,0,0,0,46,0,0,0,138,0,78,0,126,0,130,0,121,0,200,0,228,0,74,0,57,0,200,0,0,0,112,0,127,0,212,0,0,0,0,0,203,0,247,0,66,0,0,0,0,0,56,0,206,0,169,0,2,0,56,0,0,0,164,0,162,0,0,0,0,0,26,0,0,0,100,0,151,0,117,0,207,0,72,0,31,0,3,0,58,0,29,0,253,0,58,0,22,0,43,0,0,0,202,0,53,0,121,0,114,0,97,0,160,0,209,0,238,0,155,0,245,0,113,0,46,0,124,0,172,0,0,0,236,0,184,0,92,0,36,0,128,0,235,0,186,0,175,0,41,0,95,0,227,0,56,0,114,0,68,0,65,0,195,0,201,0,0,0,0,0,108,0,154,0,0,0,47,0,136,0,0,0,45,0,119,0,39,0,213,0,120,0,64,0,74,0,113,0,92,0,48,0,177,0,0,0,168,0,90,0,148,0,218,0,173,0,180,0,160,0,245,0,138,0,0,0,93,0,155,0,10,0,132,0,181,0,172,0,0,0,90,0,17,0,189,0,150,0,149,0,60,0,11,0,0,0,182,0,0,0,92,0,54,0,211,0,0,0,26,0,233,0,249,0,0,0,12,0,251,0,61,0,0,0,248,0,130,0,137,0,45,0,55,0,178,0,9,0,32,0,46,0,229,0,0,0,165,0,119,0,30,0,0,0,60,0,228,0,1,0,0,0,12,0,94,0,22,0,0,0,202,0,0,0,174,0,219,0,101,0,38,0,106,0,0,0,170,0,230,0,54,0,69,0,248,0,241,0,41,0,0,0,239,0,127,0,36,0,188,0,225,0,120,0,0,0,187,0,242,0,197,0,186,0,172,0,0,0,209,0,73,0,81,0,226,0,88,0,62,0,52,0,0,0,0,0,241,0,43,0,0,0,91,0,46,0,154,0,51,0,155,0,90,0,228,0,106,0,86,0,35,0,176,0,216,0,217,0,0,0,167,0,0,0,0,0,0,0,0,0,36,0,215,0,15,0,167,0,115,0,0,0,37,0,140,0,212,0,186,0,0,0,255,0,172,0,67,0,56,0,225,0,27,0,187,0,37,0,59,0,234,0,181,0,252,0,82,0,0,0,0,0,128,0,0,0,121,0,214,0,26,0,189,0,76,0,235,0,32,0,117,0,246,0,0,0,85,0,83,0,0,0,44,0,201,0,229,0,180,0,2,0,187,0,119,0,12,0,0,0,155,0,137,0,128,0,151,0,78,0,24,0,50,0,12,0,233,0,37,0,0,0,255,0,85,0,172,0,0,0,6,0,243,0,171,0,96,0,64,0,82,0,46,0,87,0,186,0,47,0,109,0,129,0,60,0,0,0,18,0,0,0,0,0,45,0,0,0,17,0,190,0,42,0,0,0,110,0,34,0,81,0,233,0,180,0,0,0,109,0,0,0,90,0,41,0,0,0,0,0,179,0,0,0,89,0,186,0,0,0,16,0,105,0,229,0,44,0,100,0,96,0,0,0,0,0,242,0,160,0,0,0,180,0,143,0,47,0,116,0,92,0,69,0,226,0,208,0,114,0,247,0);
signal scenario_full  : scenario_type := (95,31,185,31,174,31,174,30,92,31,109,31,241,31,85,31,48,31,38,31,141,31,213,31,42,31,150,31,196,31,254,31,160,31,252,31,252,30,190,31,108,31,56,31,56,30,21,31,185,31,137,31,87,31,87,30,46,31,179,31,138,31,131,31,122,31,236,31,147,31,147,30,78,31,249,31,42,31,33,31,216,31,225,31,226,31,98,31,247,31,247,30,71,31,98,31,198,31,49,31,186,31,79,31,79,30,112,31,67,31,81,31,4,31,156,31,47,31,237,31,88,31,88,30,88,29,94,31,161,31,82,31,163,31,170,31,170,30,170,29,117,31,175,31,254,31,63,31,58,31,209,31,254,31,254,30,254,29,131,31,76,31,72,31,104,31,242,31,72,31,191,31,115,31,225,31,155,31,155,30,155,29,70,31,117,31,69,31,164,31,87,31,136,31,9,31,9,30,129,31,9,31,9,30,122,31,122,30,122,29,122,28,122,27,17,31,138,31,76,31,135,31,123,31,123,30,225,31,225,30,179,31,50,31,146,31,193,31,188,31,78,31,179,31,158,31,52,31,52,30,83,31,162,31,59,31,184,31,23,31,155,31,118,31,193,31,148,31,122,31,122,30,14,31,6,31,38,31,11,31,194,31,151,31,151,30,106,31,106,30,229,31,47,31,47,30,122,31,29,31,172,31,241,31,195,31,137,31,31,31,31,30,229,31,41,31,243,31,165,31,71,31,45,31,122,31,68,31,125,31,5,31,125,31,125,30,125,29,232,31,6,31,154,31,154,30,154,29,5,31,242,31,242,30,29,31,29,30,104,31,188,31,188,30,243,31,43,31,24,31,24,30,2,31,11,31,184,31,110,31,110,30,94,31,8,31,7,31,117,31,77,31,62,31,31,31,204,31,129,31,66,31,88,31,133,31,133,30,82,31,82,30,82,29,48,31,97,31,97,30,124,31,215,31,215,30,136,31,232,31,232,30,232,29,137,31,217,31,1,31,99,31,231,31,218,31,222,31,53,31,137,31,180,31,25,31,54,31,250,31,147,31,181,31,178,31,76,31,76,30,231,31,12,31,240,31,240,30,240,29,252,31,245,31,7,31,168,31,24,31,24,30,32,31,25,31,204,31,53,31,134,31,216,31,40,31,141,31,239,31,239,30,74,31,123,31,87,31,215,31,149,31,160,31,49,31,8,31,8,30,224,31,105,31,105,30,15,31,15,30,15,29,102,31,164,31,113,31,149,31,60,31,36,31,12,31,12,30,157,31,149,31,130,31,249,31,57,31,216,31,183,31,183,30,81,31,29,31,29,30,50,31,138,31,191,31,191,30,16,31,210,31,210,30,129,31,165,31,165,30,165,29,134,31,134,30,241,31,108,31,76,31,78,31,191,31,194,31,209,31,32,31,32,30,32,29,32,28,125,31,229,31,158,31,25,31,105,31,86,31,247,31,247,30,119,31,81,31,228,31,125,31,190,31,171,31,228,31,228,30,11,31,112,31,77,31,93,31,124,31,124,30,10,31,180,31,61,31,218,31,191,31,176,31,176,30,176,29,73,31,39,31,191,31,191,30,45,31,38,31,38,30,38,29,204,31,253,31,37,31,234,31,132,31,81,31,117,31,117,30,103,31,183,31,148,31,148,30,133,31,133,30,133,29,241,31,144,31,44,31,126,31,66,31,20,31,20,30,20,29,240,31,240,30,46,31,46,30,138,31,78,31,126,31,130,31,121,31,200,31,228,31,74,31,57,31,200,31,200,30,112,31,127,31,212,31,212,30,212,29,203,31,247,31,66,31,66,30,66,29,56,31,206,31,169,31,2,31,56,31,56,30,164,31,162,31,162,30,162,29,26,31,26,30,100,31,151,31,117,31,207,31,72,31,31,31,3,31,58,31,29,31,253,31,58,31,22,31,43,31,43,30,202,31,53,31,121,31,114,31,97,31,160,31,209,31,238,31,155,31,245,31,113,31,46,31,124,31,172,31,172,30,236,31,184,31,92,31,36,31,128,31,235,31,186,31,175,31,41,31,95,31,227,31,56,31,114,31,68,31,65,31,195,31,201,31,201,30,201,29,108,31,154,31,154,30,47,31,136,31,136,30,45,31,119,31,39,31,213,31,120,31,64,31,74,31,113,31,92,31,48,31,177,31,177,30,168,31,90,31,148,31,218,31,173,31,180,31,160,31,245,31,138,31,138,30,93,31,155,31,10,31,132,31,181,31,172,31,172,30,90,31,17,31,189,31,150,31,149,31,60,31,11,31,11,30,182,31,182,30,92,31,54,31,211,31,211,30,26,31,233,31,249,31,249,30,12,31,251,31,61,31,61,30,248,31,130,31,137,31,45,31,55,31,178,31,9,31,32,31,46,31,229,31,229,30,165,31,119,31,30,31,30,30,60,31,228,31,1,31,1,30,12,31,94,31,22,31,22,30,202,31,202,30,174,31,219,31,101,31,38,31,106,31,106,30,170,31,230,31,54,31,69,31,248,31,241,31,41,31,41,30,239,31,127,31,36,31,188,31,225,31,120,31,120,30,187,31,242,31,197,31,186,31,172,31,172,30,209,31,73,31,81,31,226,31,88,31,62,31,52,31,52,30,52,29,241,31,43,31,43,30,91,31,46,31,154,31,51,31,155,31,90,31,228,31,106,31,86,31,35,31,176,31,216,31,217,31,217,30,167,31,167,30,167,29,167,28,167,27,36,31,215,31,15,31,167,31,115,31,115,30,37,31,140,31,212,31,186,31,186,30,255,31,172,31,67,31,56,31,225,31,27,31,187,31,37,31,59,31,234,31,181,31,252,31,82,31,82,30,82,29,128,31,128,30,121,31,214,31,26,31,189,31,76,31,235,31,32,31,117,31,246,31,246,30,85,31,83,31,83,30,44,31,201,31,229,31,180,31,2,31,187,31,119,31,12,31,12,30,155,31,137,31,128,31,151,31,78,31,24,31,50,31,12,31,233,31,37,31,37,30,255,31,85,31,172,31,172,30,6,31,243,31,171,31,96,31,64,31,82,31,46,31,87,31,186,31,47,31,109,31,129,31,60,31,60,30,18,31,18,30,18,29,45,31,45,30,17,31,190,31,42,31,42,30,110,31,34,31,81,31,233,31,180,31,180,30,109,31,109,30,90,31,41,31,41,30,41,29,179,31,179,30,89,31,186,31,186,30,16,31,105,31,229,31,44,31,100,31,96,31,96,30,96,29,242,31,160,31,160,30,180,31,143,31,47,31,116,31,92,31,69,31,226,31,208,31,114,31,247,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
