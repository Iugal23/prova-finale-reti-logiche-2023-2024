-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 477;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,111,0,206,0,75,0,23,0,197,0,0,0,102,0,137,0,88,0,93,0,233,0,143,0,0,0,3,0,56,0,0,0,190,0,190,0,188,0,71,0,168,0,114,0,0,0,0,0,230,0,230,0,54,0,0,0,146,0,195,0,92,0,88,0,82,0,129,0,111,0,172,0,155,0,75,0,49,0,118,0,101,0,72,0,206,0,84,0,0,0,186,0,188,0,242,0,94,0,170,0,97,0,128,0,0,0,188,0,102,0,236,0,197,0,0,0,55,0,122,0,81,0,181,0,168,0,161,0,56,0,0,0,41,0,211,0,32,0,141,0,182,0,178,0,106,0,35,0,211,0,45,0,184,0,200,0,209,0,131,0,0,0,0,0,100,0,186,0,232,0,25,0,170,0,237,0,109,0,174,0,138,0,0,0,62,0,180,0,163,0,245,0,28,0,30,0,151,0,65,0,0,0,235,0,63,0,66,0,239,0,253,0,109,0,192,0,28,0,229,0,50,0,218,0,214,0,204,0,57,0,9,0,9,0,108,0,226,0,0,0,118,0,131,0,0,0,253,0,0,0,122,0,5,0,196,0,197,0,240,0,118,0,64,0,158,0,0,0,235,0,0,0,53,0,197,0,253,0,153,0,29,0,254,0,144,0,0,0,70,0,201,0,0,0,46,0,138,0,95,0,136,0,238,0,200,0,80,0,8,0,0,0,122,0,0,0,50,0,132,0,26,0,64,0,69,0,240,0,128,0,122,0,84,0,13,0,35,0,238,0,165,0,197,0,231,0,208,0,21,0,78,0,159,0,0,0,239,0,239,0,107,0,0,0,18,0,55,0,17,0,94,0,140,0,165,0,172,0,0,0,223,0,114,0,91,0,244,0,0,0,0,0,47,0,254,0,160,0,199,0,0,0,12,0,7,0,0,0,150,0,177,0,197,0,72,0,195,0,139,0,102,0,141,0,119,0,53,0,0,0,211,0,53,0,164,0,167,0,109,0,231,0,53,0,194,0,63,0,0,0,151,0,126,0,135,0,40,0,252,0,72,0,0,0,13,0,83,0,0,0,19,0,181,0,0,0,59,0,0,0,78,0,101,0,169,0,66,0,132,0,0,0,164,0,0,0,197,0,235,0,205,0,191,0,0,0,236,0,206,0,75,0,111,0,99,0,30,0,194,0,195,0,0,0,0,0,223,0,187,0,100,0,200,0,12,0,190,0,141,0,131,0,188,0,66,0,0,0,246,0,103,0,89,0,187,0,193,0,74,0,0,0,0,0,48,0,57,0,146,0,148,0,45,0,216,0,61,0,93,0,110,0,213,0,214,0,117,0,0,0,0,0,46,0,176,0,0,0,246,0,97,0,207,0,238,0,88,0,0,0,235,0,218,0,114,0,202,0,209,0,110,0,0,0,0,0,249,0,32,0,229,0,0,0,144,0,8,0,225,0,98,0,0,0,246,0,207,0,40,0,230,0,189,0,221,0,46,0,108,0,188,0,0,0,64,0,0,0,0,0,0,0,0,0,50,0,31,0,248,0,21,0,251,0,0,0,1,0,208,0,40,0,67,0,217,0,206,0,155,0,38,0,142,0,17,0,0,0,0,0,101,0,180,0,141,0,84,0,0,0,0,0,89,0,0,0,112,0,0,0,117,0,231,0,196,0,104,0,0,0,174,0,0,0,13,0,0,0,126,0,38,0,253,0,54,0,253,0,49,0,73,0,142,0,178,0,75,0,178,0,0,0,177,0,220,0,239,0,0,0,58,0,0,0,10,0,120,0,7,0,137,0,0,0,66,0,0,0,121,0,241,0,0,0,150,0,207,0,209,0,75,0,87,0,0,0,88,0,32,0,103,0,196,0,214,0,180,0,0,0,132,0,26,0,253,0,43,0,182,0,73,0,140,0,59,0,24,0,0,0,88,0,149,0,0,0,8,0,185,0,215,0,30,0,0,0,26,0,51,0,88,0,191,0,0,0,234,0,211,0,210,0,238,0,0,0,0,0,0,0,200,0,82,0,89,0,86,0,186,0,0,0,90,0,241,0,0,0,34,0,0,0,61,0,80,0,187,0,0,0,0,0,1,0,0,0,0,0,170,0,123,0,205,0,0,0,42,0,114,0,204,0,59,0,0,0,126,0,173,0,0,0);
signal scenario_full  : scenario_type := (0,0,111,31,206,31,75,31,23,31,197,31,197,30,102,31,137,31,88,31,93,31,233,31,143,31,143,30,3,31,56,31,56,30,190,31,190,31,188,31,71,31,168,31,114,31,114,30,114,29,230,31,230,31,54,31,54,30,146,31,195,31,92,31,88,31,82,31,129,31,111,31,172,31,155,31,75,31,49,31,118,31,101,31,72,31,206,31,84,31,84,30,186,31,188,31,242,31,94,31,170,31,97,31,128,31,128,30,188,31,102,31,236,31,197,31,197,30,55,31,122,31,81,31,181,31,168,31,161,31,56,31,56,30,41,31,211,31,32,31,141,31,182,31,178,31,106,31,35,31,211,31,45,31,184,31,200,31,209,31,131,31,131,30,131,29,100,31,186,31,232,31,25,31,170,31,237,31,109,31,174,31,138,31,138,30,62,31,180,31,163,31,245,31,28,31,30,31,151,31,65,31,65,30,235,31,63,31,66,31,239,31,253,31,109,31,192,31,28,31,229,31,50,31,218,31,214,31,204,31,57,31,9,31,9,31,108,31,226,31,226,30,118,31,131,31,131,30,253,31,253,30,122,31,5,31,196,31,197,31,240,31,118,31,64,31,158,31,158,30,235,31,235,30,53,31,197,31,253,31,153,31,29,31,254,31,144,31,144,30,70,31,201,31,201,30,46,31,138,31,95,31,136,31,238,31,200,31,80,31,8,31,8,30,122,31,122,30,50,31,132,31,26,31,64,31,69,31,240,31,128,31,122,31,84,31,13,31,35,31,238,31,165,31,197,31,231,31,208,31,21,31,78,31,159,31,159,30,239,31,239,31,107,31,107,30,18,31,55,31,17,31,94,31,140,31,165,31,172,31,172,30,223,31,114,31,91,31,244,31,244,30,244,29,47,31,254,31,160,31,199,31,199,30,12,31,7,31,7,30,150,31,177,31,197,31,72,31,195,31,139,31,102,31,141,31,119,31,53,31,53,30,211,31,53,31,164,31,167,31,109,31,231,31,53,31,194,31,63,31,63,30,151,31,126,31,135,31,40,31,252,31,72,31,72,30,13,31,83,31,83,30,19,31,181,31,181,30,59,31,59,30,78,31,101,31,169,31,66,31,132,31,132,30,164,31,164,30,197,31,235,31,205,31,191,31,191,30,236,31,206,31,75,31,111,31,99,31,30,31,194,31,195,31,195,30,195,29,223,31,187,31,100,31,200,31,12,31,190,31,141,31,131,31,188,31,66,31,66,30,246,31,103,31,89,31,187,31,193,31,74,31,74,30,74,29,48,31,57,31,146,31,148,31,45,31,216,31,61,31,93,31,110,31,213,31,214,31,117,31,117,30,117,29,46,31,176,31,176,30,246,31,97,31,207,31,238,31,88,31,88,30,235,31,218,31,114,31,202,31,209,31,110,31,110,30,110,29,249,31,32,31,229,31,229,30,144,31,8,31,225,31,98,31,98,30,246,31,207,31,40,31,230,31,189,31,221,31,46,31,108,31,188,31,188,30,64,31,64,30,64,29,64,28,64,27,50,31,31,31,248,31,21,31,251,31,251,30,1,31,208,31,40,31,67,31,217,31,206,31,155,31,38,31,142,31,17,31,17,30,17,29,101,31,180,31,141,31,84,31,84,30,84,29,89,31,89,30,112,31,112,30,117,31,231,31,196,31,104,31,104,30,174,31,174,30,13,31,13,30,126,31,38,31,253,31,54,31,253,31,49,31,73,31,142,31,178,31,75,31,178,31,178,30,177,31,220,31,239,31,239,30,58,31,58,30,10,31,120,31,7,31,137,31,137,30,66,31,66,30,121,31,241,31,241,30,150,31,207,31,209,31,75,31,87,31,87,30,88,31,32,31,103,31,196,31,214,31,180,31,180,30,132,31,26,31,253,31,43,31,182,31,73,31,140,31,59,31,24,31,24,30,88,31,149,31,149,30,8,31,185,31,215,31,30,31,30,30,26,31,51,31,88,31,191,31,191,30,234,31,211,31,210,31,238,31,238,30,238,29,238,28,200,31,82,31,89,31,86,31,186,31,186,30,90,31,241,31,241,30,34,31,34,30,61,31,80,31,187,31,187,30,187,29,1,31,1,30,1,29,170,31,123,31,205,31,205,30,42,31,114,31,204,31,59,31,59,30,126,31,173,31,173,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
