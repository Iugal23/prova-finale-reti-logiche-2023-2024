-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 990;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (185,0,201,0,75,0,142,0,3,0,0,0,165,0,0,0,189,0,233,0,83,0,203,0,134,0,162,0,244,0,166,0,182,0,212,0,0,0,114,0,0,0,248,0,72,0,45,0,136,0,0,0,12,0,149,0,2,0,142,0,0,0,0,0,45,0,1,0,0,0,97,0,224,0,147,0,62,0,153,0,39,0,86,0,124,0,242,0,0,0,32,0,231,0,0,0,92,0,188,0,54,0,178,0,0,0,105,0,0,0,107,0,8,0,0,0,151,0,225,0,19,0,79,0,223,0,178,0,0,0,149,0,222,0,252,0,240,0,112,0,200,0,0,0,39,0,0,0,54,0,66,0,107,0,147,0,0,0,54,0,0,0,0,0,0,0,45,0,168,0,228,0,20,0,213,0,158,0,109,0,73,0,0,0,0,0,3,0,117,0,0,0,220,0,0,0,173,0,236,0,89,0,0,0,162,0,112,0,250,0,230,0,0,0,206,0,165,0,174,0,125,0,246,0,233,0,201,0,0,0,37,0,0,0,219,0,70,0,46,0,13,0,157,0,70,0,65,0,157,0,150,0,121,0,144,0,196,0,195,0,78,0,0,0,36,0,174,0,0,0,255,0,153,0,82,0,211,0,0,0,0,0,117,0,50,0,143,0,0,0,165,0,199,0,51,0,171,0,0,0,56,0,93,0,0,0,0,0,56,0,148,0,91,0,0,0,0,0,0,0,186,0,0,0,0,0,38,0,0,0,33,0,128,0,55,0,81,0,102,0,31,0,45,0,115,0,91,0,68,0,11,0,0,0,0,0,169,0,0,0,105,0,0,0,42,0,110,0,0,0,224,0,0,0,141,0,149,0,0,0,105,0,223,0,74,0,24,0,117,0,213,0,167,0,30,0,182,0,57,0,255,0,250,0,121,0,13,0,18,0,84,0,51,0,214,0,17,0,137,0,0,0,6,0,59,0,87,0,125,0,30,0,241,0,94,0,82,0,39,0,208,0,234,0,56,0,235,0,150,0,140,0,0,0,0,0,82,0,7,0,237,0,201,0,223,0,0,0,0,0,0,0,132,0,160,0,66,0,114,0,186,0,0,0,109,0,74,0,0,0,0,0,150,0,107,0,192,0,46,0,33,0,17,0,0,0,11,0,0,0,144,0,0,0,32,0,0,0,213,0,0,0,170,0,55,0,239,0,176,0,47,0,111,0,36,0,82,0,69,0,97,0,151,0,0,0,68,0,172,0,0,0,48,0,0,0,199,0,54,0,211,0,18,0,34,0,0,0,27,0,10,0,0,0,0,0,79,0,11,0,236,0,215,0,125,0,69,0,0,0,97,0,4,0,178,0,111,0,231,0,66,0,184,0,52,0,99,0,157,0,0,0,21,0,75,0,64,0,96,0,124,0,46,0,64,0,80,0,91,0,120,0,0,0,0,0,26,0,164,0,0,0,239,0,0,0,70,0,100,0,0,0,193,0,247,0,181,0,0,0,84,0,84,0,214,0,133,0,29,0,0,0,16,0,176,0,14,0,204,0,232,0,27,0,185,0,225,0,0,0,101,0,37,0,32,0,165,0,231,0,129,0,198,0,66,0,55,0,53,0,202,0,19,0,0,0,0,0,222,0,0,0,113,0,0,0,24,0,103,0,211,0,113,0,81,0,60,0,206,0,145,0,0,0,0,0,63,0,14,0,0,0,189,0,0,0,125,0,88,0,193,0,237,0,0,0,0,0,140,0,0,0,59,0,0,0,0,0,37,0,69,0,21,0,71,0,178,0,66,0,0,0,207,0,0,0,60,0,106,0,0,0,200,0,224,0,0,0,25,0,23,0,90,0,0,0,217,0,177,0,129,0,247,0,0,0,163,0,99,0,156,0,105,0,80,0,95,0,14,0,0,0,0,0,15,0,33,0,0,0,171,0,2,0,42,0,99,0,1,0,233,0,0,0,157,0,73,0,216,0,0,0,60,0,20,0,36,0,169,0,0,0,189,0,234,0,0,0,196,0,0,0,122,0,0,0,225,0,135,0,178,0,125,0,148,0,135,0,103,0,14,0,165,0,236,0,234,0,249,0,165,0,67,0,173,0,17,0,0,0,156,0,14,0,0,0,168,0,0,0,0,0,205,0,173,0,186,0,172,0,226,0,196,0,0,0,0,0,141,0,143,0,137,0,40,0,190,0,242,0,230,0,104,0,13,0,171,0,18,0,0,0,218,0,221,0,245,0,102,0,0,0,13,0,189,0,115,0,158,0,0,0,173,0,121,0,59,0,0,0,0,0,91,0,111,0,232,0,0,0,27,0,45,0,114,0,240,0,139,0,150,0,120,0,167,0,135,0,0,0,0,0,0,0,0,0,0,0,207,0,250,0,37,0,240,0,0,0,81,0,38,0,195,0,113,0,233,0,31,0,113,0,2,0,98,0,87,0,192,0,30,0,166,0,125,0,127,0,0,0,0,0,87,0,211,0,166,0,2,0,63,0,0,0,227,0,194,0,36,0,70,0,164,0,55,0,142,0,34,0,24,0,185,0,0,0,0,0,28,0,174,0,28,0,20,0,35,0,213,0,235,0,2,0,67,0,156,0,232,0,0,0,0,0,122,0,253,0,50,0,34,0,74,0,239,0,89,0,8,0,247,0,0,0,184,0,146,0,11,0,204,0,0,0,135,0,30,0,104,0,0,0,0,0,129,0,1,0,2,0,65,0,221,0,129,0,39,0,127,0,0,0,38,0,219,0,69,0,176,0,88,0,157,0,157,0,233,0,71,0,89,0,0,0,132,0,150,0,155,0,65,0,0,0,129,0,220,0,125,0,29,0,0,0,212,0,192,0,71,0,79,0,242,0,28,0,101,0,76,0,0,0,161,0,0,0,0,0,0,0,211,0,174,0,18,0,0,0,136,0,215,0,60,0,129,0,0,0,0,0,212,0,206,0,0,0,44,0,113,0,137,0,16,0,224,0,74,0,0,0,149,0,173,0,0,0,203,0,111,0,134,0,88,0,169,0,0,0,162,0,109,0,88,0,0,0,36,0,0,0,103,0,39,0,0,0,196,0,181,0,36,0,243,0,0,0,230,0,25,0,0,0,98,0,0,0,14,0,45,0,0,0,0,0,0,0,29,0,236,0,214,0,208,0,254,0,89,0,251,0,111,0,109,0,24,0,0,0,44,0,103,0,198,0,0,0,193,0,0,0,87,0,22,0,217,0,27,0,0,0,0,0,39,0,225,0,53,0,20,0,29,0,147,0,253,0,174,0,103,0,144,0,7,0,9,0,216,0,0,0,138,0,85,0,0,0,112,0,160,0,164,0,81,0,0,0,0,0,130,0,47,0,0,0,135,0,228,0,26,0,22,0,43,0,221,0,0,0,149,0,132,0,155,0,85,0,107,0,161,0,0,0,112,0,0,0,169,0,45,0,97,0,0,0,53,0,228,0,174,0,0,0,161,0,146,0,29,0,0,0,75,0,26,0,235,0,0,0,189,0,0,0,243,0,98,0,0,0,150,0,131,0,127,0,0,0,81,0,106,0,12,0,155,0,150,0,236,0,152,0,0,0,222,0,188,0,177,0,0,0,219,0,174,0,231,0,229,0,23,0,163,0,11,0,167,0,10,0,231,0,11,0,50,0,79,0,167,0,73,0,89,0,0,0,72,0,251,0,82,0,117,0,13,0,174,0,132,0,21,0,238,0,9,0,71,0,0,0,0,0,0,0,74,0,192,0,0,0,197,0,0,0,74,0,135,0,84,0,165,0,103,0,186,0,94,0,250,0,228,0,118,0,27,0,38,0,20,0,0,0,0,0,176,0,72,0,0,0,61,0,13,0,248,0,164,0,208,0,119,0,0,0,39,0,101,0,24,0,0,0,107,0,87,0,0,0,238,0,144,0,21,0,76,0,17,0,0,0,72,0,0,0,80,0,0,0,129,0,0,0,231,0,0,0,161,0,73,0,173,0,0,0,64,0,178,0,0,0,239,0,0,0,11,0,0,0,215,0,198,0,31,0,0,0,0,0,184,0,11,0,26,0,7,0,223,0,128,0,207,0,146,0,206,0,227,0,238,0,43,0,211,0,4,0,0,0,0,0,102,0,124,0,34,0,153,0,106,0,7,0,220,0,122,0,139,0,0,0,193,0,55,0,63,0,40,0,47,0,141,0,234,0,218,0,61,0,101,0,111,0,185,0,247,0,248,0,0,0,0,0,34,0,30,0,42,0,136,0,0,0,229,0,0,0,190,0,78,0,110,0,0,0,0,0,0,0,2,0,21,0,202,0,165,0,151,0,221,0,42,0,0,0,205,0,119,0,222,0,240,0,4,0,191,0,108,0,74,0,185,0,237,0,50,0,205,0,108,0,110,0,126,0,204,0,231,0,12,0,58,0,0,0,69,0,11,0,161,0,177,0,12,0,232,0,34,0,178,0,153,0,247,0,59,0,76,0,240,0,0,0);
signal scenario_full  : scenario_type := (185,31,201,31,75,31,142,31,3,31,3,30,165,31,165,30,189,31,233,31,83,31,203,31,134,31,162,31,244,31,166,31,182,31,212,31,212,30,114,31,114,30,248,31,72,31,45,31,136,31,136,30,12,31,149,31,2,31,142,31,142,30,142,29,45,31,1,31,1,30,97,31,224,31,147,31,62,31,153,31,39,31,86,31,124,31,242,31,242,30,32,31,231,31,231,30,92,31,188,31,54,31,178,31,178,30,105,31,105,30,107,31,8,31,8,30,151,31,225,31,19,31,79,31,223,31,178,31,178,30,149,31,222,31,252,31,240,31,112,31,200,31,200,30,39,31,39,30,54,31,66,31,107,31,147,31,147,30,54,31,54,30,54,29,54,28,45,31,168,31,228,31,20,31,213,31,158,31,109,31,73,31,73,30,73,29,3,31,117,31,117,30,220,31,220,30,173,31,236,31,89,31,89,30,162,31,112,31,250,31,230,31,230,30,206,31,165,31,174,31,125,31,246,31,233,31,201,31,201,30,37,31,37,30,219,31,70,31,46,31,13,31,157,31,70,31,65,31,157,31,150,31,121,31,144,31,196,31,195,31,78,31,78,30,36,31,174,31,174,30,255,31,153,31,82,31,211,31,211,30,211,29,117,31,50,31,143,31,143,30,165,31,199,31,51,31,171,31,171,30,56,31,93,31,93,30,93,29,56,31,148,31,91,31,91,30,91,29,91,28,186,31,186,30,186,29,38,31,38,30,33,31,128,31,55,31,81,31,102,31,31,31,45,31,115,31,91,31,68,31,11,31,11,30,11,29,169,31,169,30,105,31,105,30,42,31,110,31,110,30,224,31,224,30,141,31,149,31,149,30,105,31,223,31,74,31,24,31,117,31,213,31,167,31,30,31,182,31,57,31,255,31,250,31,121,31,13,31,18,31,84,31,51,31,214,31,17,31,137,31,137,30,6,31,59,31,87,31,125,31,30,31,241,31,94,31,82,31,39,31,208,31,234,31,56,31,235,31,150,31,140,31,140,30,140,29,82,31,7,31,237,31,201,31,223,31,223,30,223,29,223,28,132,31,160,31,66,31,114,31,186,31,186,30,109,31,74,31,74,30,74,29,150,31,107,31,192,31,46,31,33,31,17,31,17,30,11,31,11,30,144,31,144,30,32,31,32,30,213,31,213,30,170,31,55,31,239,31,176,31,47,31,111,31,36,31,82,31,69,31,97,31,151,31,151,30,68,31,172,31,172,30,48,31,48,30,199,31,54,31,211,31,18,31,34,31,34,30,27,31,10,31,10,30,10,29,79,31,11,31,236,31,215,31,125,31,69,31,69,30,97,31,4,31,178,31,111,31,231,31,66,31,184,31,52,31,99,31,157,31,157,30,21,31,75,31,64,31,96,31,124,31,46,31,64,31,80,31,91,31,120,31,120,30,120,29,26,31,164,31,164,30,239,31,239,30,70,31,100,31,100,30,193,31,247,31,181,31,181,30,84,31,84,31,214,31,133,31,29,31,29,30,16,31,176,31,14,31,204,31,232,31,27,31,185,31,225,31,225,30,101,31,37,31,32,31,165,31,231,31,129,31,198,31,66,31,55,31,53,31,202,31,19,31,19,30,19,29,222,31,222,30,113,31,113,30,24,31,103,31,211,31,113,31,81,31,60,31,206,31,145,31,145,30,145,29,63,31,14,31,14,30,189,31,189,30,125,31,88,31,193,31,237,31,237,30,237,29,140,31,140,30,59,31,59,30,59,29,37,31,69,31,21,31,71,31,178,31,66,31,66,30,207,31,207,30,60,31,106,31,106,30,200,31,224,31,224,30,25,31,23,31,90,31,90,30,217,31,177,31,129,31,247,31,247,30,163,31,99,31,156,31,105,31,80,31,95,31,14,31,14,30,14,29,15,31,33,31,33,30,171,31,2,31,42,31,99,31,1,31,233,31,233,30,157,31,73,31,216,31,216,30,60,31,20,31,36,31,169,31,169,30,189,31,234,31,234,30,196,31,196,30,122,31,122,30,225,31,135,31,178,31,125,31,148,31,135,31,103,31,14,31,165,31,236,31,234,31,249,31,165,31,67,31,173,31,17,31,17,30,156,31,14,31,14,30,168,31,168,30,168,29,205,31,173,31,186,31,172,31,226,31,196,31,196,30,196,29,141,31,143,31,137,31,40,31,190,31,242,31,230,31,104,31,13,31,171,31,18,31,18,30,218,31,221,31,245,31,102,31,102,30,13,31,189,31,115,31,158,31,158,30,173,31,121,31,59,31,59,30,59,29,91,31,111,31,232,31,232,30,27,31,45,31,114,31,240,31,139,31,150,31,120,31,167,31,135,31,135,30,135,29,135,28,135,27,135,26,207,31,250,31,37,31,240,31,240,30,81,31,38,31,195,31,113,31,233,31,31,31,113,31,2,31,98,31,87,31,192,31,30,31,166,31,125,31,127,31,127,30,127,29,87,31,211,31,166,31,2,31,63,31,63,30,227,31,194,31,36,31,70,31,164,31,55,31,142,31,34,31,24,31,185,31,185,30,185,29,28,31,174,31,28,31,20,31,35,31,213,31,235,31,2,31,67,31,156,31,232,31,232,30,232,29,122,31,253,31,50,31,34,31,74,31,239,31,89,31,8,31,247,31,247,30,184,31,146,31,11,31,204,31,204,30,135,31,30,31,104,31,104,30,104,29,129,31,1,31,2,31,65,31,221,31,129,31,39,31,127,31,127,30,38,31,219,31,69,31,176,31,88,31,157,31,157,31,233,31,71,31,89,31,89,30,132,31,150,31,155,31,65,31,65,30,129,31,220,31,125,31,29,31,29,30,212,31,192,31,71,31,79,31,242,31,28,31,101,31,76,31,76,30,161,31,161,30,161,29,161,28,211,31,174,31,18,31,18,30,136,31,215,31,60,31,129,31,129,30,129,29,212,31,206,31,206,30,44,31,113,31,137,31,16,31,224,31,74,31,74,30,149,31,173,31,173,30,203,31,111,31,134,31,88,31,169,31,169,30,162,31,109,31,88,31,88,30,36,31,36,30,103,31,39,31,39,30,196,31,181,31,36,31,243,31,243,30,230,31,25,31,25,30,98,31,98,30,14,31,45,31,45,30,45,29,45,28,29,31,236,31,214,31,208,31,254,31,89,31,251,31,111,31,109,31,24,31,24,30,44,31,103,31,198,31,198,30,193,31,193,30,87,31,22,31,217,31,27,31,27,30,27,29,39,31,225,31,53,31,20,31,29,31,147,31,253,31,174,31,103,31,144,31,7,31,9,31,216,31,216,30,138,31,85,31,85,30,112,31,160,31,164,31,81,31,81,30,81,29,130,31,47,31,47,30,135,31,228,31,26,31,22,31,43,31,221,31,221,30,149,31,132,31,155,31,85,31,107,31,161,31,161,30,112,31,112,30,169,31,45,31,97,31,97,30,53,31,228,31,174,31,174,30,161,31,146,31,29,31,29,30,75,31,26,31,235,31,235,30,189,31,189,30,243,31,98,31,98,30,150,31,131,31,127,31,127,30,81,31,106,31,12,31,155,31,150,31,236,31,152,31,152,30,222,31,188,31,177,31,177,30,219,31,174,31,231,31,229,31,23,31,163,31,11,31,167,31,10,31,231,31,11,31,50,31,79,31,167,31,73,31,89,31,89,30,72,31,251,31,82,31,117,31,13,31,174,31,132,31,21,31,238,31,9,31,71,31,71,30,71,29,71,28,74,31,192,31,192,30,197,31,197,30,74,31,135,31,84,31,165,31,103,31,186,31,94,31,250,31,228,31,118,31,27,31,38,31,20,31,20,30,20,29,176,31,72,31,72,30,61,31,13,31,248,31,164,31,208,31,119,31,119,30,39,31,101,31,24,31,24,30,107,31,87,31,87,30,238,31,144,31,21,31,76,31,17,31,17,30,72,31,72,30,80,31,80,30,129,31,129,30,231,31,231,30,161,31,73,31,173,31,173,30,64,31,178,31,178,30,239,31,239,30,11,31,11,30,215,31,198,31,31,31,31,30,31,29,184,31,11,31,26,31,7,31,223,31,128,31,207,31,146,31,206,31,227,31,238,31,43,31,211,31,4,31,4,30,4,29,102,31,124,31,34,31,153,31,106,31,7,31,220,31,122,31,139,31,139,30,193,31,55,31,63,31,40,31,47,31,141,31,234,31,218,31,61,31,101,31,111,31,185,31,247,31,248,31,248,30,248,29,34,31,30,31,42,31,136,31,136,30,229,31,229,30,190,31,78,31,110,31,110,30,110,29,110,28,2,31,21,31,202,31,165,31,151,31,221,31,42,31,42,30,205,31,119,31,222,31,240,31,4,31,191,31,108,31,74,31,185,31,237,31,50,31,205,31,108,31,110,31,126,31,204,31,231,31,12,31,58,31,58,30,69,31,11,31,161,31,177,31,12,31,232,31,34,31,178,31,153,31,247,31,59,31,76,31,240,31,240,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
