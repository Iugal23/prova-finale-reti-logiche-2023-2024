-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 416;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (38,0,2,0,0,0,253,0,134,0,82,0,169,0,56,0,80,0,250,0,60,0,0,0,170,0,71,0,40,0,49,0,200,0,50,0,0,0,235,0,14,0,91,0,67,0,95,0,131,0,0,0,162,0,244,0,98,0,150,0,0,0,157,0,0,0,150,0,214,0,224,0,199,0,0,0,97,0,248,0,64,0,180,0,192,0,85,0,66,0,0,0,244,0,188,0,145,0,109,0,57,0,158,0,166,0,170,0,95,0,101,0,221,0,0,0,0,0,84,0,0,0,9,0,204,0,49,0,126,0,176,0,0,0,183,0,254,0,12,0,239,0,74,0,44,0,111,0,145,0,160,0,158,0,43,0,185,0,199,0,0,0,1,0,0,0,38,0,0,0,178,0,184,0,207,0,0,0,215,0,0,0,0,0,193,0,140,0,87,0,196,0,98,0,182,0,143,0,207,0,224,0,207,0,166,0,120,0,142,0,0,0,15,0,15,0,143,0,54,0,0,0,239,0,124,0,170,0,0,0,152,0,227,0,156,0,0,0,166,0,235,0,87,0,241,0,180,0,0,0,131,0,42,0,0,0,0,0,199,0,70,0,0,0,0,0,250,0,93,0,0,0,9,0,66,0,0,0,238,0,225,0,80,0,222,0,50,0,251,0,79,0,0,0,41,0,104,0,0,0,205,0,120,0,0,0,99,0,126,0,18,0,250,0,144,0,50,0,0,0,153,0,88,0,0,0,215,0,34,0,253,0,36,0,215,0,0,0,106,0,238,0,239,0,0,0,0,0,214,0,129,0,173,0,0,0,73,0,66,0,0,0,0,0,172,0,13,0,47,0,180,0,67,0,0,0,183,0,0,0,194,0,167,0,121,0,0,0,238,0,159,0,155,0,0,0,79,0,209,0,77,0,223,0,0,0,158,0,77,0,67,0,68,0,95,0,0,0,222,0,0,0,231,0,217,0,229,0,30,0,0,0,129,0,190,0,129,0,44,0,191,0,40,0,191,0,60,0,0,0,74,0,120,0,0,0,16,0,143,0,202,0,37,0,0,0,113,0,86,0,116,0,0,0,146,0,0,0,0,0,0,0,230,0,21,0,57,0,0,0,119,0,201,0,183,0,72,0,3,0,71,0,0,0,212,0,3,0,0,0,0,0,0,0,206,0,221,0,0,0,57,0,0,0,82,0,128,0,234,0,185,0,20,0,112,0,121,0,0,0,0,0,186,0,84,0,0,0,0,0,120,0,78,0,166,0,0,0,79,0,118,0,73,0,175,0,252,0,48,0,214,0,0,0,0,0,0,0,0,0,185,0,4,0,84,0,0,0,166,0,183,0,0,0,126,0,10,0,209,0,93,0,35,0,7,0,7,0,0,0,0,0,52,0,128,0,159,0,55,0,236,0,0,0,66,0,80,0,50,0,178,0,0,0,251,0,66,0,141,0,160,0,142,0,0,0,73,0,11,0,151,0,180,0,211,0,198,0,230,0,243,0,214,0,193,0,0,0,0,0,0,0,75,0,69,0,237,0,0,0,113,0,140,0,175,0,80,0,0,0,94,0,228,0,236,0,77,0,61,0,0,0,151,0,93,0,108,0,190,0,21,0,222,0,186,0,38,0,36,0,113,0,191,0,74,0,65,0,201,0,0,0,65,0,199,0,200,0,245,0,149,0,225,0,68,0,96,0,49,0,121,0,153,0,97,0,124,0,133,0,128,0,0,0,198,0,200,0,28,0,172,0,82,0,119,0,151,0,212,0,181,0,255,0,3,0,0,0,0,0,110,0,133,0,199,0,26,0,0,0,0,0,188,0,224,0,163,0,61,0,25,0,243,0,141,0,0,0,130,0,0,0,34,0,76,0,217,0,11,0,223,0);
signal scenario_full  : scenario_type := (38,31,2,31,2,30,253,31,134,31,82,31,169,31,56,31,80,31,250,31,60,31,60,30,170,31,71,31,40,31,49,31,200,31,50,31,50,30,235,31,14,31,91,31,67,31,95,31,131,31,131,30,162,31,244,31,98,31,150,31,150,30,157,31,157,30,150,31,214,31,224,31,199,31,199,30,97,31,248,31,64,31,180,31,192,31,85,31,66,31,66,30,244,31,188,31,145,31,109,31,57,31,158,31,166,31,170,31,95,31,101,31,221,31,221,30,221,29,84,31,84,30,9,31,204,31,49,31,126,31,176,31,176,30,183,31,254,31,12,31,239,31,74,31,44,31,111,31,145,31,160,31,158,31,43,31,185,31,199,31,199,30,1,31,1,30,38,31,38,30,178,31,184,31,207,31,207,30,215,31,215,30,215,29,193,31,140,31,87,31,196,31,98,31,182,31,143,31,207,31,224,31,207,31,166,31,120,31,142,31,142,30,15,31,15,31,143,31,54,31,54,30,239,31,124,31,170,31,170,30,152,31,227,31,156,31,156,30,166,31,235,31,87,31,241,31,180,31,180,30,131,31,42,31,42,30,42,29,199,31,70,31,70,30,70,29,250,31,93,31,93,30,9,31,66,31,66,30,238,31,225,31,80,31,222,31,50,31,251,31,79,31,79,30,41,31,104,31,104,30,205,31,120,31,120,30,99,31,126,31,18,31,250,31,144,31,50,31,50,30,153,31,88,31,88,30,215,31,34,31,253,31,36,31,215,31,215,30,106,31,238,31,239,31,239,30,239,29,214,31,129,31,173,31,173,30,73,31,66,31,66,30,66,29,172,31,13,31,47,31,180,31,67,31,67,30,183,31,183,30,194,31,167,31,121,31,121,30,238,31,159,31,155,31,155,30,79,31,209,31,77,31,223,31,223,30,158,31,77,31,67,31,68,31,95,31,95,30,222,31,222,30,231,31,217,31,229,31,30,31,30,30,129,31,190,31,129,31,44,31,191,31,40,31,191,31,60,31,60,30,74,31,120,31,120,30,16,31,143,31,202,31,37,31,37,30,113,31,86,31,116,31,116,30,146,31,146,30,146,29,146,28,230,31,21,31,57,31,57,30,119,31,201,31,183,31,72,31,3,31,71,31,71,30,212,31,3,31,3,30,3,29,3,28,206,31,221,31,221,30,57,31,57,30,82,31,128,31,234,31,185,31,20,31,112,31,121,31,121,30,121,29,186,31,84,31,84,30,84,29,120,31,78,31,166,31,166,30,79,31,118,31,73,31,175,31,252,31,48,31,214,31,214,30,214,29,214,28,214,27,185,31,4,31,84,31,84,30,166,31,183,31,183,30,126,31,10,31,209,31,93,31,35,31,7,31,7,31,7,30,7,29,52,31,128,31,159,31,55,31,236,31,236,30,66,31,80,31,50,31,178,31,178,30,251,31,66,31,141,31,160,31,142,31,142,30,73,31,11,31,151,31,180,31,211,31,198,31,230,31,243,31,214,31,193,31,193,30,193,29,193,28,75,31,69,31,237,31,237,30,113,31,140,31,175,31,80,31,80,30,94,31,228,31,236,31,77,31,61,31,61,30,151,31,93,31,108,31,190,31,21,31,222,31,186,31,38,31,36,31,113,31,191,31,74,31,65,31,201,31,201,30,65,31,199,31,200,31,245,31,149,31,225,31,68,31,96,31,49,31,121,31,153,31,97,31,124,31,133,31,128,31,128,30,198,31,200,31,28,31,172,31,82,31,119,31,151,31,212,31,181,31,255,31,3,31,3,30,3,29,110,31,133,31,199,31,26,31,26,30,26,29,188,31,224,31,163,31,61,31,25,31,243,31,141,31,141,30,130,31,130,30,34,31,76,31,217,31,11,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
