-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_734 is
end project_tb_734;

architecture project_tb_arch_734 of project_tb_734 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 637;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (226,0,26,0,71,0,255,0,227,0,0,0,0,0,13,0,134,0,0,0,0,0,88,0,122,0,250,0,0,0,65,0,189,0,213,0,178,0,90,0,79,0,217,0,102,0,77,0,8,0,96,0,0,0,252,0,0,0,0,0,51,0,22,0,70,0,0,0,0,0,90,0,0,0,56,0,210,0,62,0,0,0,144,0,2,0,190,0,60,0,21,0,0,0,122,0,0,0,67,0,28,0,72,0,55,0,0,0,50,0,220,0,76,0,100,0,105,0,250,0,142,0,0,0,187,0,158,0,0,0,182,0,10,0,161,0,90,0,0,0,0,0,69,0,5,0,138,0,72,0,220,0,50,0,4,0,163,0,0,0,214,0,123,0,136,0,0,0,0,0,9,0,204,0,237,0,0,0,156,0,239,0,98,0,17,0,101,0,253,0,162,0,209,0,0,0,27,0,118,0,118,0,0,0,71,0,0,0,0,0,64,0,0,0,246,0,72,0,200,0,110,0,41,0,0,0,0,0,139,0,101,0,0,0,0,0,0,0,0,0,157,0,63,0,159,0,144,0,201,0,25,0,222,0,0,0,63,0,223,0,57,0,6,0,0,0,129,0,34,0,139,0,165,0,140,0,0,0,124,0,0,0,0,0,31,0,75,0,34,0,35,0,123,0,38,0,0,0,1,0,124,0,229,0,0,0,20,0,14,0,164,0,0,0,0,0,61,0,213,0,109,0,126,0,157,0,135,0,205,0,110,0,234,0,64,0,79,0,0,0,119,0,8,0,233,0,227,0,176,0,0,0,43,0,198,0,192,0,109,0,148,0,93,0,149,0,5,0,0,0,60,0,237,0,0,0,26,0,108,0,242,0,158,0,27,0,39,0,181,0,190,0,0,0,223,0,191,0,69,0,232,0,0,0,83,0,0,0,0,0,0,0,222,0,19,0,115,0,224,0,251,0,0,0,0,0,117,0,48,0,3,0,217,0,0,0,150,0,0,0,0,0,0,0,226,0,78,0,49,0,124,0,7,0,59,0,0,0,176,0,127,0,162,0,0,0,205,0,192,0,168,0,125,0,135,0,209,0,124,0,95,0,250,0,130,0,123,0,7,0,111,0,69,0,0,0,190,0,0,0,0,0,124,0,246,0,123,0,4,0,61,0,27,0,0,0,192,0,0,0,0,0,105,0,87,0,167,0,52,0,233,0,108,0,196,0,46,0,129,0,0,0,218,0,146,0,213,0,33,0,0,0,105,0,201,0,40,0,208,0,145,0,190,0,137,0,47,0,118,0,136,0,236,0,0,0,1,0,166,0,24,0,122,0,114,0,156,0,22,0,4,0,106,0,152,0,0,0,0,0,201,0,167,0,223,0,140,0,131,0,127,0,219,0,115,0,118,0,192,0,86,0,41,0,0,0,95,0,3,0,34,0,202,0,152,0,225,0,106,0,98,0,130,0,72,0,6,0,201,0,152,0,231,0,0,0,122,0,239,0,83,0,182,0,108,0,173,0,221,0,5,0,252,0,0,0,0,0,151,0,211,0,184,0,10,0,244,0,0,0,139,0,0,0,203,0,79,0,131,0,183,0,113,0,133,0,240,0,88,0,91,0,246,0,0,0,224,0,249,0,161,0,80,0,0,0,85,0,140,0,41,0,0,0,250,0,0,0,0,0,211,0,160,0,0,0,161,0,184,0,165,0,123,0,64,0,0,0,189,0,172,0,186,0,244,0,194,0,121,0,13,0,228,0,138,0,87,0,0,0,0,0,7,0,173,0,49,0,5,0,4,0,154,0,175,0,196,0,0,0,166,0,80,0,131,0,0,0,209,0,184,0,150,0,193,0,122,0,113,0,149,0,170,0,202,0,53,0,58,0,215,0,232,0,76,0,0,0,242,0,115,0,168,0,26,0,0,0,73,0,0,0,0,0,177,0,161,0,242,0,224,0,5,0,189,0,92,0,0,0,36,0,52,0,127,0,0,0,73,0,242,0,34,0,170,0,31,0,163,0,35,0,0,0,184,0,139,0,200,0,0,0,172,0,74,0,96,0,230,0,1,0,82,0,213,0,85,0,0,0,0,0,0,0,42,0,11,0,59,0,2,0,172,0,0,0,0,0,14,0,100,0,195,0,67,0,0,0,170,0,13,0,216,0,244,0,160,0,135,0,121,0,12,0,110,0,0,0,152,0,48,0,225,0,80,0,12,0,0,0,0,0,0,0,56,0,199,0,193,0,94,0,142,0,0,0,74,0,19,0,50,0,0,0,166,0,35,0,145,0,0,0,224,0,27,0,112,0,149,0,0,0,77,0,249,0,107,0,0,0,35,0,233,0,22,0,218,0,88,0,51,0,240,0,0,0,192,0,0,0,169,0,238,0,0,0,205,0,171,0,119,0,226,0,18,0,132,0,169,0,233,0,229,0,110,0,0,0,57,0,227,0,151,0,189,0,22,0,222,0,0,0,217,0,213,0,0,0,192,0,170,0,109,0,0,0,132,0,63,0,37,0,193,0,114,0,133,0,1,0,238,0,243,0,65,0,163,0,105,0,193,0,146,0,77,0,210,0,33,0,156,0,31,0,246,0,0,0,61,0,228,0,45,0,232,0,170,0,250,0,175,0,45,0,169,0,36,0,0,0,1,0,55,0,253,0,127,0,0,0,239,0,245,0,189,0,132,0,167,0,71,0,81,0,0,0,150,0,0,0,74,0,10,0,0,0,166,0,0,0,244,0,135,0,214,0,127,0,186,0,92,0,34,0,180,0,247,0,30,0,89,0,124,0,0,0,37,0,0,0,39,0,91,0,0,0,185,0,54,0,223,0,109,0,132,0,0,0,214,0,71,0,86,0,29,0,0,0,0,0,132,0,0,0);
signal scenario_full  : scenario_type := (226,31,26,31,71,31,255,31,227,31,227,30,227,29,13,31,134,31,134,30,134,29,88,31,122,31,250,31,250,30,65,31,189,31,213,31,178,31,90,31,79,31,217,31,102,31,77,31,8,31,96,31,96,30,252,31,252,30,252,29,51,31,22,31,70,31,70,30,70,29,90,31,90,30,56,31,210,31,62,31,62,30,144,31,2,31,190,31,60,31,21,31,21,30,122,31,122,30,67,31,28,31,72,31,55,31,55,30,50,31,220,31,76,31,100,31,105,31,250,31,142,31,142,30,187,31,158,31,158,30,182,31,10,31,161,31,90,31,90,30,90,29,69,31,5,31,138,31,72,31,220,31,50,31,4,31,163,31,163,30,214,31,123,31,136,31,136,30,136,29,9,31,204,31,237,31,237,30,156,31,239,31,98,31,17,31,101,31,253,31,162,31,209,31,209,30,27,31,118,31,118,31,118,30,71,31,71,30,71,29,64,31,64,30,246,31,72,31,200,31,110,31,41,31,41,30,41,29,139,31,101,31,101,30,101,29,101,28,101,27,157,31,63,31,159,31,144,31,201,31,25,31,222,31,222,30,63,31,223,31,57,31,6,31,6,30,129,31,34,31,139,31,165,31,140,31,140,30,124,31,124,30,124,29,31,31,75,31,34,31,35,31,123,31,38,31,38,30,1,31,124,31,229,31,229,30,20,31,14,31,164,31,164,30,164,29,61,31,213,31,109,31,126,31,157,31,135,31,205,31,110,31,234,31,64,31,79,31,79,30,119,31,8,31,233,31,227,31,176,31,176,30,43,31,198,31,192,31,109,31,148,31,93,31,149,31,5,31,5,30,60,31,237,31,237,30,26,31,108,31,242,31,158,31,27,31,39,31,181,31,190,31,190,30,223,31,191,31,69,31,232,31,232,30,83,31,83,30,83,29,83,28,222,31,19,31,115,31,224,31,251,31,251,30,251,29,117,31,48,31,3,31,217,31,217,30,150,31,150,30,150,29,150,28,226,31,78,31,49,31,124,31,7,31,59,31,59,30,176,31,127,31,162,31,162,30,205,31,192,31,168,31,125,31,135,31,209,31,124,31,95,31,250,31,130,31,123,31,7,31,111,31,69,31,69,30,190,31,190,30,190,29,124,31,246,31,123,31,4,31,61,31,27,31,27,30,192,31,192,30,192,29,105,31,87,31,167,31,52,31,233,31,108,31,196,31,46,31,129,31,129,30,218,31,146,31,213,31,33,31,33,30,105,31,201,31,40,31,208,31,145,31,190,31,137,31,47,31,118,31,136,31,236,31,236,30,1,31,166,31,24,31,122,31,114,31,156,31,22,31,4,31,106,31,152,31,152,30,152,29,201,31,167,31,223,31,140,31,131,31,127,31,219,31,115,31,118,31,192,31,86,31,41,31,41,30,95,31,3,31,34,31,202,31,152,31,225,31,106,31,98,31,130,31,72,31,6,31,201,31,152,31,231,31,231,30,122,31,239,31,83,31,182,31,108,31,173,31,221,31,5,31,252,31,252,30,252,29,151,31,211,31,184,31,10,31,244,31,244,30,139,31,139,30,203,31,79,31,131,31,183,31,113,31,133,31,240,31,88,31,91,31,246,31,246,30,224,31,249,31,161,31,80,31,80,30,85,31,140,31,41,31,41,30,250,31,250,30,250,29,211,31,160,31,160,30,161,31,184,31,165,31,123,31,64,31,64,30,189,31,172,31,186,31,244,31,194,31,121,31,13,31,228,31,138,31,87,31,87,30,87,29,7,31,173,31,49,31,5,31,4,31,154,31,175,31,196,31,196,30,166,31,80,31,131,31,131,30,209,31,184,31,150,31,193,31,122,31,113,31,149,31,170,31,202,31,53,31,58,31,215,31,232,31,76,31,76,30,242,31,115,31,168,31,26,31,26,30,73,31,73,30,73,29,177,31,161,31,242,31,224,31,5,31,189,31,92,31,92,30,36,31,52,31,127,31,127,30,73,31,242,31,34,31,170,31,31,31,163,31,35,31,35,30,184,31,139,31,200,31,200,30,172,31,74,31,96,31,230,31,1,31,82,31,213,31,85,31,85,30,85,29,85,28,42,31,11,31,59,31,2,31,172,31,172,30,172,29,14,31,100,31,195,31,67,31,67,30,170,31,13,31,216,31,244,31,160,31,135,31,121,31,12,31,110,31,110,30,152,31,48,31,225,31,80,31,12,31,12,30,12,29,12,28,56,31,199,31,193,31,94,31,142,31,142,30,74,31,19,31,50,31,50,30,166,31,35,31,145,31,145,30,224,31,27,31,112,31,149,31,149,30,77,31,249,31,107,31,107,30,35,31,233,31,22,31,218,31,88,31,51,31,240,31,240,30,192,31,192,30,169,31,238,31,238,30,205,31,171,31,119,31,226,31,18,31,132,31,169,31,233,31,229,31,110,31,110,30,57,31,227,31,151,31,189,31,22,31,222,31,222,30,217,31,213,31,213,30,192,31,170,31,109,31,109,30,132,31,63,31,37,31,193,31,114,31,133,31,1,31,238,31,243,31,65,31,163,31,105,31,193,31,146,31,77,31,210,31,33,31,156,31,31,31,246,31,246,30,61,31,228,31,45,31,232,31,170,31,250,31,175,31,45,31,169,31,36,31,36,30,1,31,55,31,253,31,127,31,127,30,239,31,245,31,189,31,132,31,167,31,71,31,81,31,81,30,150,31,150,30,74,31,10,31,10,30,166,31,166,30,244,31,135,31,214,31,127,31,186,31,92,31,34,31,180,31,247,31,30,31,89,31,124,31,124,30,37,31,37,30,39,31,91,31,91,30,185,31,54,31,223,31,109,31,132,31,132,30,214,31,71,31,86,31,29,31,29,30,29,29,132,31,132,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
