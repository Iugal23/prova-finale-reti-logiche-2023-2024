-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 651;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (141,0,210,0,174,0,69,0,75,0,61,0,207,0,104,0,0,0,0,0,151,0,80,0,181,0,0,0,0,0,247,0,0,0,172,0,146,0,159,0,76,0,183,0,166,0,21,0,74,0,172,0,236,0,91,0,0,0,183,0,73,0,3,0,178,0,159,0,54,0,7,0,76,0,0,0,130,0,58,0,168,0,139,0,0,0,239,0,246,0,234,0,88,0,203,0,45,0,75,0,132,0,0,0,207,0,0,0,91,0,217,0,253,0,3,0,128,0,129,0,0,0,21,0,236,0,142,0,144,0,170,0,0,0,151,0,141,0,0,0,113,0,0,0,8,0,147,0,208,0,0,0,58,0,0,0,115,0,249,0,155,0,21,0,26,0,0,0,136,0,95,0,144,0,81,0,0,0,139,0,0,0,244,0,222,0,33,0,212,0,0,0,101,0,139,0,185,0,127,0,45,0,142,0,113,0,0,0,242,0,156,0,89,0,76,0,40,0,126,0,203,0,1,0,148,0,117,0,162,0,110,0,0,0,158,0,160,0,0,0,104,0,66,0,120,0,22,0,97,0,91,0,127,0,129,0,172,0,0,0,129,0,21,0,109,0,181,0,78,0,154,0,0,0,51,0,239,0,239,0,27,0,6,0,36,0,146,0,92,0,81,0,0,0,47,0,248,0,14,0,230,0,181,0,0,0,118,0,242,0,63,0,124,0,139,0,244,0,185,0,247,0,207,0,126,0,180,0,76,0,23,0,246,0,150,0,158,0,128,0,227,0,56,0,172,0,17,0,205,0,214,0,0,0,0,0,43,0,87,0,0,0,72,0,28,0,119,0,42,0,118,0,203,0,55,0,231,0,79,0,177,0,77,0,218,0,18,0,161,0,236,0,0,0,134,0,49,0,171,0,73,0,0,0,106,0,126,0,16,0,0,0,0,0,45,0,72,0,72,0,65,0,0,0,134,0,17,0,104,0,142,0,124,0,195,0,220,0,46,0,179,0,94,0,0,0,0,0,14,0,110,0,195,0,0,0,40,0,186,0,109,0,101,0,53,0,188,0,146,0,41,0,36,0,249,0,138,0,15,0,10,0,100,0,46,0,254,0,0,0,129,0,81,0,82,0,26,0,105,0,159,0,4,0,0,0,91,0,71,0,45,0,159,0,192,0,136,0,0,0,97,0,154,0,0,0,118,0,77,0,168,0,254,0,81,0,3,0,0,0,1,0,79,0,0,0,39,0,138,0,80,0,43,0,93,0,248,0,0,0,21,0,196,0,0,0,71,0,55,0,0,0,223,0,82,0,238,0,229,0,64,0,79,0,40,0,215,0,0,0,1,0,254,0,33,0,176,0,245,0,65,0,164,0,104,0,0,0,40,0,120,0,65,0,138,0,173,0,0,0,207,0,160,0,65,0,28,0,0,0,76,0,163,0,113,0,179,0,96,0,120,0,27,0,32,0,51,0,23,0,160,0,133,0,0,0,109,0,0,0,241,0,0,0,0,0,0,0,0,0,77,0,120,0,0,0,224,0,57,0,72,0,0,0,0,0,255,0,0,0,226,0,146,0,160,0,0,0,210,0,179,0,58,0,194,0,0,0,92,0,197,0,107,0,113,0,253,0,0,0,92,0,155,0,0,0,25,0,178,0,130,0,49,0,25,0,0,0,0,0,116,0,42,0,1,0,132,0,78,0,0,0,28,0,129,0,189,0,77,0,6,0,0,0,187,0,132,0,32,0,0,0,211,0,108,0,3,0,0,0,146,0,194,0,0,0,20,0,224,0,98,0,216,0,0,0,0,0,0,0,210,0,171,0,154,0,182,0,91,0,0,0,0,0,212,0,181,0,206,0,190,0,213,0,0,0,49,0,225,0,27,0,163,0,74,0,67,0,166,0,31,0,173,0,154,0,238,0,0,0,253,0,0,0,216,0,6,0,177,0,36,0,159,0,107,0,111,0,160,0,157,0,0,0,0,0,0,0,0,0,45,0,52,0,0,0,108,0,0,0,0,0,207,0,0,0,102,0,216,0,169,0,0,0,241,0,95,0,79,0,174,0,0,0,0,0,0,0,167,0,160,0,154,0,105,0,44,0,0,0,35,0,117,0,65,0,31,0,0,0,193,0,97,0,132,0,155,0,128,0,212,0,223,0,3,0,3,0,235,0,133,0,129,0,79,0,0,0,49,0,47,0,58,0,35,0,214,0,204,0,175,0,128,0,164,0,79,0,113,0,57,0,196,0,253,0,197,0,75,0,0,0,176,0,0,0,213,0,218,0,0,0,1,0,8,0,0,0,115,0,0,0,0,0,251,0,0,0,112,0,221,0,183,0,250,0,19,0,130,0,7,0,156,0,0,0,205,0,251,0,223,0,62,0,87,0,36,0,248,0,0,0,15,0,128,0,244,0,213,0,81,0,209,0,9,0,0,0,62,0,245,0,172,0,0,0,17,0,0,0,207,0,119,0,0,0,0,0,12,0,0,0,72,0,121,0,0,0,66,0,0,0,222,0,33,0,226,0,226,0,208,0,57,0,0,0,183,0,251,0,76,0,249,0,71,0,0,0,0,0,69,0,212,0,0,0,122,0,0,0,174,0,0,0,84,0,0,0,96,0,207,0,24,0,51,0,0,0,22,0,0,0,89,0,0,0,61,0,168,0,117,0,216,0,106,0,72,0,110,0,63,0,6,0,35,0,71,0,220,0,48,0,0,0,143,0,106,0,0,0,160,0,245,0,176,0,186,0,105,0,74,0,0,0,246,0,170,0,58,0,230,0,220,0,248,0,14,0,11,0,22,0,132,0,0,0,33,0,164,0,0,0,0,0,162,0,0,0,57,0,20,0,151,0,16,0,227,0,216,0,208,0,103,0,136,0,107,0,237,0,180,0,86,0,185,0,242,0,15,0,142,0,25,0,1,0,0,0,0,0,188,0);
signal scenario_full  : scenario_type := (141,31,210,31,174,31,69,31,75,31,61,31,207,31,104,31,104,30,104,29,151,31,80,31,181,31,181,30,181,29,247,31,247,30,172,31,146,31,159,31,76,31,183,31,166,31,21,31,74,31,172,31,236,31,91,31,91,30,183,31,73,31,3,31,178,31,159,31,54,31,7,31,76,31,76,30,130,31,58,31,168,31,139,31,139,30,239,31,246,31,234,31,88,31,203,31,45,31,75,31,132,31,132,30,207,31,207,30,91,31,217,31,253,31,3,31,128,31,129,31,129,30,21,31,236,31,142,31,144,31,170,31,170,30,151,31,141,31,141,30,113,31,113,30,8,31,147,31,208,31,208,30,58,31,58,30,115,31,249,31,155,31,21,31,26,31,26,30,136,31,95,31,144,31,81,31,81,30,139,31,139,30,244,31,222,31,33,31,212,31,212,30,101,31,139,31,185,31,127,31,45,31,142,31,113,31,113,30,242,31,156,31,89,31,76,31,40,31,126,31,203,31,1,31,148,31,117,31,162,31,110,31,110,30,158,31,160,31,160,30,104,31,66,31,120,31,22,31,97,31,91,31,127,31,129,31,172,31,172,30,129,31,21,31,109,31,181,31,78,31,154,31,154,30,51,31,239,31,239,31,27,31,6,31,36,31,146,31,92,31,81,31,81,30,47,31,248,31,14,31,230,31,181,31,181,30,118,31,242,31,63,31,124,31,139,31,244,31,185,31,247,31,207,31,126,31,180,31,76,31,23,31,246,31,150,31,158,31,128,31,227,31,56,31,172,31,17,31,205,31,214,31,214,30,214,29,43,31,87,31,87,30,72,31,28,31,119,31,42,31,118,31,203,31,55,31,231,31,79,31,177,31,77,31,218,31,18,31,161,31,236,31,236,30,134,31,49,31,171,31,73,31,73,30,106,31,126,31,16,31,16,30,16,29,45,31,72,31,72,31,65,31,65,30,134,31,17,31,104,31,142,31,124,31,195,31,220,31,46,31,179,31,94,31,94,30,94,29,14,31,110,31,195,31,195,30,40,31,186,31,109,31,101,31,53,31,188,31,146,31,41,31,36,31,249,31,138,31,15,31,10,31,100,31,46,31,254,31,254,30,129,31,81,31,82,31,26,31,105,31,159,31,4,31,4,30,91,31,71,31,45,31,159,31,192,31,136,31,136,30,97,31,154,31,154,30,118,31,77,31,168,31,254,31,81,31,3,31,3,30,1,31,79,31,79,30,39,31,138,31,80,31,43,31,93,31,248,31,248,30,21,31,196,31,196,30,71,31,55,31,55,30,223,31,82,31,238,31,229,31,64,31,79,31,40,31,215,31,215,30,1,31,254,31,33,31,176,31,245,31,65,31,164,31,104,31,104,30,40,31,120,31,65,31,138,31,173,31,173,30,207,31,160,31,65,31,28,31,28,30,76,31,163,31,113,31,179,31,96,31,120,31,27,31,32,31,51,31,23,31,160,31,133,31,133,30,109,31,109,30,241,31,241,30,241,29,241,28,241,27,77,31,120,31,120,30,224,31,57,31,72,31,72,30,72,29,255,31,255,30,226,31,146,31,160,31,160,30,210,31,179,31,58,31,194,31,194,30,92,31,197,31,107,31,113,31,253,31,253,30,92,31,155,31,155,30,25,31,178,31,130,31,49,31,25,31,25,30,25,29,116,31,42,31,1,31,132,31,78,31,78,30,28,31,129,31,189,31,77,31,6,31,6,30,187,31,132,31,32,31,32,30,211,31,108,31,3,31,3,30,146,31,194,31,194,30,20,31,224,31,98,31,216,31,216,30,216,29,216,28,210,31,171,31,154,31,182,31,91,31,91,30,91,29,212,31,181,31,206,31,190,31,213,31,213,30,49,31,225,31,27,31,163,31,74,31,67,31,166,31,31,31,173,31,154,31,238,31,238,30,253,31,253,30,216,31,6,31,177,31,36,31,159,31,107,31,111,31,160,31,157,31,157,30,157,29,157,28,157,27,45,31,52,31,52,30,108,31,108,30,108,29,207,31,207,30,102,31,216,31,169,31,169,30,241,31,95,31,79,31,174,31,174,30,174,29,174,28,167,31,160,31,154,31,105,31,44,31,44,30,35,31,117,31,65,31,31,31,31,30,193,31,97,31,132,31,155,31,128,31,212,31,223,31,3,31,3,31,235,31,133,31,129,31,79,31,79,30,49,31,47,31,58,31,35,31,214,31,204,31,175,31,128,31,164,31,79,31,113,31,57,31,196,31,253,31,197,31,75,31,75,30,176,31,176,30,213,31,218,31,218,30,1,31,8,31,8,30,115,31,115,30,115,29,251,31,251,30,112,31,221,31,183,31,250,31,19,31,130,31,7,31,156,31,156,30,205,31,251,31,223,31,62,31,87,31,36,31,248,31,248,30,15,31,128,31,244,31,213,31,81,31,209,31,9,31,9,30,62,31,245,31,172,31,172,30,17,31,17,30,207,31,119,31,119,30,119,29,12,31,12,30,72,31,121,31,121,30,66,31,66,30,222,31,33,31,226,31,226,31,208,31,57,31,57,30,183,31,251,31,76,31,249,31,71,31,71,30,71,29,69,31,212,31,212,30,122,31,122,30,174,31,174,30,84,31,84,30,96,31,207,31,24,31,51,31,51,30,22,31,22,30,89,31,89,30,61,31,168,31,117,31,216,31,106,31,72,31,110,31,63,31,6,31,35,31,71,31,220,31,48,31,48,30,143,31,106,31,106,30,160,31,245,31,176,31,186,31,105,31,74,31,74,30,246,31,170,31,58,31,230,31,220,31,248,31,14,31,11,31,22,31,132,31,132,30,33,31,164,31,164,30,164,29,162,31,162,30,57,31,20,31,151,31,16,31,227,31,216,31,208,31,103,31,136,31,107,31,237,31,180,31,86,31,185,31,242,31,15,31,142,31,25,31,1,31,1,30,1,29,188,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
