-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_99 is
end project_tb_99;

architecture project_tb_arch_99 of project_tb_99 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 586;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,10,0,0,0,145,0,29,0,0,0,141,0,226,0,0,0,225,0,239,0,90,0,171,0,86,0,159,0,79,0,156,0,190,0,99,0,171,0,0,0,0,0,54,0,148,0,32,0,22,0,228,0,255,0,75,0,0,0,0,0,148,0,74,0,92,0,179,0,53,0,13,0,254,0,102,0,56,0,57,0,240,0,125,0,124,0,0,0,0,0,132,0,10,0,13,0,191,0,214,0,197,0,0,0,241,0,70,0,79,0,151,0,101,0,241,0,25,0,30,0,13,0,0,0,219,0,228,0,255,0,161,0,143,0,79,0,0,0,149,0,15,0,53,0,133,0,92,0,156,0,227,0,185,0,0,0,72,0,215,0,174,0,134,0,118,0,0,0,102,0,0,0,33,0,156,0,41,0,41,0,178,0,214,0,0,0,182,0,242,0,18,0,201,0,222,0,186,0,0,0,172,0,61,0,143,0,0,0,115,0,7,0,67,0,2,0,217,0,91,0,0,0,0,0,183,0,215,0,70,0,243,0,42,0,32,0,52,0,248,0,85,0,27,0,99,0,0,0,201,0,89,0,220,0,0,0,2,0,253,0,180,0,255,0,3,0,0,0,71,0,116,0,242,0,62,0,63,0,0,0,234,0,32,0,128,0,0,0,10,0,145,0,148,0,255,0,159,0,4,0,0,0,0,0,53,0,144,0,176,0,118,0,6,0,60,0,237,0,124,0,231,0,96,0,65,0,252,0,188,0,87,0,233,0,57,0,227,0,232,0,29,0,119,0,190,0,111,0,47,0,0,0,14,0,254,0,0,0,41,0,0,0,253,0,50,0,197,0,211,0,208,0,0,0,227,0,35,0,21,0,252,0,150,0,242,0,0,0,0,0,25,0,221,0,113,0,254,0,224,0,252,0,0,0,39,0,0,0,0,0,59,0,184,0,95,0,166,0,184,0,109,0,3,0,244,0,222,0,89,0,85,0,232,0,159,0,79,0,164,0,0,0,6,0,32,0,10,0,237,0,0,0,119,0,121,0,80,0,84,0,71,0,218,0,21,0,99,0,0,0,149,0,189,0,245,0,171,0,159,0,120,0,251,0,228,0,81,0,78,0,3,0,49,0,246,0,0,0,181,0,114,0,136,0,187,0,141,0,0,0,125,0,227,0,127,0,241,0,0,0,125,0,210,0,233,0,193,0,37,0,158,0,17,0,0,0,117,0,222,0,151,0,202,0,202,0,0,0,59,0,0,0,37,0,248,0,0,0,19,0,153,0,0,0,200,0,187,0,89,0,176,0,174,0,166,0,149,0,23,0,79,0,188,0,82,0,160,0,141,0,1,0,170,0,106,0,65,0,212,0,71,0,98,0,104,0,0,0,106,0,219,0,178,0,216,0,106,0,16,0,39,0,170,0,181,0,85,0,0,0,186,0,251,0,0,0,35,0,12,0,104,0,4,0,0,0,64,0,0,0,169,0,0,0,55,0,73,0,229,0,157,0,41,0,0,0,0,0,0,0,0,0,0,0,29,0,0,0,0,0,56,0,69,0,93,0,222,0,211,0,0,0,0,0,198,0,123,0,199,0,232,0,0,0,165,0,205,0,157,0,120,0,217,0,25,0,175,0,113,0,182,0,75,0,0,0,64,0,241,0,0,0,0,0,0,0,46,0,72,0,96,0,137,0,181,0,0,0,119,0,67,0,0,0,65,0,0,0,235,0,70,0,244,0,84,0,231,0,0,0,0,0,0,0,195,0,240,0,176,0,240,0,117,0,217,0,134,0,131,0,61,0,252,0,85,0,46,0,17,0,47,0,2,0,0,0,138,0,190,0,127,0,203,0,1,0,156,0,29,0,0,0,108,0,0,0,84,0,0,0,0,0,75,0,0,0,68,0,218,0,100,0,204,0,132,0,5,0,240,0,247,0,33,0,212,0,8,0,230,0,132,0,181,0,53,0,60,0,0,0,0,0,51,0,138,0,46,0,0,0,0,0,82,0,0,0,112,0,0,0,87,0,44,0,171,0,213,0,172,0,168,0,0,0,213,0,254,0,68,0,203,0,128,0,151,0,0,0,216,0,0,0,65,0,0,0,57,0,204,0,159,0,0,0,0,0,168,0,141,0,213,0,0,0,0,0,0,0,154,0,52,0,109,0,129,0,7,0,50,0,45,0,231,0,22,0,202,0,85,0,139,0,167,0,0,0,0,0,89,0,121,0,193,0,55,0,78,0,44,0,76,0,0,0,0,0,0,0,119,0,0,0,166,0,0,0,164,0,40,0,110,0,181,0,188,0,255,0,133,0,33,0,5,0,108,0,152,0,242,0,81,0,87,0,221,0,95,0,231,0,159,0,0,0,122,0,228,0,93,0,189,0,10,0,154,0,194,0,0,0,195,0,0,0,0,0,0,0,108,0,75,0,0,0,219,0,0,0,92,0,135,0,19,0,0,0,77,0,138,0,235,0,132,0,176,0,107,0,235,0,0,0,219,0,27,0,205,0,141,0,220,0,238,0,85,0,191,0,121,0,148,0,188,0,0,0,0,0,126,0,0,0,57,0,102,0,122,0,158,0,62,0,6,0,106,0,241,0,97,0,0,0,250,0,145,0,247,0,244,0,4,0,247,0,13,0,13,0,248,0);
signal scenario_full  : scenario_type := (0,0,10,31,10,30,145,31,29,31,29,30,141,31,226,31,226,30,225,31,239,31,90,31,171,31,86,31,159,31,79,31,156,31,190,31,99,31,171,31,171,30,171,29,54,31,148,31,32,31,22,31,228,31,255,31,75,31,75,30,75,29,148,31,74,31,92,31,179,31,53,31,13,31,254,31,102,31,56,31,57,31,240,31,125,31,124,31,124,30,124,29,132,31,10,31,13,31,191,31,214,31,197,31,197,30,241,31,70,31,79,31,151,31,101,31,241,31,25,31,30,31,13,31,13,30,219,31,228,31,255,31,161,31,143,31,79,31,79,30,149,31,15,31,53,31,133,31,92,31,156,31,227,31,185,31,185,30,72,31,215,31,174,31,134,31,118,31,118,30,102,31,102,30,33,31,156,31,41,31,41,31,178,31,214,31,214,30,182,31,242,31,18,31,201,31,222,31,186,31,186,30,172,31,61,31,143,31,143,30,115,31,7,31,67,31,2,31,217,31,91,31,91,30,91,29,183,31,215,31,70,31,243,31,42,31,32,31,52,31,248,31,85,31,27,31,99,31,99,30,201,31,89,31,220,31,220,30,2,31,253,31,180,31,255,31,3,31,3,30,71,31,116,31,242,31,62,31,63,31,63,30,234,31,32,31,128,31,128,30,10,31,145,31,148,31,255,31,159,31,4,31,4,30,4,29,53,31,144,31,176,31,118,31,6,31,60,31,237,31,124,31,231,31,96,31,65,31,252,31,188,31,87,31,233,31,57,31,227,31,232,31,29,31,119,31,190,31,111,31,47,31,47,30,14,31,254,31,254,30,41,31,41,30,253,31,50,31,197,31,211,31,208,31,208,30,227,31,35,31,21,31,252,31,150,31,242,31,242,30,242,29,25,31,221,31,113,31,254,31,224,31,252,31,252,30,39,31,39,30,39,29,59,31,184,31,95,31,166,31,184,31,109,31,3,31,244,31,222,31,89,31,85,31,232,31,159,31,79,31,164,31,164,30,6,31,32,31,10,31,237,31,237,30,119,31,121,31,80,31,84,31,71,31,218,31,21,31,99,31,99,30,149,31,189,31,245,31,171,31,159,31,120,31,251,31,228,31,81,31,78,31,3,31,49,31,246,31,246,30,181,31,114,31,136,31,187,31,141,31,141,30,125,31,227,31,127,31,241,31,241,30,125,31,210,31,233,31,193,31,37,31,158,31,17,31,17,30,117,31,222,31,151,31,202,31,202,31,202,30,59,31,59,30,37,31,248,31,248,30,19,31,153,31,153,30,200,31,187,31,89,31,176,31,174,31,166,31,149,31,23,31,79,31,188,31,82,31,160,31,141,31,1,31,170,31,106,31,65,31,212,31,71,31,98,31,104,31,104,30,106,31,219,31,178,31,216,31,106,31,16,31,39,31,170,31,181,31,85,31,85,30,186,31,251,31,251,30,35,31,12,31,104,31,4,31,4,30,64,31,64,30,169,31,169,30,55,31,73,31,229,31,157,31,41,31,41,30,41,29,41,28,41,27,41,26,29,31,29,30,29,29,56,31,69,31,93,31,222,31,211,31,211,30,211,29,198,31,123,31,199,31,232,31,232,30,165,31,205,31,157,31,120,31,217,31,25,31,175,31,113,31,182,31,75,31,75,30,64,31,241,31,241,30,241,29,241,28,46,31,72,31,96,31,137,31,181,31,181,30,119,31,67,31,67,30,65,31,65,30,235,31,70,31,244,31,84,31,231,31,231,30,231,29,231,28,195,31,240,31,176,31,240,31,117,31,217,31,134,31,131,31,61,31,252,31,85,31,46,31,17,31,47,31,2,31,2,30,138,31,190,31,127,31,203,31,1,31,156,31,29,31,29,30,108,31,108,30,84,31,84,30,84,29,75,31,75,30,68,31,218,31,100,31,204,31,132,31,5,31,240,31,247,31,33,31,212,31,8,31,230,31,132,31,181,31,53,31,60,31,60,30,60,29,51,31,138,31,46,31,46,30,46,29,82,31,82,30,112,31,112,30,87,31,44,31,171,31,213,31,172,31,168,31,168,30,213,31,254,31,68,31,203,31,128,31,151,31,151,30,216,31,216,30,65,31,65,30,57,31,204,31,159,31,159,30,159,29,168,31,141,31,213,31,213,30,213,29,213,28,154,31,52,31,109,31,129,31,7,31,50,31,45,31,231,31,22,31,202,31,85,31,139,31,167,31,167,30,167,29,89,31,121,31,193,31,55,31,78,31,44,31,76,31,76,30,76,29,76,28,119,31,119,30,166,31,166,30,164,31,40,31,110,31,181,31,188,31,255,31,133,31,33,31,5,31,108,31,152,31,242,31,81,31,87,31,221,31,95,31,231,31,159,31,159,30,122,31,228,31,93,31,189,31,10,31,154,31,194,31,194,30,195,31,195,30,195,29,195,28,108,31,75,31,75,30,219,31,219,30,92,31,135,31,19,31,19,30,77,31,138,31,235,31,132,31,176,31,107,31,235,31,235,30,219,31,27,31,205,31,141,31,220,31,238,31,85,31,191,31,121,31,148,31,188,31,188,30,188,29,126,31,126,30,57,31,102,31,122,31,158,31,62,31,6,31,106,31,241,31,97,31,97,30,250,31,145,31,247,31,244,31,4,31,247,31,13,31,13,31,248,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
