-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 326;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (174,0,151,0,205,0,18,0,59,0,164,0,0,0,0,0,219,0,0,0,0,0,0,0,61,0,176,0,73,0,0,0,184,0,0,0,0,0,130,0,181,0,0,0,175,0,0,0,135,0,245,0,78,0,251,0,161,0,0,0,224,0,238,0,0,0,0,0,2,0,78,0,166,0,235,0,233,0,211,0,0,0,107,0,231,0,83,0,45,0,0,0,161,0,0,0,216,0,54,0,25,0,196,0,142,0,0,0,236,0,144,0,203,0,190,0,0,0,235,0,0,0,0,0,207,0,176,0,241,0,203,0,228,0,88,0,92,0,250,0,92,0,12,0,170,0,20,0,99,0,114,0,132,0,22,0,23,0,123,0,171,0,115,0,150,0,0,0,24,0,221,0,0,0,10,0,86,0,172,0,49,0,39,0,50,0,0,0,36,0,200,0,192,0,237,0,59,0,137,0,0,0,196,0,246,0,168,0,177,0,11,0,92,0,150,0,0,0,82,0,79,0,150,0,222,0,155,0,246,0,0,0,0,0,140,0,0,0,0,0,183,0,118,0,115,0,222,0,12,0,20,0,0,0,8,0,37,0,126,0,0,0,78,0,57,0,0,0,125,0,66,0,226,0,11,0,143,0,19,0,2,0,188,0,0,0,244,0,24,0,203,0,0,0,176,0,117,0,37,0,231,0,173,0,44,0,58,0,4,0,250,0,0,0,30,0,165,0,81,0,201,0,0,0,241,0,91,0,93,0,35,0,42,0,132,0,124,0,59,0,88,0,75,0,0,0,197,0,0,0,85,0,142,0,48,0,208,0,0,0,84,0,199,0,61,0,27,0,0,0,110,0,0,0,0,0,237,0,97,0,236,0,149,0,0,0,1,0,28,0,3,0,40,0,143,0,11,0,163,0,58,0,86,0,81,0,161,0,110,0,215,0,0,0,217,0,0,0,0,0,161,0,0,0,113,0,146,0,121,0,37,0,92,0,203,0,142,0,221,0,155,0,0,0,0,0,188,0,47,0,0,0,0,0,122,0,110,0,0,0,207,0,204,0,117,0,109,0,0,0,136,0,68,0,97,0,1,0,195,0,0,0,214,0,115,0,91,0,0,0,247,0,67,0,60,0,0,0,201,0,0,0,70,0,10,0,229,0,0,0,123,0,245,0,129,0,0,0,117,0,0,0,90,0,95,0,0,0,136,0,249,0,0,0,82,0,141,0,202,0,96,0,237,0,0,0,95,0,0,0,173,0,232,0,53,0,82,0,189,0,246,0,24,0,0,0,0,0,182,0,0,0,3,0,0,0,132,0,76,0,17,0,0,0,0,0,171,0,111,0,227,0,213,0,103,0,161,0,0,0,21,0,67,0,64,0,246,0,0,0,100,0,0,0,144,0,16,0,171,0,64,0,223,0,112,0,167,0,0,0,13,0,0,0,240,0,55,0,116,0,216,0,116,0,68,0,240,0,0,0,202,0);
signal scenario_full  : scenario_type := (174,31,151,31,205,31,18,31,59,31,164,31,164,30,164,29,219,31,219,30,219,29,219,28,61,31,176,31,73,31,73,30,184,31,184,30,184,29,130,31,181,31,181,30,175,31,175,30,135,31,245,31,78,31,251,31,161,31,161,30,224,31,238,31,238,30,238,29,2,31,78,31,166,31,235,31,233,31,211,31,211,30,107,31,231,31,83,31,45,31,45,30,161,31,161,30,216,31,54,31,25,31,196,31,142,31,142,30,236,31,144,31,203,31,190,31,190,30,235,31,235,30,235,29,207,31,176,31,241,31,203,31,228,31,88,31,92,31,250,31,92,31,12,31,170,31,20,31,99,31,114,31,132,31,22,31,23,31,123,31,171,31,115,31,150,31,150,30,24,31,221,31,221,30,10,31,86,31,172,31,49,31,39,31,50,31,50,30,36,31,200,31,192,31,237,31,59,31,137,31,137,30,196,31,246,31,168,31,177,31,11,31,92,31,150,31,150,30,82,31,79,31,150,31,222,31,155,31,246,31,246,30,246,29,140,31,140,30,140,29,183,31,118,31,115,31,222,31,12,31,20,31,20,30,8,31,37,31,126,31,126,30,78,31,57,31,57,30,125,31,66,31,226,31,11,31,143,31,19,31,2,31,188,31,188,30,244,31,24,31,203,31,203,30,176,31,117,31,37,31,231,31,173,31,44,31,58,31,4,31,250,31,250,30,30,31,165,31,81,31,201,31,201,30,241,31,91,31,93,31,35,31,42,31,132,31,124,31,59,31,88,31,75,31,75,30,197,31,197,30,85,31,142,31,48,31,208,31,208,30,84,31,199,31,61,31,27,31,27,30,110,31,110,30,110,29,237,31,97,31,236,31,149,31,149,30,1,31,28,31,3,31,40,31,143,31,11,31,163,31,58,31,86,31,81,31,161,31,110,31,215,31,215,30,217,31,217,30,217,29,161,31,161,30,113,31,146,31,121,31,37,31,92,31,203,31,142,31,221,31,155,31,155,30,155,29,188,31,47,31,47,30,47,29,122,31,110,31,110,30,207,31,204,31,117,31,109,31,109,30,136,31,68,31,97,31,1,31,195,31,195,30,214,31,115,31,91,31,91,30,247,31,67,31,60,31,60,30,201,31,201,30,70,31,10,31,229,31,229,30,123,31,245,31,129,31,129,30,117,31,117,30,90,31,95,31,95,30,136,31,249,31,249,30,82,31,141,31,202,31,96,31,237,31,237,30,95,31,95,30,173,31,232,31,53,31,82,31,189,31,246,31,24,31,24,30,24,29,182,31,182,30,3,31,3,30,132,31,76,31,17,31,17,30,17,29,171,31,111,31,227,31,213,31,103,31,161,31,161,30,21,31,67,31,64,31,246,31,246,30,100,31,100,30,144,31,16,31,171,31,64,31,223,31,112,31,167,31,167,30,13,31,13,30,240,31,55,31,116,31,216,31,116,31,68,31,240,31,240,30,202,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
