-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_187 is
end project_tb_187;

architecture project_tb_arch_187 of project_tb_187 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 372;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (241,0,252,0,131,0,170,0,86,0,0,0,22,0,217,0,18,0,94,0,209,0,2,0,0,0,0,0,123,0,0,0,117,0,95,0,0,0,5,0,217,0,82,0,87,0,28,0,160,0,0,0,184,0,0,0,67,0,0,0,112,0,89,0,205,0,87,0,13,0,0,0,189,0,97,0,175,0,219,0,128,0,72,0,159,0,95,0,56,0,154,0,214,0,128,0,0,0,208,0,222,0,0,0,76,0,0,0,0,0,57,0,249,0,91,0,0,0,186,0,0,0,79,0,208,0,182,0,0,0,75,0,216,0,0,0,141,0,165,0,111,0,27,0,0,0,52,0,0,0,72,0,240,0,15,0,19,0,44,0,45,0,165,0,155,0,158,0,0,0,175,0,118,0,255,0,75,0,72,0,218,0,175,0,38,0,0,0,61,0,91,0,44,0,190,0,145,0,0,0,117,0,56,0,48,0,248,0,21,0,98,0,0,0,0,0,160,0,1,0,224,0,31,0,28,0,0,0,180,0,115,0,0,0,0,0,52,0,145,0,19,0,53,0,51,0,40,0,136,0,241,0,102,0,0,0,0,0,154,0,94,0,151,0,41,0,67,0,111,0,117,0,163,0,241,0,0,0,128,0,76,0,88,0,182,0,228,0,0,0,128,0,169,0,97,0,46,0,85,0,16,0,231,0,177,0,163,0,97,0,0,0,236,0,0,0,34,0,57,0,196,0,154,0,140,0,0,0,237,0,162,0,221,0,0,0,205,0,0,0,184,0,40,0,114,0,231,0,67,0,0,0,0,0,121,0,18,0,53,0,194,0,163,0,7,0,0,0,153,0,241,0,56,0,135,0,247,0,61,0,41,0,106,0,193,0,0,0,153,0,74,0,201,0,43,0,131,0,186,0,210,0,246,0,17,0,79,0,180,0,0,0,198,0,0,0,27,0,217,0,0,0,2,0,132,0,210,0,0,0,0,0,0,0,154,0,25,0,64,0,151,0,0,0,250,0,186,0,241,0,176,0,0,0,101,0,65,0,147,0,138,0,156,0,202,0,185,0,247,0,158,0,177,0,0,0,104,0,16,0,218,0,0,0,19,0,0,0,12,0,245,0,142,0,0,0,164,0,227,0,124,0,224,0,0,0,132,0,154,0,49,0,190,0,219,0,117,0,38,0,0,0,162,0,151,0,255,0,76,0,139,0,114,0,0,0,165,0,87,0,72,0,188,0,19,0,0,0,170,0,208,0,96,0,6,0,0,0,36,0,170,0,157,0,0,0,44,0,107,0,188,0,138,0,0,0,32,0,185,0,143,0,0,0,0,0,147,0,50,0,188,0,0,0,123,0,14,0,0,0,105,0,0,0,155,0,0,0,0,0,207,0,134,0,0,0,243,0,150,0,41,0,0,0,0,0,100,0,32,0,0,0,214,0,157,0,8,0,2,0,39,0,46,0,0,0,120,0,219,0,243,0,0,0,131,0,76,0,204,0,101,0,0,0,148,0,232,0,49,0,0,0,214,0,0,0,0,0,70,0,114,0,69,0,29,0,148,0,158,0,27,0,0,0,18,0,0,0,138,0,155,0,0,0,190,0,15,0,152,0,183,0,0,0,0,0,32,0,67,0,219,0,79,0,150,0,220,0,172,0,0,0,101,0,202,0,0,0,173,0,0,0,0,0);
signal scenario_full  : scenario_type := (241,31,252,31,131,31,170,31,86,31,86,30,22,31,217,31,18,31,94,31,209,31,2,31,2,30,2,29,123,31,123,30,117,31,95,31,95,30,5,31,217,31,82,31,87,31,28,31,160,31,160,30,184,31,184,30,67,31,67,30,112,31,89,31,205,31,87,31,13,31,13,30,189,31,97,31,175,31,219,31,128,31,72,31,159,31,95,31,56,31,154,31,214,31,128,31,128,30,208,31,222,31,222,30,76,31,76,30,76,29,57,31,249,31,91,31,91,30,186,31,186,30,79,31,208,31,182,31,182,30,75,31,216,31,216,30,141,31,165,31,111,31,27,31,27,30,52,31,52,30,72,31,240,31,15,31,19,31,44,31,45,31,165,31,155,31,158,31,158,30,175,31,118,31,255,31,75,31,72,31,218,31,175,31,38,31,38,30,61,31,91,31,44,31,190,31,145,31,145,30,117,31,56,31,48,31,248,31,21,31,98,31,98,30,98,29,160,31,1,31,224,31,31,31,28,31,28,30,180,31,115,31,115,30,115,29,52,31,145,31,19,31,53,31,51,31,40,31,136,31,241,31,102,31,102,30,102,29,154,31,94,31,151,31,41,31,67,31,111,31,117,31,163,31,241,31,241,30,128,31,76,31,88,31,182,31,228,31,228,30,128,31,169,31,97,31,46,31,85,31,16,31,231,31,177,31,163,31,97,31,97,30,236,31,236,30,34,31,57,31,196,31,154,31,140,31,140,30,237,31,162,31,221,31,221,30,205,31,205,30,184,31,40,31,114,31,231,31,67,31,67,30,67,29,121,31,18,31,53,31,194,31,163,31,7,31,7,30,153,31,241,31,56,31,135,31,247,31,61,31,41,31,106,31,193,31,193,30,153,31,74,31,201,31,43,31,131,31,186,31,210,31,246,31,17,31,79,31,180,31,180,30,198,31,198,30,27,31,217,31,217,30,2,31,132,31,210,31,210,30,210,29,210,28,154,31,25,31,64,31,151,31,151,30,250,31,186,31,241,31,176,31,176,30,101,31,65,31,147,31,138,31,156,31,202,31,185,31,247,31,158,31,177,31,177,30,104,31,16,31,218,31,218,30,19,31,19,30,12,31,245,31,142,31,142,30,164,31,227,31,124,31,224,31,224,30,132,31,154,31,49,31,190,31,219,31,117,31,38,31,38,30,162,31,151,31,255,31,76,31,139,31,114,31,114,30,165,31,87,31,72,31,188,31,19,31,19,30,170,31,208,31,96,31,6,31,6,30,36,31,170,31,157,31,157,30,44,31,107,31,188,31,138,31,138,30,32,31,185,31,143,31,143,30,143,29,147,31,50,31,188,31,188,30,123,31,14,31,14,30,105,31,105,30,155,31,155,30,155,29,207,31,134,31,134,30,243,31,150,31,41,31,41,30,41,29,100,31,32,31,32,30,214,31,157,31,8,31,2,31,39,31,46,31,46,30,120,31,219,31,243,31,243,30,131,31,76,31,204,31,101,31,101,30,148,31,232,31,49,31,49,30,214,31,214,30,214,29,70,31,114,31,69,31,29,31,148,31,158,31,27,31,27,30,18,31,18,30,138,31,155,31,155,30,190,31,15,31,152,31,183,31,183,30,183,29,32,31,67,31,219,31,79,31,150,31,220,31,172,31,172,30,101,31,202,31,202,30,173,31,173,30,173,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
