-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_705 is
end project_tb_705;

architecture project_tb_arch_705 of project_tb_705 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 842;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,244,0,99,0,154,0,219,0,198,0,142,0,239,0,166,0,0,0,26,0,156,0,84,0,239,0,92,0,0,0,0,0,6,0,176,0,234,0,0,0,7,0,0,0,203,0,244,0,180,0,88,0,0,0,21,0,0,0,0,0,56,0,67,0,156,0,0,0,0,0,0,0,222,0,0,0,181,0,154,0,115,0,0,0,160,0,155,0,7,0,156,0,199,0,72,0,168,0,182,0,72,0,192,0,103,0,240,0,96,0,95,0,162,0,199,0,73,0,225,0,216,0,110,0,61,0,99,0,53,0,0,0,78,0,165,0,149,0,120,0,165,0,0,0,0,0,253,0,254,0,86,0,238,0,95,0,20,0,231,0,0,0,0,0,208,0,0,0,239,0,171,0,177,0,81,0,71,0,137,0,163,0,0,0,6,0,0,0,162,0,171,0,204,0,125,0,0,0,140,0,0,0,77,0,41,0,174,0,152,0,116,0,193,0,226,0,0,0,243,0,233,0,159,0,188,0,210,0,0,0,0,0,3,0,218,0,242,0,14,0,236,0,91,0,103,0,70,0,251,0,242,0,218,0,19,0,102,0,0,0,253,0,11,0,148,0,175,0,50,0,44,0,112,0,229,0,0,0,0,0,0,0,61,0,211,0,201,0,22,0,8,0,0,0,56,0,30,0,130,0,151,0,179,0,14,0,109,0,0,0,60,0,12,0,104,0,78,0,64,0,70,0,0,0,125,0,233,0,105,0,89,0,156,0,84,0,32,0,99,0,130,0,0,0,185,0,200,0,161,0,211,0,203,0,57,0,84,0,120,0,0,0,23,0,241,0,126,0,74,0,198,0,0,0,164,0,46,0,235,0,187,0,120,0,170,0,214,0,248,0,226,0,177,0,223,0,164,0,20,0,12,0,12,0,155,0,0,0,181,0,10,0,115,0,125,0,180,0,0,0,57,0,159,0,0,0,112,0,194,0,150,0,157,0,230,0,143,0,68,0,203,0,0,0,182,0,36,0,0,0,0,0,201,0,136,0,156,0,0,0,122,0,0,0,155,0,225,0,0,0,0,0,58,0,0,0,198,0,79,0,0,0,0,0,189,0,152,0,0,0,142,0,149,0,232,0,225,0,228,0,209,0,45,0,0,0,12,0,0,0,27,0,56,0,0,0,52,0,29,0,142,0,219,0,167,0,194,0,47,0,205,0,204,0,177,0,19,0,0,0,60,0,161,0,143,0,51,0,112,0,165,0,109,0,239,0,91,0,107,0,81,0,158,0,224,0,0,0,163,0,61,0,159,0,127,0,133,0,6,0,173,0,119,0,237,0,51,0,67,0,71,0,20,0,226,0,60,0,218,0,0,0,81,0,153,0,61,0,79,0,104,0,158,0,43,0,38,0,146,0,173,0,6,0,0,0,111,0,96,0,224,0,0,0,142,0,69,0,0,0,25,0,47,0,213,0,251,0,53,0,0,0,46,0,132,0,69,0,168,0,216,0,0,0,0,0,160,0,140,0,248,0,240,0,86,0,27,0,61,0,176,0,206,0,0,0,0,0,0,0,0,0,248,0,76,0,26,0,105,0,122,0,156,0,205,0,141,0,56,0,217,0,235,0,0,0,0,0,0,0,199,0,175,0,248,0,68,0,98,0,252,0,0,0,34,0,0,0,0,0,0,0,58,0,0,0,0,0,81,0,94,0,162,0,1,0,0,0,20,0,99,0,17,0,252,0,242,0,97,0,22,0,193,0,61,0,135,0,0,0,121,0,69,0,247,0,188,0,226,0,143,0,93,0,47,0,34,0,68,0,130,0,0,0,0,0,40,0,177,0,158,0,139,0,21,0,122,0,163,0,178,0,66,0,46,0,34,0,0,0,12,0,79,0,3,0,230,0,157,0,17,0,143,0,219,0,250,0,129,0,81,0,31,0,209,0,0,0,143,0,28,0,155,0,0,0,62,0,0,0,103,0,35,0,0,0,0,0,79,0,161,0,61,0,172,0,54,0,0,0,110,0,167,0,193,0,19,0,209,0,111,0,233,0,0,0,93,0,59,0,0,0,124,0,176,0,0,0,0,0,30,0,85,0,141,0,103,0,162,0,232,0,219,0,154,0,158,0,252,0,88,0,15,0,102,0,133,0,57,0,154,0,22,0,37,0,255,0,0,0,250,0,170,0,0,0,254,0,0,0,124,0,0,0,0,0,14,0,172,0,43,0,109,0,98,0,241,0,111,0,159,0,6,0,0,0,0,0,174,0,78,0,34,0,17,0,0,0,33,0,0,0,192,0,0,0,126,0,4,0,207,0,196,0,0,0,177,0,8,0,0,0,0,0,130,0,215,0,60,0,233,0,0,0,174,0,17,0,170,0,172,0,0,0,178,0,0,0,18,0,111,0,82,0,197,0,134,0,0,0,0,0,188,0,0,0,83,0,0,0,0,0,92,0,22,0,64,0,50,0,16,0,215,0,99,0,59,0,134,0,231,0,163,0,0,0,250,0,0,0,193,0,230,0,244,0,0,0,61,0,70,0,0,0,64,0,154,0,238,0,182,0,0,0,160,0,219,0,223,0,200,0,213,0,21,0,244,0,248,0,0,0,72,0,240,0,86,0,203,0,95,0,117,0,0,0,185,0,59,0,240,0,35,0,0,0,111,0,96,0,44,0,192,0,209,0,0,0,0,0,0,0,27,0,63,0,121,0,187,0,217,0,234,0,102,0,81,0,0,0,52,0,15,0,246,0,126,0,189,0,93,0,68,0,0,0,0,0,81,0,162,0,0,0,0,0,100,0,185,0,0,0,135,0,185,0,198,0,0,0,133,0,0,0,18,0,62,0,0,0,13,0,0,0,27,0,4,0,191,0,0,0,0,0,119,0,219,0,36,0,0,0,167,0,0,0,19,0,251,0,28,0,35,0,241,0,57,0,0,0,182,0,174,0,0,0,190,0,72,0,52,0,0,0,247,0,180,0,160,0,201,0,24,0,0,0,0,0,113,0,134,0,0,0,0,0,139,0,31,0,0,0,230,0,114,0,204,0,8,0,29,0,0,0,0,0,0,0,59,0,243,0,111,0,218,0,136,0,85,0,139,0,82,0,0,0,67,0,119,0,20,0,89,0,150,0,194,0,61,0,0,0,0,0,248,0,173,0,0,0,118,0,191,0,189,0,0,0,143,0,109,0,137,0,39,0,197,0,131,0,2,0,39,0,0,0,0,0,24,0,0,0,63,0,179,0,108,0,116,0,217,0,175,0,231,0,139,0,249,0,11,0,0,0,20,0,7,0,18,0,41,0,235,0,70,0,190,0,85,0,200,0,101,0,30,0,193,0,189,0,53,0,0,0,47,0,199,0,0,0,0,0,0,0,186,0,225,0,109,0,174,0,56,0,0,0,68,0,115,0,242,0,107,0,137,0,12,0,161,0,136,0,10,0,171,0,62,0,171,0,75,0,157,0,169,0,119,0,140,0,176,0,57,0,243,0,21,0,109,0,38,0,0,0,135,0,4,0,9,0,89,0,188,0,0,0,0,0,203,0,149,0,209,0,234,0,208,0,38,0,0,0,125,0,185,0,108,0,55,0,236,0,118,0,104,0,0,0,205,0,95,0,70,0,223,0,121,0,119,0,190,0,253,0,218,0,27,0,113,0,0,0,132,0,0,0,215,0,209,0,91,0,6,0,10,0,17,0,192,0,240,0,231,0,0,0,0,0,0,0,45,0,230,0,0,0,161,0,68,0,85,0,39,0,185,0,0,0,6,0,97,0,142,0,0,0,13,0,169,0,49,0);
signal scenario_full  : scenario_type := (214,31,244,31,99,31,154,31,219,31,198,31,142,31,239,31,166,31,166,30,26,31,156,31,84,31,239,31,92,31,92,30,92,29,6,31,176,31,234,31,234,30,7,31,7,30,203,31,244,31,180,31,88,31,88,30,21,31,21,30,21,29,56,31,67,31,156,31,156,30,156,29,156,28,222,31,222,30,181,31,154,31,115,31,115,30,160,31,155,31,7,31,156,31,199,31,72,31,168,31,182,31,72,31,192,31,103,31,240,31,96,31,95,31,162,31,199,31,73,31,225,31,216,31,110,31,61,31,99,31,53,31,53,30,78,31,165,31,149,31,120,31,165,31,165,30,165,29,253,31,254,31,86,31,238,31,95,31,20,31,231,31,231,30,231,29,208,31,208,30,239,31,171,31,177,31,81,31,71,31,137,31,163,31,163,30,6,31,6,30,162,31,171,31,204,31,125,31,125,30,140,31,140,30,77,31,41,31,174,31,152,31,116,31,193,31,226,31,226,30,243,31,233,31,159,31,188,31,210,31,210,30,210,29,3,31,218,31,242,31,14,31,236,31,91,31,103,31,70,31,251,31,242,31,218,31,19,31,102,31,102,30,253,31,11,31,148,31,175,31,50,31,44,31,112,31,229,31,229,30,229,29,229,28,61,31,211,31,201,31,22,31,8,31,8,30,56,31,30,31,130,31,151,31,179,31,14,31,109,31,109,30,60,31,12,31,104,31,78,31,64,31,70,31,70,30,125,31,233,31,105,31,89,31,156,31,84,31,32,31,99,31,130,31,130,30,185,31,200,31,161,31,211,31,203,31,57,31,84,31,120,31,120,30,23,31,241,31,126,31,74,31,198,31,198,30,164,31,46,31,235,31,187,31,120,31,170,31,214,31,248,31,226,31,177,31,223,31,164,31,20,31,12,31,12,31,155,31,155,30,181,31,10,31,115,31,125,31,180,31,180,30,57,31,159,31,159,30,112,31,194,31,150,31,157,31,230,31,143,31,68,31,203,31,203,30,182,31,36,31,36,30,36,29,201,31,136,31,156,31,156,30,122,31,122,30,155,31,225,31,225,30,225,29,58,31,58,30,198,31,79,31,79,30,79,29,189,31,152,31,152,30,142,31,149,31,232,31,225,31,228,31,209,31,45,31,45,30,12,31,12,30,27,31,56,31,56,30,52,31,29,31,142,31,219,31,167,31,194,31,47,31,205,31,204,31,177,31,19,31,19,30,60,31,161,31,143,31,51,31,112,31,165,31,109,31,239,31,91,31,107,31,81,31,158,31,224,31,224,30,163,31,61,31,159,31,127,31,133,31,6,31,173,31,119,31,237,31,51,31,67,31,71,31,20,31,226,31,60,31,218,31,218,30,81,31,153,31,61,31,79,31,104,31,158,31,43,31,38,31,146,31,173,31,6,31,6,30,111,31,96,31,224,31,224,30,142,31,69,31,69,30,25,31,47,31,213,31,251,31,53,31,53,30,46,31,132,31,69,31,168,31,216,31,216,30,216,29,160,31,140,31,248,31,240,31,86,31,27,31,61,31,176,31,206,31,206,30,206,29,206,28,206,27,248,31,76,31,26,31,105,31,122,31,156,31,205,31,141,31,56,31,217,31,235,31,235,30,235,29,235,28,199,31,175,31,248,31,68,31,98,31,252,31,252,30,34,31,34,30,34,29,34,28,58,31,58,30,58,29,81,31,94,31,162,31,1,31,1,30,20,31,99,31,17,31,252,31,242,31,97,31,22,31,193,31,61,31,135,31,135,30,121,31,69,31,247,31,188,31,226,31,143,31,93,31,47,31,34,31,68,31,130,31,130,30,130,29,40,31,177,31,158,31,139,31,21,31,122,31,163,31,178,31,66,31,46,31,34,31,34,30,12,31,79,31,3,31,230,31,157,31,17,31,143,31,219,31,250,31,129,31,81,31,31,31,209,31,209,30,143,31,28,31,155,31,155,30,62,31,62,30,103,31,35,31,35,30,35,29,79,31,161,31,61,31,172,31,54,31,54,30,110,31,167,31,193,31,19,31,209,31,111,31,233,31,233,30,93,31,59,31,59,30,124,31,176,31,176,30,176,29,30,31,85,31,141,31,103,31,162,31,232,31,219,31,154,31,158,31,252,31,88,31,15,31,102,31,133,31,57,31,154,31,22,31,37,31,255,31,255,30,250,31,170,31,170,30,254,31,254,30,124,31,124,30,124,29,14,31,172,31,43,31,109,31,98,31,241,31,111,31,159,31,6,31,6,30,6,29,174,31,78,31,34,31,17,31,17,30,33,31,33,30,192,31,192,30,126,31,4,31,207,31,196,31,196,30,177,31,8,31,8,30,8,29,130,31,215,31,60,31,233,31,233,30,174,31,17,31,170,31,172,31,172,30,178,31,178,30,18,31,111,31,82,31,197,31,134,31,134,30,134,29,188,31,188,30,83,31,83,30,83,29,92,31,22,31,64,31,50,31,16,31,215,31,99,31,59,31,134,31,231,31,163,31,163,30,250,31,250,30,193,31,230,31,244,31,244,30,61,31,70,31,70,30,64,31,154,31,238,31,182,31,182,30,160,31,219,31,223,31,200,31,213,31,21,31,244,31,248,31,248,30,72,31,240,31,86,31,203,31,95,31,117,31,117,30,185,31,59,31,240,31,35,31,35,30,111,31,96,31,44,31,192,31,209,31,209,30,209,29,209,28,27,31,63,31,121,31,187,31,217,31,234,31,102,31,81,31,81,30,52,31,15,31,246,31,126,31,189,31,93,31,68,31,68,30,68,29,81,31,162,31,162,30,162,29,100,31,185,31,185,30,135,31,185,31,198,31,198,30,133,31,133,30,18,31,62,31,62,30,13,31,13,30,27,31,4,31,191,31,191,30,191,29,119,31,219,31,36,31,36,30,167,31,167,30,19,31,251,31,28,31,35,31,241,31,57,31,57,30,182,31,174,31,174,30,190,31,72,31,52,31,52,30,247,31,180,31,160,31,201,31,24,31,24,30,24,29,113,31,134,31,134,30,134,29,139,31,31,31,31,30,230,31,114,31,204,31,8,31,29,31,29,30,29,29,29,28,59,31,243,31,111,31,218,31,136,31,85,31,139,31,82,31,82,30,67,31,119,31,20,31,89,31,150,31,194,31,61,31,61,30,61,29,248,31,173,31,173,30,118,31,191,31,189,31,189,30,143,31,109,31,137,31,39,31,197,31,131,31,2,31,39,31,39,30,39,29,24,31,24,30,63,31,179,31,108,31,116,31,217,31,175,31,231,31,139,31,249,31,11,31,11,30,20,31,7,31,18,31,41,31,235,31,70,31,190,31,85,31,200,31,101,31,30,31,193,31,189,31,53,31,53,30,47,31,199,31,199,30,199,29,199,28,186,31,225,31,109,31,174,31,56,31,56,30,68,31,115,31,242,31,107,31,137,31,12,31,161,31,136,31,10,31,171,31,62,31,171,31,75,31,157,31,169,31,119,31,140,31,176,31,57,31,243,31,21,31,109,31,38,31,38,30,135,31,4,31,9,31,89,31,188,31,188,30,188,29,203,31,149,31,209,31,234,31,208,31,38,31,38,30,125,31,185,31,108,31,55,31,236,31,118,31,104,31,104,30,205,31,95,31,70,31,223,31,121,31,119,31,190,31,253,31,218,31,27,31,113,31,113,30,132,31,132,30,215,31,209,31,91,31,6,31,10,31,17,31,192,31,240,31,231,31,231,30,231,29,231,28,45,31,230,31,230,30,161,31,68,31,85,31,39,31,185,31,185,30,6,31,97,31,142,31,142,30,13,31,169,31,49,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
