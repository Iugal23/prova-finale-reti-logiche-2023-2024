-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_680 is
end project_tb_680;

architecture project_tb_arch_680 of project_tb_680 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 867;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (96,0,0,0,216,0,196,0,175,0,244,0,108,0,111,0,124,0,0,0,12,0,83,0,222,0,23,0,241,0,202,0,159,0,136,0,162,0,0,0,140,0,244,0,4,0,117,0,101,0,203,0,0,0,141,0,199,0,194,0,0,0,236,0,226,0,1,0,83,0,0,0,101,0,0,0,224,0,0,0,45,0,164,0,0,0,101,0,140,0,174,0,189,0,0,0,202,0,198,0,98,0,159,0,51,0,0,0,26,0,235,0,0,0,230,0,136,0,0,0,0,0,231,0,181,0,194,0,95,0,31,0,109,0,208,0,95,0,178,0,138,0,132,0,213,0,0,0,109,0,0,0,0,0,19,0,158,0,193,0,0,0,203,0,173,0,213,0,82,0,113,0,59,0,0,0,0,0,36,0,249,0,0,0,40,0,100,0,0,0,0,0,212,0,105,0,125,0,207,0,222,0,88,0,0,0,122,0,177,0,76,0,0,0,0,0,0,0,97,0,117,0,163,0,0,0,102,0,0,0,156,0,45,0,6,0,27,0,252,0,250,0,138,0,0,0,55,0,219,0,127,0,37,0,214,0,182,0,0,0,0,0,200,0,202,0,0,0,5,0,3,0,246,0,57,0,202,0,86,0,0,0,0,0,0,0,231,0,0,0,42,0,244,0,106,0,63,0,0,0,186,0,210,0,13,0,96,0,0,0,231,0,211,0,0,0,192,0,155,0,150,0,138,0,112,0,130,0,97,0,68,0,96,0,240,0,44,0,190,0,227,0,254,0,168,0,171,0,224,0,0,0,13,0,13,0,78,0,54,0,175,0,23,0,0,0,17,0,183,0,209,0,53,0,167,0,42,0,105,0,133,0,242,0,254,0,53,0,219,0,2,0,182,0,128,0,68,0,105,0,72,0,170,0,164,0,136,0,244,0,0,0,144,0,248,0,2,0,72,0,0,0,35,0,0,0,0,0,174,0,193,0,153,0,180,0,208,0,243,0,176,0,0,0,201,0,0,0,240,0,0,0,6,0,99,0,206,0,227,0,193,0,124,0,0,0,43,0,0,0,75,0,0,0,0,0,25,0,236,0,22,0,36,0,222,0,115,0,0,0,58,0,158,0,43,0,0,0,74,0,0,0,50,0,38,0,0,0,105,0,44,0,168,0,165,0,175,0,181,0,245,0,160,0,103,0,6,0,170,0,0,0,219,0,0,0,138,0,219,0,115,0,28,0,231,0,190,0,99,0,144,0,137,0,29,0,119,0,180,0,55,0,0,0,3,0,249,0,62,0,71,0,0,0,46,0,121,0,233,0,166,0,73,0,124,0,52,0,107,0,0,0,86,0,0,0,152,0,234,0,58,0,37,0,156,0,48,0,141,0,84,0,29,0,5,0,249,0,98,0,195,0,121,0,0,0,243,0,0,0,153,0,0,0,69,0,222,0,62,0,169,0,248,0,89,0,0,0,241,0,204,0,119,0,171,0,248,0,41,0,55,0,63,0,128,0,82,0,62,0,109,0,100,0,168,0,82,0,180,0,66,0,205,0,60,0,122,0,158,0,146,0,36,0,176,0,203,0,222,0,104,0,226,0,210,0,48,0,0,0,0,0,233,0,19,0,71,0,70,0,244,0,236,0,1,0,137,0,159,0,165,0,235,0,156,0,0,0,0,0,103,0,34,0,182,0,24,0,0,0,0,0,20,0,39,0,165,0,99,0,122,0,158,0,0,0,162,0,89,0,155,0,207,0,126,0,185,0,39,0,0,0,0,0,94,0,7,0,38,0,0,0,103,0,209,0,196,0,0,0,54,0,154,0,119,0,196,0,59,0,0,0,184,0,19,0,21,0,13,0,189,0,34,0,33,0,93,0,88,0,0,0,0,0,128,0,5,0,0,0,0,0,243,0,37,0,229,0,229,0,161,0,33,0,0,0,37,0,235,0,197,0,28,0,0,0,179,0,113,0,138,0,0,0,98,0,197,0,192,0,10,0,148,0,35,0,153,0,101,0,0,0,6,0,249,0,29,0,90,0,27,0,58,0,211,0,0,0,199,0,0,0,44,0,121,0,154,0,54,0,216,0,96,0,214,0,154,0,75,0,74,0,150,0,106,0,65,0,43,0,145,0,0,0,0,0,194,0,205,0,152,0,100,0,214,0,244,0,108,0,0,0,0,0,49,0,178,0,117,0,34,0,16,0,127,0,191,0,46,0,243,0,194,0,240,0,196,0,179,0,148,0,42,0,180,0,211,0,0,0,0,0,171,0,238,0,188,0,110,0,72,0,0,0,159,0,223,0,104,0,111,0,255,0,173,0,241,0,117,0,128,0,0,0,123,0,20,0,142,0,0,0,176,0,20,0,217,0,181,0,235,0,168,0,0,0,157,0,0,0,134,0,226,0,18,0,0,0,125,0,0,0,154,0,224,0,137,0,119,0,135,0,0,0,215,0,235,0,159,0,0,0,0,0,160,0,117,0,175,0,19,0,41,0,0,0,0,0,249,0,0,0,194,0,81,0,225,0,226,0,0,0,244,0,0,0,58,0,73,0,104,0,183,0,0,0,0,0,0,0,0,0,22,0,0,0,0,0,0,0,151,0,87,0,25,0,0,0,117,0,0,0,0,0,232,0,162,0,173,0,217,0,174,0,69,0,111,0,0,0,0,0,181,0,170,0,9,0,29,0,57,0,17,0,110,0,40,0,47,0,31,0,0,0,0,0,110,0,117,0,178,0,0,0,157,0,98,0,72,0,0,0,225,0,108,0,13,0,152,0,0,0,66,0,132,0,0,0,236,0,212,0,0,0,162,0,95,0,46,0,22,0,175,0,220,0,213,0,0,0,11,0,113,0,76,0,94,0,119,0,124,0,155,0,181,0,181,0,0,0,0,0,0,0,189,0,69,0,169,0,11,0,0,0,82,0,238,0,5,0,14,0,0,0,205,0,141,0,23,0,33,0,196,0,140,0,41,0,49,0,45,0,83,0,192,0,0,0,224,0,0,0,171,0,109,0,164,0,0,0,207,0,198,0,60,0,0,0,31,0,0,0,80,0,203,0,235,0,17,0,47,0,0,0,0,0,169,0,0,0,249,0,98,0,26,0,68,0,150,0,0,0,49,0,0,0,8,0,160,0,237,0,132,0,189,0,220,0,69,0,45,0,216,0,47,0,1,0,132,0,0,0,0,0,29,0,127,0,225,0,235,0,168,0,184,0,67,0,146,0,0,0,249,0,0,0,246,0,54,0,60,0,220,0,5,0,70,0,155,0,188,0,241,0,233,0,59,0,77,0,145,0,0,0,0,0,56,0,8,0,138,0,161,0,225,0,252,0,184,0,78,0,114,0,168,0,163,0,0,0,195,0,119,0,0,0,98,0,42,0,0,0,225,0,232,0,0,0,193,0,19,0,0,0,0,0,119,0,191,0,91,0,0,0,0,0,0,0,67,0,201,0,223,0,97,0,165,0,0,0,249,0,111,0,152,0,193,0,191,0,0,0,212,0,102,0,177,0,158,0,127,0,0,0,34,0,111,0,56,0,0,0,54,0,203,0,57,0,100,0,139,0,0,0,1,0,62,0,45,0,0,0,35,0,0,0,0,0,84,0,253,0,95,0,0,0,229,0,0,0,122,0,60,0,201,0,234,0,217,0,2,0,223,0,249,0,250,0,128,0,91,0,119,0,255,0,0,0,0,0,43,0,255,0,211,0,187,0,30,0,229,0,43,0,24,0,253,0,10,0,223,0,74,0,124,0,165,0,97,0,0,0,241,0,0,0,30,0,33,0,0,0,148,0,0,0,222,0,6,0,14,0,151,0,147,0,148,0,151,0,0,0,207,0,62,0,218,0,90,0,0,0,79,0,75,0,11,0,52,0,211,0,162,0,50,0,56,0,231,0,16,0,14,0);
signal scenario_full  : scenario_type := (96,31,96,30,216,31,196,31,175,31,244,31,108,31,111,31,124,31,124,30,12,31,83,31,222,31,23,31,241,31,202,31,159,31,136,31,162,31,162,30,140,31,244,31,4,31,117,31,101,31,203,31,203,30,141,31,199,31,194,31,194,30,236,31,226,31,1,31,83,31,83,30,101,31,101,30,224,31,224,30,45,31,164,31,164,30,101,31,140,31,174,31,189,31,189,30,202,31,198,31,98,31,159,31,51,31,51,30,26,31,235,31,235,30,230,31,136,31,136,30,136,29,231,31,181,31,194,31,95,31,31,31,109,31,208,31,95,31,178,31,138,31,132,31,213,31,213,30,109,31,109,30,109,29,19,31,158,31,193,31,193,30,203,31,173,31,213,31,82,31,113,31,59,31,59,30,59,29,36,31,249,31,249,30,40,31,100,31,100,30,100,29,212,31,105,31,125,31,207,31,222,31,88,31,88,30,122,31,177,31,76,31,76,30,76,29,76,28,97,31,117,31,163,31,163,30,102,31,102,30,156,31,45,31,6,31,27,31,252,31,250,31,138,31,138,30,55,31,219,31,127,31,37,31,214,31,182,31,182,30,182,29,200,31,202,31,202,30,5,31,3,31,246,31,57,31,202,31,86,31,86,30,86,29,86,28,231,31,231,30,42,31,244,31,106,31,63,31,63,30,186,31,210,31,13,31,96,31,96,30,231,31,211,31,211,30,192,31,155,31,150,31,138,31,112,31,130,31,97,31,68,31,96,31,240,31,44,31,190,31,227,31,254,31,168,31,171,31,224,31,224,30,13,31,13,31,78,31,54,31,175,31,23,31,23,30,17,31,183,31,209,31,53,31,167,31,42,31,105,31,133,31,242,31,254,31,53,31,219,31,2,31,182,31,128,31,68,31,105,31,72,31,170,31,164,31,136,31,244,31,244,30,144,31,248,31,2,31,72,31,72,30,35,31,35,30,35,29,174,31,193,31,153,31,180,31,208,31,243,31,176,31,176,30,201,31,201,30,240,31,240,30,6,31,99,31,206,31,227,31,193,31,124,31,124,30,43,31,43,30,75,31,75,30,75,29,25,31,236,31,22,31,36,31,222,31,115,31,115,30,58,31,158,31,43,31,43,30,74,31,74,30,50,31,38,31,38,30,105,31,44,31,168,31,165,31,175,31,181,31,245,31,160,31,103,31,6,31,170,31,170,30,219,31,219,30,138,31,219,31,115,31,28,31,231,31,190,31,99,31,144,31,137,31,29,31,119,31,180,31,55,31,55,30,3,31,249,31,62,31,71,31,71,30,46,31,121,31,233,31,166,31,73,31,124,31,52,31,107,31,107,30,86,31,86,30,152,31,234,31,58,31,37,31,156,31,48,31,141,31,84,31,29,31,5,31,249,31,98,31,195,31,121,31,121,30,243,31,243,30,153,31,153,30,69,31,222,31,62,31,169,31,248,31,89,31,89,30,241,31,204,31,119,31,171,31,248,31,41,31,55,31,63,31,128,31,82,31,62,31,109,31,100,31,168,31,82,31,180,31,66,31,205,31,60,31,122,31,158,31,146,31,36,31,176,31,203,31,222,31,104,31,226,31,210,31,48,31,48,30,48,29,233,31,19,31,71,31,70,31,244,31,236,31,1,31,137,31,159,31,165,31,235,31,156,31,156,30,156,29,103,31,34,31,182,31,24,31,24,30,24,29,20,31,39,31,165,31,99,31,122,31,158,31,158,30,162,31,89,31,155,31,207,31,126,31,185,31,39,31,39,30,39,29,94,31,7,31,38,31,38,30,103,31,209,31,196,31,196,30,54,31,154,31,119,31,196,31,59,31,59,30,184,31,19,31,21,31,13,31,189,31,34,31,33,31,93,31,88,31,88,30,88,29,128,31,5,31,5,30,5,29,243,31,37,31,229,31,229,31,161,31,33,31,33,30,37,31,235,31,197,31,28,31,28,30,179,31,113,31,138,31,138,30,98,31,197,31,192,31,10,31,148,31,35,31,153,31,101,31,101,30,6,31,249,31,29,31,90,31,27,31,58,31,211,31,211,30,199,31,199,30,44,31,121,31,154,31,54,31,216,31,96,31,214,31,154,31,75,31,74,31,150,31,106,31,65,31,43,31,145,31,145,30,145,29,194,31,205,31,152,31,100,31,214,31,244,31,108,31,108,30,108,29,49,31,178,31,117,31,34,31,16,31,127,31,191,31,46,31,243,31,194,31,240,31,196,31,179,31,148,31,42,31,180,31,211,31,211,30,211,29,171,31,238,31,188,31,110,31,72,31,72,30,159,31,223,31,104,31,111,31,255,31,173,31,241,31,117,31,128,31,128,30,123,31,20,31,142,31,142,30,176,31,20,31,217,31,181,31,235,31,168,31,168,30,157,31,157,30,134,31,226,31,18,31,18,30,125,31,125,30,154,31,224,31,137,31,119,31,135,31,135,30,215,31,235,31,159,31,159,30,159,29,160,31,117,31,175,31,19,31,41,31,41,30,41,29,249,31,249,30,194,31,81,31,225,31,226,31,226,30,244,31,244,30,58,31,73,31,104,31,183,31,183,30,183,29,183,28,183,27,22,31,22,30,22,29,22,28,151,31,87,31,25,31,25,30,117,31,117,30,117,29,232,31,162,31,173,31,217,31,174,31,69,31,111,31,111,30,111,29,181,31,170,31,9,31,29,31,57,31,17,31,110,31,40,31,47,31,31,31,31,30,31,29,110,31,117,31,178,31,178,30,157,31,98,31,72,31,72,30,225,31,108,31,13,31,152,31,152,30,66,31,132,31,132,30,236,31,212,31,212,30,162,31,95,31,46,31,22,31,175,31,220,31,213,31,213,30,11,31,113,31,76,31,94,31,119,31,124,31,155,31,181,31,181,31,181,30,181,29,181,28,189,31,69,31,169,31,11,31,11,30,82,31,238,31,5,31,14,31,14,30,205,31,141,31,23,31,33,31,196,31,140,31,41,31,49,31,45,31,83,31,192,31,192,30,224,31,224,30,171,31,109,31,164,31,164,30,207,31,198,31,60,31,60,30,31,31,31,30,80,31,203,31,235,31,17,31,47,31,47,30,47,29,169,31,169,30,249,31,98,31,26,31,68,31,150,31,150,30,49,31,49,30,8,31,160,31,237,31,132,31,189,31,220,31,69,31,45,31,216,31,47,31,1,31,132,31,132,30,132,29,29,31,127,31,225,31,235,31,168,31,184,31,67,31,146,31,146,30,249,31,249,30,246,31,54,31,60,31,220,31,5,31,70,31,155,31,188,31,241,31,233,31,59,31,77,31,145,31,145,30,145,29,56,31,8,31,138,31,161,31,225,31,252,31,184,31,78,31,114,31,168,31,163,31,163,30,195,31,119,31,119,30,98,31,42,31,42,30,225,31,232,31,232,30,193,31,19,31,19,30,19,29,119,31,191,31,91,31,91,30,91,29,91,28,67,31,201,31,223,31,97,31,165,31,165,30,249,31,111,31,152,31,193,31,191,31,191,30,212,31,102,31,177,31,158,31,127,31,127,30,34,31,111,31,56,31,56,30,54,31,203,31,57,31,100,31,139,31,139,30,1,31,62,31,45,31,45,30,35,31,35,30,35,29,84,31,253,31,95,31,95,30,229,31,229,30,122,31,60,31,201,31,234,31,217,31,2,31,223,31,249,31,250,31,128,31,91,31,119,31,255,31,255,30,255,29,43,31,255,31,211,31,187,31,30,31,229,31,43,31,24,31,253,31,10,31,223,31,74,31,124,31,165,31,97,31,97,30,241,31,241,30,30,31,33,31,33,30,148,31,148,30,222,31,6,31,14,31,151,31,147,31,148,31,151,31,151,30,207,31,62,31,218,31,90,31,90,30,79,31,75,31,11,31,52,31,211,31,162,31,50,31,56,31,231,31,16,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
