-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 887;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (81,0,214,0,198,0,0,0,153,0,227,0,96,0,180,0,203,0,0,0,164,0,39,0,247,0,62,0,68,0,250,0,135,0,28,0,170,0,49,0,190,0,0,0,0,0,244,0,88,0,109,0,158,0,230,0,187,0,123,0,219,0,202,0,0,0,253,0,175,0,161,0,0,0,169,0,140,0,32,0,101,0,229,0,0,0,0,0,152,0,0,0,89,0,40,0,59,0,218,0,198,0,104,0,65,0,44,0,182,0,59,0,40,0,179,0,249,0,44,0,96,0,137,0,194,0,193,0,249,0,110,0,114,0,149,0,0,0,0,0,247,0,109,0,55,0,15,0,98,0,0,0,0,0,97,0,0,0,89,0,37,0,178,0,0,0,248,0,5,0,58,0,195,0,17,0,198,0,56,0,0,0,0,0,16,0,178,0,46,0,36,0,125,0,240,0,68,0,255,0,106,0,24,0,21,0,203,0,157,0,24,0,234,0,64,0,98,0,76,0,126,0,0,0,0,0,47,0,0,0,209,0,184,0,176,0,205,0,185,0,0,0,31,0,63,0,158,0,187,0,29,0,58,0,213,0,118,0,0,0,0,0,26,0,102,0,0,0,32,0,0,0,54,0,0,0,76,0,0,0,201,0,0,0,0,0,187,0,210,0,0,0,82,0,250,0,29,0,91,0,126,0,160,0,37,0,126,0,3,0,88,0,111,0,97,0,252,0,230,0,245,0,90,0,0,0,0,0,0,0,64,0,0,0,239,0,0,0,232,0,116,0,206,0,226,0,212,0,0,0,0,0,51,0,0,0,85,0,184,0,112,0,100,0,0,0,89,0,0,0,0,0,90,0,238,0,163,0,245,0,119,0,34,0,12,0,0,0,10,0,175,0,0,0,45,0,34,0,165,0,167,0,246,0,0,0,0,0,172,0,157,0,75,0,0,0,80,0,219,0,71,0,121,0,241,0,66,0,127,0,0,0,222,0,108,0,137,0,51,0,0,0,137,0,130,0,7,0,66,0,31,0,148,0,255,0,45,0,15,0,167,0,44,0,255,0,205,0,67,0,41,0,96,0,14,0,93,0,0,0,132,0,94,0,135,0,138,0,247,0,229,0,73,0,58,0,0,0,112,0,77,0,114,0,186,0,8,0,0,0,3,0,88,0,37,0,14,0,105,0,7,0,39,0,88,0,0,0,0,0,77,0,201,0,70,0,224,0,92,0,152,0,0,0,0,0,28,0,216,0,0,0,0,0,121,0,245,0,132,0,158,0,153,0,178,0,0,0,0,0,194,0,111,0,230,0,105,0,35,0,0,0,220,0,176,0,0,0,233,0,242,0,48,0,77,0,0,0,222,0,0,0,138,0,223,0,0,0,251,0,197,0,103,0,0,0,103,0,187,0,42,0,202,0,36,0,40,0,248,0,134,0,206,0,233,0,231,0,44,0,100,0,0,0,108,0,62,0,0,0,208,0,180,0,18,0,74,0,225,0,234,0,197,0,235,0,78,0,165,0,190,0,0,0,93,0,102,0,0,0,0,0,253,0,132,0,39,0,231,0,39,0,25,0,68,0,107,0,0,0,130,0,38,0,81,0,233,0,70,0,28,0,119,0,200,0,78,0,0,0,152,0,87,0,0,0,73,0,99,0,226,0,0,0,174,0,133,0,21,0,144,0,5,0,0,0,162,0,188,0,55,0,155,0,183,0,0,0,22,0,29,0,143,0,223,0,201,0,245,0,202,0,0,0,0,0,216,0,200,0,35,0,158,0,163,0,13,0,21,0,33,0,150,0,239,0,201,0,165,0,195,0,44,0,198,0,225,0,215,0,146,0,141,0,129,0,36,0,213,0,37,0,251,0,53,0,0,0,15,0,160,0,0,0,0,0,0,0,76,0,0,0,0,0,0,0,241,0,183,0,0,0,28,0,160,0,0,0,33,0,0,0,0,0,217,0,0,0,190,0,148,0,83,0,161,0,220,0,114,0,11,0,43,0,0,0,181,0,229,0,0,0,230,0,0,0,0,0,117,0,95,0,0,0,0,0,205,0,108,0,0,0,177,0,0,0,85,0,193,0,0,0,209,0,14,0,140,0,0,0,0,0,91,0,57,0,254,0,0,0,130,0,180,0,54,0,110,0,13,0,0,0,238,0,244,0,126,0,0,0,94,0,0,0,233,0,13,0,36,0,0,0,49,0,194,0,31,0,62,0,0,0,101,0,172,0,146,0,75,0,223,0,247,0,178,0,177,0,136,0,224,0,140,0,219,0,73,0,174,0,169,0,115,0,45,0,109,0,0,0,23,0,0,0,32,0,135,0,52,0,251,0,34,0,0,0,0,0,114,0,4,0,16,0,153,0,193,0,70,0,33,0,213,0,1,0,0,0,45,0,0,0,91,0,148,0,218,0,41,0,239,0,0,0,2,0,0,0,20,0,190,0,192,0,66,0,75,0,171,0,98,0,173,0,0,0,112,0,32,0,86,0,109,0,239,0,0,0,81,0,91,0,0,0,10,0,231,0,92,0,220,0,0,0,215,0,123,0,0,0,183,0,63,0,218,0,166,0,243,0,59,0,164,0,7,0,0,0,35,0,0,0,191,0,254,0,0,0,96,0,0,0,205,0,84,0,105,0,0,0,227,0,124,0,192,0,91,0,0,0,0,0,138,0,246,0,35,0,175,0,242,0,49,0,110,0,109,0,233,0,113,0,168,0,86,0,0,0,104,0,229,0,0,0,74,0,43,0,74,0,126,0,150,0,86,0,0,0,139,0,18,0,89,0,55,0,0,0,0,0,7,0,0,0,0,0,4,0,0,0,111,0,220,0,137,0,124,0,239,0,198,0,56,0,223,0,151,0,27,0,220,0,200,0,187,0,118,0,0,0,24,0,0,0,173,0,121,0,52,0,118,0,101,0,206,0,0,0,20,0,165,0,0,0,140,0,49,0,0,0,241,0,128,0,0,0,126,0,96,0,29,0,169,0,93,0,54,0,249,0,160,0,118,0,51,0,178,0,0,0,156,0,203,0,75,0,37,0,73,0,211,0,160,0,0,0,45,0,130,0,0,0,0,0,0,0,184,0,131,0,167,0,30,0,193,0,131,0,38,0,118,0,0,0,87,0,43,0,2,0,0,0,0,0,80,0,0,0,78,0,23,0,236,0,179,0,102,0,2,0,85,0,226,0,0,0,171,0,0,0,8,0,0,0,0,0,193,0,232,0,231,0,7,0,0,0,50,0,83,0,175,0,0,0,69,0,25,0,238,0,28,0,0,0,103,0,70,0,0,0,172,0,130,0,0,0,15,0,103,0,105,0,24,0,122,0,0,0,11,0,214,0,17,0,97,0,92,0,0,0,175,0,27,0,105,0,95,0,247,0,0,0,0,0,0,0,216,0,0,0,165,0,0,0,3,0,57,0,107,0,150,0,70,0,152,0,54,0,164,0,43,0,79,0,131,0,46,0,19,0,133,0,0,0,236,0,88,0,172,0,160,0,16,0,104,0,0,0,79,0,190,0,0,0,11,0,85,0,242,0,0,0,220,0,36,0,181,0,96,0,79,0,189,0,0,0,145,0,0,0,172,0,121,0,50,0,70,0,20,0,229,0,194,0,0,0,196,0,78,0,171,0,151,0,193,0,0,0,18,0,197,0,214,0,221,0,122,0,91,0,44,0,233,0,142,0,246,0,25,0,218,0,243,0,103,0,11,0,144,0,0,0,198,0,184,0,94,0,142,0,226,0,83,0,52,0,187,0,59,0,64,0,226,0,105,0,68,0,181,0,165,0,209,0,134,0,156,0,0,0,41,0,0,0,83,0,240,0,157,0,250,0,39,0,254,0,196,0,120,0,77,0,76,0,0,0,157,0,0,0,0,0,227,0,203,0,48,0,25,0,250,0,205,0,183,0,0,0,151,0,0,0,70,0,234,0,66,0,31,0,109,0,0,0,26,0,29,0,0,0,98,0,20,0,62,0,254,0,0,0,0,0,141,0);
signal scenario_full  : scenario_type := (81,31,214,31,198,31,198,30,153,31,227,31,96,31,180,31,203,31,203,30,164,31,39,31,247,31,62,31,68,31,250,31,135,31,28,31,170,31,49,31,190,31,190,30,190,29,244,31,88,31,109,31,158,31,230,31,187,31,123,31,219,31,202,31,202,30,253,31,175,31,161,31,161,30,169,31,140,31,32,31,101,31,229,31,229,30,229,29,152,31,152,30,89,31,40,31,59,31,218,31,198,31,104,31,65,31,44,31,182,31,59,31,40,31,179,31,249,31,44,31,96,31,137,31,194,31,193,31,249,31,110,31,114,31,149,31,149,30,149,29,247,31,109,31,55,31,15,31,98,31,98,30,98,29,97,31,97,30,89,31,37,31,178,31,178,30,248,31,5,31,58,31,195,31,17,31,198,31,56,31,56,30,56,29,16,31,178,31,46,31,36,31,125,31,240,31,68,31,255,31,106,31,24,31,21,31,203,31,157,31,24,31,234,31,64,31,98,31,76,31,126,31,126,30,126,29,47,31,47,30,209,31,184,31,176,31,205,31,185,31,185,30,31,31,63,31,158,31,187,31,29,31,58,31,213,31,118,31,118,30,118,29,26,31,102,31,102,30,32,31,32,30,54,31,54,30,76,31,76,30,201,31,201,30,201,29,187,31,210,31,210,30,82,31,250,31,29,31,91,31,126,31,160,31,37,31,126,31,3,31,88,31,111,31,97,31,252,31,230,31,245,31,90,31,90,30,90,29,90,28,64,31,64,30,239,31,239,30,232,31,116,31,206,31,226,31,212,31,212,30,212,29,51,31,51,30,85,31,184,31,112,31,100,31,100,30,89,31,89,30,89,29,90,31,238,31,163,31,245,31,119,31,34,31,12,31,12,30,10,31,175,31,175,30,45,31,34,31,165,31,167,31,246,31,246,30,246,29,172,31,157,31,75,31,75,30,80,31,219,31,71,31,121,31,241,31,66,31,127,31,127,30,222,31,108,31,137,31,51,31,51,30,137,31,130,31,7,31,66,31,31,31,148,31,255,31,45,31,15,31,167,31,44,31,255,31,205,31,67,31,41,31,96,31,14,31,93,31,93,30,132,31,94,31,135,31,138,31,247,31,229,31,73,31,58,31,58,30,112,31,77,31,114,31,186,31,8,31,8,30,3,31,88,31,37,31,14,31,105,31,7,31,39,31,88,31,88,30,88,29,77,31,201,31,70,31,224,31,92,31,152,31,152,30,152,29,28,31,216,31,216,30,216,29,121,31,245,31,132,31,158,31,153,31,178,31,178,30,178,29,194,31,111,31,230,31,105,31,35,31,35,30,220,31,176,31,176,30,233,31,242,31,48,31,77,31,77,30,222,31,222,30,138,31,223,31,223,30,251,31,197,31,103,31,103,30,103,31,187,31,42,31,202,31,36,31,40,31,248,31,134,31,206,31,233,31,231,31,44,31,100,31,100,30,108,31,62,31,62,30,208,31,180,31,18,31,74,31,225,31,234,31,197,31,235,31,78,31,165,31,190,31,190,30,93,31,102,31,102,30,102,29,253,31,132,31,39,31,231,31,39,31,25,31,68,31,107,31,107,30,130,31,38,31,81,31,233,31,70,31,28,31,119,31,200,31,78,31,78,30,152,31,87,31,87,30,73,31,99,31,226,31,226,30,174,31,133,31,21,31,144,31,5,31,5,30,162,31,188,31,55,31,155,31,183,31,183,30,22,31,29,31,143,31,223,31,201,31,245,31,202,31,202,30,202,29,216,31,200,31,35,31,158,31,163,31,13,31,21,31,33,31,150,31,239,31,201,31,165,31,195,31,44,31,198,31,225,31,215,31,146,31,141,31,129,31,36,31,213,31,37,31,251,31,53,31,53,30,15,31,160,31,160,30,160,29,160,28,76,31,76,30,76,29,76,28,241,31,183,31,183,30,28,31,160,31,160,30,33,31,33,30,33,29,217,31,217,30,190,31,148,31,83,31,161,31,220,31,114,31,11,31,43,31,43,30,181,31,229,31,229,30,230,31,230,30,230,29,117,31,95,31,95,30,95,29,205,31,108,31,108,30,177,31,177,30,85,31,193,31,193,30,209,31,14,31,140,31,140,30,140,29,91,31,57,31,254,31,254,30,130,31,180,31,54,31,110,31,13,31,13,30,238,31,244,31,126,31,126,30,94,31,94,30,233,31,13,31,36,31,36,30,49,31,194,31,31,31,62,31,62,30,101,31,172,31,146,31,75,31,223,31,247,31,178,31,177,31,136,31,224,31,140,31,219,31,73,31,174,31,169,31,115,31,45,31,109,31,109,30,23,31,23,30,32,31,135,31,52,31,251,31,34,31,34,30,34,29,114,31,4,31,16,31,153,31,193,31,70,31,33,31,213,31,1,31,1,30,45,31,45,30,91,31,148,31,218,31,41,31,239,31,239,30,2,31,2,30,20,31,190,31,192,31,66,31,75,31,171,31,98,31,173,31,173,30,112,31,32,31,86,31,109,31,239,31,239,30,81,31,91,31,91,30,10,31,231,31,92,31,220,31,220,30,215,31,123,31,123,30,183,31,63,31,218,31,166,31,243,31,59,31,164,31,7,31,7,30,35,31,35,30,191,31,254,31,254,30,96,31,96,30,205,31,84,31,105,31,105,30,227,31,124,31,192,31,91,31,91,30,91,29,138,31,246,31,35,31,175,31,242,31,49,31,110,31,109,31,233,31,113,31,168,31,86,31,86,30,104,31,229,31,229,30,74,31,43,31,74,31,126,31,150,31,86,31,86,30,139,31,18,31,89,31,55,31,55,30,55,29,7,31,7,30,7,29,4,31,4,30,111,31,220,31,137,31,124,31,239,31,198,31,56,31,223,31,151,31,27,31,220,31,200,31,187,31,118,31,118,30,24,31,24,30,173,31,121,31,52,31,118,31,101,31,206,31,206,30,20,31,165,31,165,30,140,31,49,31,49,30,241,31,128,31,128,30,126,31,96,31,29,31,169,31,93,31,54,31,249,31,160,31,118,31,51,31,178,31,178,30,156,31,203,31,75,31,37,31,73,31,211,31,160,31,160,30,45,31,130,31,130,30,130,29,130,28,184,31,131,31,167,31,30,31,193,31,131,31,38,31,118,31,118,30,87,31,43,31,2,31,2,30,2,29,80,31,80,30,78,31,23,31,236,31,179,31,102,31,2,31,85,31,226,31,226,30,171,31,171,30,8,31,8,30,8,29,193,31,232,31,231,31,7,31,7,30,50,31,83,31,175,31,175,30,69,31,25,31,238,31,28,31,28,30,103,31,70,31,70,30,172,31,130,31,130,30,15,31,103,31,105,31,24,31,122,31,122,30,11,31,214,31,17,31,97,31,92,31,92,30,175,31,27,31,105,31,95,31,247,31,247,30,247,29,247,28,216,31,216,30,165,31,165,30,3,31,57,31,107,31,150,31,70,31,152,31,54,31,164,31,43,31,79,31,131,31,46,31,19,31,133,31,133,30,236,31,88,31,172,31,160,31,16,31,104,31,104,30,79,31,190,31,190,30,11,31,85,31,242,31,242,30,220,31,36,31,181,31,96,31,79,31,189,31,189,30,145,31,145,30,172,31,121,31,50,31,70,31,20,31,229,31,194,31,194,30,196,31,78,31,171,31,151,31,193,31,193,30,18,31,197,31,214,31,221,31,122,31,91,31,44,31,233,31,142,31,246,31,25,31,218,31,243,31,103,31,11,31,144,31,144,30,198,31,184,31,94,31,142,31,226,31,83,31,52,31,187,31,59,31,64,31,226,31,105,31,68,31,181,31,165,31,209,31,134,31,156,31,156,30,41,31,41,30,83,31,240,31,157,31,250,31,39,31,254,31,196,31,120,31,77,31,76,31,76,30,157,31,157,30,157,29,227,31,203,31,48,31,25,31,250,31,205,31,183,31,183,30,151,31,151,30,70,31,234,31,66,31,31,31,109,31,109,30,26,31,29,31,29,30,98,31,20,31,62,31,254,31,254,30,254,29,141,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
