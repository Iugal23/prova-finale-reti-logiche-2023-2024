-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 954;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,162,0,0,0,0,0,0,0,112,0,210,0,222,0,222,0,242,0,2,0,217,0,92,0,207,0,33,0,89,0,193,0,159,0,117,0,148,0,1,0,213,0,117,0,53,0,0,0,175,0,127,0,109,0,0,0,42,0,0,0,93,0,0,0,55,0,0,0,45,0,107,0,69,0,0,0,87,0,37,0,0,0,241,0,148,0,239,0,226,0,250,0,210,0,0,0,82,0,52,0,118,0,194,0,158,0,253,0,0,0,112,0,120,0,229,0,58,0,0,0,93,0,0,0,1,0,26,0,52,0,0,0,192,0,200,0,59,0,161,0,180,0,0,0,192,0,0,0,85,0,230,0,187,0,61,0,92,0,209,0,0,0,16,0,174,0,140,0,175,0,0,0,216,0,224,0,0,0,159,0,58,0,96,0,0,0,235,0,0,0,0,0,202,0,127,0,244,0,102,0,230,0,129,0,36,0,245,0,177,0,96,0,220,0,216,0,61,0,0,0,0,0,0,0,0,0,127,0,83,0,24,0,16,0,43,0,135,0,223,0,3,0,116,0,207,0,83,0,79,0,228,0,158,0,0,0,0,0,121,0,111,0,70,0,37,0,203,0,189,0,227,0,247,0,89,0,120,0,0,0,224,0,235,0,180,0,0,0,68,0,41,0,252,0,218,0,7,0,154,0,144,0,47,0,106,0,228,0,50,0,253,0,87,0,45,0,148,0,131,0,137,0,169,0,0,0,142,0,148,0,238,0,224,0,245,0,77,0,0,0,4,0,126,0,55,0,247,0,0,0,226,0,110,0,10,0,124,0,15,0,202,0,230,0,142,0,82,0,128,0,0,0,195,0,0,0,31,0,129,0,34,0,0,0,216,0,0,0,40,0,226,0,225,0,72,0,0,0,238,0,167,0,0,0,93,0,66,0,117,0,58,0,139,0,0,0,197,0,158,0,206,0,148,0,204,0,200,0,0,0,0,0,117,0,100,0,216,0,189,0,233,0,112,0,128,0,158,0,47,0,231,0,193,0,28,0,166,0,182,0,0,0,68,0,89,0,207,0,0,0,0,0,168,0,138,0,94,0,0,0,205,0,0,0,164,0,49,0,182,0,3,0,57,0,0,0,49,0,232,0,0,0,0,0,111,0,244,0,112,0,209,0,85,0,7,0,238,0,65,0,0,0,216,0,0,0,30,0,82,0,50,0,12,0,42,0,25,0,0,0,0,0,7,0,102,0,46,0,128,0,0,0,0,0,205,0,247,0,11,0,181,0,0,0,126,0,155,0,156,0,244,0,174,0,149,0,56,0,111,0,141,0,89,0,238,0,30,0,251,0,186,0,129,0,252,0,29,0,155,0,65,0,181,0,49,0,58,0,227,0,0,0,61,0,27,0,0,0,1,0,155,0,144,0,192,0,6,0,0,0,203,0,26,0,0,0,208,0,20,0,176,0,245,0,13,0,160,0,0,0,84,0,71,0,0,0,0,0,0,0,237,0,87,0,0,0,123,0,0,0,213,0,0,0,225,0,72,0,123,0,197,0,1,0,212,0,14,0,134,0,74,0,140,0,168,0,0,0,209,0,62,0,0,0,127,0,95,0,10,0,181,0,235,0,26,0,93,0,0,0,228,0,0,0,131,0,0,0,18,0,5,0,0,0,171,0,208,0,143,0,131,0,135,0,192,0,0,0,0,0,61,0,205,0,117,0,141,0,0,0,103,0,18,0,0,0,0,0,175,0,0,0,0,0,129,0,193,0,195,0,0,0,168,0,193,0,230,0,144,0,194,0,13,0,95,0,98,0,53,0,0,0,111,0,207,0,157,0,0,0,22,0,85,0,187,0,67,0,176,0,16,0,0,0,136,0,138,0,79,0,0,0,2,0,0,0,240,0,3,0,62,0,156,0,98,0,183,0,131,0,131,0,155,0,149,0,168,0,22,0,27,0,17,0,187,0,92,0,199,0,0,0,230,0,133,0,79,0,228,0,62,0,0,0,0,0,18,0,43,0,0,0,166,0,193,0,0,0,0,0,219,0,66,0,207,0,255,0,187,0,219,0,27,0,56,0,146,0,151,0,235,0,207,0,0,0,161,0,76,0,76,0,0,0,0,0,50,0,200,0,212,0,221,0,184,0,181,0,85,0,157,0,226,0,76,0,68,0,77,0,153,0,254,0,0,0,0,0,160,0,90,0,109,0,231,0,140,0,19,0,0,0,0,0,155,0,138,0,143,0,209,0,230,0,0,0,231,0,159,0,111,0,116,0,81,0,21,0,42,0,218,0,40,0,14,0,4,0,0,0,149,0,229,0,230,0,139,0,16,0,93,0,0,0,126,0,230,0,37,0,0,0,0,0,0,0,96,0,0,0,0,0,40,0,182,0,30,0,0,0,7,0,121,0,148,0,205,0,0,0,80,0,0,0,18,0,195,0,103,0,221,0,122,0,58,0,0,0,230,0,180,0,180,0,104,0,245,0,40,0,117,0,89,0,68,0,190,0,138,0,244,0,115,0,243,0,173,0,132,0,0,0,197,0,8,0,0,0,97,0,189,0,18,0,172,0,108,0,189,0,178,0,0,0,133,0,0,0,0,0,103,0,200,0,89,0,0,0,135,0,239,0,0,0,0,0,217,0,226,0,228,0,179,0,222,0,0,0,0,0,65,0,11,0,173,0,0,0,16,0,138,0,8,0,73,0,0,0,130,0,158,0,176,0,124,0,75,0,12,0,103,0,85,0,61,0,70,0,7,0,140,0,63,0,214,0,221,0,228,0,125,0,0,0,154,0,0,0,50,0,0,0,204,0,110,0,157,0,10,0,53,0,192,0,80,0,210,0,43,0,107,0,0,0,131,0,103,0,159,0,123,0,128,0,0,0,3,0,191,0,129,0,161,0,252,0,139,0,97,0,0,0,0,0,5,0,0,0,73,0,1,0,98,0,15,0,213,0,247,0,78,0,140,0,162,0,55,0,6,0,165,0,169,0,239,0,0,0,244,0,0,0,116,0,171,0,28,0,20,0,188,0,202,0,0,0,32,0,14,0,116,0,208,0,242,0,116,0,120,0,168,0,0,0,0,0,0,0,128,0,130,0,107,0,1,0,148,0,172,0,0,0,145,0,5,0,204,0,90,0,0,0,94,0,187,0,111,0,16,0,59,0,155,0,75,0,108,0,65,0,244,0,136,0,70,0,45,0,114,0,41,0,199,0,29,0,193,0,0,0,164,0,87,0,210,0,90,0,115,0,0,0,224,0,2,0,134,0,74,0,73,0,0,0,10,0,0,0,0,0,47,0,0,0,198,0,21,0,0,0,134,0,37,0,70,0,204,0,107,0,231,0,151,0,12,0,0,0,186,0,195,0,162,0,240,0,97,0,139,0,71,0,200,0,0,0,0,0,117,0,29,0,0,0,165,0,138,0,130,0,0,0,0,0,0,0,164,0,158,0,0,0,0,0,202,0,120,0,197,0,185,0,193,0,0,0,117,0,0,0,0,0,72,0,25,0,231,0,0,0,133,0,91,0,36,0,96,0,191,0,212,0,78,0,135,0,92,0,0,0,213,0,223,0,7,0,235,0,0,0,128,0,0,0,66,0,0,0,150,0,89,0,136,0,199,0,127,0,191,0,0,0,0,0,39,0,191,0,0,0,11,0,233,0,43,0,206,0,140,0,224,0,11,0,224,0,166,0,241,0,183,0,95,0,196,0,98,0,35,0,133,0,42,0,101,0,118,0,249,0,70,0,173,0,0,0,135,0,0,0,189,0,85,0,180,0,10,0,153,0,127,0,0,0,78,0,135,0,0,0,172,0,0,0,0,0,104,0,0,0,15,0,0,0,70,0,0,0,0,0,201,0,182,0,28,0,0,0,148,0,103,0,0,0,30,0,88,0,23,0,0,0,45,0,62,0,17,0,99,0,0,0,0,0,0,0,104,0,210,0,0,0,83,0,0,0,235,0,62,0,3,0,251,0,172,0,235,0,36,0,77,0,27,0,30,0,111,0,49,0,70,0,191,0,15,0,197,0,144,0,156,0,107,0,181,0,82,0,134,0,0,0,253,0,221,0,84,0,10,0,153,0,179,0,250,0,0,0,66,0,27,0,229,0,25,0,108,0,0,0,22,0,143,0,16,0,66,0,0,0,0,0,155,0,0,0,179,0,210,0,58,0,85,0,0,0,0,0,177,0,10,0,229,0,0,0,240,0,249,0,6,0,129,0,39,0,52,0,143,0,226,0,227,0,142,0,123,0,192,0,49,0,104,0,16,0,0,0,0,0,0,0,0,0,127,0);
signal scenario_full  : scenario_type := (195,31,162,31,162,30,162,29,162,28,112,31,210,31,222,31,222,31,242,31,2,31,217,31,92,31,207,31,33,31,89,31,193,31,159,31,117,31,148,31,1,31,213,31,117,31,53,31,53,30,175,31,127,31,109,31,109,30,42,31,42,30,93,31,93,30,55,31,55,30,45,31,107,31,69,31,69,30,87,31,37,31,37,30,241,31,148,31,239,31,226,31,250,31,210,31,210,30,82,31,52,31,118,31,194,31,158,31,253,31,253,30,112,31,120,31,229,31,58,31,58,30,93,31,93,30,1,31,26,31,52,31,52,30,192,31,200,31,59,31,161,31,180,31,180,30,192,31,192,30,85,31,230,31,187,31,61,31,92,31,209,31,209,30,16,31,174,31,140,31,175,31,175,30,216,31,224,31,224,30,159,31,58,31,96,31,96,30,235,31,235,30,235,29,202,31,127,31,244,31,102,31,230,31,129,31,36,31,245,31,177,31,96,31,220,31,216,31,61,31,61,30,61,29,61,28,61,27,127,31,83,31,24,31,16,31,43,31,135,31,223,31,3,31,116,31,207,31,83,31,79,31,228,31,158,31,158,30,158,29,121,31,111,31,70,31,37,31,203,31,189,31,227,31,247,31,89,31,120,31,120,30,224,31,235,31,180,31,180,30,68,31,41,31,252,31,218,31,7,31,154,31,144,31,47,31,106,31,228,31,50,31,253,31,87,31,45,31,148,31,131,31,137,31,169,31,169,30,142,31,148,31,238,31,224,31,245,31,77,31,77,30,4,31,126,31,55,31,247,31,247,30,226,31,110,31,10,31,124,31,15,31,202,31,230,31,142,31,82,31,128,31,128,30,195,31,195,30,31,31,129,31,34,31,34,30,216,31,216,30,40,31,226,31,225,31,72,31,72,30,238,31,167,31,167,30,93,31,66,31,117,31,58,31,139,31,139,30,197,31,158,31,206,31,148,31,204,31,200,31,200,30,200,29,117,31,100,31,216,31,189,31,233,31,112,31,128,31,158,31,47,31,231,31,193,31,28,31,166,31,182,31,182,30,68,31,89,31,207,31,207,30,207,29,168,31,138,31,94,31,94,30,205,31,205,30,164,31,49,31,182,31,3,31,57,31,57,30,49,31,232,31,232,30,232,29,111,31,244,31,112,31,209,31,85,31,7,31,238,31,65,31,65,30,216,31,216,30,30,31,82,31,50,31,12,31,42,31,25,31,25,30,25,29,7,31,102,31,46,31,128,31,128,30,128,29,205,31,247,31,11,31,181,31,181,30,126,31,155,31,156,31,244,31,174,31,149,31,56,31,111,31,141,31,89,31,238,31,30,31,251,31,186,31,129,31,252,31,29,31,155,31,65,31,181,31,49,31,58,31,227,31,227,30,61,31,27,31,27,30,1,31,155,31,144,31,192,31,6,31,6,30,203,31,26,31,26,30,208,31,20,31,176,31,245,31,13,31,160,31,160,30,84,31,71,31,71,30,71,29,71,28,237,31,87,31,87,30,123,31,123,30,213,31,213,30,225,31,72,31,123,31,197,31,1,31,212,31,14,31,134,31,74,31,140,31,168,31,168,30,209,31,62,31,62,30,127,31,95,31,10,31,181,31,235,31,26,31,93,31,93,30,228,31,228,30,131,31,131,30,18,31,5,31,5,30,171,31,208,31,143,31,131,31,135,31,192,31,192,30,192,29,61,31,205,31,117,31,141,31,141,30,103,31,18,31,18,30,18,29,175,31,175,30,175,29,129,31,193,31,195,31,195,30,168,31,193,31,230,31,144,31,194,31,13,31,95,31,98,31,53,31,53,30,111,31,207,31,157,31,157,30,22,31,85,31,187,31,67,31,176,31,16,31,16,30,136,31,138,31,79,31,79,30,2,31,2,30,240,31,3,31,62,31,156,31,98,31,183,31,131,31,131,31,155,31,149,31,168,31,22,31,27,31,17,31,187,31,92,31,199,31,199,30,230,31,133,31,79,31,228,31,62,31,62,30,62,29,18,31,43,31,43,30,166,31,193,31,193,30,193,29,219,31,66,31,207,31,255,31,187,31,219,31,27,31,56,31,146,31,151,31,235,31,207,31,207,30,161,31,76,31,76,31,76,30,76,29,50,31,200,31,212,31,221,31,184,31,181,31,85,31,157,31,226,31,76,31,68,31,77,31,153,31,254,31,254,30,254,29,160,31,90,31,109,31,231,31,140,31,19,31,19,30,19,29,155,31,138,31,143,31,209,31,230,31,230,30,231,31,159,31,111,31,116,31,81,31,21,31,42,31,218,31,40,31,14,31,4,31,4,30,149,31,229,31,230,31,139,31,16,31,93,31,93,30,126,31,230,31,37,31,37,30,37,29,37,28,96,31,96,30,96,29,40,31,182,31,30,31,30,30,7,31,121,31,148,31,205,31,205,30,80,31,80,30,18,31,195,31,103,31,221,31,122,31,58,31,58,30,230,31,180,31,180,31,104,31,245,31,40,31,117,31,89,31,68,31,190,31,138,31,244,31,115,31,243,31,173,31,132,31,132,30,197,31,8,31,8,30,97,31,189,31,18,31,172,31,108,31,189,31,178,31,178,30,133,31,133,30,133,29,103,31,200,31,89,31,89,30,135,31,239,31,239,30,239,29,217,31,226,31,228,31,179,31,222,31,222,30,222,29,65,31,11,31,173,31,173,30,16,31,138,31,8,31,73,31,73,30,130,31,158,31,176,31,124,31,75,31,12,31,103,31,85,31,61,31,70,31,7,31,140,31,63,31,214,31,221,31,228,31,125,31,125,30,154,31,154,30,50,31,50,30,204,31,110,31,157,31,10,31,53,31,192,31,80,31,210,31,43,31,107,31,107,30,131,31,103,31,159,31,123,31,128,31,128,30,3,31,191,31,129,31,161,31,252,31,139,31,97,31,97,30,97,29,5,31,5,30,73,31,1,31,98,31,15,31,213,31,247,31,78,31,140,31,162,31,55,31,6,31,165,31,169,31,239,31,239,30,244,31,244,30,116,31,171,31,28,31,20,31,188,31,202,31,202,30,32,31,14,31,116,31,208,31,242,31,116,31,120,31,168,31,168,30,168,29,168,28,128,31,130,31,107,31,1,31,148,31,172,31,172,30,145,31,5,31,204,31,90,31,90,30,94,31,187,31,111,31,16,31,59,31,155,31,75,31,108,31,65,31,244,31,136,31,70,31,45,31,114,31,41,31,199,31,29,31,193,31,193,30,164,31,87,31,210,31,90,31,115,31,115,30,224,31,2,31,134,31,74,31,73,31,73,30,10,31,10,30,10,29,47,31,47,30,198,31,21,31,21,30,134,31,37,31,70,31,204,31,107,31,231,31,151,31,12,31,12,30,186,31,195,31,162,31,240,31,97,31,139,31,71,31,200,31,200,30,200,29,117,31,29,31,29,30,165,31,138,31,130,31,130,30,130,29,130,28,164,31,158,31,158,30,158,29,202,31,120,31,197,31,185,31,193,31,193,30,117,31,117,30,117,29,72,31,25,31,231,31,231,30,133,31,91,31,36,31,96,31,191,31,212,31,78,31,135,31,92,31,92,30,213,31,223,31,7,31,235,31,235,30,128,31,128,30,66,31,66,30,150,31,89,31,136,31,199,31,127,31,191,31,191,30,191,29,39,31,191,31,191,30,11,31,233,31,43,31,206,31,140,31,224,31,11,31,224,31,166,31,241,31,183,31,95,31,196,31,98,31,35,31,133,31,42,31,101,31,118,31,249,31,70,31,173,31,173,30,135,31,135,30,189,31,85,31,180,31,10,31,153,31,127,31,127,30,78,31,135,31,135,30,172,31,172,30,172,29,104,31,104,30,15,31,15,30,70,31,70,30,70,29,201,31,182,31,28,31,28,30,148,31,103,31,103,30,30,31,88,31,23,31,23,30,45,31,62,31,17,31,99,31,99,30,99,29,99,28,104,31,210,31,210,30,83,31,83,30,235,31,62,31,3,31,251,31,172,31,235,31,36,31,77,31,27,31,30,31,111,31,49,31,70,31,191,31,15,31,197,31,144,31,156,31,107,31,181,31,82,31,134,31,134,30,253,31,221,31,84,31,10,31,153,31,179,31,250,31,250,30,66,31,27,31,229,31,25,31,108,31,108,30,22,31,143,31,16,31,66,31,66,30,66,29,155,31,155,30,179,31,210,31,58,31,85,31,85,30,85,29,177,31,10,31,229,31,229,30,240,31,249,31,6,31,129,31,39,31,52,31,143,31,226,31,227,31,142,31,123,31,192,31,49,31,104,31,16,31,16,30,16,29,16,28,16,27,127,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
