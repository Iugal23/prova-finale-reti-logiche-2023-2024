-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 864;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (29,0,85,0,0,0,54,0,86,0,178,0,221,0,232,0,19,0,93,0,215,0,170,0,220,0,53,0,81,0,0,0,192,0,0,0,0,0,172,0,26,0,229,0,0,0,0,0,150,0,238,0,156,0,118,0,13,0,202,0,94,0,115,0,192,0,48,0,138,0,23,0,224,0,164,0,194,0,114,0,0,0,34,0,139,0,241,0,215,0,38,0,103,0,226,0,36,0,26,0,113,0,240,0,245,0,144,0,52,0,145,0,246,0,94,0,44,0,247,0,0,0,0,0,182,0,10,0,215,0,105,0,123,0,90,0,191,0,238,0,198,0,147,0,54,0,0,0,83,0,234,0,0,0,215,0,138,0,0,0,0,0,191,0,141,0,142,0,73,0,95,0,0,0,109,0,141,0,248,0,91,0,216,0,0,0,15,0,222,0,204,0,45,0,92,0,16,0,29,0,177,0,18,0,0,0,0,0,24,0,122,0,228,0,173,0,95,0,0,0,82,0,69,0,29,0,133,0,89,0,0,0,193,0,213,0,226,0,0,0,249,0,222,0,107,0,98,0,134,0,5,0,246,0,66,0,96,0,250,0,216,0,233,0,190,0,5,0,239,0,0,0,149,0,205,0,177,0,71,0,111,0,0,0,134,0,24,0,121,0,160,0,231,0,0,0,195,0,235,0,214,0,183,0,190,0,250,0,74,0,174,0,60,0,0,0,225,0,147,0,108,0,250,0,238,0,0,0,0,0,192,0,51,0,0,0,175,0,237,0,96,0,179,0,219,0,198,0,226,0,184,0,41,0,43,0,137,0,160,0,95,0,232,0,211,0,233,0,118,0,215,0,80,0,0,0,0,0,14,0,182,0,55,0,247,0,136,0,113,0,95,0,0,0,64,0,130,0,110,0,192,0,216,0,85,0,209,0,113,0,203,0,188,0,191,0,104,0,0,0,0,0,255,0,86,0,0,0,0,0,121,0,150,0,37,0,55,0,88,0,81,0,93,0,29,0,108,0,61,0,141,0,97,0,90,0,0,0,95,0,51,0,24,0,225,0,68,0,0,0,7,0,11,0,66,0,168,0,30,0,0,0,165,0,62,0,77,0,74,0,0,0,82,0,179,0,195,0,254,0,120,0,200,0,253,0,0,0,34,0,0,0,104,0,171,0,143,0,162,0,0,0,180,0,195,0,66,0,182,0,252,0,186,0,137,0,116,0,71,0,119,0,138,0,242,0,99,0,0,0,200,0,65,0,181,0,182,0,0,0,216,0,0,0,127,0,0,0,39,0,217,0,0,0,48,0,0,0,171,0,3,0,0,0,19,0,57,0,48,0,202,0,0,0,194,0,185,0,0,0,233,0,8,0,128,0,0,0,0,0,21,0,231,0,1,0,149,0,183,0,192,0,0,0,0,0,93,0,10,0,252,0,91,0,114,0,91,0,0,0,214,0,214,0,107,0,176,0,60,0,13,0,175,0,157,0,235,0,49,0,254,0,0,0,132,0,0,0,114,0,98,0,171,0,105,0,0,0,118,0,69,0,0,0,220,0,176,0,101,0,37,0,242,0,120,0,197,0,59,0,61,0,46,0,79,0,0,0,206,0,112,0,0,0,161,0,222,0,156,0,0,0,254,0,209,0,30,0,0,0,167,0,110,0,97,0,128,0,73,0,0,0,151,0,147,0,204,0,217,0,159,0,227,0,50,0,16,0,121,0,9,0,0,0,208,0,114,0,135,0,194,0,169,0,62,0,187,0,227,0,78,0,151,0,239,0,96,0,213,0,191,0,21,0,127,0,9,0,183,0,121,0,0,0,98,0,0,0,254,0,64,0,187,0,71,0,215,0,217,0,53,0,58,0,67,0,86,0,207,0,0,0,0,0,240,0,0,0,0,0,0,0,0,0,0,0,205,0,0,0,160,0,105,0,109,0,35,0,0,0,81,0,28,0,0,0,176,0,147,0,33,0,56,0,140,0,24,0,208,0,252,0,241,0,176,0,0,0,215,0,226,0,150,0,185,0,153,0,227,0,178,0,0,0,205,0,0,0,0,0,243,0,112,0,0,0,212,0,80,0,181,0,0,0,115,0,222,0,211,0,200,0,206,0,9,0,18,0,251,0,97,0,0,0,170,0,0,0,232,0,17,0,19,0,1,0,221,0,0,0,170,0,24,0,0,0,82,0,40,0,92,0,147,0,43,0,80,0,0,0,183,0,191,0,0,0,250,0,221,0,127,0,0,0,149,0,182,0,17,0,181,0,22,0,0,0,0,0,101,0,254,0,168,0,144,0,102,0,245,0,181,0,131,0,0,0,87,0,75,0,97,0,42,0,211,0,220,0,55,0,53,0,44,0,173,0,0,0,216,0,0,0,172,0,241,0,202,0,0,0,189,0,0,0,62,0,228,0,179,0,195,0,174,0,78,0,0,0,40,0,50,0,0,0,243,0,120,0,95,0,0,0,213,0,38,0,139,0,131,0,213,0,146,0,33,0,105,0,0,0,176,0,105,0,81,0,31,0,227,0,93,0,155,0,12,0,132,0,0,0,1,0,93,0,0,0,144,0,0,0,159,0,253,0,126,0,108,0,188,0,151,0,93,0,0,0,50,0,251,0,99,0,105,0,246,0,10,0,44,0,149,0,9,0,247,0,153,0,27,0,128,0,20,0,78,0,7,0,221,0,209,0,168,0,0,0,66,0,0,0,207,0,220,0,113,0,227,0,114,0,73,0,62,0,208,0,0,0,0,0,72,0,207,0,239,0,253,0,16,0,152,0,20,0,185,0,202,0,193,0,195,0,0,0,0,0,89,0,156,0,138,0,206,0,89,0,12,0,10,0,99,0,201,0,201,0,208,0,220,0,215,0,101,0,102,0,94,0,151,0,57,0,88,0,214,0,21,0,2,0,156,0,253,0,169,0,67,0,55,0,0,0,16,0,0,0,188,0,252,0,242,0,50,0,231,0,0,0,0,0,90,0,0,0,177,0,0,0,201,0,0,0,6,0,38,0,145,0,174,0,0,0,228,0,57,0,28,0,233,0,168,0,102,0,246,0,217,0,0,0,59,0,25,0,226,0,189,0,194,0,229,0,184,0,0,0,238,0,63,0,55,0,99,0,130,0,0,0,0,0,0,0,113,0,246,0,193,0,100,0,228,0,0,0,198,0,40,0,236,0,0,0,7,0,177,0,200,0,252,0,31,0,204,0,12,0,120,0,0,0,17,0,101,0,0,0,124,0,62,0,11,0,236,0,16,0,72,0,104,0,0,0,14,0,244,0,138,0,0,0,197,0,115,0,22,0,42,0,116,0,0,0,126,0,187,0,218,0,3,0,37,0,0,0,215,0,147,0,96,0,254,0,107,0,238,0,188,0,220,0,161,0,118,0,133,0,71,0,237,0,239,0,91,0,188,0,153,0,0,0,141,0,228,0,19,0,103,0,230,0,37,0,96,0,134,0,194,0,252,0,80,0,184,0,162,0,227,0,142,0,0,0,0,0,120,0,10,0,238,0,25,0,139,0,212,0,176,0,86,0,116,0,243,0,0,0,0,0,40,0,0,0,0,0,0,0,248,0,217,0,36,0,118,0,0,0,64,0,13,0,0,0,216,0,17,0,163,0,60,0,39,0,0,0,135,0,197,0,0,0,21,0,89,0,0,0,195,0,92,0,178,0,196,0,240,0,178,0,49,0,122,0,167,0,45,0,0,0,0,0,210,0,196,0,241,0,80,0,167,0,0,0,49,0,196,0,147,0,0,0,150,0,68,0,13,0,122,0,37,0,27,0,116,0,187,0,212,0,247,0,1,0,62,0,216,0,208,0,0,0,190,0,56,0,64,0,0,0,68,0,220,0,58,0,0,0,56,0,11,0,0,0,0,0,210,0,56,0);
signal scenario_full  : scenario_type := (29,31,85,31,85,30,54,31,86,31,178,31,221,31,232,31,19,31,93,31,215,31,170,31,220,31,53,31,81,31,81,30,192,31,192,30,192,29,172,31,26,31,229,31,229,30,229,29,150,31,238,31,156,31,118,31,13,31,202,31,94,31,115,31,192,31,48,31,138,31,23,31,224,31,164,31,194,31,114,31,114,30,34,31,139,31,241,31,215,31,38,31,103,31,226,31,36,31,26,31,113,31,240,31,245,31,144,31,52,31,145,31,246,31,94,31,44,31,247,31,247,30,247,29,182,31,10,31,215,31,105,31,123,31,90,31,191,31,238,31,198,31,147,31,54,31,54,30,83,31,234,31,234,30,215,31,138,31,138,30,138,29,191,31,141,31,142,31,73,31,95,31,95,30,109,31,141,31,248,31,91,31,216,31,216,30,15,31,222,31,204,31,45,31,92,31,16,31,29,31,177,31,18,31,18,30,18,29,24,31,122,31,228,31,173,31,95,31,95,30,82,31,69,31,29,31,133,31,89,31,89,30,193,31,213,31,226,31,226,30,249,31,222,31,107,31,98,31,134,31,5,31,246,31,66,31,96,31,250,31,216,31,233,31,190,31,5,31,239,31,239,30,149,31,205,31,177,31,71,31,111,31,111,30,134,31,24,31,121,31,160,31,231,31,231,30,195,31,235,31,214,31,183,31,190,31,250,31,74,31,174,31,60,31,60,30,225,31,147,31,108,31,250,31,238,31,238,30,238,29,192,31,51,31,51,30,175,31,237,31,96,31,179,31,219,31,198,31,226,31,184,31,41,31,43,31,137,31,160,31,95,31,232,31,211,31,233,31,118,31,215,31,80,31,80,30,80,29,14,31,182,31,55,31,247,31,136,31,113,31,95,31,95,30,64,31,130,31,110,31,192,31,216,31,85,31,209,31,113,31,203,31,188,31,191,31,104,31,104,30,104,29,255,31,86,31,86,30,86,29,121,31,150,31,37,31,55,31,88,31,81,31,93,31,29,31,108,31,61,31,141,31,97,31,90,31,90,30,95,31,51,31,24,31,225,31,68,31,68,30,7,31,11,31,66,31,168,31,30,31,30,30,165,31,62,31,77,31,74,31,74,30,82,31,179,31,195,31,254,31,120,31,200,31,253,31,253,30,34,31,34,30,104,31,171,31,143,31,162,31,162,30,180,31,195,31,66,31,182,31,252,31,186,31,137,31,116,31,71,31,119,31,138,31,242,31,99,31,99,30,200,31,65,31,181,31,182,31,182,30,216,31,216,30,127,31,127,30,39,31,217,31,217,30,48,31,48,30,171,31,3,31,3,30,19,31,57,31,48,31,202,31,202,30,194,31,185,31,185,30,233,31,8,31,128,31,128,30,128,29,21,31,231,31,1,31,149,31,183,31,192,31,192,30,192,29,93,31,10,31,252,31,91,31,114,31,91,31,91,30,214,31,214,31,107,31,176,31,60,31,13,31,175,31,157,31,235,31,49,31,254,31,254,30,132,31,132,30,114,31,98,31,171,31,105,31,105,30,118,31,69,31,69,30,220,31,176,31,101,31,37,31,242,31,120,31,197,31,59,31,61,31,46,31,79,31,79,30,206,31,112,31,112,30,161,31,222,31,156,31,156,30,254,31,209,31,30,31,30,30,167,31,110,31,97,31,128,31,73,31,73,30,151,31,147,31,204,31,217,31,159,31,227,31,50,31,16,31,121,31,9,31,9,30,208,31,114,31,135,31,194,31,169,31,62,31,187,31,227,31,78,31,151,31,239,31,96,31,213,31,191,31,21,31,127,31,9,31,183,31,121,31,121,30,98,31,98,30,254,31,64,31,187,31,71,31,215,31,217,31,53,31,58,31,67,31,86,31,207,31,207,30,207,29,240,31,240,30,240,29,240,28,240,27,240,26,205,31,205,30,160,31,105,31,109,31,35,31,35,30,81,31,28,31,28,30,176,31,147,31,33,31,56,31,140,31,24,31,208,31,252,31,241,31,176,31,176,30,215,31,226,31,150,31,185,31,153,31,227,31,178,31,178,30,205,31,205,30,205,29,243,31,112,31,112,30,212,31,80,31,181,31,181,30,115,31,222,31,211,31,200,31,206,31,9,31,18,31,251,31,97,31,97,30,170,31,170,30,232,31,17,31,19,31,1,31,221,31,221,30,170,31,24,31,24,30,82,31,40,31,92,31,147,31,43,31,80,31,80,30,183,31,191,31,191,30,250,31,221,31,127,31,127,30,149,31,182,31,17,31,181,31,22,31,22,30,22,29,101,31,254,31,168,31,144,31,102,31,245,31,181,31,131,31,131,30,87,31,75,31,97,31,42,31,211,31,220,31,55,31,53,31,44,31,173,31,173,30,216,31,216,30,172,31,241,31,202,31,202,30,189,31,189,30,62,31,228,31,179,31,195,31,174,31,78,31,78,30,40,31,50,31,50,30,243,31,120,31,95,31,95,30,213,31,38,31,139,31,131,31,213,31,146,31,33,31,105,31,105,30,176,31,105,31,81,31,31,31,227,31,93,31,155,31,12,31,132,31,132,30,1,31,93,31,93,30,144,31,144,30,159,31,253,31,126,31,108,31,188,31,151,31,93,31,93,30,50,31,251,31,99,31,105,31,246,31,10,31,44,31,149,31,9,31,247,31,153,31,27,31,128,31,20,31,78,31,7,31,221,31,209,31,168,31,168,30,66,31,66,30,207,31,220,31,113,31,227,31,114,31,73,31,62,31,208,31,208,30,208,29,72,31,207,31,239,31,253,31,16,31,152,31,20,31,185,31,202,31,193,31,195,31,195,30,195,29,89,31,156,31,138,31,206,31,89,31,12,31,10,31,99,31,201,31,201,31,208,31,220,31,215,31,101,31,102,31,94,31,151,31,57,31,88,31,214,31,21,31,2,31,156,31,253,31,169,31,67,31,55,31,55,30,16,31,16,30,188,31,252,31,242,31,50,31,231,31,231,30,231,29,90,31,90,30,177,31,177,30,201,31,201,30,6,31,38,31,145,31,174,31,174,30,228,31,57,31,28,31,233,31,168,31,102,31,246,31,217,31,217,30,59,31,25,31,226,31,189,31,194,31,229,31,184,31,184,30,238,31,63,31,55,31,99,31,130,31,130,30,130,29,130,28,113,31,246,31,193,31,100,31,228,31,228,30,198,31,40,31,236,31,236,30,7,31,177,31,200,31,252,31,31,31,204,31,12,31,120,31,120,30,17,31,101,31,101,30,124,31,62,31,11,31,236,31,16,31,72,31,104,31,104,30,14,31,244,31,138,31,138,30,197,31,115,31,22,31,42,31,116,31,116,30,126,31,187,31,218,31,3,31,37,31,37,30,215,31,147,31,96,31,254,31,107,31,238,31,188,31,220,31,161,31,118,31,133,31,71,31,237,31,239,31,91,31,188,31,153,31,153,30,141,31,228,31,19,31,103,31,230,31,37,31,96,31,134,31,194,31,252,31,80,31,184,31,162,31,227,31,142,31,142,30,142,29,120,31,10,31,238,31,25,31,139,31,212,31,176,31,86,31,116,31,243,31,243,30,243,29,40,31,40,30,40,29,40,28,248,31,217,31,36,31,118,31,118,30,64,31,13,31,13,30,216,31,17,31,163,31,60,31,39,31,39,30,135,31,197,31,197,30,21,31,89,31,89,30,195,31,92,31,178,31,196,31,240,31,178,31,49,31,122,31,167,31,45,31,45,30,45,29,210,31,196,31,241,31,80,31,167,31,167,30,49,31,196,31,147,31,147,30,150,31,68,31,13,31,122,31,37,31,27,31,116,31,187,31,212,31,247,31,1,31,62,31,216,31,208,31,208,30,190,31,56,31,64,31,64,30,68,31,220,31,58,31,58,30,56,31,11,31,11,30,11,29,210,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
