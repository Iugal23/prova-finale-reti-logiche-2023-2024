-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 992;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (94,0,30,0,169,0,181,0,0,0,106,0,255,0,55,0,0,0,221,0,0,0,233,0,69,0,21,0,89,0,0,0,130,0,21,0,30,0,46,0,170,0,153,0,0,0,94,0,39,0,150,0,144,0,98,0,172,0,26,0,112,0,239,0,81,0,0,0,0,0,152,0,205,0,33,0,64,0,92,0,8,0,61,0,3,0,0,0,111,0,7,0,184,0,177,0,183,0,49,0,190,0,86,0,134,0,85,0,111,0,209,0,83,0,111,0,236,0,161,0,204,0,155,0,33,0,159,0,234,0,229,0,151,0,207,0,208,0,0,0,0,0,9,0,39,0,137,0,218,0,85,0,130,0,149,0,81,0,17,0,90,0,0,0,82,0,202,0,158,0,228,0,155,0,0,0,0,0,0,0,216,0,36,0,137,0,59,0,0,0,3,0,122,0,179,0,0,0,87,0,109,0,169,0,239,0,187,0,0,0,46,0,179,0,0,0,73,0,0,0,169,0,255,0,77,0,157,0,74,0,0,0,49,0,192,0,0,0,39,0,202,0,0,0,115,0,33,0,0,0,56,0,16,0,204,0,0,0,94,0,209,0,0,0,206,0,55,0,175,0,85,0,178,0,214,0,227,0,46,0,81,0,168,0,84,0,70,0,248,0,0,0,119,0,216,0,0,0,235,0,107,0,86,0,81,0,0,0,210,0,173,0,14,0,144,0,168,0,36,0,118,0,0,0,154,0,31,0,240,0,80,0,30,0,146,0,84,0,214,0,63,0,0,0,205,0,0,0,0,0,0,0,0,0,76,0,0,0,0,0,88,0,205,0,89,0,0,0,26,0,114,0,71,0,30,0,95,0,77,0,89,0,0,0,180,0,138,0,80,0,176,0,240,0,47,0,6,0,205,0,190,0,0,0,0,0,111,0,0,0,93,0,235,0,254,0,175,0,0,0,77,0,31,0,86,0,131,0,0,0,21,0,237,0,247,0,197,0,127,0,43,0,176,0,240,0,232,0,0,0,142,0,118,0,151,0,173,0,0,0,176,0,0,0,136,0,5,0,229,0,80,0,156,0,14,0,241,0,175,0,243,0,37,0,137,0,170,0,201,0,110,0,251,0,75,0,72,0,145,0,187,0,118,0,0,0,167,0,152,0,0,0,20,0,6,0,0,0,136,0,223,0,65,0,75,0,67,0,196,0,118,0,96,0,0,0,115,0,180,0,239,0,0,0,193,0,0,0,238,0,113,0,75,0,214,0,193,0,0,0,141,0,0,0,0,0,0,0,143,0,54,0,75,0,174,0,202,0,34,0,0,0,154,0,22,0,71,0,76,0,113,0,0,0,90,0,128,0,49,0,0,0,87,0,226,0,89,0,0,0,0,0,182,0,87,0,171,0,36,0,110,0,198,0,135,0,143,0,12,0,80,0,103,0,240,0,140,0,0,0,227,0,248,0,1,0,227,0,0,0,187,0,52,0,32,0,108,0,63,0,189,0,68,0,221,0,126,0,0,0,74,0,138,0,0,0,191,0,251,0,0,0,234,0,223,0,0,0,25,0,194,0,0,0,80,0,4,0,0,0,219,0,235,0,189,0,121,0,17,0,63,0,189,0,11,0,43,0,144,0,33,0,0,0,32,0,123,0,24,0,129,0,111,0,116,0,103,0,72,0,28,0,124,0,1,0,192,0,0,0,253,0,0,0,20,0,95,0,187,0,192,0,68,0,218,0,107,0,107,0,138,0,2,0,63,0,59,0,0,0,157,0,22,0,105,0,7,0,191,0,209,0,57,0,140,0,0,0,0,0,22,0,209,0,0,0,114,0,0,0,0,0,204,0,247,0,81,0,77,0,189,0,124,0,215,0,179,0,10,0,113,0,15,0,78,0,32,0,101,0,133,0,0,0,24,0,237,0,99,0,35,0,53,0,18,0,62,0,157,0,66,0,96,0,0,0,83,0,37,0,0,0,183,0,22,0,0,0,181,0,0,0,196,0,91,0,17,0,64,0,0,0,0,0,213,0,0,0,231,0,13,0,160,0,77,0,0,0,78,0,0,0,79,0,0,0,124,0,0,0,68,0,5,0,0,0,140,0,230,0,0,0,221,0,98,0,150,0,230,0,35,0,147,0,12,0,192,0,155,0,227,0,0,0,27,0,229,0,129,0,137,0,113,0,8,0,0,0,75,0,161,0,56,0,2,0,47,0,194,0,0,0,108,0,209,0,232,0,0,0,186,0,0,0,0,0,125,0,62,0,117,0,228,0,0,0,0,0,55,0,142,0,89,0,234,0,194,0,100,0,5,0,220,0,240,0,112,0,0,0,237,0,0,0,0,0,185,0,0,0,0,0,195,0,116,0,107,0,220,0,44,0,74,0,181,0,221,0,0,0,0,0,211,0,228,0,254,0,224,0,235,0,195,0,38,0,27,0,159,0,202,0,151,0,24,0,66,0,85,0,109,0,103,0,106,0,76,0,32,0,2,0,191,0,121,0,143,0,154,0,246,0,226,0,19,0,12,0,0,0,21,0,124,0,156,0,4,0,150,0,129,0,232,0,69,0,8,0,53,0,119,0,198,0,58,0,188,0,115,0,222,0,160,0,57,0,18,0,40,0,0,0,0,0,154,0,20,0,147,0,6,0,91,0,80,0,115,0,0,0,115,0,146,0,0,0,232,0,213,0,85,0,48,0,53,0,210,0,68,0,110,0,99,0,207,0,14,0,157,0,12,0,174,0,0,0,76,0,123,0,182,0,16,0,19,0,167,0,43,0,0,0,152,0,27,0,196,0,122,0,0,0,0,0,121,0,0,0,229,0,73,0,26,0,130,0,185,0,0,0,0,0,97,0,108,0,0,0,0,0,0,0,0,0,235,0,166,0,32,0,0,0,0,0,11,0,242,0,0,0,77,0,41,0,170,0,0,0,163,0,175,0,114,0,132,0,197,0,0,0,94,0,26,0,107,0,0,0,74,0,102,0,49,0,48,0,231,0,0,0,2,0,0,0,97,0,84,0,229,0,147,0,50,0,0,0,73,0,222,0,116,0,87,0,9,0,111,0,4,0,85,0,26,0,250,0,0,0,68,0,154,0,246,0,0,0,43,0,175,0,242,0,116,0,238,0,32,0,57,0,118,0,0,0,10,0,215,0,0,0,0,0,60,0,189,0,68,0,5,0,20,0,0,0,208,0,57,0,108,0,42,0,181,0,3,0,188,0,150,0,150,0,181,0,171,0,226,0,0,0,67,0,218,0,223,0,173,0,97,0,0,0,150,0,115,0,45,0,151,0,41,0,64,0,127,0,1,0,85,0,0,0,0,0,115,0,7,0,47,0,23,0,71,0,9,0,59,0,0,0,190,0,243,0,126,0,105,0,110,0,192,0,0,0,195,0,197,0,181,0,217,0,216,0,97,0,78,0,83,0,83,0,205,0,67,0,192,0,10,0,13,0,0,0,0,0,0,0,144,0,232,0,72,0,62,0,228,0,26,0,230,0,0,0,90,0,184,0,0,0,188,0,27,0,46,0,0,0,204,0,224,0,0,0,107,0,240,0,48,0,119,0,125,0,30,0,158,0,223,0,3,0,90,0,70,0,92,0,117,0,26,0,18,0,0,0,158,0,74,0,0,0,15,0,16,0,0,0,44,0,216,0,0,0,171,0,218,0,0,0,164,0,177,0,79,0,132,0,107,0,202,0,12,0,0,0,20,0,93,0,187,0,30,0,252,0,254,0,0,0,107,0,38,0,249,0,164,0,149,0,0,0,4,0,198,0,119,0,27,0,192,0,237,0,71,0,0,0,240,0,38,0,178,0,2,0,170,0,0,0,174,0,168,0,0,0,6,0,93,0,90,0,0,0,41,0,7,0,218,0,0,0,248,0,121,0,214,0,22,0,204,0,66,0,0,0,143,0,153,0,0,0,167,0,0,0,157,0,19,0,0,0,153,0,0,0,113,0,40,0,194,0,0,0,71,0,11,0,10,0,212,0,0,0,228,0,120,0,30,0,0,0,0,0,147,0,145,0,68,0,217,0,89,0,0,0,241,0,0,0,0,0,187,0,22,0,144,0,192,0,0,0,173,0,134,0,25,0,141,0,192,0,0,0,239,0,192,0,237,0,91,0,26,0,23,0,97,0,63,0,180,0,55,0,165,0,131,0,208,0,0,0,0,0,155,0,26,0,117,0,53,0,114,0,164,0,0,0,7,0,19,0,76,0,114,0,178,0,119,0,141,0,8,0,201,0,0,0,189,0,0,0,84,0,100,0,0,0,229,0,165,0,109,0,0,0,79,0,0,0,0,0,98,0,174,0,109,0,132,0,0,0,207,0,72,0,18,0,196,0,55,0,0,0,172,0,219,0,0,0,68,0,0,0,50,0,88,0,9,0,221,0,61,0,0,0,28,0,111,0,9,0,42,0,24,0,202,0,239,0,0,0,0,0,255,0,109,0,173,0,217,0,0,0);
signal scenario_full  : scenario_type := (94,31,30,31,169,31,181,31,181,30,106,31,255,31,55,31,55,30,221,31,221,30,233,31,69,31,21,31,89,31,89,30,130,31,21,31,30,31,46,31,170,31,153,31,153,30,94,31,39,31,150,31,144,31,98,31,172,31,26,31,112,31,239,31,81,31,81,30,81,29,152,31,205,31,33,31,64,31,92,31,8,31,61,31,3,31,3,30,111,31,7,31,184,31,177,31,183,31,49,31,190,31,86,31,134,31,85,31,111,31,209,31,83,31,111,31,236,31,161,31,204,31,155,31,33,31,159,31,234,31,229,31,151,31,207,31,208,31,208,30,208,29,9,31,39,31,137,31,218,31,85,31,130,31,149,31,81,31,17,31,90,31,90,30,82,31,202,31,158,31,228,31,155,31,155,30,155,29,155,28,216,31,36,31,137,31,59,31,59,30,3,31,122,31,179,31,179,30,87,31,109,31,169,31,239,31,187,31,187,30,46,31,179,31,179,30,73,31,73,30,169,31,255,31,77,31,157,31,74,31,74,30,49,31,192,31,192,30,39,31,202,31,202,30,115,31,33,31,33,30,56,31,16,31,204,31,204,30,94,31,209,31,209,30,206,31,55,31,175,31,85,31,178,31,214,31,227,31,46,31,81,31,168,31,84,31,70,31,248,31,248,30,119,31,216,31,216,30,235,31,107,31,86,31,81,31,81,30,210,31,173,31,14,31,144,31,168,31,36,31,118,31,118,30,154,31,31,31,240,31,80,31,30,31,146,31,84,31,214,31,63,31,63,30,205,31,205,30,205,29,205,28,205,27,76,31,76,30,76,29,88,31,205,31,89,31,89,30,26,31,114,31,71,31,30,31,95,31,77,31,89,31,89,30,180,31,138,31,80,31,176,31,240,31,47,31,6,31,205,31,190,31,190,30,190,29,111,31,111,30,93,31,235,31,254,31,175,31,175,30,77,31,31,31,86,31,131,31,131,30,21,31,237,31,247,31,197,31,127,31,43,31,176,31,240,31,232,31,232,30,142,31,118,31,151,31,173,31,173,30,176,31,176,30,136,31,5,31,229,31,80,31,156,31,14,31,241,31,175,31,243,31,37,31,137,31,170,31,201,31,110,31,251,31,75,31,72,31,145,31,187,31,118,31,118,30,167,31,152,31,152,30,20,31,6,31,6,30,136,31,223,31,65,31,75,31,67,31,196,31,118,31,96,31,96,30,115,31,180,31,239,31,239,30,193,31,193,30,238,31,113,31,75,31,214,31,193,31,193,30,141,31,141,30,141,29,141,28,143,31,54,31,75,31,174,31,202,31,34,31,34,30,154,31,22,31,71,31,76,31,113,31,113,30,90,31,128,31,49,31,49,30,87,31,226,31,89,31,89,30,89,29,182,31,87,31,171,31,36,31,110,31,198,31,135,31,143,31,12,31,80,31,103,31,240,31,140,31,140,30,227,31,248,31,1,31,227,31,227,30,187,31,52,31,32,31,108,31,63,31,189,31,68,31,221,31,126,31,126,30,74,31,138,31,138,30,191,31,251,31,251,30,234,31,223,31,223,30,25,31,194,31,194,30,80,31,4,31,4,30,219,31,235,31,189,31,121,31,17,31,63,31,189,31,11,31,43,31,144,31,33,31,33,30,32,31,123,31,24,31,129,31,111,31,116,31,103,31,72,31,28,31,124,31,1,31,192,31,192,30,253,31,253,30,20,31,95,31,187,31,192,31,68,31,218,31,107,31,107,31,138,31,2,31,63,31,59,31,59,30,157,31,22,31,105,31,7,31,191,31,209,31,57,31,140,31,140,30,140,29,22,31,209,31,209,30,114,31,114,30,114,29,204,31,247,31,81,31,77,31,189,31,124,31,215,31,179,31,10,31,113,31,15,31,78,31,32,31,101,31,133,31,133,30,24,31,237,31,99,31,35,31,53,31,18,31,62,31,157,31,66,31,96,31,96,30,83,31,37,31,37,30,183,31,22,31,22,30,181,31,181,30,196,31,91,31,17,31,64,31,64,30,64,29,213,31,213,30,231,31,13,31,160,31,77,31,77,30,78,31,78,30,79,31,79,30,124,31,124,30,68,31,5,31,5,30,140,31,230,31,230,30,221,31,98,31,150,31,230,31,35,31,147,31,12,31,192,31,155,31,227,31,227,30,27,31,229,31,129,31,137,31,113,31,8,31,8,30,75,31,161,31,56,31,2,31,47,31,194,31,194,30,108,31,209,31,232,31,232,30,186,31,186,30,186,29,125,31,62,31,117,31,228,31,228,30,228,29,55,31,142,31,89,31,234,31,194,31,100,31,5,31,220,31,240,31,112,31,112,30,237,31,237,30,237,29,185,31,185,30,185,29,195,31,116,31,107,31,220,31,44,31,74,31,181,31,221,31,221,30,221,29,211,31,228,31,254,31,224,31,235,31,195,31,38,31,27,31,159,31,202,31,151,31,24,31,66,31,85,31,109,31,103,31,106,31,76,31,32,31,2,31,191,31,121,31,143,31,154,31,246,31,226,31,19,31,12,31,12,30,21,31,124,31,156,31,4,31,150,31,129,31,232,31,69,31,8,31,53,31,119,31,198,31,58,31,188,31,115,31,222,31,160,31,57,31,18,31,40,31,40,30,40,29,154,31,20,31,147,31,6,31,91,31,80,31,115,31,115,30,115,31,146,31,146,30,232,31,213,31,85,31,48,31,53,31,210,31,68,31,110,31,99,31,207,31,14,31,157,31,12,31,174,31,174,30,76,31,123,31,182,31,16,31,19,31,167,31,43,31,43,30,152,31,27,31,196,31,122,31,122,30,122,29,121,31,121,30,229,31,73,31,26,31,130,31,185,31,185,30,185,29,97,31,108,31,108,30,108,29,108,28,108,27,235,31,166,31,32,31,32,30,32,29,11,31,242,31,242,30,77,31,41,31,170,31,170,30,163,31,175,31,114,31,132,31,197,31,197,30,94,31,26,31,107,31,107,30,74,31,102,31,49,31,48,31,231,31,231,30,2,31,2,30,97,31,84,31,229,31,147,31,50,31,50,30,73,31,222,31,116,31,87,31,9,31,111,31,4,31,85,31,26,31,250,31,250,30,68,31,154,31,246,31,246,30,43,31,175,31,242,31,116,31,238,31,32,31,57,31,118,31,118,30,10,31,215,31,215,30,215,29,60,31,189,31,68,31,5,31,20,31,20,30,208,31,57,31,108,31,42,31,181,31,3,31,188,31,150,31,150,31,181,31,171,31,226,31,226,30,67,31,218,31,223,31,173,31,97,31,97,30,150,31,115,31,45,31,151,31,41,31,64,31,127,31,1,31,85,31,85,30,85,29,115,31,7,31,47,31,23,31,71,31,9,31,59,31,59,30,190,31,243,31,126,31,105,31,110,31,192,31,192,30,195,31,197,31,181,31,217,31,216,31,97,31,78,31,83,31,83,31,205,31,67,31,192,31,10,31,13,31,13,30,13,29,13,28,144,31,232,31,72,31,62,31,228,31,26,31,230,31,230,30,90,31,184,31,184,30,188,31,27,31,46,31,46,30,204,31,224,31,224,30,107,31,240,31,48,31,119,31,125,31,30,31,158,31,223,31,3,31,90,31,70,31,92,31,117,31,26,31,18,31,18,30,158,31,74,31,74,30,15,31,16,31,16,30,44,31,216,31,216,30,171,31,218,31,218,30,164,31,177,31,79,31,132,31,107,31,202,31,12,31,12,30,20,31,93,31,187,31,30,31,252,31,254,31,254,30,107,31,38,31,249,31,164,31,149,31,149,30,4,31,198,31,119,31,27,31,192,31,237,31,71,31,71,30,240,31,38,31,178,31,2,31,170,31,170,30,174,31,168,31,168,30,6,31,93,31,90,31,90,30,41,31,7,31,218,31,218,30,248,31,121,31,214,31,22,31,204,31,66,31,66,30,143,31,153,31,153,30,167,31,167,30,157,31,19,31,19,30,153,31,153,30,113,31,40,31,194,31,194,30,71,31,11,31,10,31,212,31,212,30,228,31,120,31,30,31,30,30,30,29,147,31,145,31,68,31,217,31,89,31,89,30,241,31,241,30,241,29,187,31,22,31,144,31,192,31,192,30,173,31,134,31,25,31,141,31,192,31,192,30,239,31,192,31,237,31,91,31,26,31,23,31,97,31,63,31,180,31,55,31,165,31,131,31,208,31,208,30,208,29,155,31,26,31,117,31,53,31,114,31,164,31,164,30,7,31,19,31,76,31,114,31,178,31,119,31,141,31,8,31,201,31,201,30,189,31,189,30,84,31,100,31,100,30,229,31,165,31,109,31,109,30,79,31,79,30,79,29,98,31,174,31,109,31,132,31,132,30,207,31,72,31,18,31,196,31,55,31,55,30,172,31,219,31,219,30,68,31,68,30,50,31,88,31,9,31,221,31,61,31,61,30,28,31,111,31,9,31,42,31,24,31,202,31,239,31,239,30,239,29,255,31,109,31,173,31,217,31,217,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
