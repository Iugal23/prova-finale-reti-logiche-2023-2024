-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_812 is
end project_tb_812;

architecture project_tb_arch_812 of project_tb_812 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 607;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,198,0,154,0,0,0,36,0,36,0,170,0,30,0,0,0,142,0,234,0,157,0,158,0,10,0,123,0,227,0,181,0,220,0,140,0,209,0,0,0,0,0,42,0,57,0,249,0,0,0,0,0,0,0,39,0,65,0,76,0,217,0,0,0,173,0,0,0,135,0,0,0,0,0,188,0,209,0,142,0,242,0,202,0,0,0,14,0,235,0,141,0,0,0,181,0,0,0,89,0,53,0,132,0,196,0,46,0,0,0,94,0,0,0,102,0,5,0,129,0,171,0,25,0,151,0,165,0,34,0,64,0,0,0,11,0,17,0,207,0,0,0,43,0,183,0,89,0,198,0,186,0,116,0,235,0,44,0,72,0,0,0,165,0,71,0,87,0,253,0,0,0,83,0,127,0,57,0,205,0,25,0,95,0,192,0,159,0,197,0,0,0,157,0,47,0,84,0,153,0,91,0,9,0,214,0,89,0,108,0,0,0,197,0,50,0,50,0,81,0,146,0,248,0,0,0,92,0,118,0,79,0,106,0,38,0,184,0,0,0,24,0,0,0,102,0,74,0,35,0,254,0,200,0,66,0,190,0,0,0,27,0,170,0,50,0,0,0,175,0,0,0,238,0,0,0,150,0,184,0,14,0,0,0,73,0,239,0,232,0,0,0,67,0,90,0,186,0,0,0,0,0,0,0,59,0,98,0,129,0,114,0,62,0,133,0,146,0,151,0,100,0,0,0,0,0,41,0,0,0,85,0,0,0,0,0,208,0,0,0,98,0,199,0,0,0,103,0,38,0,0,0,199,0,252,0,78,0,104,0,194,0,100,0,0,0,188,0,187,0,93,0,255,0,0,0,50,0,208,0,77,0,4,0,173,0,205,0,140,0,131,0,209,0,0,0,226,0,30,0,91,0,188,0,229,0,0,0,0,0,190,0,126,0,0,0,4,0,125,0,0,0,0,0,86,0,108,0,197,0,0,0,210,0,0,0,0,0,135,0,0,0,0,0,136,0,16,0,77,0,143,0,0,0,196,0,0,0,0,0,0,0,0,0,237,0,180,0,223,0,131,0,0,0,205,0,0,0,114,0,0,0,147,0,125,0,217,0,0,0,167,0,0,0,142,0,100,0,2,0,162,0,0,0,47,0,237,0,9,0,30,0,0,0,52,0,195,0,0,0,127,0,153,0,159,0,224,0,0,0,130,0,0,0,0,0,0,0,0,0,0,0,207,0,0,0,118,0,78,0,30,0,175,0,161,0,122,0,7,0,0,0,17,0,0,0,255,0,0,0,72,0,232,0,178,0,155,0,116,0,0,0,0,0,0,0,47,0,152,0,202,0,147,0,0,0,0,0,67,0,179,0,47,0,97,0,231,0,0,0,53,0,0,0,15,0,0,0,42,0,9,0,0,0,60,0,0,0,200,0,0,0,229,0,15,0,229,0,0,0,76,0,184,0,11,0,144,0,0,0,130,0,0,0,196,0,0,0,0,0,128,0,205,0,188,0,199,0,95,0,49,0,198,0,0,0,71,0,150,0,0,0,206,0,132,0,79,0,185,0,17,0,4,0,1,0,6,0,13,0,114,0,0,0,0,0,44,0,166,0,0,0,2,0,157,0,40,0,135,0,47,0,28,0,53,0,0,0,121,0,178,0,227,0,228,0,131,0,20,0,219,0,32,0,207,0,29,0,108,0,0,0,88,0,0,0,165,0,0,0,0,0,31,0,51,0,238,0,11,0,210,0,0,0,0,0,18,0,64,0,255,0,88,0,33,0,177,0,100,0,63,0,156,0,246,0,119,0,0,0,101,0,28,0,163,0,48,0,250,0,214,0,240,0,6,0,116,0,211,0,52,0,0,0,249,0,75,0,0,0,25,0,0,0,14,0,25,0,0,0,0,0,0,0,64,0,65,0,179,0,101,0,67,0,0,0,0,0,0,0,158,0,9,0,148,0,0,0,42,0,96,0,154,0,34,0,234,0,148,0,122,0,206,0,212,0,18,0,167,0,206,0,184,0,0,0,0,0,0,0,121,0,230,0,47,0,0,0,108,0,73,0,3,0,0,0,133,0,0,0,83,0,0,0,0,0,105,0,240,0,198,0,178,0,70,0,222,0,49,0,104,0,85,0,17,0,83,0,0,0,71,0,249,0,167,0,133,0,0,0,242,0,131,0,23,0,180,0,109,0,161,0,93,0,122,0,201,0,95,0,144,0,161,0,46,0,222,0,36,0,170,0,111,0,0,0,113,0,131,0,35,0,46,0,119,0,0,0,255,0,0,0,220,0,243,0,0,0,68,0,33,0,72,0,192,0,0,0,79,0,29,0,62,0,50,0,89,0,133,0,0,0,45,0,252,0,0,0,131,0,154,0,248,0,165,0,0,0,161,0,60,0,0,0,0,0,3,0,148,0,166,0,0,0,0,0,197,0,0,0,0,0,218,0,216,0,0,0,0,0,0,0,122,0,3,0,0,0,0,0,0,0,191,0,188,0,169,0,227,0,0,0,248,0,200,0,134,0,99,0,52,0,191,0,88,0,10,0,0,0,63,0,201,0,0,0,54,0,114,0,152,0,14,0,37,0,228,0,0,0,254,0,0,0,0,0,231,0,229,0,205,0,14,0,73,0,42,0,0,0,0,0,204,0,196,0,91,0,0,0,59,0,126,0,69,0,102,0,1,0,77,0,47,0,0,0,166,0,0,0,81,0,215,0,83,0,194,0,8,0,224,0);
signal scenario_full  : scenario_type := (0,0,198,31,154,31,154,30,36,31,36,31,170,31,30,31,30,30,142,31,234,31,157,31,158,31,10,31,123,31,227,31,181,31,220,31,140,31,209,31,209,30,209,29,42,31,57,31,249,31,249,30,249,29,249,28,39,31,65,31,76,31,217,31,217,30,173,31,173,30,135,31,135,30,135,29,188,31,209,31,142,31,242,31,202,31,202,30,14,31,235,31,141,31,141,30,181,31,181,30,89,31,53,31,132,31,196,31,46,31,46,30,94,31,94,30,102,31,5,31,129,31,171,31,25,31,151,31,165,31,34,31,64,31,64,30,11,31,17,31,207,31,207,30,43,31,183,31,89,31,198,31,186,31,116,31,235,31,44,31,72,31,72,30,165,31,71,31,87,31,253,31,253,30,83,31,127,31,57,31,205,31,25,31,95,31,192,31,159,31,197,31,197,30,157,31,47,31,84,31,153,31,91,31,9,31,214,31,89,31,108,31,108,30,197,31,50,31,50,31,81,31,146,31,248,31,248,30,92,31,118,31,79,31,106,31,38,31,184,31,184,30,24,31,24,30,102,31,74,31,35,31,254,31,200,31,66,31,190,31,190,30,27,31,170,31,50,31,50,30,175,31,175,30,238,31,238,30,150,31,184,31,14,31,14,30,73,31,239,31,232,31,232,30,67,31,90,31,186,31,186,30,186,29,186,28,59,31,98,31,129,31,114,31,62,31,133,31,146,31,151,31,100,31,100,30,100,29,41,31,41,30,85,31,85,30,85,29,208,31,208,30,98,31,199,31,199,30,103,31,38,31,38,30,199,31,252,31,78,31,104,31,194,31,100,31,100,30,188,31,187,31,93,31,255,31,255,30,50,31,208,31,77,31,4,31,173,31,205,31,140,31,131,31,209,31,209,30,226,31,30,31,91,31,188,31,229,31,229,30,229,29,190,31,126,31,126,30,4,31,125,31,125,30,125,29,86,31,108,31,197,31,197,30,210,31,210,30,210,29,135,31,135,30,135,29,136,31,16,31,77,31,143,31,143,30,196,31,196,30,196,29,196,28,196,27,237,31,180,31,223,31,131,31,131,30,205,31,205,30,114,31,114,30,147,31,125,31,217,31,217,30,167,31,167,30,142,31,100,31,2,31,162,31,162,30,47,31,237,31,9,31,30,31,30,30,52,31,195,31,195,30,127,31,153,31,159,31,224,31,224,30,130,31,130,30,130,29,130,28,130,27,130,26,207,31,207,30,118,31,78,31,30,31,175,31,161,31,122,31,7,31,7,30,17,31,17,30,255,31,255,30,72,31,232,31,178,31,155,31,116,31,116,30,116,29,116,28,47,31,152,31,202,31,147,31,147,30,147,29,67,31,179,31,47,31,97,31,231,31,231,30,53,31,53,30,15,31,15,30,42,31,9,31,9,30,60,31,60,30,200,31,200,30,229,31,15,31,229,31,229,30,76,31,184,31,11,31,144,31,144,30,130,31,130,30,196,31,196,30,196,29,128,31,205,31,188,31,199,31,95,31,49,31,198,31,198,30,71,31,150,31,150,30,206,31,132,31,79,31,185,31,17,31,4,31,1,31,6,31,13,31,114,31,114,30,114,29,44,31,166,31,166,30,2,31,157,31,40,31,135,31,47,31,28,31,53,31,53,30,121,31,178,31,227,31,228,31,131,31,20,31,219,31,32,31,207,31,29,31,108,31,108,30,88,31,88,30,165,31,165,30,165,29,31,31,51,31,238,31,11,31,210,31,210,30,210,29,18,31,64,31,255,31,88,31,33,31,177,31,100,31,63,31,156,31,246,31,119,31,119,30,101,31,28,31,163,31,48,31,250,31,214,31,240,31,6,31,116,31,211,31,52,31,52,30,249,31,75,31,75,30,25,31,25,30,14,31,25,31,25,30,25,29,25,28,64,31,65,31,179,31,101,31,67,31,67,30,67,29,67,28,158,31,9,31,148,31,148,30,42,31,96,31,154,31,34,31,234,31,148,31,122,31,206,31,212,31,18,31,167,31,206,31,184,31,184,30,184,29,184,28,121,31,230,31,47,31,47,30,108,31,73,31,3,31,3,30,133,31,133,30,83,31,83,30,83,29,105,31,240,31,198,31,178,31,70,31,222,31,49,31,104,31,85,31,17,31,83,31,83,30,71,31,249,31,167,31,133,31,133,30,242,31,131,31,23,31,180,31,109,31,161,31,93,31,122,31,201,31,95,31,144,31,161,31,46,31,222,31,36,31,170,31,111,31,111,30,113,31,131,31,35,31,46,31,119,31,119,30,255,31,255,30,220,31,243,31,243,30,68,31,33,31,72,31,192,31,192,30,79,31,29,31,62,31,50,31,89,31,133,31,133,30,45,31,252,31,252,30,131,31,154,31,248,31,165,31,165,30,161,31,60,31,60,30,60,29,3,31,148,31,166,31,166,30,166,29,197,31,197,30,197,29,218,31,216,31,216,30,216,29,216,28,122,31,3,31,3,30,3,29,3,28,191,31,188,31,169,31,227,31,227,30,248,31,200,31,134,31,99,31,52,31,191,31,88,31,10,31,10,30,63,31,201,31,201,30,54,31,114,31,152,31,14,31,37,31,228,31,228,30,254,31,254,30,254,29,231,31,229,31,205,31,14,31,73,31,42,31,42,30,42,29,204,31,196,31,91,31,91,30,59,31,126,31,69,31,102,31,1,31,77,31,47,31,47,30,166,31,166,30,81,31,215,31,83,31,194,31,8,31,224,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
