-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_679 is
end project_tb_679;

architecture project_tb_arch_679 of project_tb_679 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 873;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,162,0,146,0,248,0,19,0,0,0,132,0,170,0,180,0,224,0,0,0,66,0,185,0,97,0,162,0,138,0,34,0,133,0,0,0,175,0,97,0,15,0,0,0,41,0,19,0,42,0,95,0,175,0,148,0,241,0,220,0,0,0,102,0,91,0,0,0,252,0,183,0,174,0,37,0,0,0,251,0,121,0,230,0,0,0,196,0,214,0,11,0,182,0,0,0,138,0,186,0,0,0,0,0,97,0,0,0,146,0,163,0,154,0,134,0,36,0,104,0,50,0,111,0,0,0,177,0,238,0,0,0,156,0,0,0,59,0,138,0,60,0,0,0,0,0,59,0,0,0,57,0,124,0,123,0,92,0,137,0,0,0,132,0,20,0,85,0,123,0,0,0,0,0,12,0,63,0,144,0,154,0,134,0,206,0,0,0,0,0,0,0,0,0,0,0,46,0,250,0,192,0,137,0,224,0,106,0,154,0,0,0,68,0,161,0,105,0,93,0,56,0,0,0,0,0,1,0,196,0,0,0,0,0,228,0,112,0,167,0,0,0,159,0,225,0,49,0,62,0,191,0,235,0,0,0,206,0,189,0,209,0,63,0,0,0,0,0,170,0,0,0,31,0,164,0,0,0,230,0,171,0,71,0,0,0,9,0,119,0,0,0,251,0,40,0,105,0,80,0,58,0,10,0,0,0,46,0,235,0,221,0,195,0,82,0,154,0,0,0,0,0,171,0,183,0,222,0,0,0,141,0,173,0,209,0,162,0,36,0,144,0,136,0,140,0,0,0,0,0,95,0,229,0,177,0,194,0,219,0,0,0,0,0,105,0,68,0,0,0,30,0,0,0,171,0,28,0,48,0,86,0,159,0,217,0,38,0,118,0,0,0,109,0,7,0,139,0,0,0,41,0,105,0,0,0,113,0,111,0,107,0,1,0,142,0,0,0,214,0,0,0,186,0,131,0,82,0,234,0,71,0,0,0,0,0,0,0,216,0,139,0,125,0,219,0,0,0,184,0,0,0,150,0,0,0,55,0,0,0,76,0,2,0,86,0,126,0,74,0,184,0,44,0,154,0,133,0,0,0,137,0,119,0,104,0,205,0,199,0,205,0,205,0,23,0,232,0,137,0,58,0,234,0,71,0,93,0,68,0,184,0,220,0,98,0,29,0,39,0,7,0,26,0,69,0,0,0,103,0,194,0,165,0,147,0,0,0,57,0,74,0,58,0,84,0,0,0,45,0,101,0,0,0,181,0,12,0,0,0,0,0,136,0,175,0,131,0,33,0,0,0,0,0,75,0,0,0,115,0,120,0,89,0,106,0,12,0,213,0,73,0,27,0,129,0,47,0,0,0,158,0,109,0,76,0,24,0,193,0,41,0,0,0,154,0,248,0,24,0,249,0,33,0,107,0,244,0,151,0,21,0,229,0,46,0,37,0,0,0,0,0,0,0,167,0,232,0,244,0,153,0,16,0,184,0,0,0,33,0,0,0,216,0,0,0,0,0,145,0,40,0,0,0,122,0,39,0,0,0,34,0,38,0,0,0,224,0,122,0,0,0,103,0,98,0,197,0,0,0,61,0,24,0,0,0,41,0,233,0,210,0,200,0,119,0,160,0,201,0,149,0,1,0,136,0,99,0,244,0,159,0,28,0,55,0,85,0,0,0,75,0,161,0,0,0,123,0,104,0,0,0,163,0,225,0,128,0,0,0,43,0,250,0,0,0,125,0,217,0,12,0,52,0,247,0,0,0,170,0,48,0,100,0,119,0,67,0,62,0,0,0,106,0,131,0,0,0,63,0,221,0,6,0,128,0,236,0,246,0,175,0,0,0,45,0,213,0,0,0,0,0,206,0,112,0,0,0,13,0,36,0,0,0,96,0,218,0,205,0,174,0,95,0,163,0,29,0,219,0,0,0,179,0,192,0,0,0,0,0,28,0,174,0,237,0,169,0,138,0,5,0,131,0,3,0,157,0,68,0,32,0,207,0,52,0,182,0,0,0,0,0,233,0,188,0,137,0,34,0,0,0,20,0,187,0,0,0,159,0,150,0,0,0,209,0,58,0,162,0,172,0,8,0,255,0,39,0,189,0,82,0,213,0,101,0,47,0,160,0,152,0,0,0,212,0,231,0,158,0,100,0,0,0,72,0,208,0,255,0,92,0,144,0,171,0,109,0,129,0,1,0,252,0,11,0,68,0,0,0,254,0,191,0,114,0,210,0,98,0,153,0,161,0,0,0,23,0,174,0,5,0,146,0,222,0,116,0,109,0,30,0,139,0,249,0,210,0,40,0,0,0,191,0,246,0,49,0,136,0,109,0,59,0,91,0,23,0,6,0,78,0,131,0,31,0,150,0,80,0,232,0,191,0,0,0,0,0,0,0,166,0,82,0,0,0,97,0,212,0,54,0,0,0,0,0,180,0,157,0,223,0,0,0,207,0,222,0,45,0,176,0,0,0,41,0,114,0,167,0,102,0,0,0,108,0,0,0,79,0,138,0,53,0,42,0,56,0,130,0,231,0,0,0,204,0,214,0,198,0,119,0,88,0,248,0,0,0,224,0,0,0,51,0,232,0,245,0,154,0,16,0,0,0,239,0,104,0,0,0,182,0,148,0,107,0,120,0,195,0,245,0,110,0,152,0,0,0,113,0,0,0,133,0,0,0,218,0,94,0,108,0,110,0,192,0,26,0,152,0,0,0,0,0,255,0,0,0,218,0,39,0,241,0,44,0,115,0,124,0,0,0,247,0,86,0,85,0,0,0,0,0,68,0,7,0,221,0,0,0,137,0,243,0,250,0,94,0,120,0,38,0,42,0,0,0,151,0,82,0,65,0,224,0,196,0,138,0,14,0,42,0,1,0,153,0,213,0,115,0,5,0,74,0,0,0,0,0,0,0,183,0,42,0,85,0,222,0,94,0,20,0,28,0,57,0,0,0,0,0,250,0,224,0,7,0,247,0,0,0,197,0,0,0,156,0,4,0,0,0,131,0,195,0,24,0,0,0,72,0,214,0,33,0,59,0,127,0,0,0,0,0,70,0,0,0,0,0,32,0,114,0,35,0,131,0,144,0,252,0,0,0,186,0,98,0,166,0,21,0,29,0,148,0,108,0,225,0,200,0,109,0,37,0,239,0,0,0,207,0,100,0,163,0,187,0,130,0,0,0,0,0,0,0,174,0,17,0,238,0,217,0,58,0,3,0,48,0,4,0,177,0,88,0,93,0,0,0,0,0,200,0,0,0,13,0,0,0,68,0,51,0,27,0,0,0,226,0,78,0,0,0,11,0,245,0,0,0,172,0,167,0,0,0,0,0,0,0,17,0,0,0,129,0,27,0,172,0,49,0,133,0,187,0,125,0,141,0,237,0,126,0,217,0,34,0,150,0,0,0,0,0,204,0,254,0,0,0,11,0,225,0,0,0,0,0,5,0,8,0,0,0,33,0,106,0,40,0,24,0,0,0,33,0,0,0,0,0,0,0,39,0,194,0,149,0,213,0,239,0,166,0,216,0,134,0,74,0,0,0,0,0,207,0,92,0,215,0,169,0,0,0,0,0,151,0,49,0,98,0,0,0,84,0,0,0,0,0,175,0,12,0,51,0,131,0,9,0,124,0,186,0,230,0,168,0,165,0,0,0,155,0,255,0,227,0,123,0,242,0,68,0,0,0,12,0,0,0,9,0,86,0,145,0,101,0,128,0,0,0,209,0,118,0,179,0,77,0,0,0,0,0,58,0,199,0,27,0,0,0,79,0,227,0,77,0,0,0,94,0,246,0,187,0,121,0,65,0,111,0,91,0,62,0,0,0,230,0,159,0,55,0,125,0,185,0,122,0,0,0,252,0,106,0,132,0,245,0,0,0,105,0,164,0,0,0,2,0,170,0,0,0,126,0,0,0,0,0,132,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,162,31,146,31,248,31,19,31,19,30,132,31,170,31,180,31,224,31,224,30,66,31,185,31,97,31,162,31,138,31,34,31,133,31,133,30,175,31,97,31,15,31,15,30,41,31,19,31,42,31,95,31,175,31,148,31,241,31,220,31,220,30,102,31,91,31,91,30,252,31,183,31,174,31,37,31,37,30,251,31,121,31,230,31,230,30,196,31,214,31,11,31,182,31,182,30,138,31,186,31,186,30,186,29,97,31,97,30,146,31,163,31,154,31,134,31,36,31,104,31,50,31,111,31,111,30,177,31,238,31,238,30,156,31,156,30,59,31,138,31,60,31,60,30,60,29,59,31,59,30,57,31,124,31,123,31,92,31,137,31,137,30,132,31,20,31,85,31,123,31,123,30,123,29,12,31,63,31,144,31,154,31,134,31,206,31,206,30,206,29,206,28,206,27,206,26,46,31,250,31,192,31,137,31,224,31,106,31,154,31,154,30,68,31,161,31,105,31,93,31,56,31,56,30,56,29,1,31,196,31,196,30,196,29,228,31,112,31,167,31,167,30,159,31,225,31,49,31,62,31,191,31,235,31,235,30,206,31,189,31,209,31,63,31,63,30,63,29,170,31,170,30,31,31,164,31,164,30,230,31,171,31,71,31,71,30,9,31,119,31,119,30,251,31,40,31,105,31,80,31,58,31,10,31,10,30,46,31,235,31,221,31,195,31,82,31,154,31,154,30,154,29,171,31,183,31,222,31,222,30,141,31,173,31,209,31,162,31,36,31,144,31,136,31,140,31,140,30,140,29,95,31,229,31,177,31,194,31,219,31,219,30,219,29,105,31,68,31,68,30,30,31,30,30,171,31,28,31,48,31,86,31,159,31,217,31,38,31,118,31,118,30,109,31,7,31,139,31,139,30,41,31,105,31,105,30,113,31,111,31,107,31,1,31,142,31,142,30,214,31,214,30,186,31,131,31,82,31,234,31,71,31,71,30,71,29,71,28,216,31,139,31,125,31,219,31,219,30,184,31,184,30,150,31,150,30,55,31,55,30,76,31,2,31,86,31,126,31,74,31,184,31,44,31,154,31,133,31,133,30,137,31,119,31,104,31,205,31,199,31,205,31,205,31,23,31,232,31,137,31,58,31,234,31,71,31,93,31,68,31,184,31,220,31,98,31,29,31,39,31,7,31,26,31,69,31,69,30,103,31,194,31,165,31,147,31,147,30,57,31,74,31,58,31,84,31,84,30,45,31,101,31,101,30,181,31,12,31,12,30,12,29,136,31,175,31,131,31,33,31,33,30,33,29,75,31,75,30,115,31,120,31,89,31,106,31,12,31,213,31,73,31,27,31,129,31,47,31,47,30,158,31,109,31,76,31,24,31,193,31,41,31,41,30,154,31,248,31,24,31,249,31,33,31,107,31,244,31,151,31,21,31,229,31,46,31,37,31,37,30,37,29,37,28,167,31,232,31,244,31,153,31,16,31,184,31,184,30,33,31,33,30,216,31,216,30,216,29,145,31,40,31,40,30,122,31,39,31,39,30,34,31,38,31,38,30,224,31,122,31,122,30,103,31,98,31,197,31,197,30,61,31,24,31,24,30,41,31,233,31,210,31,200,31,119,31,160,31,201,31,149,31,1,31,136,31,99,31,244,31,159,31,28,31,55,31,85,31,85,30,75,31,161,31,161,30,123,31,104,31,104,30,163,31,225,31,128,31,128,30,43,31,250,31,250,30,125,31,217,31,12,31,52,31,247,31,247,30,170,31,48,31,100,31,119,31,67,31,62,31,62,30,106,31,131,31,131,30,63,31,221,31,6,31,128,31,236,31,246,31,175,31,175,30,45,31,213,31,213,30,213,29,206,31,112,31,112,30,13,31,36,31,36,30,96,31,218,31,205,31,174,31,95,31,163,31,29,31,219,31,219,30,179,31,192,31,192,30,192,29,28,31,174,31,237,31,169,31,138,31,5,31,131,31,3,31,157,31,68,31,32,31,207,31,52,31,182,31,182,30,182,29,233,31,188,31,137,31,34,31,34,30,20,31,187,31,187,30,159,31,150,31,150,30,209,31,58,31,162,31,172,31,8,31,255,31,39,31,189,31,82,31,213,31,101,31,47,31,160,31,152,31,152,30,212,31,231,31,158,31,100,31,100,30,72,31,208,31,255,31,92,31,144,31,171,31,109,31,129,31,1,31,252,31,11,31,68,31,68,30,254,31,191,31,114,31,210,31,98,31,153,31,161,31,161,30,23,31,174,31,5,31,146,31,222,31,116,31,109,31,30,31,139,31,249,31,210,31,40,31,40,30,191,31,246,31,49,31,136,31,109,31,59,31,91,31,23,31,6,31,78,31,131,31,31,31,150,31,80,31,232,31,191,31,191,30,191,29,191,28,166,31,82,31,82,30,97,31,212,31,54,31,54,30,54,29,180,31,157,31,223,31,223,30,207,31,222,31,45,31,176,31,176,30,41,31,114,31,167,31,102,31,102,30,108,31,108,30,79,31,138,31,53,31,42,31,56,31,130,31,231,31,231,30,204,31,214,31,198,31,119,31,88,31,248,31,248,30,224,31,224,30,51,31,232,31,245,31,154,31,16,31,16,30,239,31,104,31,104,30,182,31,148,31,107,31,120,31,195,31,245,31,110,31,152,31,152,30,113,31,113,30,133,31,133,30,218,31,94,31,108,31,110,31,192,31,26,31,152,31,152,30,152,29,255,31,255,30,218,31,39,31,241,31,44,31,115,31,124,31,124,30,247,31,86,31,85,31,85,30,85,29,68,31,7,31,221,31,221,30,137,31,243,31,250,31,94,31,120,31,38,31,42,31,42,30,151,31,82,31,65,31,224,31,196,31,138,31,14,31,42,31,1,31,153,31,213,31,115,31,5,31,74,31,74,30,74,29,74,28,183,31,42,31,85,31,222,31,94,31,20,31,28,31,57,31,57,30,57,29,250,31,224,31,7,31,247,31,247,30,197,31,197,30,156,31,4,31,4,30,131,31,195,31,24,31,24,30,72,31,214,31,33,31,59,31,127,31,127,30,127,29,70,31,70,30,70,29,32,31,114,31,35,31,131,31,144,31,252,31,252,30,186,31,98,31,166,31,21,31,29,31,148,31,108,31,225,31,200,31,109,31,37,31,239,31,239,30,207,31,100,31,163,31,187,31,130,31,130,30,130,29,130,28,174,31,17,31,238,31,217,31,58,31,3,31,48,31,4,31,177,31,88,31,93,31,93,30,93,29,200,31,200,30,13,31,13,30,68,31,51,31,27,31,27,30,226,31,78,31,78,30,11,31,245,31,245,30,172,31,167,31,167,30,167,29,167,28,17,31,17,30,129,31,27,31,172,31,49,31,133,31,187,31,125,31,141,31,237,31,126,31,217,31,34,31,150,31,150,30,150,29,204,31,254,31,254,30,11,31,225,31,225,30,225,29,5,31,8,31,8,30,33,31,106,31,40,31,24,31,24,30,33,31,33,30,33,29,33,28,39,31,194,31,149,31,213,31,239,31,166,31,216,31,134,31,74,31,74,30,74,29,207,31,92,31,215,31,169,31,169,30,169,29,151,31,49,31,98,31,98,30,84,31,84,30,84,29,175,31,12,31,51,31,131,31,9,31,124,31,186,31,230,31,168,31,165,31,165,30,155,31,255,31,227,31,123,31,242,31,68,31,68,30,12,31,12,30,9,31,86,31,145,31,101,31,128,31,128,30,209,31,118,31,179,31,77,31,77,30,77,29,58,31,199,31,27,31,27,30,79,31,227,31,77,31,77,30,94,31,246,31,187,31,121,31,65,31,111,31,91,31,62,31,62,30,230,31,159,31,55,31,125,31,185,31,122,31,122,30,252,31,106,31,132,31,245,31,245,30,105,31,164,31,164,30,2,31,170,31,170,30,126,31,126,30,126,29,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
