-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 825;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (54,0,73,0,213,0,22,0,168,0,24,0,60,0,0,0,249,0,240,0,125,0,172,0,138,0,0,0,165,0,191,0,204,0,36,0,28,0,177,0,193,0,153,0,234,0,11,0,0,0,80,0,29,0,193,0,88,0,0,0,138,0,124,0,225,0,231,0,15,0,219,0,0,0,0,0,202,0,137,0,151,0,25,0,210,0,30,0,98,0,36,0,0,0,244,0,162,0,44,0,0,0,47,0,141,0,65,0,103,0,196,0,0,0,56,0,6,0,0,0,178,0,180,0,76,0,102,0,230,0,0,0,18,0,240,0,20,0,235,0,170,0,21,0,4,0,128,0,111,0,198,0,1,0,164,0,23,0,96,0,100,0,145,0,81,0,0,0,0,0,11,0,142,0,0,0,224,0,164,0,55,0,34,0,72,0,37,0,125,0,0,0,0,0,54,0,207,0,0,0,128,0,210,0,7,0,63,0,0,0,17,0,0,0,173,0,99,0,200,0,0,0,178,0,240,0,80,0,216,0,0,0,73,0,0,0,15,0,255,0,0,0,197,0,0,0,56,0,72,0,0,0,53,0,138,0,194,0,0,0,65,0,180,0,2,0,68,0,119,0,0,0,88,0,132,0,45,0,0,0,54,0,151,0,182,0,120,0,51,0,124,0,0,0,0,0,89,0,91,0,164,0,186,0,0,0,82,0,0,0,202,0,0,0,251,0,124,0,91,0,0,0,36,0,0,0,0,0,199,0,31,0,155,0,0,0,87,0,198,0,153,0,50,0,75,0,135,0,32,0,19,0,194,0,113,0,210,0,145,0,233,0,129,0,0,0,151,0,232,0,120,0,0,0,0,0,26,0,195,0,98,0,4,0,0,0,0,0,35,0,0,0,0,0,0,0,0,0,53,0,39,0,23,0,63,0,174,0,126,0,149,0,90,0,0,0,106,0,24,0,158,0,33,0,167,0,0,0,148,0,0,0,49,0,252,0,188,0,141,0,54,0,247,0,53,0,164,0,112,0,28,0,247,0,175,0,0,0,84,0,0,0,186,0,187,0,140,0,0,0,153,0,0,0,87,0,117,0,0,0,87,0,16,0,197,0,132,0,177,0,213,0,29,0,184,0,147,0,0,0,232,0,156,0,102,0,91,0,229,0,20,0,91,0,80,0,0,0,211,0,218,0,17,0,233,0,252,0,49,0,0,0,81,0,0,0,0,0,78,0,0,0,32,0,252,0,156,0,245,0,0,0,0,0,106,0,184,0,255,0,215,0,133,0,0,0,30,0,191,0,17,0,251,0,131,0,0,0,232,0,0,0,204,0,114,0,159,0,198,0,135,0,40,0,183,0,92,0,111,0,0,0,196,0,192,0,82,0,25,0,38,0,101,0,188,0,88,0,175,0,57,0,171,0,0,0,99,0,93,0,100,0,84,0,22,0,62,0,67,0,0,0,241,0,181,0,242,0,61,0,29,0,0,0,0,0,201,0,22,0,186,0,252,0,14,0,180,0,0,0,74,0,205,0,145,0,0,0,208,0,0,0,93,0,0,0,74,0,59,0,208,0,0,0,71,0,150,0,244,0,126,0,120,0,0,0,161,0,159,0,199,0,0,0,182,0,190,0,0,0,0,0,21,0,0,0,141,0,0,0,254,0,0,0,0,0,152,0,195,0,0,0,234,0,0,0,37,0,83,0,0,0,191,0,26,0,230,0,198,0,240,0,0,0,102,0,15,0,0,0,0,0,157,0,59,0,99,0,98,0,153,0,85,0,117,0,113,0,24,0,162,0,131,0,172,0,16,0,9,0,35,0,198,0,248,0,248,0,0,0,0,0,227,0,0,0,169,0,164,0,174,0,152,0,64,0,147,0,242,0,59,0,198,0,0,0,91,0,215,0,44,0,135,0,190,0,0,0,49,0,33,0,0,0,9,0,71,0,0,0,119,0,12,0,136,0,34,0,78,0,79,0,86,0,145,0,180,0,0,0,0,0,237,0,52,0,53,0,0,0,0,0,0,0,186,0,152,0,145,0,0,0,204,0,81,0,22,0,112,0,140,0,178,0,205,0,14,0,50,0,21,0,83,0,19,0,0,0,23,0,236,0,212,0,74,0,0,0,221,0,160,0,182,0,208,0,0,0,19,0,33,0,197,0,0,0,146,0,0,0,25,0,199,0,64,0,67,0,47,0,202,0,0,0,0,0,244,0,0,0,123,0,145,0,0,0,0,0,67,0,0,0,140,0,0,0,160,0,134,0,236,0,166,0,65,0,55,0,154,0,227,0,158,0,62,0,31,0,226,0,69,0,98,0,98,0,0,0,89,0,0,0,70,0,36,0,198,0,199,0,41,0,59,0,0,0,221,0,0,0,249,0,138,0,141,0,210,0,130,0,174,0,147,0,0,0,199,0,172,0,254,0,173,0,241,0,82,0,0,0,30,0,64,0,22,0,45,0,211,0,0,0,225,0,0,0,195,0,192,0,171,0,0,0,202,0,143,0,81,0,106,0,0,0,128,0,59,0,2,0,33,0,184,0,238,0,117,0,30,0,1,0,164,0,217,0,75,0,35,0,93,0,44,0,202,0,172,0,56,0,4,0,210,0,38,0,70,0,28,0,0,0,147,0,107,0,108,0,0,0,140,0,117,0,54,0,0,0,138,0,217,0,161,0,235,0,252,0,12,0,0,0,215,0,103,0,149,0,0,0,0,0,0,0,0,0,246,0,0,0,106,0,194,0,80,0,0,0,81,0,0,0,36,0,56,0,0,0,233,0,239,0,51,0,179,0,0,0,180,0,221,0,143,0,196,0,0,0,56,0,189,0,175,0,75,0,210,0,3,0,55,0,0,0,112,0,217,0,1,0,133,0,216,0,0,0,0,0,239,0,99,0,0,0,70,0,40,0,0,0,113,0,225,0,0,0,33,0,103,0,125,0,251,0,211,0,236,0,243,0,173,0,0,0,162,0,62,0,30,0,254,0,149,0,20,0,223,0,143,0,37,0,217,0,107,0,62,0,216,0,34,0,248,0,0,0,0,0,37,0,64,0,245,0,80,0,121,0,0,0,91,0,250,0,159,0,100,0,91,0,15,0,71,0,167,0,47,0,76,0,0,0,250,0,0,0,0,0,0,0,7,0,12,0,0,0,74,0,5,0,0,0,77,0,224,0,123,0,105,0,0,0,113,0,0,0,15,0,80,0,122,0,85,0,233,0,44,0,205,0,99,0,193,0,0,0,54,0,0,0,0,0,36,0,0,0,0,0,157,0,146,0,140,0,5,0,2,0,14,0,209,0,18,0,249,0,0,0,196,0,103,0,136,0,153,0,125,0,0,0,98,0,145,0,90,0,53,0,20,0,223,0,6,0,202,0,247,0,128,0,161,0,32,0,62,0,186,0,32,0,52,0,116,0,0,0,163,0,0,0,240,0,37,0,251,0,0,0,235,0,0,0,8,0,69,0,239,0,222,0,96,0,140,0,0,0,0,0,246,0,139,0,0,0,0,0,22,0,251,0,145,0,66,0,100,0,132,0,90,0,0,0,4,0,244,0,0,0,102,0,36,0,255,0,55,0,20,0,170,0,0,0,180,0,161,0,136,0,208,0,0,0,220,0,6,0,225,0,0,0,41,0,139,0,12,0,27,0,53,0,7,0,124,0,206,0,46,0,0,0,95,0,66,0,93,0,0,0,39,0,255,0,187,0,79,0,0,0,16,0);
signal scenario_full  : scenario_type := (54,31,73,31,213,31,22,31,168,31,24,31,60,31,60,30,249,31,240,31,125,31,172,31,138,31,138,30,165,31,191,31,204,31,36,31,28,31,177,31,193,31,153,31,234,31,11,31,11,30,80,31,29,31,193,31,88,31,88,30,138,31,124,31,225,31,231,31,15,31,219,31,219,30,219,29,202,31,137,31,151,31,25,31,210,31,30,31,98,31,36,31,36,30,244,31,162,31,44,31,44,30,47,31,141,31,65,31,103,31,196,31,196,30,56,31,6,31,6,30,178,31,180,31,76,31,102,31,230,31,230,30,18,31,240,31,20,31,235,31,170,31,21,31,4,31,128,31,111,31,198,31,1,31,164,31,23,31,96,31,100,31,145,31,81,31,81,30,81,29,11,31,142,31,142,30,224,31,164,31,55,31,34,31,72,31,37,31,125,31,125,30,125,29,54,31,207,31,207,30,128,31,210,31,7,31,63,31,63,30,17,31,17,30,173,31,99,31,200,31,200,30,178,31,240,31,80,31,216,31,216,30,73,31,73,30,15,31,255,31,255,30,197,31,197,30,56,31,72,31,72,30,53,31,138,31,194,31,194,30,65,31,180,31,2,31,68,31,119,31,119,30,88,31,132,31,45,31,45,30,54,31,151,31,182,31,120,31,51,31,124,31,124,30,124,29,89,31,91,31,164,31,186,31,186,30,82,31,82,30,202,31,202,30,251,31,124,31,91,31,91,30,36,31,36,30,36,29,199,31,31,31,155,31,155,30,87,31,198,31,153,31,50,31,75,31,135,31,32,31,19,31,194,31,113,31,210,31,145,31,233,31,129,31,129,30,151,31,232,31,120,31,120,30,120,29,26,31,195,31,98,31,4,31,4,30,4,29,35,31,35,30,35,29,35,28,35,27,53,31,39,31,23,31,63,31,174,31,126,31,149,31,90,31,90,30,106,31,24,31,158,31,33,31,167,31,167,30,148,31,148,30,49,31,252,31,188,31,141,31,54,31,247,31,53,31,164,31,112,31,28,31,247,31,175,31,175,30,84,31,84,30,186,31,187,31,140,31,140,30,153,31,153,30,87,31,117,31,117,30,87,31,16,31,197,31,132,31,177,31,213,31,29,31,184,31,147,31,147,30,232,31,156,31,102,31,91,31,229,31,20,31,91,31,80,31,80,30,211,31,218,31,17,31,233,31,252,31,49,31,49,30,81,31,81,30,81,29,78,31,78,30,32,31,252,31,156,31,245,31,245,30,245,29,106,31,184,31,255,31,215,31,133,31,133,30,30,31,191,31,17,31,251,31,131,31,131,30,232,31,232,30,204,31,114,31,159,31,198,31,135,31,40,31,183,31,92,31,111,31,111,30,196,31,192,31,82,31,25,31,38,31,101,31,188,31,88,31,175,31,57,31,171,31,171,30,99,31,93,31,100,31,84,31,22,31,62,31,67,31,67,30,241,31,181,31,242,31,61,31,29,31,29,30,29,29,201,31,22,31,186,31,252,31,14,31,180,31,180,30,74,31,205,31,145,31,145,30,208,31,208,30,93,31,93,30,74,31,59,31,208,31,208,30,71,31,150,31,244,31,126,31,120,31,120,30,161,31,159,31,199,31,199,30,182,31,190,31,190,30,190,29,21,31,21,30,141,31,141,30,254,31,254,30,254,29,152,31,195,31,195,30,234,31,234,30,37,31,83,31,83,30,191,31,26,31,230,31,198,31,240,31,240,30,102,31,15,31,15,30,15,29,157,31,59,31,99,31,98,31,153,31,85,31,117,31,113,31,24,31,162,31,131,31,172,31,16,31,9,31,35,31,198,31,248,31,248,31,248,30,248,29,227,31,227,30,169,31,164,31,174,31,152,31,64,31,147,31,242,31,59,31,198,31,198,30,91,31,215,31,44,31,135,31,190,31,190,30,49,31,33,31,33,30,9,31,71,31,71,30,119,31,12,31,136,31,34,31,78,31,79,31,86,31,145,31,180,31,180,30,180,29,237,31,52,31,53,31,53,30,53,29,53,28,186,31,152,31,145,31,145,30,204,31,81,31,22,31,112,31,140,31,178,31,205,31,14,31,50,31,21,31,83,31,19,31,19,30,23,31,236,31,212,31,74,31,74,30,221,31,160,31,182,31,208,31,208,30,19,31,33,31,197,31,197,30,146,31,146,30,25,31,199,31,64,31,67,31,47,31,202,31,202,30,202,29,244,31,244,30,123,31,145,31,145,30,145,29,67,31,67,30,140,31,140,30,160,31,134,31,236,31,166,31,65,31,55,31,154,31,227,31,158,31,62,31,31,31,226,31,69,31,98,31,98,31,98,30,89,31,89,30,70,31,36,31,198,31,199,31,41,31,59,31,59,30,221,31,221,30,249,31,138,31,141,31,210,31,130,31,174,31,147,31,147,30,199,31,172,31,254,31,173,31,241,31,82,31,82,30,30,31,64,31,22,31,45,31,211,31,211,30,225,31,225,30,195,31,192,31,171,31,171,30,202,31,143,31,81,31,106,31,106,30,128,31,59,31,2,31,33,31,184,31,238,31,117,31,30,31,1,31,164,31,217,31,75,31,35,31,93,31,44,31,202,31,172,31,56,31,4,31,210,31,38,31,70,31,28,31,28,30,147,31,107,31,108,31,108,30,140,31,117,31,54,31,54,30,138,31,217,31,161,31,235,31,252,31,12,31,12,30,215,31,103,31,149,31,149,30,149,29,149,28,149,27,246,31,246,30,106,31,194,31,80,31,80,30,81,31,81,30,36,31,56,31,56,30,233,31,239,31,51,31,179,31,179,30,180,31,221,31,143,31,196,31,196,30,56,31,189,31,175,31,75,31,210,31,3,31,55,31,55,30,112,31,217,31,1,31,133,31,216,31,216,30,216,29,239,31,99,31,99,30,70,31,40,31,40,30,113,31,225,31,225,30,33,31,103,31,125,31,251,31,211,31,236,31,243,31,173,31,173,30,162,31,62,31,30,31,254,31,149,31,20,31,223,31,143,31,37,31,217,31,107,31,62,31,216,31,34,31,248,31,248,30,248,29,37,31,64,31,245,31,80,31,121,31,121,30,91,31,250,31,159,31,100,31,91,31,15,31,71,31,167,31,47,31,76,31,76,30,250,31,250,30,250,29,250,28,7,31,12,31,12,30,74,31,5,31,5,30,77,31,224,31,123,31,105,31,105,30,113,31,113,30,15,31,80,31,122,31,85,31,233,31,44,31,205,31,99,31,193,31,193,30,54,31,54,30,54,29,36,31,36,30,36,29,157,31,146,31,140,31,5,31,2,31,14,31,209,31,18,31,249,31,249,30,196,31,103,31,136,31,153,31,125,31,125,30,98,31,145,31,90,31,53,31,20,31,223,31,6,31,202,31,247,31,128,31,161,31,32,31,62,31,186,31,32,31,52,31,116,31,116,30,163,31,163,30,240,31,37,31,251,31,251,30,235,31,235,30,8,31,69,31,239,31,222,31,96,31,140,31,140,30,140,29,246,31,139,31,139,30,139,29,22,31,251,31,145,31,66,31,100,31,132,31,90,31,90,30,4,31,244,31,244,30,102,31,36,31,255,31,55,31,20,31,170,31,170,30,180,31,161,31,136,31,208,31,208,30,220,31,6,31,225,31,225,30,41,31,139,31,12,31,27,31,53,31,7,31,124,31,206,31,46,31,46,30,95,31,66,31,93,31,93,30,39,31,255,31,187,31,79,31,79,30,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
