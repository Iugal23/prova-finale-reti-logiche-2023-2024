-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_469 is
end project_tb_469;

architecture project_tb_arch_469 of project_tb_469 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 807;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,181,0,0,0,155,0,67,0,172,0,12,0,69,0,250,0,167,0,180,0,66,0,74,0,21,0,11,0,0,0,144,0,0,0,118,0,236,0,127,0,48,0,36,0,163,0,179,0,100,0,158,0,40,0,92,0,105,0,0,0,245,0,158,0,0,0,35,0,51,0,0,0,0,0,246,0,246,0,209,0,145,0,244,0,193,0,14,0,29,0,0,0,0,0,181,0,200,0,58,0,160,0,0,0,24,0,72,0,0,0,232,0,0,0,198,0,210,0,179,0,91,0,249,0,105,0,67,0,230,0,81,0,251,0,82,0,222,0,79,0,28,0,97,0,14,0,157,0,70,0,14,0,242,0,0,0,0,0,22,0,0,0,53,0,153,0,101,0,69,0,61,0,0,0,140,0,4,0,235,0,239,0,19,0,36,0,81,0,15,0,24,0,120,0,0,0,251,0,95,0,105,0,253,0,0,0,147,0,251,0,222,0,25,0,165,0,15,0,0,0,193,0,148,0,213,0,252,0,37,0,88,0,16,0,77,0,20,0,85,0,144,0,0,0,0,0,73,0,58,0,81,0,159,0,182,0,199,0,98,0,33,0,76,0,0,0,242,0,219,0,226,0,3,0,250,0,31,0,0,0,65,0,99,0,79,0,227,0,247,0,0,0,0,0,69,0,0,0,0,0,54,0,147,0,249,0,158,0,0,0,68,0,250,0,0,0,233,0,200,0,0,0,234,0,30,0,14,0,248,0,106,0,76,0,77,0,113,0,0,0,54,0,198,0,58,0,125,0,0,0,176,0,179,0,139,0,125,0,0,0,15,0,62,0,140,0,0,0,228,0,0,0,0,0,131,0,0,0,105,0,238,0,33,0,0,0,59,0,99,0,200,0,66,0,2,0,37,0,179,0,157,0,29,0,161,0,171,0,206,0,141,0,10,0,0,0,2,0,37,0,246,0,180,0,208,0,253,0,119,0,57,0,197,0,116,0,136,0,206,0,170,0,24,0,56,0,181,0,147,0,115,0,102,0,76,0,0,0,58,0,212,0,113,0,94,0,156,0,11,0,71,0,48,0,94,0,60,0,227,0,29,0,0,0,244,0,125,0,0,0,58,0,5,0,37,0,15,0,243,0,151,0,252,0,0,0,99,0,80,0,145,0,13,0,11,0,126,0,97,0,45,0,18,0,77,0,67,0,188,0,8,0,97,0,234,0,213,0,187,0,92,0,200,0,0,0,0,0,5,0,0,0,81,0,79,0,113,0,112,0,211,0,37,0,0,0,18,0,95,0,198,0,193,0,190,0,233,0,0,0,0,0,89,0,247,0,43,0,111,0,235,0,0,0,115,0,0,0,134,0,179,0,18,0,78,0,172,0,0,0,63,0,109,0,49,0,135,0,160,0,107,0,183,0,109,0,0,0,0,0,138,0,0,0,0,0,245,0,159,0,0,0,6,0,141,0,247,0,252,0,55,0,62,0,0,0,25,0,0,0,45,0,76,0,67,0,0,0,0,0,138,0,0,0,0,0,237,0,244,0,80,0,148,0,117,0,0,0,56,0,88,0,140,0,105,0,27,0,0,0,215,0,127,0,154,0,159,0,77,0,13,0,194,0,57,0,74,0,183,0,146,0,0,0,51,0,217,0,208,0,0,0,130,0,0,0,115,0,176,0,76,0,0,0,83,0,134,0,35,0,169,0,47,0,96,0,100,0,222,0,76,0,161,0,37,0,163,0,166,0,218,0,0,0,125,0,188,0,0,0,0,0,3,0,172,0,101,0,203,0,148,0,0,0,178,0,54,0,190,0,0,0,81,0,34,0,225,0,161,0,125,0,42,0,254,0,189,0,109,0,0,0,138,0,40,0,0,0,17,0,18,0,20,0,250,0,43,0,176,0,135,0,196,0,96,0,40,0,45,0,58,0,0,0,244,0,113,0,133,0,0,0,0,0,69,0,8,0,175,0,156,0,99,0,236,0,150,0,129,0,192,0,0,0,105,0,94,0,92,0,37,0,0,0,147,0,62,0,249,0,75,0,0,0,147,0,30,0,153,0,71,0,29,0,0,0,46,0,0,0,21,0,92,0,198,0,51,0,249,0,37,0,234,0,0,0,42,0,43,0,141,0,56,0,108,0,172,0,87,0,12,0,249,0,122,0,0,0,95,0,0,0,133,0,29,0,121,0,132,0,0,0,153,0,154,0,174,0,118,0,200,0,17,0,0,0,191,0,106,0,0,0,3,0,34,0,74,0,244,0,52,0,242,0,0,0,0,0,145,0,0,0,129,0,121,0,231,0,0,0,184,0,236,0,147,0,45,0,199,0,57,0,172,0,0,0,62,0,31,0,122,0,64,0,214,0,41,0,69,0,195,0,0,0,26,0,186,0,152,0,0,0,252,0,185,0,128,0,119,0,0,0,167,0,199,0,95,0,249,0,5,0,30,0,241,0,116,0,234,0,222,0,238,0,139,0,183,0,132,0,0,0,150,0,149,0,0,0,207,0,204,0,244,0,0,0,238,0,168,0,94,0,171,0,202,0,0,0,28,0,0,0,131,0,253,0,0,0,34,0,134,0,61,0,227,0,247,0,243,0,84,0,250,0,68,0,165,0,240,0,165,0,103,0,36,0,78,0,160,0,36,0,247,0,251,0,0,0,197,0,197,0,8,0,208,0,0,0,247,0,255,0,120,0,92,0,195,0,26,0,0,0,89,0,0,0,135,0,206,0,3,0,183,0,146,0,74,0,43,0,99,0,128,0,0,0,67,0,0,0,0,0,180,0,60,0,117,0,67,0,255,0,12,0,23,0,0,0,194,0,0,0,2,0,0,0,0,0,48,0,84,0,207,0,40,0,49,0,0,0,200,0,245,0,212,0,2,0,177,0,113,0,0,0,0,0,220,0,0,0,238,0,150,0,132,0,0,0,10,0,124,0,252,0,219,0,250,0,251,0,44,0,76,0,105,0,161,0,151,0,33,0,168,0,0,0,46,0,109,0,0,0,66,0,241,0,138,0,0,0,9,0,42,0,111,0,125,0,0,0,3,0,54,0,226,0,103,0,255,0,0,0,80,0,0,0,0,0,103,0,15,0,52,0,158,0,155,0,118,0,213,0,116,0,255,0,0,0,0,0,168,0,74,0,105,0,0,0,26,0,187,0,178,0,180,0,112,0,22,0,0,0,128,0,20,0,221,0,184,0,96,0,0,0,18,0,0,0,204,0,159,0,0,0,59,0,19,0,245,0,252,0,215,0,178,0,95,0,161,0,122,0,217,0,0,0,5,0,0,0,2,0,50,0,113,0,139,0,31,0,58,0,235,0,0,0,0,0,2,0,156,0,61,0,57,0,0,0,167,0,0,0,138,0,217,0,255,0,68,0,161,0,60,0,0,0,0,0,57,0,89,0,0,0,0,0,33,0,0,0,0,0,101,0,0,0,0,0,221,0,149,0,246,0,185,0,48,0,173,0,0,0,0,0,212,0,60,0,118,0,0,0,0,0,137,0,20,0,0,0,0,0,235,0,50,0,32,0,139,0,127,0,251,0,47,0,240,0,233,0,204,0,0,0,112,0,246,0,158,0,59,0,151,0,0,0,0,0,0,0,26,0,127,0,9,0,207,0,126,0,0,0);
signal scenario_full  : scenario_type := (0,0,181,31,181,30,155,31,67,31,172,31,12,31,69,31,250,31,167,31,180,31,66,31,74,31,21,31,11,31,11,30,144,31,144,30,118,31,236,31,127,31,48,31,36,31,163,31,179,31,100,31,158,31,40,31,92,31,105,31,105,30,245,31,158,31,158,30,35,31,51,31,51,30,51,29,246,31,246,31,209,31,145,31,244,31,193,31,14,31,29,31,29,30,29,29,181,31,200,31,58,31,160,31,160,30,24,31,72,31,72,30,232,31,232,30,198,31,210,31,179,31,91,31,249,31,105,31,67,31,230,31,81,31,251,31,82,31,222,31,79,31,28,31,97,31,14,31,157,31,70,31,14,31,242,31,242,30,242,29,22,31,22,30,53,31,153,31,101,31,69,31,61,31,61,30,140,31,4,31,235,31,239,31,19,31,36,31,81,31,15,31,24,31,120,31,120,30,251,31,95,31,105,31,253,31,253,30,147,31,251,31,222,31,25,31,165,31,15,31,15,30,193,31,148,31,213,31,252,31,37,31,88,31,16,31,77,31,20,31,85,31,144,31,144,30,144,29,73,31,58,31,81,31,159,31,182,31,199,31,98,31,33,31,76,31,76,30,242,31,219,31,226,31,3,31,250,31,31,31,31,30,65,31,99,31,79,31,227,31,247,31,247,30,247,29,69,31,69,30,69,29,54,31,147,31,249,31,158,31,158,30,68,31,250,31,250,30,233,31,200,31,200,30,234,31,30,31,14,31,248,31,106,31,76,31,77,31,113,31,113,30,54,31,198,31,58,31,125,31,125,30,176,31,179,31,139,31,125,31,125,30,15,31,62,31,140,31,140,30,228,31,228,30,228,29,131,31,131,30,105,31,238,31,33,31,33,30,59,31,99,31,200,31,66,31,2,31,37,31,179,31,157,31,29,31,161,31,171,31,206,31,141,31,10,31,10,30,2,31,37,31,246,31,180,31,208,31,253,31,119,31,57,31,197,31,116,31,136,31,206,31,170,31,24,31,56,31,181,31,147,31,115,31,102,31,76,31,76,30,58,31,212,31,113,31,94,31,156,31,11,31,71,31,48,31,94,31,60,31,227,31,29,31,29,30,244,31,125,31,125,30,58,31,5,31,37,31,15,31,243,31,151,31,252,31,252,30,99,31,80,31,145,31,13,31,11,31,126,31,97,31,45,31,18,31,77,31,67,31,188,31,8,31,97,31,234,31,213,31,187,31,92,31,200,31,200,30,200,29,5,31,5,30,81,31,79,31,113,31,112,31,211,31,37,31,37,30,18,31,95,31,198,31,193,31,190,31,233,31,233,30,233,29,89,31,247,31,43,31,111,31,235,31,235,30,115,31,115,30,134,31,179,31,18,31,78,31,172,31,172,30,63,31,109,31,49,31,135,31,160,31,107,31,183,31,109,31,109,30,109,29,138,31,138,30,138,29,245,31,159,31,159,30,6,31,141,31,247,31,252,31,55,31,62,31,62,30,25,31,25,30,45,31,76,31,67,31,67,30,67,29,138,31,138,30,138,29,237,31,244,31,80,31,148,31,117,31,117,30,56,31,88,31,140,31,105,31,27,31,27,30,215,31,127,31,154,31,159,31,77,31,13,31,194,31,57,31,74,31,183,31,146,31,146,30,51,31,217,31,208,31,208,30,130,31,130,30,115,31,176,31,76,31,76,30,83,31,134,31,35,31,169,31,47,31,96,31,100,31,222,31,76,31,161,31,37,31,163,31,166,31,218,31,218,30,125,31,188,31,188,30,188,29,3,31,172,31,101,31,203,31,148,31,148,30,178,31,54,31,190,31,190,30,81,31,34,31,225,31,161,31,125,31,42,31,254,31,189,31,109,31,109,30,138,31,40,31,40,30,17,31,18,31,20,31,250,31,43,31,176,31,135,31,196,31,96,31,40,31,45,31,58,31,58,30,244,31,113,31,133,31,133,30,133,29,69,31,8,31,175,31,156,31,99,31,236,31,150,31,129,31,192,31,192,30,105,31,94,31,92,31,37,31,37,30,147,31,62,31,249,31,75,31,75,30,147,31,30,31,153,31,71,31,29,31,29,30,46,31,46,30,21,31,92,31,198,31,51,31,249,31,37,31,234,31,234,30,42,31,43,31,141,31,56,31,108,31,172,31,87,31,12,31,249,31,122,31,122,30,95,31,95,30,133,31,29,31,121,31,132,31,132,30,153,31,154,31,174,31,118,31,200,31,17,31,17,30,191,31,106,31,106,30,3,31,34,31,74,31,244,31,52,31,242,31,242,30,242,29,145,31,145,30,129,31,121,31,231,31,231,30,184,31,236,31,147,31,45,31,199,31,57,31,172,31,172,30,62,31,31,31,122,31,64,31,214,31,41,31,69,31,195,31,195,30,26,31,186,31,152,31,152,30,252,31,185,31,128,31,119,31,119,30,167,31,199,31,95,31,249,31,5,31,30,31,241,31,116,31,234,31,222,31,238,31,139,31,183,31,132,31,132,30,150,31,149,31,149,30,207,31,204,31,244,31,244,30,238,31,168,31,94,31,171,31,202,31,202,30,28,31,28,30,131,31,253,31,253,30,34,31,134,31,61,31,227,31,247,31,243,31,84,31,250,31,68,31,165,31,240,31,165,31,103,31,36,31,78,31,160,31,36,31,247,31,251,31,251,30,197,31,197,31,8,31,208,31,208,30,247,31,255,31,120,31,92,31,195,31,26,31,26,30,89,31,89,30,135,31,206,31,3,31,183,31,146,31,74,31,43,31,99,31,128,31,128,30,67,31,67,30,67,29,180,31,60,31,117,31,67,31,255,31,12,31,23,31,23,30,194,31,194,30,2,31,2,30,2,29,48,31,84,31,207,31,40,31,49,31,49,30,200,31,245,31,212,31,2,31,177,31,113,31,113,30,113,29,220,31,220,30,238,31,150,31,132,31,132,30,10,31,124,31,252,31,219,31,250,31,251,31,44,31,76,31,105,31,161,31,151,31,33,31,168,31,168,30,46,31,109,31,109,30,66,31,241,31,138,31,138,30,9,31,42,31,111,31,125,31,125,30,3,31,54,31,226,31,103,31,255,31,255,30,80,31,80,30,80,29,103,31,15,31,52,31,158,31,155,31,118,31,213,31,116,31,255,31,255,30,255,29,168,31,74,31,105,31,105,30,26,31,187,31,178,31,180,31,112,31,22,31,22,30,128,31,20,31,221,31,184,31,96,31,96,30,18,31,18,30,204,31,159,31,159,30,59,31,19,31,245,31,252,31,215,31,178,31,95,31,161,31,122,31,217,31,217,30,5,31,5,30,2,31,50,31,113,31,139,31,31,31,58,31,235,31,235,30,235,29,2,31,156,31,61,31,57,31,57,30,167,31,167,30,138,31,217,31,255,31,68,31,161,31,60,31,60,30,60,29,57,31,89,31,89,30,89,29,33,31,33,30,33,29,101,31,101,30,101,29,221,31,149,31,246,31,185,31,48,31,173,31,173,30,173,29,212,31,60,31,118,31,118,30,118,29,137,31,20,31,20,30,20,29,235,31,50,31,32,31,139,31,127,31,251,31,47,31,240,31,233,31,204,31,204,30,112,31,246,31,158,31,59,31,151,31,151,30,151,29,151,28,26,31,127,31,9,31,207,31,126,31,126,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
