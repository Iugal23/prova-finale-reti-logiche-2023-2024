-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_208 is
end project_tb_208;

architecture project_tb_arch_208 of project_tb_208 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1023;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (130,0,5,0,0,0,31,0,0,0,175,0,0,0,63,0,16,0,94,0,79,0,143,0,229,0,56,0,103,0,191,0,138,0,58,0,184,0,4,0,203,0,251,0,181,0,0,0,251,0,135,0,23,0,107,0,95,0,14,0,0,0,35,0,4,0,40,0,0,0,85,0,70,0,238,0,113,0,57,0,215,0,136,0,45,0,153,0,217,0,90,0,27,0,89,0,0,0,203,0,217,0,86,0,0,0,204,0,36,0,206,0,0,0,32,0,49,0,191,0,147,0,0,0,83,0,53,0,207,0,30,0,23,0,83,0,3,0,200,0,137,0,0,0,87,0,2,0,244,0,0,0,0,0,0,0,177,0,0,0,204,0,0,0,64,0,0,0,80,0,136,0,97,0,46,0,188,0,215,0,0,0,215,0,0,0,0,0,0,0,0,0,167,0,139,0,188,0,0,0,72,0,239,0,74,0,28,0,136,0,39,0,0,0,191,0,82,0,171,0,0,0,252,0,106,0,0,0,229,0,242,0,173,0,169,0,0,0,7,0,26,0,0,0,64,0,103,0,9,0,8,0,177,0,126,0,179,0,40,0,0,0,135,0,215,0,103,0,55,0,250,0,19,0,139,0,239,0,38,0,246,0,0,0,86,0,0,0,175,0,168,0,115,0,0,0,137,0,82,0,179,0,13,0,243,0,119,0,123,0,43,0,9,0,141,0,2,0,100,0,238,0,0,0,93,0,2,0,53,0,235,0,145,0,95,0,99,0,169,0,254,0,183,0,179,0,0,0,19,0,150,0,58,0,203,0,216,0,228,0,250,0,160,0,7,0,9,0,61,0,113,0,179,0,0,0,247,0,0,0,0,0,131,0,228,0,217,0,0,0,166,0,33,0,51,0,221,0,0,0,232,0,0,0,0,0,0,0,137,0,0,0,0,0,107,0,0,0,78,0,240,0,218,0,115,0,0,0,242,0,252,0,131,0,148,0,133,0,92,0,41,0,63,0,210,0,154,0,131,0,18,0,138,0,0,0,0,0,69,0,30,0,240,0,80,0,161,0,72,0,47,0,0,0,127,0,63,0,108,0,71,0,0,0,24,0,31,0,201,0,18,0,0,0,125,0,123,0,208,0,0,0,15,0,139,0,14,0,51,0,82,0,105,0,188,0,16,0,120,0,48,0,177,0,0,0,63,0,144,0,120,0,215,0,26,0,149,0,49,0,192,0,233,0,0,0,115,0,167,0,0,0,0,0,0,0,34,0,0,0,126,0,66,0,193,0,18,0,0,0,139,0,136,0,96,0,121,0,0,0,0,0,65,0,184,0,0,0,109,0,16,0,108,0,6,0,89,0,184,0,35,0,0,0,210,0,0,0,0,0,225,0,191,0,193,0,196,0,204,0,0,0,138,0,53,0,101,0,216,0,0,0,156,0,0,0,32,0,234,0,0,0,65,0,210,0,80,0,92,0,153,0,57,0,31,0,218,0,187,0,92,0,46,0,113,0,0,0,97,0,0,0,63,0,0,0,0,0,0,0,12,0,53,0,132,0,151,0,58,0,157,0,255,0,225,0,155,0,131,0,34,0,23,0,40,0,0,0,159,0,102,0,25,0,0,0,101,0,134,0,158,0,0,0,101,0,1,0,0,0,188,0,53,0,29,0,0,0,67,0,133,0,137,0,216,0,110,0,157,0,24,0,253,0,135,0,12,0,9,0,141,0,238,0,131,0,172,0,137,0,0,0,217,0,146,0,47,0,0,0,101,0,148,0,223,0,213,0,0,0,0,0,120,0,0,0,176,0,179,0,0,0,150,0,61,0,211,0,0,0,0,0,33,0,215,0,96,0,0,0,113,0,229,0,178,0,187,0,0,0,222,0,15,0,110,0,0,0,5,0,223,0,155,0,46,0,181,0,0,0,15,0,187,0,141,0,0,0,235,0,223,0,29,0,81,0,0,0,66,0,0,0,0,0,9,0,13,0,113,0,41,0,166,0,53,0,0,0,24,0,129,0,161,0,102,0,199,0,152,0,55,0,19,0,139,0,135,0,209,0,6,0,0,0,3,0,0,0,0,0,0,0,0,0,18,0,170,0,170,0,114,0,60,0,33,0,217,0,0,0,251,0,184,0,228,0,100,0,168,0,0,0,199,0,36,0,183,0,174,0,0,0,113,0,224,0,238,0,240,0,52,0,0,0,131,0,0,0,0,0,250,0,219,0,243,0,178,0,0,0,214,0,221,0,0,0,31,0,0,0,178,0,129,0,0,0,0,0,0,0,0,0,58,0,238,0,142,0,126,0,31,0,112,0,127,0,127,0,2,0,0,0,0,0,242,0,238,0,154,0,0,0,0,0,193,0,45,0,121,0,43,0,27,0,17,0,232,0,0,0,147,0,0,0,185,0,86,0,88,0,205,0,5,0,70,0,146,0,5,0,0,0,0,0,0,0,220,0,243,0,181,0,29,0,0,0,92,0,0,0,36,0,0,0,168,0,0,0,0,0,33,0,189,0,0,0,0,0,244,0,107,0,170,0,15,0,186,0,121,0,224,0,175,0,31,0,170,0,65,0,54,0,194,0,15,0,157,0,0,0,104,0,217,0,118,0,1,0,249,0,141,0,0,0,111,0,0,0,20,0,83,0,59,0,0,0,213,0,1,0,158,0,0,0,83,0,41,0,175,0,0,0,19,0,172,0,32,0,108,0,115,0,0,0,199,0,56,0,91,0,72,0,250,0,3,0,209,0,0,0,5,0,243,0,0,0,154,0,90,0,248,0,0,0,133,0,207,0,231,0,111,0,0,0,55,0,52,0,130,0,133,0,0,0,206,0,122,0,161,0,91,0,171,0,41,0,170,0,247,0,0,0,201,0,11,0,139,0,0,0,165,0,0,0,35,0,63,0,68,0,15,0,248,0,49,0,157,0,0,0,231,0,21,0,125,0,0,0,175,0,0,0,46,0,198,0,141,0,14,0,0,0,101,0,0,0,236,0,164,0,0,0,31,0,0,0,0,0,84,0,157,0,26,0,8,0,11,0,196,0,0,0,202,0,37,0,115,0,249,0,0,0,0,0,65,0,166,0,90,0,0,0,142,0,163,0,0,0,194,0,106,0,198,0,16,0,239,0,107,0,19,0,171,0,246,0,0,0,0,0,83,0,0,0,116,0,189,0,162,0,5,0,49,0,93,0,56,0,92,0,214,0,48,0,66,0,0,0,0,0,229,0,225,0,78,0,39,0,111,0,248,0,5,0,115,0,175,0,67,0,36,0,0,0,66,0,120,0,119,0,253,0,0,0,87,0,41,0,12,0,145,0,57,0,7,0,0,0,241,0,75,0,6,0,162,0,0,0,250,0,162,0,231,0,127,0,77,0,123,0,7,0,119,0,34,0,63,0,209,0,0,0,0,0,0,0,96,0,47,0,0,0,29,0,191,0,135,0,57,0,231,0,225,0,246,0,23,0,0,0,1,0,0,0,166,0,86,0,122,0,185,0,253,0,220,0,52,0,180,0,136,0,80,0,197,0,71,0,60,0,154,0,217,0,83,0,20,0,79,0,11,0,46,0,39,0,227,0,226,0,0,0,115,0,134,0,0,0,97,0,0,0,0,0,62,0,71,0,46,0,185,0,182,0,111,0,146,0,44,0,0,0,134,0,0,0,24,0,11,0,35,0,70,0,243,0,222,0,169,0,197,0,23,0,8,0,253,0,196,0,0,0,147,0,228,0,24,0,0,0,166,0,0,0,94,0,11,0,0,0,247,0,239,0,101,0,149,0,19,0,123,0,168,0,0,0,217,0,37,0,0,0,148,0,5,0,13,0,56,0,0,0,120,0,104,0,71,0,217,0,62,0,0,0,97,0,0,0,10,0,32,0,172,0,52,0,214,0,102,0,57,0,128,0,169,0,25,0,22,0,0,0,78,0,0,0,205,0,61,0,98,0,234,0,125,0,134,0,28,0,225,0,195,0,0,0,248,0,41,0,146,0,40,0,97,0,82,0,207,0,224,0,182,0,18,0,76,0,156,0,139,0,45,0,0,0,0,0,50,0,199,0,98,0,9,0,0,0,31,0,80,0,69,0,0,0,253,0,198,0,26,0,0,0,95,0,65,0,0,0,27,0,162,0,41,0,104,0,0,0,0,0,46,0,153,0,39,0,0,0,182,0,136,0,166,0,164,0,229,0,220,0,43,0,122,0,0,0,83,0,201,0,55,0,181,0,181,0,205,0,177,0,0,0,0,0,7,0,198,0,104,0,167,0,169,0,226,0,235,0,17,0,163,0,0,0,0,0,142,0,154,0,67,0,104,0,184,0,0,0,0,0,224,0,144,0,0,0,0,0,0,0,62,0,190,0,0,0,107,0,0,0,168,0,222,0,0,0,99,0,191,0,214,0,32,0,185,0,237,0,20,0,0,0,0,0,199,0,24,0,229,0,0,0,140,0,138,0,94,0,192,0,92,0,132,0,23,0,147,0,13,0,87,0,116,0,45,0,0,0,176,0,163,0,186,0,118,0,0,0,236,0,0,0,0,0,61,0,142,0,208,0,170,0,224,0,0,0,89,0,129,0,113,0,25,0,166,0,198,0,218,0,210,0,254,0);
signal scenario_full  : scenario_type := (130,31,5,31,5,30,31,31,31,30,175,31,175,30,63,31,16,31,94,31,79,31,143,31,229,31,56,31,103,31,191,31,138,31,58,31,184,31,4,31,203,31,251,31,181,31,181,30,251,31,135,31,23,31,107,31,95,31,14,31,14,30,35,31,4,31,40,31,40,30,85,31,70,31,238,31,113,31,57,31,215,31,136,31,45,31,153,31,217,31,90,31,27,31,89,31,89,30,203,31,217,31,86,31,86,30,204,31,36,31,206,31,206,30,32,31,49,31,191,31,147,31,147,30,83,31,53,31,207,31,30,31,23,31,83,31,3,31,200,31,137,31,137,30,87,31,2,31,244,31,244,30,244,29,244,28,177,31,177,30,204,31,204,30,64,31,64,30,80,31,136,31,97,31,46,31,188,31,215,31,215,30,215,31,215,30,215,29,215,28,215,27,167,31,139,31,188,31,188,30,72,31,239,31,74,31,28,31,136,31,39,31,39,30,191,31,82,31,171,31,171,30,252,31,106,31,106,30,229,31,242,31,173,31,169,31,169,30,7,31,26,31,26,30,64,31,103,31,9,31,8,31,177,31,126,31,179,31,40,31,40,30,135,31,215,31,103,31,55,31,250,31,19,31,139,31,239,31,38,31,246,31,246,30,86,31,86,30,175,31,168,31,115,31,115,30,137,31,82,31,179,31,13,31,243,31,119,31,123,31,43,31,9,31,141,31,2,31,100,31,238,31,238,30,93,31,2,31,53,31,235,31,145,31,95,31,99,31,169,31,254,31,183,31,179,31,179,30,19,31,150,31,58,31,203,31,216,31,228,31,250,31,160,31,7,31,9,31,61,31,113,31,179,31,179,30,247,31,247,30,247,29,131,31,228,31,217,31,217,30,166,31,33,31,51,31,221,31,221,30,232,31,232,30,232,29,232,28,137,31,137,30,137,29,107,31,107,30,78,31,240,31,218,31,115,31,115,30,242,31,252,31,131,31,148,31,133,31,92,31,41,31,63,31,210,31,154,31,131,31,18,31,138,31,138,30,138,29,69,31,30,31,240,31,80,31,161,31,72,31,47,31,47,30,127,31,63,31,108,31,71,31,71,30,24,31,31,31,201,31,18,31,18,30,125,31,123,31,208,31,208,30,15,31,139,31,14,31,51,31,82,31,105,31,188,31,16,31,120,31,48,31,177,31,177,30,63,31,144,31,120,31,215,31,26,31,149,31,49,31,192,31,233,31,233,30,115,31,167,31,167,30,167,29,167,28,34,31,34,30,126,31,66,31,193,31,18,31,18,30,139,31,136,31,96,31,121,31,121,30,121,29,65,31,184,31,184,30,109,31,16,31,108,31,6,31,89,31,184,31,35,31,35,30,210,31,210,30,210,29,225,31,191,31,193,31,196,31,204,31,204,30,138,31,53,31,101,31,216,31,216,30,156,31,156,30,32,31,234,31,234,30,65,31,210,31,80,31,92,31,153,31,57,31,31,31,218,31,187,31,92,31,46,31,113,31,113,30,97,31,97,30,63,31,63,30,63,29,63,28,12,31,53,31,132,31,151,31,58,31,157,31,255,31,225,31,155,31,131,31,34,31,23,31,40,31,40,30,159,31,102,31,25,31,25,30,101,31,134,31,158,31,158,30,101,31,1,31,1,30,188,31,53,31,29,31,29,30,67,31,133,31,137,31,216,31,110,31,157,31,24,31,253,31,135,31,12,31,9,31,141,31,238,31,131,31,172,31,137,31,137,30,217,31,146,31,47,31,47,30,101,31,148,31,223,31,213,31,213,30,213,29,120,31,120,30,176,31,179,31,179,30,150,31,61,31,211,31,211,30,211,29,33,31,215,31,96,31,96,30,113,31,229,31,178,31,187,31,187,30,222,31,15,31,110,31,110,30,5,31,223,31,155,31,46,31,181,31,181,30,15,31,187,31,141,31,141,30,235,31,223,31,29,31,81,31,81,30,66,31,66,30,66,29,9,31,13,31,113,31,41,31,166,31,53,31,53,30,24,31,129,31,161,31,102,31,199,31,152,31,55,31,19,31,139,31,135,31,209,31,6,31,6,30,3,31,3,30,3,29,3,28,3,27,18,31,170,31,170,31,114,31,60,31,33,31,217,31,217,30,251,31,184,31,228,31,100,31,168,31,168,30,199,31,36,31,183,31,174,31,174,30,113,31,224,31,238,31,240,31,52,31,52,30,131,31,131,30,131,29,250,31,219,31,243,31,178,31,178,30,214,31,221,31,221,30,31,31,31,30,178,31,129,31,129,30,129,29,129,28,129,27,58,31,238,31,142,31,126,31,31,31,112,31,127,31,127,31,2,31,2,30,2,29,242,31,238,31,154,31,154,30,154,29,193,31,45,31,121,31,43,31,27,31,17,31,232,31,232,30,147,31,147,30,185,31,86,31,88,31,205,31,5,31,70,31,146,31,5,31,5,30,5,29,5,28,220,31,243,31,181,31,29,31,29,30,92,31,92,30,36,31,36,30,168,31,168,30,168,29,33,31,189,31,189,30,189,29,244,31,107,31,170,31,15,31,186,31,121,31,224,31,175,31,31,31,170,31,65,31,54,31,194,31,15,31,157,31,157,30,104,31,217,31,118,31,1,31,249,31,141,31,141,30,111,31,111,30,20,31,83,31,59,31,59,30,213,31,1,31,158,31,158,30,83,31,41,31,175,31,175,30,19,31,172,31,32,31,108,31,115,31,115,30,199,31,56,31,91,31,72,31,250,31,3,31,209,31,209,30,5,31,243,31,243,30,154,31,90,31,248,31,248,30,133,31,207,31,231,31,111,31,111,30,55,31,52,31,130,31,133,31,133,30,206,31,122,31,161,31,91,31,171,31,41,31,170,31,247,31,247,30,201,31,11,31,139,31,139,30,165,31,165,30,35,31,63,31,68,31,15,31,248,31,49,31,157,31,157,30,231,31,21,31,125,31,125,30,175,31,175,30,46,31,198,31,141,31,14,31,14,30,101,31,101,30,236,31,164,31,164,30,31,31,31,30,31,29,84,31,157,31,26,31,8,31,11,31,196,31,196,30,202,31,37,31,115,31,249,31,249,30,249,29,65,31,166,31,90,31,90,30,142,31,163,31,163,30,194,31,106,31,198,31,16,31,239,31,107,31,19,31,171,31,246,31,246,30,246,29,83,31,83,30,116,31,189,31,162,31,5,31,49,31,93,31,56,31,92,31,214,31,48,31,66,31,66,30,66,29,229,31,225,31,78,31,39,31,111,31,248,31,5,31,115,31,175,31,67,31,36,31,36,30,66,31,120,31,119,31,253,31,253,30,87,31,41,31,12,31,145,31,57,31,7,31,7,30,241,31,75,31,6,31,162,31,162,30,250,31,162,31,231,31,127,31,77,31,123,31,7,31,119,31,34,31,63,31,209,31,209,30,209,29,209,28,96,31,47,31,47,30,29,31,191,31,135,31,57,31,231,31,225,31,246,31,23,31,23,30,1,31,1,30,166,31,86,31,122,31,185,31,253,31,220,31,52,31,180,31,136,31,80,31,197,31,71,31,60,31,154,31,217,31,83,31,20,31,79,31,11,31,46,31,39,31,227,31,226,31,226,30,115,31,134,31,134,30,97,31,97,30,97,29,62,31,71,31,46,31,185,31,182,31,111,31,146,31,44,31,44,30,134,31,134,30,24,31,11,31,35,31,70,31,243,31,222,31,169,31,197,31,23,31,8,31,253,31,196,31,196,30,147,31,228,31,24,31,24,30,166,31,166,30,94,31,11,31,11,30,247,31,239,31,101,31,149,31,19,31,123,31,168,31,168,30,217,31,37,31,37,30,148,31,5,31,13,31,56,31,56,30,120,31,104,31,71,31,217,31,62,31,62,30,97,31,97,30,10,31,32,31,172,31,52,31,214,31,102,31,57,31,128,31,169,31,25,31,22,31,22,30,78,31,78,30,205,31,61,31,98,31,234,31,125,31,134,31,28,31,225,31,195,31,195,30,248,31,41,31,146,31,40,31,97,31,82,31,207,31,224,31,182,31,18,31,76,31,156,31,139,31,45,31,45,30,45,29,50,31,199,31,98,31,9,31,9,30,31,31,80,31,69,31,69,30,253,31,198,31,26,31,26,30,95,31,65,31,65,30,27,31,162,31,41,31,104,31,104,30,104,29,46,31,153,31,39,31,39,30,182,31,136,31,166,31,164,31,229,31,220,31,43,31,122,31,122,30,83,31,201,31,55,31,181,31,181,31,205,31,177,31,177,30,177,29,7,31,198,31,104,31,167,31,169,31,226,31,235,31,17,31,163,31,163,30,163,29,142,31,154,31,67,31,104,31,184,31,184,30,184,29,224,31,144,31,144,30,144,29,144,28,62,31,190,31,190,30,107,31,107,30,168,31,222,31,222,30,99,31,191,31,214,31,32,31,185,31,237,31,20,31,20,30,20,29,199,31,24,31,229,31,229,30,140,31,138,31,94,31,192,31,92,31,132,31,23,31,147,31,13,31,87,31,116,31,45,31,45,30,176,31,163,31,186,31,118,31,118,30,236,31,236,30,236,29,61,31,142,31,208,31,170,31,224,31,224,30,89,31,129,31,113,31,25,31,166,31,198,31,218,31,210,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
