-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_925 is
end project_tb_925;

architecture project_tb_arch_925 of project_tb_925 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 670;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (38,0,173,0,224,0,105,0,75,0,238,0,180,0,0,0,0,0,193,0,0,0,94,0,3,0,132,0,183,0,15,0,15,0,80,0,0,0,126,0,207,0,0,0,0,0,88,0,58,0,32,0,73,0,146,0,12,0,94,0,0,0,78,0,232,0,155,0,99,0,86,0,154,0,178,0,0,0,33,0,174,0,83,0,136,0,110,0,147,0,223,0,197,0,65,0,26,0,65,0,162,0,18,0,82,0,219,0,244,0,75,0,0,0,133,0,29,0,110,0,75,0,0,0,206,0,0,0,0,0,56,0,35,0,254,0,69,0,100,0,191,0,69,0,145,0,0,0,42,0,62,0,0,0,71,0,49,0,184,0,99,0,0,0,175,0,179,0,251,0,85,0,225,0,9,0,134,0,240,0,137,0,73,0,176,0,28,0,125,0,49,0,210,0,192,0,101,0,51,0,182,0,180,0,191,0,165,0,0,0,118,0,253,0,0,0,3,0,89,0,118,0,135,0,136,0,230,0,0,0,5,0,137,0,202,0,85,0,140,0,0,0,2,0,165,0,0,0,0,0,248,0,0,0,37,0,0,0,126,0,0,0,0,0,83,0,18,0,226,0,204,0,3,0,59,0,76,0,87,0,0,0,160,0,69,0,0,0,0,0,108,0,0,0,98,0,240,0,183,0,0,0,87,0,90,0,207,0,53,0,124,0,0,0,183,0,139,0,129,0,0,0,56,0,50,0,142,0,163,0,173,0,169,0,172,0,200,0,0,0,43,0,213,0,0,0,143,0,162,0,0,0,229,0,95,0,157,0,0,0,225,0,228,0,116,0,243,0,171,0,148,0,162,0,249,0,81,0,195,0,226,0,0,0,0,0,4,0,0,0,26,0,251,0,153,0,32,0,166,0,0,0,114,0,7,0,34,0,31,0,113,0,30,0,127,0,124,0,231,0,23,0,63,0,5,0,0,0,102,0,88,0,62,0,0,0,52,0,41,0,0,0,0,0,186,0,164,0,26,0,0,0,125,0,150,0,226,0,0,0,244,0,127,0,120,0,198,0,0,0,0,0,141,0,0,0,98,0,230,0,26,0,208,0,211,0,0,0,119,0,0,0,127,0,224,0,219,0,151,0,108,0,225,0,0,0,44,0,229,0,221,0,29,0,225,0,0,0,0,0,30,0,0,0,76,0,0,0,96,0,130,0,81,0,2,0,136,0,0,0,138,0,151,0,244,0,242,0,63,0,0,0,78,0,0,0,197,0,242,0,92,0,111,0,157,0,219,0,139,0,0,0,227,0,17,0,0,0,209,0,0,0,174,0,192,0,24,0,155,0,110,0,223,0,0,0,89,0,193,0,252,0,61,0,206,0,195,0,175,0,231,0,0,0,245,0,163,0,106,0,239,0,204,0,229,0,212,0,18,0,233,0,241,0,95,0,95,0,142,0,0,0,0,0,131,0,116,0,71,0,0,0,237,0,82,0,156,0,210,0,182,0,246,0,193,0,222,0,126,0,134,0,251,0,156,0,68,0,243,0,133,0,0,0,111,0,118,0,237,0,251,0,203,0,203,0,222,0,47,0,132,0,0,0,198,0,138,0,239,0,93,0,163,0,176,0,145,0,101,0,147,0,0,0,38,0,14,0,144,0,0,0,78,0,90,0,187,0,251,0,147,0,0,0,131,0,110,0,0,0,70,0,0,0,20,0,209,0,0,0,141,0,37,0,76,0,53,0,241,0,0,0,122,0,230,0,0,0,60,0,0,0,0,0,112,0,74,0,238,0,36,0,2,0,20,0,59,0,0,0,206,0,0,0,138,0,0,0,46,0,0,0,59,0,229,0,236,0,19,0,57,0,158,0,0,0,51,0,71,0,2,0,142,0,3,0,0,0,71,0,181,0,68,0,240,0,253,0,0,0,245,0,60,0,41,0,207,0,150,0,229,0,205,0,0,0,0,0,56,0,168,0,248,0,120,0,196,0,150,0,146,0,181,0,118,0,196,0,42,0,145,0,18,0,213,0,11,0,161,0,0,0,99,0,201,0,204,0,0,0,227,0,209,0,128,0,1,0,0,0,0,0,131,0,203,0,0,0,227,0,0,0,0,0,209,0,0,0,89,0,255,0,211,0,18,0,33,0,81,0,151,0,195,0,72,0,225,0,214,0,248,0,0,0,188,0,0,0,144,0,0,0,0,0,191,0,10,0,91,0,177,0,26,0,61,0,124,0,152,0,0,0,226,0,161,0,171,0,40,0,139,0,9,0,145,0,85,0,10,0,155,0,0,0,8,0,185,0,48,0,111,0,183,0,116,0,0,0,53,0,63,0,0,0,71,0,48,0,185,0,145,0,0,0,64,0,235,0,248,0,182,0,0,0,209,0,195,0,181,0,145,0,219,0,220,0,53,0,155,0,22,0,47,0,128,0,0,0,186,0,66,0,243,0,214,0,172,0,203,0,57,0,84,0,0,0,42,0,40,0,108,0,0,0,195,0,0,0,202,0,10,0,41,0,201,0,38,0,247,0,247,0,128,0,180,0,114,0,33,0,0,0,35,0,197,0,158,0,168,0,55,0,0,0,0,0,0,0,46,0,86,0,239,0,72,0,216,0,0,0,164,0,138,0,209,0,23,0,113,0,8,0,227,0,42,0,4,0,0,0,171,0,0,0,0,0,254,0,139,0,225,0,95,0,32,0,117,0,246,0,205,0,155,0,38,0,161,0,0,0,183,0,0,0,131,0,113,0,97,0,0,0,0,0,227,0,47,0,224,0,47,0,57,0,0,0,81,0,0,0,119,0,40,0,186,0,0,0,224,0,126,0,245,0,209,0,122,0,89,0,79,0,192,0,248,0,145,0,0,0,0,0,49,0,0,0,120,0,132,0,236,0,87,0,160,0,58,0,6,0,0,0,196,0,220,0,112,0,241,0,237,0,0,0,155,0,144,0,191,0,0,0,72,0,105,0,174,0,188,0,182,0,54,0,219,0,0,0,136,0,11,0,0,0,0,0,209,0,206,0);
signal scenario_full  : scenario_type := (38,31,173,31,224,31,105,31,75,31,238,31,180,31,180,30,180,29,193,31,193,30,94,31,3,31,132,31,183,31,15,31,15,31,80,31,80,30,126,31,207,31,207,30,207,29,88,31,58,31,32,31,73,31,146,31,12,31,94,31,94,30,78,31,232,31,155,31,99,31,86,31,154,31,178,31,178,30,33,31,174,31,83,31,136,31,110,31,147,31,223,31,197,31,65,31,26,31,65,31,162,31,18,31,82,31,219,31,244,31,75,31,75,30,133,31,29,31,110,31,75,31,75,30,206,31,206,30,206,29,56,31,35,31,254,31,69,31,100,31,191,31,69,31,145,31,145,30,42,31,62,31,62,30,71,31,49,31,184,31,99,31,99,30,175,31,179,31,251,31,85,31,225,31,9,31,134,31,240,31,137,31,73,31,176,31,28,31,125,31,49,31,210,31,192,31,101,31,51,31,182,31,180,31,191,31,165,31,165,30,118,31,253,31,253,30,3,31,89,31,118,31,135,31,136,31,230,31,230,30,5,31,137,31,202,31,85,31,140,31,140,30,2,31,165,31,165,30,165,29,248,31,248,30,37,31,37,30,126,31,126,30,126,29,83,31,18,31,226,31,204,31,3,31,59,31,76,31,87,31,87,30,160,31,69,31,69,30,69,29,108,31,108,30,98,31,240,31,183,31,183,30,87,31,90,31,207,31,53,31,124,31,124,30,183,31,139,31,129,31,129,30,56,31,50,31,142,31,163,31,173,31,169,31,172,31,200,31,200,30,43,31,213,31,213,30,143,31,162,31,162,30,229,31,95,31,157,31,157,30,225,31,228,31,116,31,243,31,171,31,148,31,162,31,249,31,81,31,195,31,226,31,226,30,226,29,4,31,4,30,26,31,251,31,153,31,32,31,166,31,166,30,114,31,7,31,34,31,31,31,113,31,30,31,127,31,124,31,231,31,23,31,63,31,5,31,5,30,102,31,88,31,62,31,62,30,52,31,41,31,41,30,41,29,186,31,164,31,26,31,26,30,125,31,150,31,226,31,226,30,244,31,127,31,120,31,198,31,198,30,198,29,141,31,141,30,98,31,230,31,26,31,208,31,211,31,211,30,119,31,119,30,127,31,224,31,219,31,151,31,108,31,225,31,225,30,44,31,229,31,221,31,29,31,225,31,225,30,225,29,30,31,30,30,76,31,76,30,96,31,130,31,81,31,2,31,136,31,136,30,138,31,151,31,244,31,242,31,63,31,63,30,78,31,78,30,197,31,242,31,92,31,111,31,157,31,219,31,139,31,139,30,227,31,17,31,17,30,209,31,209,30,174,31,192,31,24,31,155,31,110,31,223,31,223,30,89,31,193,31,252,31,61,31,206,31,195,31,175,31,231,31,231,30,245,31,163,31,106,31,239,31,204,31,229,31,212,31,18,31,233,31,241,31,95,31,95,31,142,31,142,30,142,29,131,31,116,31,71,31,71,30,237,31,82,31,156,31,210,31,182,31,246,31,193,31,222,31,126,31,134,31,251,31,156,31,68,31,243,31,133,31,133,30,111,31,118,31,237,31,251,31,203,31,203,31,222,31,47,31,132,31,132,30,198,31,138,31,239,31,93,31,163,31,176,31,145,31,101,31,147,31,147,30,38,31,14,31,144,31,144,30,78,31,90,31,187,31,251,31,147,31,147,30,131,31,110,31,110,30,70,31,70,30,20,31,209,31,209,30,141,31,37,31,76,31,53,31,241,31,241,30,122,31,230,31,230,30,60,31,60,30,60,29,112,31,74,31,238,31,36,31,2,31,20,31,59,31,59,30,206,31,206,30,138,31,138,30,46,31,46,30,59,31,229,31,236,31,19,31,57,31,158,31,158,30,51,31,71,31,2,31,142,31,3,31,3,30,71,31,181,31,68,31,240,31,253,31,253,30,245,31,60,31,41,31,207,31,150,31,229,31,205,31,205,30,205,29,56,31,168,31,248,31,120,31,196,31,150,31,146,31,181,31,118,31,196,31,42,31,145,31,18,31,213,31,11,31,161,31,161,30,99,31,201,31,204,31,204,30,227,31,209,31,128,31,1,31,1,30,1,29,131,31,203,31,203,30,227,31,227,30,227,29,209,31,209,30,89,31,255,31,211,31,18,31,33,31,81,31,151,31,195,31,72,31,225,31,214,31,248,31,248,30,188,31,188,30,144,31,144,30,144,29,191,31,10,31,91,31,177,31,26,31,61,31,124,31,152,31,152,30,226,31,161,31,171,31,40,31,139,31,9,31,145,31,85,31,10,31,155,31,155,30,8,31,185,31,48,31,111,31,183,31,116,31,116,30,53,31,63,31,63,30,71,31,48,31,185,31,145,31,145,30,64,31,235,31,248,31,182,31,182,30,209,31,195,31,181,31,145,31,219,31,220,31,53,31,155,31,22,31,47,31,128,31,128,30,186,31,66,31,243,31,214,31,172,31,203,31,57,31,84,31,84,30,42,31,40,31,108,31,108,30,195,31,195,30,202,31,10,31,41,31,201,31,38,31,247,31,247,31,128,31,180,31,114,31,33,31,33,30,35,31,197,31,158,31,168,31,55,31,55,30,55,29,55,28,46,31,86,31,239,31,72,31,216,31,216,30,164,31,138,31,209,31,23,31,113,31,8,31,227,31,42,31,4,31,4,30,171,31,171,30,171,29,254,31,139,31,225,31,95,31,32,31,117,31,246,31,205,31,155,31,38,31,161,31,161,30,183,31,183,30,131,31,113,31,97,31,97,30,97,29,227,31,47,31,224,31,47,31,57,31,57,30,81,31,81,30,119,31,40,31,186,31,186,30,224,31,126,31,245,31,209,31,122,31,89,31,79,31,192,31,248,31,145,31,145,30,145,29,49,31,49,30,120,31,132,31,236,31,87,31,160,31,58,31,6,31,6,30,196,31,220,31,112,31,241,31,237,31,237,30,155,31,144,31,191,31,191,30,72,31,105,31,174,31,188,31,182,31,54,31,219,31,219,30,136,31,11,31,11,30,11,29,209,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
