-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 894;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,0,0,228,0,221,0,203,0,228,0,78,0,0,0,40,0,0,0,97,0,8,0,80,0,7,0,91,0,181,0,20,0,166,0,111,0,107,0,64,0,215,0,199,0,42,0,229,0,0,0,0,0,111,0,213,0,87,0,152,0,231,0,75,0,0,0,146,0,0,0,0,0,62,0,90,0,89,0,232,0,94,0,37,0,0,0,142,0,179,0,136,0,0,0,186,0,0,0,47,0,99,0,36,0,120,0,47,0,132,0,37,0,0,0,241,0,0,0,102,0,83,0,0,0,143,0,84,0,155,0,240,0,180,0,189,0,24,0,17,0,184,0,61,0,231,0,0,0,57,0,187,0,158,0,212,0,0,0,164,0,0,0,90,0,17,0,199,0,223,0,106,0,136,0,0,0,0,0,37,0,157,0,233,0,0,0,233,0,92,0,255,0,87,0,2,0,152,0,102,0,82,0,169,0,0,0,169,0,6,0,168,0,158,0,0,0,234,0,99,0,61,0,177,0,0,0,177,0,246,0,0,0,139,0,1,0,43,0,170,0,155,0,38,0,72,0,0,0,214,0,0,0,191,0,163,0,101,0,199,0,154,0,69,0,35,0,43,0,45,0,0,0,0,0,0,0,0,0,117,0,0,0,209,0,168,0,188,0,148,0,0,0,134,0,225,0,136,0,0,0,29,0,226,0,240,0,229,0,148,0,178,0,48,0,79,0,194,0,0,0,184,0,0,0,46,0,99,0,91,0,238,0,0,0,172,0,42,0,31,0,160,0,205,0,86,0,188,0,0,0,187,0,149,0,0,0,216,0,132,0,28,0,15,0,84,0,118,0,195,0,99,0,190,0,213,0,16,0,144,0,3,0,133,0,210,0,0,0,43,0,101,0,42,0,114,0,23,0,53,0,228,0,214,0,159,0,0,0,133,0,0,0,58,0,0,0,38,0,36,0,17,0,0,0,0,0,157,0,58,0,0,0,107,0,51,0,15,0,200,0,241,0,0,0,62,0,0,0,27,0,0,0,19,0,222,0,136,0,0,0,155,0,96,0,171,0,155,0,163,0,0,0,16,0,24,0,141,0,0,0,0,0,143,0,33,0,50,0,101,0,54,0,82,0,211,0,182,0,249,0,206,0,109,0,221,0,69,0,115,0,18,0,204,0,0,0,232,0,121,0,251,0,176,0,37,0,0,0,26,0,183,0,129,0,73,0,190,0,195,0,201,0,102,0,0,0,254,0,0,0,82,0,73,0,23,0,71,0,223,0,0,0,0,0,30,0,150,0,113,0,195,0,3,0,70,0,242,0,79,0,41,0,238,0,0,0,35,0,218,0,57,0,138,0,213,0,0,0,8,0,0,0,239,0,66,0,0,0,106,0,149,0,170,0,10,0,147,0,53,0,26,0,234,0,102,0,52,0,80,0,5,0,191,0,116,0,209,0,154,0,98,0,198,0,152,0,213,0,175,0,64,0,160,0,110,0,249,0,104,0,248,0,9,0,0,0,0,0,219,0,104,0,0,0,135,0,131,0,241,0,81,0,0,0,57,0,26,0,151,0,161,0,101,0,242,0,55,0,90,0,0,0,154,0,0,0,0,0,101,0,25,0,0,0,142,0,224,0,134,0,192,0,220,0,129,0,252,0,22,0,142,0,230,0,192,0,192,0,63,0,166,0,57,0,0,0,0,0,24,0,0,0,230,0,105,0,152,0,248,0,76,0,187,0,244,0,213,0,201,0,164,0,47,0,0,0,188,0,98,0,120,0,241,0,0,0,230,0,71,0,162,0,9,0,93,0,9,0,95,0,0,0,100,0,0,0,55,0,217,0,39,0,37,0,0,0,0,0,108,0,0,0,224,0,59,0,49,0,23,0,13,0,0,0,21,0,9,0,100,0,56,0,195,0,223,0,122,0,35,0,228,0,0,0,105,0,74,0,248,0,0,0,0,0,71,0,67,0,226,0,32,0,130,0,160,0,0,0,0,0,0,0,154,0,0,0,0,0,0,0,166,0,155,0,82,0,0,0,0,0,219,0,0,0,0,0,17,0,69,0,58,0,0,0,118,0,187,0,168,0,14,0,87,0,164,0,137,0,113,0,141,0,247,0,0,0,100,0,232,0,150,0,4,0,243,0,208,0,61,0,0,0,45,0,251,0,102,0,192,0,95,0,151,0,0,0,183,0,13,0,49,0,181,0,179,0,167,0,238,0,0,0,251,0,0,0,77,0,195,0,135,0,225,0,75,0,243,0,162,0,22,0,174,0,23,0,117,0,216,0,239,0,132,0,178,0,0,0,64,0,77,0,48,0,113,0,54,0,136,0,112,0,0,0,77,0,101,0,1,0,0,0,200,0,177,0,133,0,231,0,5,0,225,0,10,0,13,0,68,0,201,0,215,0,254,0,0,0,0,0,0,0,132,0,94,0,241,0,165,0,153,0,193,0,115,0,223,0,73,0,117,0,167,0,0,0,0,0,80,0,249,0,165,0,61,0,103,0,151,0,157,0,59,0,0,0,56,0,24,0,43,0,13,0,187,0,82,0,47,0,59,0,197,0,156,0,0,0,199,0,114,0,135,0,216,0,148,0,223,0,162,0,0,0,9,0,221,0,204,0,97,0,10,0,0,0,224,0,0,0,27,0,0,0,220,0,87,0,134,0,247,0,0,0,28,0,239,0,114,0,28,0,8,0,37,0,105,0,161,0,201,0,72,0,139,0,255,0,0,0,133,0,211,0,250,0,79,0,219,0,0,0,239,0,227,0,83,0,249,0,222,0,0,0,72,0,0,0,0,0,0,0,138,0,115,0,56,0,0,0,43,0,65,0,155,0,206,0,0,0,106,0,243,0,240,0,90,0,195,0,0,0,40,0,151,0,225,0,138,0,0,0,13,0,173,0,148,0,101,0,222,0,144,0,23,0,0,0,0,0,192,0,0,0,221,0,254,0,111,0,25,0,0,0,12,0,221,0,211,0,37,0,183,0,43,0,194,0,83,0,0,0,118,0,199,0,5,0,0,0,212,0,181,0,13,0,225,0,79,0,106,0,253,0,96,0,0,0,233,0,192,0,41,0,144,0,71,0,48,0,51,0,199,0,10,0,122,0,44,0,49,0,0,0,167,0,177,0,213,0,176,0,88,0,0,0,200,0,133,0,170,0,22,0,214,0,175,0,78,0,226,0,0,0,0,0,39,0,209,0,143,0,57,0,33,0,240,0,193,0,20,0,165,0,0,0,188,0,153,0,88,0,0,0,5,0,9,0,178,0,32,0,167,0,102,0,235,0,136,0,0,0,73,0,28,0,49,0,201,0,222,0,0,0,87,0,67,0,219,0,0,0,56,0,138,0,254,0,143,0,119,0,180,0,0,0,4,0,55,0,0,0,231,0,231,0,212,0,85,0,83,0,188,0,117,0,205,0,0,0,105,0,0,0,157,0,0,0,0,0,62,0,114,0,72,0,0,0,180,0,213,0,105,0,211,0,0,0,246,0,117,0,135,0,160,0,0,0,246,0,0,0,228,0,69,0,188,0,0,0,223,0,62,0,83,0,219,0,0,0,39,0,127,0,0,0,0,0,50,0,239,0,0,0,0,0,229,0,53,0,115,0,144,0,108,0,187,0,254,0,0,0,0,0,63,0,182,0,0,0,68,0,0,0,19,0,240,0,49,0,0,0,109,0,106,0,171,0,0,0,38,0,9,0,203,0,0,0,222,0,137,0,55,0,15,0,77,0,93,0,0,0,128,0,168,0,89,0,38,0,141,0,179,0,0,0,0,0,136,0,246,0,7,0,179,0,157,0,102,0,152,0,180,0,23,0,39,0,4,0,0,0,0,0,144,0,174,0,61,0,70,0,0,0,205,0,193,0,87,0,178,0,193,0,18,0,173,0,158,0,0,0,188,0,38,0,159,0,234,0,17,0,137,0,214,0,198,0,249,0,0,0,0,0,236,0,51,0,187,0,38,0,129,0,162,0,152,0,77,0,0,0,0,0,145,0,0,0,0,0,0,0,249,0,56,0);
signal scenario_full  : scenario_type := (232,31,232,30,228,31,221,31,203,31,228,31,78,31,78,30,40,31,40,30,97,31,8,31,80,31,7,31,91,31,181,31,20,31,166,31,111,31,107,31,64,31,215,31,199,31,42,31,229,31,229,30,229,29,111,31,213,31,87,31,152,31,231,31,75,31,75,30,146,31,146,30,146,29,62,31,90,31,89,31,232,31,94,31,37,31,37,30,142,31,179,31,136,31,136,30,186,31,186,30,47,31,99,31,36,31,120,31,47,31,132,31,37,31,37,30,241,31,241,30,102,31,83,31,83,30,143,31,84,31,155,31,240,31,180,31,189,31,24,31,17,31,184,31,61,31,231,31,231,30,57,31,187,31,158,31,212,31,212,30,164,31,164,30,90,31,17,31,199,31,223,31,106,31,136,31,136,30,136,29,37,31,157,31,233,31,233,30,233,31,92,31,255,31,87,31,2,31,152,31,102,31,82,31,169,31,169,30,169,31,6,31,168,31,158,31,158,30,234,31,99,31,61,31,177,31,177,30,177,31,246,31,246,30,139,31,1,31,43,31,170,31,155,31,38,31,72,31,72,30,214,31,214,30,191,31,163,31,101,31,199,31,154,31,69,31,35,31,43,31,45,31,45,30,45,29,45,28,45,27,117,31,117,30,209,31,168,31,188,31,148,31,148,30,134,31,225,31,136,31,136,30,29,31,226,31,240,31,229,31,148,31,178,31,48,31,79,31,194,31,194,30,184,31,184,30,46,31,99,31,91,31,238,31,238,30,172,31,42,31,31,31,160,31,205,31,86,31,188,31,188,30,187,31,149,31,149,30,216,31,132,31,28,31,15,31,84,31,118,31,195,31,99,31,190,31,213,31,16,31,144,31,3,31,133,31,210,31,210,30,43,31,101,31,42,31,114,31,23,31,53,31,228,31,214,31,159,31,159,30,133,31,133,30,58,31,58,30,38,31,36,31,17,31,17,30,17,29,157,31,58,31,58,30,107,31,51,31,15,31,200,31,241,31,241,30,62,31,62,30,27,31,27,30,19,31,222,31,136,31,136,30,155,31,96,31,171,31,155,31,163,31,163,30,16,31,24,31,141,31,141,30,141,29,143,31,33,31,50,31,101,31,54,31,82,31,211,31,182,31,249,31,206,31,109,31,221,31,69,31,115,31,18,31,204,31,204,30,232,31,121,31,251,31,176,31,37,31,37,30,26,31,183,31,129,31,73,31,190,31,195,31,201,31,102,31,102,30,254,31,254,30,82,31,73,31,23,31,71,31,223,31,223,30,223,29,30,31,150,31,113,31,195,31,3,31,70,31,242,31,79,31,41,31,238,31,238,30,35,31,218,31,57,31,138,31,213,31,213,30,8,31,8,30,239,31,66,31,66,30,106,31,149,31,170,31,10,31,147,31,53,31,26,31,234,31,102,31,52,31,80,31,5,31,191,31,116,31,209,31,154,31,98,31,198,31,152,31,213,31,175,31,64,31,160,31,110,31,249,31,104,31,248,31,9,31,9,30,9,29,219,31,104,31,104,30,135,31,131,31,241,31,81,31,81,30,57,31,26,31,151,31,161,31,101,31,242,31,55,31,90,31,90,30,154,31,154,30,154,29,101,31,25,31,25,30,142,31,224,31,134,31,192,31,220,31,129,31,252,31,22,31,142,31,230,31,192,31,192,31,63,31,166,31,57,31,57,30,57,29,24,31,24,30,230,31,105,31,152,31,248,31,76,31,187,31,244,31,213,31,201,31,164,31,47,31,47,30,188,31,98,31,120,31,241,31,241,30,230,31,71,31,162,31,9,31,93,31,9,31,95,31,95,30,100,31,100,30,55,31,217,31,39,31,37,31,37,30,37,29,108,31,108,30,224,31,59,31,49,31,23,31,13,31,13,30,21,31,9,31,100,31,56,31,195,31,223,31,122,31,35,31,228,31,228,30,105,31,74,31,248,31,248,30,248,29,71,31,67,31,226,31,32,31,130,31,160,31,160,30,160,29,160,28,154,31,154,30,154,29,154,28,166,31,155,31,82,31,82,30,82,29,219,31,219,30,219,29,17,31,69,31,58,31,58,30,118,31,187,31,168,31,14,31,87,31,164,31,137,31,113,31,141,31,247,31,247,30,100,31,232,31,150,31,4,31,243,31,208,31,61,31,61,30,45,31,251,31,102,31,192,31,95,31,151,31,151,30,183,31,13,31,49,31,181,31,179,31,167,31,238,31,238,30,251,31,251,30,77,31,195,31,135,31,225,31,75,31,243,31,162,31,22,31,174,31,23,31,117,31,216,31,239,31,132,31,178,31,178,30,64,31,77,31,48,31,113,31,54,31,136,31,112,31,112,30,77,31,101,31,1,31,1,30,200,31,177,31,133,31,231,31,5,31,225,31,10,31,13,31,68,31,201,31,215,31,254,31,254,30,254,29,254,28,132,31,94,31,241,31,165,31,153,31,193,31,115,31,223,31,73,31,117,31,167,31,167,30,167,29,80,31,249,31,165,31,61,31,103,31,151,31,157,31,59,31,59,30,56,31,24,31,43,31,13,31,187,31,82,31,47,31,59,31,197,31,156,31,156,30,199,31,114,31,135,31,216,31,148,31,223,31,162,31,162,30,9,31,221,31,204,31,97,31,10,31,10,30,224,31,224,30,27,31,27,30,220,31,87,31,134,31,247,31,247,30,28,31,239,31,114,31,28,31,8,31,37,31,105,31,161,31,201,31,72,31,139,31,255,31,255,30,133,31,211,31,250,31,79,31,219,31,219,30,239,31,227,31,83,31,249,31,222,31,222,30,72,31,72,30,72,29,72,28,138,31,115,31,56,31,56,30,43,31,65,31,155,31,206,31,206,30,106,31,243,31,240,31,90,31,195,31,195,30,40,31,151,31,225,31,138,31,138,30,13,31,173,31,148,31,101,31,222,31,144,31,23,31,23,30,23,29,192,31,192,30,221,31,254,31,111,31,25,31,25,30,12,31,221,31,211,31,37,31,183,31,43,31,194,31,83,31,83,30,118,31,199,31,5,31,5,30,212,31,181,31,13,31,225,31,79,31,106,31,253,31,96,31,96,30,233,31,192,31,41,31,144,31,71,31,48,31,51,31,199,31,10,31,122,31,44,31,49,31,49,30,167,31,177,31,213,31,176,31,88,31,88,30,200,31,133,31,170,31,22,31,214,31,175,31,78,31,226,31,226,30,226,29,39,31,209,31,143,31,57,31,33,31,240,31,193,31,20,31,165,31,165,30,188,31,153,31,88,31,88,30,5,31,9,31,178,31,32,31,167,31,102,31,235,31,136,31,136,30,73,31,28,31,49,31,201,31,222,31,222,30,87,31,67,31,219,31,219,30,56,31,138,31,254,31,143,31,119,31,180,31,180,30,4,31,55,31,55,30,231,31,231,31,212,31,85,31,83,31,188,31,117,31,205,31,205,30,105,31,105,30,157,31,157,30,157,29,62,31,114,31,72,31,72,30,180,31,213,31,105,31,211,31,211,30,246,31,117,31,135,31,160,31,160,30,246,31,246,30,228,31,69,31,188,31,188,30,223,31,62,31,83,31,219,31,219,30,39,31,127,31,127,30,127,29,50,31,239,31,239,30,239,29,229,31,53,31,115,31,144,31,108,31,187,31,254,31,254,30,254,29,63,31,182,31,182,30,68,31,68,30,19,31,240,31,49,31,49,30,109,31,106,31,171,31,171,30,38,31,9,31,203,31,203,30,222,31,137,31,55,31,15,31,77,31,93,31,93,30,128,31,168,31,89,31,38,31,141,31,179,31,179,30,179,29,136,31,246,31,7,31,179,31,157,31,102,31,152,31,180,31,23,31,39,31,4,31,4,30,4,29,144,31,174,31,61,31,70,31,70,30,205,31,193,31,87,31,178,31,193,31,18,31,173,31,158,31,158,30,188,31,38,31,159,31,234,31,17,31,137,31,214,31,198,31,249,31,249,30,249,29,236,31,51,31,187,31,38,31,129,31,162,31,152,31,77,31,77,30,77,29,145,31,145,30,145,29,145,28,249,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
