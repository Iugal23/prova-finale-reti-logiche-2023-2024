-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_260 is
end project_tb_260;

architecture project_tb_arch_260 of project_tb_260 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 627;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (33,0,197,0,115,0,83,0,56,0,210,0,0,0,90,0,0,0,122,0,154,0,243,0,121,0,235,0,0,0,26,0,0,0,67,0,116,0,0,0,0,0,131,0,32,0,133,0,65,0,206,0,87,0,0,0,63,0,7,0,124,0,42,0,210,0,152,0,58,0,0,0,139,0,44,0,6,0,45,0,164,0,103,0,0,0,152,0,54,0,0,0,69,0,91,0,152,0,206,0,36,0,0,0,171,0,0,0,53,0,195,0,177,0,177,0,158,0,0,0,0,0,0,0,210,0,192,0,211,0,0,0,235,0,91,0,149,0,115,0,180,0,242,0,3,0,206,0,218,0,22,0,179,0,211,0,0,0,116,0,170,0,229,0,0,0,156,0,166,0,165,0,108,0,148,0,166,0,32,0,152,0,82,0,17,0,161,0,165,0,0,0,0,0,0,0,112,0,163,0,235,0,254,0,27,0,0,0,0,0,62,0,190,0,199,0,177,0,177,0,179,0,0,0,87,0,0,0,13,0,246,0,210,0,254,0,83,0,220,0,136,0,97,0,47,0,21,0,145,0,48,0,34,0,8,0,0,0,0,0,242,0,22,0,0,0,84,0,35,0,214,0,194,0,162,0,115,0,243,0,50,0,69,0,194,0,177,0,237,0,167,0,0,0,41,0,0,0,146,0,163,0,216,0,195,0,252,0,46,0,241,0,118,0,19,0,73,0,233,0,232,0,138,0,0,0,26,0,218,0,163,0,38,0,217,0,159,0,111,0,54,0,59,0,246,0,220,0,125,0,0,0,88,0,79,0,127,0,118,0,0,0,0,0,149,0,70,0,0,0,186,0,0,0,202,0,105,0,80,0,30,0,241,0,0,0,94,0,21,0,7,0,0,0,0,0,136,0,99,0,249,0,152,0,181,0,65,0,248,0,0,0,86,0,0,0,106,0,44,0,53,0,221,0,95,0,49,0,139,0,0,0,154,0,122,0,9,0,117,0,149,0,174,0,180,0,0,0,253,0,127,0,16,0,132,0,174,0,0,0,127,0,179,0,148,0,20,0,19,0,120,0,229,0,0,0,57,0,26,0,200,0,201,0,133,0,0,0,0,0,218,0,2,0,105,0,44,0,0,0,149,0,125,0,25,0,0,0,80,0,173,0,0,0,151,0,0,0,217,0,0,0,153,0,138,0,0,0,48,0,0,0,20,0,215,0,64,0,0,0,234,0,0,0,245,0,172,0,9,0,142,0,0,0,69,0,0,0,0,0,111,0,154,0,0,0,50,0,131,0,109,0,0,0,138,0,0,0,228,0,0,0,0,0,6,0,234,0,92,0,116,0,160,0,0,0,117,0,0,0,25,0,174,0,238,0,179,0,118,0,115,0,133,0,252,0,8,0,174,0,27,0,77,0,222,0,91,0,0,0,125,0,69,0,0,0,170,0,75,0,220,0,0,0,101,0,174,0,88,0,95,0,122,0,56,0,8,0,188,0,226,0,123,0,81,0,180,0,194,0,0,0,104,0,183,0,0,0,10,0,67,0,54,0,106,0,0,0,125,0,91,0,2,0,111,0,203,0,200,0,59,0,108,0,94,0,57,0,88,0,155,0,127,0,9,0,88,0,215,0,207,0,132,0,11,0,215,0,30,0,62,0,100,0,187,0,0,0,145,0,187,0,198,0,0,0,6,0,50,0,134,0,0,0,184,0,67,0,173,0,30,0,226,0,240,0,50,0,192,0,84,0,54,0,16,0,97,0,81,0,31,0,220,0,208,0,96,0,188,0,182,0,195,0,67,0,0,0,186,0,0,0,112,0,0,0,0,0,138,0,142,0,0,0,146,0,0,0,49,0,4,0,0,0,228,0,0,0,88,0,2,0,58,0,153,0,30,0,102,0,231,0,195,0,10,0,106,0,2,0,10,0,102,0,110,0,206,0,63,0,154,0,15,0,0,0,0,0,0,0,223,0,208,0,113,0,41,0,180,0,119,0,210,0,233,0,2,0,54,0,52,0,135,0,52,0,22,0,52,0,226,0,104,0,136,0,189,0,0,0,0,0,72,0,0,0,62,0,120,0,124,0,37,0,99,0,0,0,0,0,68,0,212,0,79,0,201,0,72,0,0,0,0,0,110,0,86,0,0,0,172,0,219,0,236,0,154,0,64,0,226,0,244,0,0,0,201,0,141,0,138,0,0,0,195,0,0,0,224,0,0,0,39,0,115,0,66,0,0,0,76,0,139,0,105,0,122,0,0,0,96,0,122,0,214,0,78,0,227,0,252,0,85,0,21,0,17,0,0,0,71,0,131,0,233,0,61,0,126,0,70,0,45,0,0,0,183,0,0,0,216,0,155,0,0,0,100,0,64,0,207,0,43,0,0,0,217,0,0,0,25,0,181,0,0,0,109,0,1,0,129,0,23,0,102,0,98,0,0,0,99,0,101,0,0,0,0,0,76,0,229,0,0,0,226,0,99,0,198,0,0,0,254,0,204,0,54,0,182,0,238,0,0,0,103,0,16,0,255,0,121,0,239,0,225,0,188,0,0,0,190,0,17,0,41,0,211,0,197,0,0,0,159,0,234,0,221,0,0,0,0,0,108,0,0,0,196,0,21,0,0,0,0,0,0,0,116,0,219,0,207,0,0,0,56,0,46,0,145,0,229,0,1,0,71,0,142,0,0,0,195,0,78,0,1,0,111,0,0,0,132,0,98,0,84,0,185,0,109,0,237,0,255,0,111,0,82,0,147,0,167,0,82,0,98,0,252,0,74,0,18,0,91,0,134,0,25,0,255,0,88,0,59,0,231,0,73,0,119,0,115,0,0,0);
signal scenario_full  : scenario_type := (33,31,197,31,115,31,83,31,56,31,210,31,210,30,90,31,90,30,122,31,154,31,243,31,121,31,235,31,235,30,26,31,26,30,67,31,116,31,116,30,116,29,131,31,32,31,133,31,65,31,206,31,87,31,87,30,63,31,7,31,124,31,42,31,210,31,152,31,58,31,58,30,139,31,44,31,6,31,45,31,164,31,103,31,103,30,152,31,54,31,54,30,69,31,91,31,152,31,206,31,36,31,36,30,171,31,171,30,53,31,195,31,177,31,177,31,158,31,158,30,158,29,158,28,210,31,192,31,211,31,211,30,235,31,91,31,149,31,115,31,180,31,242,31,3,31,206,31,218,31,22,31,179,31,211,31,211,30,116,31,170,31,229,31,229,30,156,31,166,31,165,31,108,31,148,31,166,31,32,31,152,31,82,31,17,31,161,31,165,31,165,30,165,29,165,28,112,31,163,31,235,31,254,31,27,31,27,30,27,29,62,31,190,31,199,31,177,31,177,31,179,31,179,30,87,31,87,30,13,31,246,31,210,31,254,31,83,31,220,31,136,31,97,31,47,31,21,31,145,31,48,31,34,31,8,31,8,30,8,29,242,31,22,31,22,30,84,31,35,31,214,31,194,31,162,31,115,31,243,31,50,31,69,31,194,31,177,31,237,31,167,31,167,30,41,31,41,30,146,31,163,31,216,31,195,31,252,31,46,31,241,31,118,31,19,31,73,31,233,31,232,31,138,31,138,30,26,31,218,31,163,31,38,31,217,31,159,31,111,31,54,31,59,31,246,31,220,31,125,31,125,30,88,31,79,31,127,31,118,31,118,30,118,29,149,31,70,31,70,30,186,31,186,30,202,31,105,31,80,31,30,31,241,31,241,30,94,31,21,31,7,31,7,30,7,29,136,31,99,31,249,31,152,31,181,31,65,31,248,31,248,30,86,31,86,30,106,31,44,31,53,31,221,31,95,31,49,31,139,31,139,30,154,31,122,31,9,31,117,31,149,31,174,31,180,31,180,30,253,31,127,31,16,31,132,31,174,31,174,30,127,31,179,31,148,31,20,31,19,31,120,31,229,31,229,30,57,31,26,31,200,31,201,31,133,31,133,30,133,29,218,31,2,31,105,31,44,31,44,30,149,31,125,31,25,31,25,30,80,31,173,31,173,30,151,31,151,30,217,31,217,30,153,31,138,31,138,30,48,31,48,30,20,31,215,31,64,31,64,30,234,31,234,30,245,31,172,31,9,31,142,31,142,30,69,31,69,30,69,29,111,31,154,31,154,30,50,31,131,31,109,31,109,30,138,31,138,30,228,31,228,30,228,29,6,31,234,31,92,31,116,31,160,31,160,30,117,31,117,30,25,31,174,31,238,31,179,31,118,31,115,31,133,31,252,31,8,31,174,31,27,31,77,31,222,31,91,31,91,30,125,31,69,31,69,30,170,31,75,31,220,31,220,30,101,31,174,31,88,31,95,31,122,31,56,31,8,31,188,31,226,31,123,31,81,31,180,31,194,31,194,30,104,31,183,31,183,30,10,31,67,31,54,31,106,31,106,30,125,31,91,31,2,31,111,31,203,31,200,31,59,31,108,31,94,31,57,31,88,31,155,31,127,31,9,31,88,31,215,31,207,31,132,31,11,31,215,31,30,31,62,31,100,31,187,31,187,30,145,31,187,31,198,31,198,30,6,31,50,31,134,31,134,30,184,31,67,31,173,31,30,31,226,31,240,31,50,31,192,31,84,31,54,31,16,31,97,31,81,31,31,31,220,31,208,31,96,31,188,31,182,31,195,31,67,31,67,30,186,31,186,30,112,31,112,30,112,29,138,31,142,31,142,30,146,31,146,30,49,31,4,31,4,30,228,31,228,30,88,31,2,31,58,31,153,31,30,31,102,31,231,31,195,31,10,31,106,31,2,31,10,31,102,31,110,31,206,31,63,31,154,31,15,31,15,30,15,29,15,28,223,31,208,31,113,31,41,31,180,31,119,31,210,31,233,31,2,31,54,31,52,31,135,31,52,31,22,31,52,31,226,31,104,31,136,31,189,31,189,30,189,29,72,31,72,30,62,31,120,31,124,31,37,31,99,31,99,30,99,29,68,31,212,31,79,31,201,31,72,31,72,30,72,29,110,31,86,31,86,30,172,31,219,31,236,31,154,31,64,31,226,31,244,31,244,30,201,31,141,31,138,31,138,30,195,31,195,30,224,31,224,30,39,31,115,31,66,31,66,30,76,31,139,31,105,31,122,31,122,30,96,31,122,31,214,31,78,31,227,31,252,31,85,31,21,31,17,31,17,30,71,31,131,31,233,31,61,31,126,31,70,31,45,31,45,30,183,31,183,30,216,31,155,31,155,30,100,31,64,31,207,31,43,31,43,30,217,31,217,30,25,31,181,31,181,30,109,31,1,31,129,31,23,31,102,31,98,31,98,30,99,31,101,31,101,30,101,29,76,31,229,31,229,30,226,31,99,31,198,31,198,30,254,31,204,31,54,31,182,31,238,31,238,30,103,31,16,31,255,31,121,31,239,31,225,31,188,31,188,30,190,31,17,31,41,31,211,31,197,31,197,30,159,31,234,31,221,31,221,30,221,29,108,31,108,30,196,31,21,31,21,30,21,29,21,28,116,31,219,31,207,31,207,30,56,31,46,31,145,31,229,31,1,31,71,31,142,31,142,30,195,31,78,31,1,31,111,31,111,30,132,31,98,31,84,31,185,31,109,31,237,31,255,31,111,31,82,31,147,31,167,31,82,31,98,31,252,31,74,31,18,31,91,31,134,31,25,31,255,31,88,31,59,31,231,31,73,31,119,31,115,31,115,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
