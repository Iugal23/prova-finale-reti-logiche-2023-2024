-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 993;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,143,0,200,0,0,0,49,0,188,0,31,0,50,0,0,0,94,0,113,0,0,0,116,0,99,0,38,0,20,0,11,0,0,0,165,0,0,0,138,0,192,0,181,0,205,0,0,0,44,0,0,0,229,0,170,0,68,0,16,0,187,0,4,0,0,0,209,0,181,0,0,0,36,0,0,0,112,0,108,0,202,0,221,0,243,0,0,0,0,0,35,0,0,0,106,0,203,0,0,0,63,0,15,0,4,0,66,0,0,0,134,0,0,0,69,0,245,0,60,0,90,0,152,0,163,0,165,0,68,0,154,0,0,0,0,0,20,0,20,0,0,0,0,0,0,0,0,0,156,0,94,0,90,0,0,0,127,0,95,0,50,0,170,0,110,0,0,0,0,0,244,0,175,0,123,0,110,0,138,0,155,0,140,0,0,0,244,0,218,0,0,0,207,0,0,0,197,0,4,0,0,0,0,0,190,0,139,0,239,0,36,0,164,0,0,0,0,0,209,0,26,0,85,0,172,0,0,0,62,0,26,0,129,0,114,0,225,0,243,0,93,0,159,0,100,0,214,0,236,0,0,0,0,0,0,0,88,0,196,0,178,0,208,0,22,0,132,0,226,0,0,0,51,0,16,0,230,0,76,0,0,0,134,0,20,0,243,0,181,0,207,0,115,0,131,0,197,0,0,0,167,0,7,0,0,0,171,0,229,0,0,0,201,0,15,0,210,0,0,0,180,0,244,0,208,0,94,0,0,0,178,0,0,0,3,0,204,0,3,0,136,0,123,0,128,0,210,0,0,0,0,0,0,0,0,0,143,0,231,0,55,0,60,0,52,0,65,0,121,0,0,0,167,0,0,0,122,0,159,0,122,0,178,0,253,0,118,0,108,0,0,0,187,0,132,0,24,0,0,0,225,0,122,0,186,0,122,0,57,0,0,0,210,0,0,0,48,0,134,0,89,0,177,0,242,0,111,0,215,0,0,0,243,0,249,0,71,0,158,0,20,0,0,0,189,0,36,0,132,0,69,0,183,0,72,0,0,0,222,0,171,0,233,0,112,0,110,0,195,0,0,0,0,0,0,0,223,0,5,0,89,0,212,0,48,0,29,0,167,0,121,0,0,0,82,0,160,0,117,0,196,0,254,0,0,0,180,0,40,0,177,0,181,0,100,0,166,0,115,0,134,0,129,0,131,0,0,0,15,0,0,0,137,0,67,0,206,0,0,0,73,0,25,0,5,0,0,0,39,0,107,0,80,0,117,0,255,0,47,0,0,0,126,0,23,0,220,0,81,0,16,0,214,0,74,0,226,0,36,0,104,0,0,0,50,0,201,0,0,0,193,0,131,0,240,0,0,0,72,0,98,0,157,0,37,0,124,0,233,0,231,0,29,0,101,0,120,0,82,0,0,0,202,0,182,0,150,0,0,0,175,0,32,0,0,0,235,0,187,0,98,0,94,0,77,0,196,0,60,0,0,0,185,0,40,0,0,0,0,0,191,0,253,0,78,0,75,0,59,0,66,0,102,0,217,0,90,0,79,0,178,0,0,0,0,0,142,0,53,0,96,0,106,0,63,0,73,0,166,0,0,0,133,0,0,0,194,0,186,0,4,0,111,0,0,0,231,0,146,0,0,0,0,0,0,0,0,0,194,0,102,0,0,0,208,0,0,0,238,0,146,0,70,0,76,0,198,0,248,0,63,0,0,0,5,0,34,0,141,0,245,0,187,0,252,0,228,0,117,0,0,0,172,0,64,0,33,0,0,0,135,0,38,0,0,0,247,0,44,0,204,0,70,0,0,0,91,0,119,0,146,0,0,0,97,0,41,0,214,0,0,0,94,0,135,0,147,0,239,0,2,0,232,0,61,0,175,0,0,0,0,0,222,0,0,0,212,0,15,0,74,0,0,0,28,0,216,0,183,0,217,0,95,0,80,0,179,0,248,0,62,0,117,0,0,0,165,0,8,0,0,0,7,0,238,0,235,0,2,0,0,0,39,0,37,0,240,0,120,0,0,0,216,0,119,0,156,0,0,0,0,0,122,0,96,0,87,0,112,0,123,0,0,0,229,0,65,0,116,0,189,0,17,0,178,0,168,0,0,0,10,0,56,0,58,0,117,0,33,0,149,0,17,0,0,0,5,0,54,0,0,0,37,0,223,0,20,0,159,0,0,0,220,0,220,0,200,0,0,0,149,0,60,0,33,0,189,0,0,0,91,0,18,0,124,0,227,0,7,0,107,0,0,0,179,0,47,0,120,0,183,0,126,0,40,0,101,0,111,0,197,0,69,0,152,0,0,0,0,0,156,0,0,0,192,0,229,0,193,0,218,0,63,0,217,0,0,0,0,0,92,0,79,0,117,0,210,0,241,0,50,0,32,0,86,0,179,0,61,0,192,0,117,0,3,0,177,0,63,0,191,0,175,0,85,0,141,0,0,0,209,0,0,0,178,0,50,0,33,0,33,0,8,0,0,0,0,0,254,0,117,0,0,0,245,0,202,0,107,0,68,0,10,0,218,0,248,0,146,0,65,0,17,0,41,0,0,0,37,0,121,0,0,0,75,0,0,0,248,0,0,0,224,0,108,0,8,0,22,0,62,0,74,0,133,0,161,0,218,0,0,0,0,0,158,0,223,0,184,0,38,0,29,0,0,0,250,0,154,0,251,0,75,0,156,0,18,0,112,0,134,0,0,0,63,0,90,0,149,0,152,0,0,0,234,0,194,0,172,0,0,0,0,0,6,0,83,0,0,0,186,0,121,0,0,0,175,0,88,0,34,0,78,0,53,0,11,0,157,0,184,0,4,0,195,0,0,0,168,0,80,0,0,0,212,0,0,0,0,0,0,0,19,0,194,0,83,0,0,0,85,0,30,0,19,0,201,0,251,0,15,0,0,0,124,0,200,0,93,0,0,0,77,0,165,0,176,0,104,0,80,0,253,0,32,0,195,0,55,0,101,0,177,0,0,0,29,0,196,0,0,0,0,0,151,0,61,0,0,0,17,0,0,0,121,0,174,0,47,0,0,0,29,0,0,0,0,0,57,0,178,0,92,0,0,0,95,0,0,0,193,0,45,0,87,0,196,0,46,0,108,0,0,0,125,0,226,0,0,0,221,0,127,0,68,0,231,0,41,0,142,0,0,0,225,0,118,0,0,0,0,0,14,0,0,0,0,0,248,0,216,0,201,0,153,0,0,0,0,0,36,0,25,0,120,0,105,0,78,0,190,0,149,0,136,0,118,0,242,0,158,0,0,0,83,0,163,0,223,0,211,0,214,0,156,0,0,0,0,0,189,0,14,0,254,0,0,0,63,0,138,0,56,0,0,0,220,0,0,0,88,0,99,0,96,0,163,0,20,0,0,0,0,0,0,0,124,0,0,0,0,0,0,0,231,0,0,0,126,0,34,0,199,0,134,0,0,0,220,0,64,0,202,0,192,0,0,0,128,0,155,0,215,0,5,0,97,0,76,0,191,0,50,0,0,0,0,0,121,0,88,0,0,0,251,0,58,0,167,0,159,0,121,0,163,0,175,0,0,0,51,0,0,0,0,0,0,0,146,0,173,0,80,0,165,0,15,0,47,0,24,0,134,0,180,0,81,0,41,0,229,0,168,0,0,0,95,0,22,0,62,0,85,0,12,0,13,0,221,0,242,0,0,0,0,0,20,0,57,0,42,0,241,0,57,0,84,0,51,0,92,0,63,0,119,0,251,0,4,0,50,0,152,0,77,0,241,0,69,0,50,0,196,0,0,0,144,0,234,0,238,0,0,0,157,0,228,0,68,0,128,0,52,0,42,0,9,0,152,0,208,0,2,0,3,0,0,0,0,0,91,0,49,0,185,0,65,0,177,0,0,0,60,0,97,0,180,0,115,0,221,0,212,0,185,0,27,0,71,0,201,0,175,0,0,0,0,0,36,0,244,0,0,0,248,0,0,0,218,0,156,0,151,0,139,0,57,0,44,0,167,0,189,0,54,0,99,0,0,0,19,0,23,0,109,0,191,0,111,0,84,0,0,0,175,0,69,0,192,0,0,0,144,0,93,0,0,0,30,0,150,0,133,0,148,0,161,0,0,0,38,0,214,0,155,0,81,0,155,0,73,0,114,0,170,0,167,0,248,0,39,0,204,0,76,0,177,0,0,0,174,0,147,0,0,0,0,0,239,0,221,0,126,0,146,0,18,0,44,0,138,0,79,0,255,0,202,0,129,0,32,0,204,0,204,0,217,0,19,0,0,0,229,0,189,0,74,0,212,0,0,0,215,0,166,0,208,0,213,0,0,0,102,0,59,0,0,0,222,0,252,0,89,0,201,0,0,0,154,0,170,0,250,0,250,0,16,0,0,0,239,0,114,0,0,0,228,0,43,0,0,0,111,0,156,0,0,0,106,0,217,0,0,0,103,0,188,0,103,0,248,0,159,0,0,0,0,0,0,0,0,0,142,0,236,0,18,0,34,0,0,0,88,0);
signal scenario_full  : scenario_type := (87,31,143,31,200,31,200,30,49,31,188,31,31,31,50,31,50,30,94,31,113,31,113,30,116,31,99,31,38,31,20,31,11,31,11,30,165,31,165,30,138,31,192,31,181,31,205,31,205,30,44,31,44,30,229,31,170,31,68,31,16,31,187,31,4,31,4,30,209,31,181,31,181,30,36,31,36,30,112,31,108,31,202,31,221,31,243,31,243,30,243,29,35,31,35,30,106,31,203,31,203,30,63,31,15,31,4,31,66,31,66,30,134,31,134,30,69,31,245,31,60,31,90,31,152,31,163,31,165,31,68,31,154,31,154,30,154,29,20,31,20,31,20,30,20,29,20,28,20,27,156,31,94,31,90,31,90,30,127,31,95,31,50,31,170,31,110,31,110,30,110,29,244,31,175,31,123,31,110,31,138,31,155,31,140,31,140,30,244,31,218,31,218,30,207,31,207,30,197,31,4,31,4,30,4,29,190,31,139,31,239,31,36,31,164,31,164,30,164,29,209,31,26,31,85,31,172,31,172,30,62,31,26,31,129,31,114,31,225,31,243,31,93,31,159,31,100,31,214,31,236,31,236,30,236,29,236,28,88,31,196,31,178,31,208,31,22,31,132,31,226,31,226,30,51,31,16,31,230,31,76,31,76,30,134,31,20,31,243,31,181,31,207,31,115,31,131,31,197,31,197,30,167,31,7,31,7,30,171,31,229,31,229,30,201,31,15,31,210,31,210,30,180,31,244,31,208,31,94,31,94,30,178,31,178,30,3,31,204,31,3,31,136,31,123,31,128,31,210,31,210,30,210,29,210,28,210,27,143,31,231,31,55,31,60,31,52,31,65,31,121,31,121,30,167,31,167,30,122,31,159,31,122,31,178,31,253,31,118,31,108,31,108,30,187,31,132,31,24,31,24,30,225,31,122,31,186,31,122,31,57,31,57,30,210,31,210,30,48,31,134,31,89,31,177,31,242,31,111,31,215,31,215,30,243,31,249,31,71,31,158,31,20,31,20,30,189,31,36,31,132,31,69,31,183,31,72,31,72,30,222,31,171,31,233,31,112,31,110,31,195,31,195,30,195,29,195,28,223,31,5,31,89,31,212,31,48,31,29,31,167,31,121,31,121,30,82,31,160,31,117,31,196,31,254,31,254,30,180,31,40,31,177,31,181,31,100,31,166,31,115,31,134,31,129,31,131,31,131,30,15,31,15,30,137,31,67,31,206,31,206,30,73,31,25,31,5,31,5,30,39,31,107,31,80,31,117,31,255,31,47,31,47,30,126,31,23,31,220,31,81,31,16,31,214,31,74,31,226,31,36,31,104,31,104,30,50,31,201,31,201,30,193,31,131,31,240,31,240,30,72,31,98,31,157,31,37,31,124,31,233,31,231,31,29,31,101,31,120,31,82,31,82,30,202,31,182,31,150,31,150,30,175,31,32,31,32,30,235,31,187,31,98,31,94,31,77,31,196,31,60,31,60,30,185,31,40,31,40,30,40,29,191,31,253,31,78,31,75,31,59,31,66,31,102,31,217,31,90,31,79,31,178,31,178,30,178,29,142,31,53,31,96,31,106,31,63,31,73,31,166,31,166,30,133,31,133,30,194,31,186,31,4,31,111,31,111,30,231,31,146,31,146,30,146,29,146,28,146,27,194,31,102,31,102,30,208,31,208,30,238,31,146,31,70,31,76,31,198,31,248,31,63,31,63,30,5,31,34,31,141,31,245,31,187,31,252,31,228,31,117,31,117,30,172,31,64,31,33,31,33,30,135,31,38,31,38,30,247,31,44,31,204,31,70,31,70,30,91,31,119,31,146,31,146,30,97,31,41,31,214,31,214,30,94,31,135,31,147,31,239,31,2,31,232,31,61,31,175,31,175,30,175,29,222,31,222,30,212,31,15,31,74,31,74,30,28,31,216,31,183,31,217,31,95,31,80,31,179,31,248,31,62,31,117,31,117,30,165,31,8,31,8,30,7,31,238,31,235,31,2,31,2,30,39,31,37,31,240,31,120,31,120,30,216,31,119,31,156,31,156,30,156,29,122,31,96,31,87,31,112,31,123,31,123,30,229,31,65,31,116,31,189,31,17,31,178,31,168,31,168,30,10,31,56,31,58,31,117,31,33,31,149,31,17,31,17,30,5,31,54,31,54,30,37,31,223,31,20,31,159,31,159,30,220,31,220,31,200,31,200,30,149,31,60,31,33,31,189,31,189,30,91,31,18,31,124,31,227,31,7,31,107,31,107,30,179,31,47,31,120,31,183,31,126,31,40,31,101,31,111,31,197,31,69,31,152,31,152,30,152,29,156,31,156,30,192,31,229,31,193,31,218,31,63,31,217,31,217,30,217,29,92,31,79,31,117,31,210,31,241,31,50,31,32,31,86,31,179,31,61,31,192,31,117,31,3,31,177,31,63,31,191,31,175,31,85,31,141,31,141,30,209,31,209,30,178,31,50,31,33,31,33,31,8,31,8,30,8,29,254,31,117,31,117,30,245,31,202,31,107,31,68,31,10,31,218,31,248,31,146,31,65,31,17,31,41,31,41,30,37,31,121,31,121,30,75,31,75,30,248,31,248,30,224,31,108,31,8,31,22,31,62,31,74,31,133,31,161,31,218,31,218,30,218,29,158,31,223,31,184,31,38,31,29,31,29,30,250,31,154,31,251,31,75,31,156,31,18,31,112,31,134,31,134,30,63,31,90,31,149,31,152,31,152,30,234,31,194,31,172,31,172,30,172,29,6,31,83,31,83,30,186,31,121,31,121,30,175,31,88,31,34,31,78,31,53,31,11,31,157,31,184,31,4,31,195,31,195,30,168,31,80,31,80,30,212,31,212,30,212,29,212,28,19,31,194,31,83,31,83,30,85,31,30,31,19,31,201,31,251,31,15,31,15,30,124,31,200,31,93,31,93,30,77,31,165,31,176,31,104,31,80,31,253,31,32,31,195,31,55,31,101,31,177,31,177,30,29,31,196,31,196,30,196,29,151,31,61,31,61,30,17,31,17,30,121,31,174,31,47,31,47,30,29,31,29,30,29,29,57,31,178,31,92,31,92,30,95,31,95,30,193,31,45,31,87,31,196,31,46,31,108,31,108,30,125,31,226,31,226,30,221,31,127,31,68,31,231,31,41,31,142,31,142,30,225,31,118,31,118,30,118,29,14,31,14,30,14,29,248,31,216,31,201,31,153,31,153,30,153,29,36,31,25,31,120,31,105,31,78,31,190,31,149,31,136,31,118,31,242,31,158,31,158,30,83,31,163,31,223,31,211,31,214,31,156,31,156,30,156,29,189,31,14,31,254,31,254,30,63,31,138,31,56,31,56,30,220,31,220,30,88,31,99,31,96,31,163,31,20,31,20,30,20,29,20,28,124,31,124,30,124,29,124,28,231,31,231,30,126,31,34,31,199,31,134,31,134,30,220,31,64,31,202,31,192,31,192,30,128,31,155,31,215,31,5,31,97,31,76,31,191,31,50,31,50,30,50,29,121,31,88,31,88,30,251,31,58,31,167,31,159,31,121,31,163,31,175,31,175,30,51,31,51,30,51,29,51,28,146,31,173,31,80,31,165,31,15,31,47,31,24,31,134,31,180,31,81,31,41,31,229,31,168,31,168,30,95,31,22,31,62,31,85,31,12,31,13,31,221,31,242,31,242,30,242,29,20,31,57,31,42,31,241,31,57,31,84,31,51,31,92,31,63,31,119,31,251,31,4,31,50,31,152,31,77,31,241,31,69,31,50,31,196,31,196,30,144,31,234,31,238,31,238,30,157,31,228,31,68,31,128,31,52,31,42,31,9,31,152,31,208,31,2,31,3,31,3,30,3,29,91,31,49,31,185,31,65,31,177,31,177,30,60,31,97,31,180,31,115,31,221,31,212,31,185,31,27,31,71,31,201,31,175,31,175,30,175,29,36,31,244,31,244,30,248,31,248,30,218,31,156,31,151,31,139,31,57,31,44,31,167,31,189,31,54,31,99,31,99,30,19,31,23,31,109,31,191,31,111,31,84,31,84,30,175,31,69,31,192,31,192,30,144,31,93,31,93,30,30,31,150,31,133,31,148,31,161,31,161,30,38,31,214,31,155,31,81,31,155,31,73,31,114,31,170,31,167,31,248,31,39,31,204,31,76,31,177,31,177,30,174,31,147,31,147,30,147,29,239,31,221,31,126,31,146,31,18,31,44,31,138,31,79,31,255,31,202,31,129,31,32,31,204,31,204,31,217,31,19,31,19,30,229,31,189,31,74,31,212,31,212,30,215,31,166,31,208,31,213,31,213,30,102,31,59,31,59,30,222,31,252,31,89,31,201,31,201,30,154,31,170,31,250,31,250,31,16,31,16,30,239,31,114,31,114,30,228,31,43,31,43,30,111,31,156,31,156,30,106,31,217,31,217,30,103,31,188,31,103,31,248,31,159,31,159,30,159,29,159,28,159,27,142,31,236,31,18,31,34,31,34,30,88,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
