-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 307;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (52,0,138,0,73,0,52,0,225,0,96,0,113,0,200,0,158,0,85,0,17,0,159,0,64,0,194,0,92,0,161,0,37,0,156,0,160,0,153,0,0,0,119,0,61,0,182,0,66,0,136,0,185,0,62,0,1,0,0,0,0,0,89,0,74,0,0,0,213,0,0,0,193,0,15,0,0,0,232,0,164,0,72,0,168,0,139,0,204,0,0,0,91,0,0,0,34,0,116,0,0,0,147,0,0,0,0,0,89,0,112,0,29,0,167,0,19,0,149,0,134,0,252,0,147,0,205,0,21,0,245,0,75,0,227,0,122,0,190,0,147,0,0,0,0,0,84,0,135,0,0,0,89,0,0,0,248,0,101,0,248,0,0,0,103,0,13,0,33,0,188,0,148,0,112,0,201,0,0,0,0,0,200,0,234,0,27,0,110,0,0,0,95,0,117,0,0,0,131,0,205,0,0,0,109,0,252,0,130,0,68,0,41,0,229,0,68,0,94,0,128,0,110,0,0,0,78,0,250,0,0,0,117,0,82,0,0,0,253,0,0,0,0,0,211,0,58,0,27,0,206,0,56,0,0,0,181,0,142,0,12,0,94,0,160,0,158,0,169,0,0,0,230,0,0,0,0,0,147,0,13,0,0,0,105,0,78,0,201,0,55,0,226,0,47,0,117,0,208,0,43,0,57,0,0,0,44,0,0,0,153,0,0,0,0,0,219,0,34,0,0,0,169,0,113,0,161,0,132,0,0,0,127,0,134,0,0,0,81,0,151,0,50,0,192,0,206,0,178,0,0,0,184,0,95,0,101,0,218,0,0,0,183,0,179,0,75,0,124,0,129,0,10,0,153,0,99,0,62,0,108,0,236,0,0,0,40,0,17,0,127,0,178,0,127,0,190,0,106,0,11,0,52,0,73,0,222,0,118,0,16,0,25,0,166,0,128,0,141,0,76,0,175,0,62,0,196,0,86,0,0,0,129,0,184,0,67,0,0,0,23,0,108,0,84,0,166,0,172,0,214,0,0,0,0,0,73,0,107,0,213,0,122,0,205,0,0,0,209,0,217,0,0,0,0,0,167,0,0,0,48,0,197,0,50,0,36,0,215,0,0,0,0,0,195,0,74,0,228,0,214,0,59,0,0,0,185,0,235,0,7,0,96,0,118,0,238,0,213,0,231,0,100,0,150,0,18,0,51,0,0,0,0,0,0,0,233,0,77,0,188,0,0,0,105,0,217,0,6,0,0,0,92,0,23,0,185,0,67,0,15,0,255,0,66,0,164,0,97,0,197,0,69,0,64,0,176,0,214,0,78,0,195,0,49,0,222,0,0,0,159,0,170,0,2,0,0,0,84,0,109,0,10,0,223,0,13,0,15,0,117,0,254,0);
signal scenario_full  : scenario_type := (52,31,138,31,73,31,52,31,225,31,96,31,113,31,200,31,158,31,85,31,17,31,159,31,64,31,194,31,92,31,161,31,37,31,156,31,160,31,153,31,153,30,119,31,61,31,182,31,66,31,136,31,185,31,62,31,1,31,1,30,1,29,89,31,74,31,74,30,213,31,213,30,193,31,15,31,15,30,232,31,164,31,72,31,168,31,139,31,204,31,204,30,91,31,91,30,34,31,116,31,116,30,147,31,147,30,147,29,89,31,112,31,29,31,167,31,19,31,149,31,134,31,252,31,147,31,205,31,21,31,245,31,75,31,227,31,122,31,190,31,147,31,147,30,147,29,84,31,135,31,135,30,89,31,89,30,248,31,101,31,248,31,248,30,103,31,13,31,33,31,188,31,148,31,112,31,201,31,201,30,201,29,200,31,234,31,27,31,110,31,110,30,95,31,117,31,117,30,131,31,205,31,205,30,109,31,252,31,130,31,68,31,41,31,229,31,68,31,94,31,128,31,110,31,110,30,78,31,250,31,250,30,117,31,82,31,82,30,253,31,253,30,253,29,211,31,58,31,27,31,206,31,56,31,56,30,181,31,142,31,12,31,94,31,160,31,158,31,169,31,169,30,230,31,230,30,230,29,147,31,13,31,13,30,105,31,78,31,201,31,55,31,226,31,47,31,117,31,208,31,43,31,57,31,57,30,44,31,44,30,153,31,153,30,153,29,219,31,34,31,34,30,169,31,113,31,161,31,132,31,132,30,127,31,134,31,134,30,81,31,151,31,50,31,192,31,206,31,178,31,178,30,184,31,95,31,101,31,218,31,218,30,183,31,179,31,75,31,124,31,129,31,10,31,153,31,99,31,62,31,108,31,236,31,236,30,40,31,17,31,127,31,178,31,127,31,190,31,106,31,11,31,52,31,73,31,222,31,118,31,16,31,25,31,166,31,128,31,141,31,76,31,175,31,62,31,196,31,86,31,86,30,129,31,184,31,67,31,67,30,23,31,108,31,84,31,166,31,172,31,214,31,214,30,214,29,73,31,107,31,213,31,122,31,205,31,205,30,209,31,217,31,217,30,217,29,167,31,167,30,48,31,197,31,50,31,36,31,215,31,215,30,215,29,195,31,74,31,228,31,214,31,59,31,59,30,185,31,235,31,7,31,96,31,118,31,238,31,213,31,231,31,100,31,150,31,18,31,51,31,51,30,51,29,51,28,233,31,77,31,188,31,188,30,105,31,217,31,6,31,6,30,92,31,23,31,185,31,67,31,15,31,255,31,66,31,164,31,97,31,197,31,69,31,64,31,176,31,214,31,78,31,195,31,49,31,222,31,222,30,159,31,170,31,2,31,2,30,84,31,109,31,10,31,223,31,13,31,15,31,117,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
