-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 534;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,0,0,41,0,12,0,239,0,96,0,209,0,48,0,109,0,88,0,254,0,131,0,253,0,12,0,0,0,0,0,0,0,52,0,132,0,14,0,50,0,52,0,59,0,0,0,216,0,211,0,0,0,3,0,169,0,170,0,68,0,85,0,102,0,22,0,184,0,0,0,151,0,42,0,6,0,19,0,126,0,236,0,187,0,181,0,154,0,239,0,27,0,250,0,10,0,111,0,7,0,71,0,218,0,48,0,203,0,70,0,0,0,66,0,236,0,66,0,216,0,114,0,156,0,210,0,183,0,0,0,89,0,10,0,93,0,238,0,244,0,10,0,0,0,143,0,4,0,172,0,11,0,73,0,114,0,62,0,20,0,135,0,19,0,66,0,168,0,97,0,194,0,0,0,144,0,0,0,63,0,162,0,207,0,190,0,160,0,161,0,79,0,0,0,194,0,106,0,206,0,81,0,206,0,61,0,229,0,169,0,164,0,0,0,15,0,139,0,33,0,0,0,247,0,177,0,233,0,227,0,0,0,203,0,172,0,180,0,71,0,215,0,8,0,120,0,100,0,31,0,84,0,0,0,252,0,0,0,227,0,84,0,195,0,0,0,111,0,112,0,170,0,217,0,191,0,123,0,42,0,0,0,119,0,202,0,97,0,181,0,112,0,148,0,166,0,133,0,16,0,0,0,0,0,62,0,88,0,0,0,135,0,179,0,123,0,178,0,80,0,0,0,144,0,103,0,9,0,215,0,0,0,105,0,125,0,219,0,238,0,92,0,156,0,237,0,116,0,93,0,49,0,0,0,107,0,35,0,3,0,112,0,0,0,178,0,0,0,233,0,95,0,122,0,133,0,31,0,227,0,0,0,212,0,176,0,228,0,224,0,226,0,174,0,197,0,0,0,0,0,218,0,0,0,62,0,34,0,84,0,0,0,0,0,0,0,98,0,0,0,0,0,191,0,0,0,13,0,216,0,89,0,103,0,55,0,179,0,107,0,4,0,0,0,56,0,165,0,228,0,113,0,0,0,0,0,237,0,0,0,147,0,120,0,214,0,96,0,228,0,244,0,17,0,137,0,195,0,109,0,191,0,87,0,234,0,239,0,131,0,158,0,24,0,0,0,190,0,88,0,65,0,37,0,7,0,0,0,15,0,0,0,182,0,128,0,23,0,69,0,0,0,124,0,8,0,185,0,194,0,0,0,0,0,0,0,33,0,0,0,21,0,20,0,162,0,11,0,48,0,48,0,80,0,0,0,53,0,230,0,0,0,0,0,52,0,157,0,128,0,49,0,0,0,2,0,0,0,0,0,227,0,52,0,190,0,210,0,158,0,237,0,21,0,0,0,196,0,0,0,210,0,160,0,15,0,134,0,157,0,37,0,45,0,135,0,182,0,108,0,238,0,0,0,54,0,242,0,244,0,75,0,236,0,108,0,69,0,197,0,0,0,72,0,188,0,12,0,0,0,21,0,0,0,0,0,58,0,243,0,92,0,60,0,237,0,82,0,251,0,28,0,0,0,160,0,0,0,41,0,6,0,41,0,70,0,0,0,47,0,131,0,145,0,189,0,68,0,0,0,188,0,0,0,249,0,248,0,51,0,78,0,52,0,113,0,90,0,0,0,0,0,59,0,0,0,153,0,0,0,6,0,0,0,6,0,40,0,0,0,0,0,123,0,231,0,208,0,0,0,0,0,43,0,52,0,107,0,57,0,96,0,49,0,203,0,161,0,244,0,193,0,0,0,90,0,236,0,176,0,0,0,0,0,0,0,0,0,0,0,140,0,63,0,5,0,86,0,0,0,105,0,133,0,123,0,241,0,82,0,198,0,121,0,0,0,0,0,217,0,0,0,0,0,209,0,42,0,7,0,238,0,227,0,160,0,51,0,0,0,231,0,0,0,51,0,163,0,156,0,0,0,73,0,231,0,27,0,0,0,217,0,138,0,55,0,201,0,101,0,156,0,188,0,71,0,249,0,202,0,0,0,18,0,207,0,38,0,19,0,0,0,131,0,106,0,0,0,146,0,0,0,0,0,53,0,81,0,0,0,5,0,0,0,120,0,0,0,0,0,0,0,69,0,0,0,26,0,182,0,100,0,177,0,186,0,130,0,0,0,157,0,131,0,254,0,232,0,125,0,239,0,104,0,20,0,0,0,252,0,44,0,29,0,30,0,99,0,101,0,167,0,137,0,0,0,36,0,108,0,164,0,83,0,5,0,69,0,190,0,139,0,0,0,0,0,254,0,241,0,225,0,210,0,108,0,0,0,133,0,159,0,0,0,129,0,64,0,41,0,242,0,179,0,59,0,80,0,86,0,225,0,0,0,94,0,0,0,18,0,234,0,45,0,86,0,91,0,88,0,0,0,0,0,19,0,63,0,0,0,101,0,74,0,202,0);
signal scenario_full  : scenario_type := (24,31,24,30,41,31,12,31,239,31,96,31,209,31,48,31,109,31,88,31,254,31,131,31,253,31,12,31,12,30,12,29,12,28,52,31,132,31,14,31,50,31,52,31,59,31,59,30,216,31,211,31,211,30,3,31,169,31,170,31,68,31,85,31,102,31,22,31,184,31,184,30,151,31,42,31,6,31,19,31,126,31,236,31,187,31,181,31,154,31,239,31,27,31,250,31,10,31,111,31,7,31,71,31,218,31,48,31,203,31,70,31,70,30,66,31,236,31,66,31,216,31,114,31,156,31,210,31,183,31,183,30,89,31,10,31,93,31,238,31,244,31,10,31,10,30,143,31,4,31,172,31,11,31,73,31,114,31,62,31,20,31,135,31,19,31,66,31,168,31,97,31,194,31,194,30,144,31,144,30,63,31,162,31,207,31,190,31,160,31,161,31,79,31,79,30,194,31,106,31,206,31,81,31,206,31,61,31,229,31,169,31,164,31,164,30,15,31,139,31,33,31,33,30,247,31,177,31,233,31,227,31,227,30,203,31,172,31,180,31,71,31,215,31,8,31,120,31,100,31,31,31,84,31,84,30,252,31,252,30,227,31,84,31,195,31,195,30,111,31,112,31,170,31,217,31,191,31,123,31,42,31,42,30,119,31,202,31,97,31,181,31,112,31,148,31,166,31,133,31,16,31,16,30,16,29,62,31,88,31,88,30,135,31,179,31,123,31,178,31,80,31,80,30,144,31,103,31,9,31,215,31,215,30,105,31,125,31,219,31,238,31,92,31,156,31,237,31,116,31,93,31,49,31,49,30,107,31,35,31,3,31,112,31,112,30,178,31,178,30,233,31,95,31,122,31,133,31,31,31,227,31,227,30,212,31,176,31,228,31,224,31,226,31,174,31,197,31,197,30,197,29,218,31,218,30,62,31,34,31,84,31,84,30,84,29,84,28,98,31,98,30,98,29,191,31,191,30,13,31,216,31,89,31,103,31,55,31,179,31,107,31,4,31,4,30,56,31,165,31,228,31,113,31,113,30,113,29,237,31,237,30,147,31,120,31,214,31,96,31,228,31,244,31,17,31,137,31,195,31,109,31,191,31,87,31,234,31,239,31,131,31,158,31,24,31,24,30,190,31,88,31,65,31,37,31,7,31,7,30,15,31,15,30,182,31,128,31,23,31,69,31,69,30,124,31,8,31,185,31,194,31,194,30,194,29,194,28,33,31,33,30,21,31,20,31,162,31,11,31,48,31,48,31,80,31,80,30,53,31,230,31,230,30,230,29,52,31,157,31,128,31,49,31,49,30,2,31,2,30,2,29,227,31,52,31,190,31,210,31,158,31,237,31,21,31,21,30,196,31,196,30,210,31,160,31,15,31,134,31,157,31,37,31,45,31,135,31,182,31,108,31,238,31,238,30,54,31,242,31,244,31,75,31,236,31,108,31,69,31,197,31,197,30,72,31,188,31,12,31,12,30,21,31,21,30,21,29,58,31,243,31,92,31,60,31,237,31,82,31,251,31,28,31,28,30,160,31,160,30,41,31,6,31,41,31,70,31,70,30,47,31,131,31,145,31,189,31,68,31,68,30,188,31,188,30,249,31,248,31,51,31,78,31,52,31,113,31,90,31,90,30,90,29,59,31,59,30,153,31,153,30,6,31,6,30,6,31,40,31,40,30,40,29,123,31,231,31,208,31,208,30,208,29,43,31,52,31,107,31,57,31,96,31,49,31,203,31,161,31,244,31,193,31,193,30,90,31,236,31,176,31,176,30,176,29,176,28,176,27,176,26,140,31,63,31,5,31,86,31,86,30,105,31,133,31,123,31,241,31,82,31,198,31,121,31,121,30,121,29,217,31,217,30,217,29,209,31,42,31,7,31,238,31,227,31,160,31,51,31,51,30,231,31,231,30,51,31,163,31,156,31,156,30,73,31,231,31,27,31,27,30,217,31,138,31,55,31,201,31,101,31,156,31,188,31,71,31,249,31,202,31,202,30,18,31,207,31,38,31,19,31,19,30,131,31,106,31,106,30,146,31,146,30,146,29,53,31,81,31,81,30,5,31,5,30,120,31,120,30,120,29,120,28,69,31,69,30,26,31,182,31,100,31,177,31,186,31,130,31,130,30,157,31,131,31,254,31,232,31,125,31,239,31,104,31,20,31,20,30,252,31,44,31,29,31,30,31,99,31,101,31,167,31,137,31,137,30,36,31,108,31,164,31,83,31,5,31,69,31,190,31,139,31,139,30,139,29,254,31,241,31,225,31,210,31,108,31,108,30,133,31,159,31,159,30,129,31,64,31,41,31,242,31,179,31,59,31,80,31,86,31,225,31,225,30,94,31,94,30,18,31,234,31,45,31,86,31,91,31,88,31,88,30,88,29,19,31,63,31,63,30,101,31,74,31,202,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
