-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_41 is
end project_tb_41;

architecture project_tb_arch_41 of project_tb_41 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 630;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (43,0,69,0,26,0,144,0,159,0,46,0,240,0,0,0,223,0,171,0,127,0,91,0,246,0,201,0,220,0,64,0,0,0,26,0,21,0,0,0,121,0,102,0,227,0,0,0,42,0,10,0,19,0,50,0,234,0,136,0,40,0,152,0,137,0,49,0,0,0,101,0,217,0,0,0,77,0,182,0,0,0,143,0,207,0,121,0,26,0,99,0,243,0,79,0,103,0,156,0,0,0,216,0,0,0,27,0,6,0,253,0,84,0,0,0,120,0,185,0,87,0,0,0,13,0,167,0,0,0,206,0,183,0,241,0,222,0,193,0,230,0,18,0,38,0,102,0,220,0,109,0,7,0,51,0,110,0,210,0,245,0,0,0,74,0,0,0,196,0,0,0,168,0,0,0,68,0,37,0,0,0,81,0,193,0,146,0,112,0,189,0,60,0,189,0,239,0,33,0,226,0,0,0,13,0,221,0,159,0,0,0,122,0,42,0,0,0,226,0,14,0,158,0,204,0,129,0,253,0,254,0,200,0,50,0,38,0,8,0,2,0,111,0,150,0,72,0,4,0,0,0,154,0,159,0,91,0,33,0,138,0,56,0,10,0,10,0,127,0,235,0,184,0,218,0,18,0,134,0,57,0,113,0,57,0,39,0,229,0,166,0,185,0,0,0,167,0,208,0,206,0,94,0,45,0,115,0,189,0,199,0,0,0,95,0,96,0,13,0,135,0,237,0,26,0,90,0,193,0,156,0,38,0,242,0,0,0,197,0,150,0,152,0,0,0,0,0,0,0,168,0,91,0,43,0,19,0,0,0,0,0,0,0,128,0,18,0,174,0,78,0,179,0,142,0,115,0,11,0,0,0,195,0,62,0,236,0,33,0,142,0,202,0,97,0,171,0,61,0,160,0,200,0,219,0,135,0,105,0,166,0,0,0,0,0,189,0,212,0,76,0,209,0,73,0,205,0,0,0,0,0,16,0,210,0,0,0,239,0,27,0,217,0,16,0,155,0,247,0,0,0,70,0,97,0,69,0,79,0,69,0,25,0,95,0,0,0,31,0,0,0,51,0,49,0,0,0,115,0,172,0,199,0,161,0,189,0,22,0,0,0,231,0,246,0,35,0,0,0,174,0,188,0,0,0,67,0,40,0,130,0,11,0,171,0,243,0,67,0,109,0,0,0,52,0,149,0,251,0,60,0,193,0,19,0,67,0,0,0,222,0,248,0,16,0,17,0,86,0,117,0,143,0,42,0,225,0,231,0,0,0,38,0,5,0,0,0,113,0,122,0,0,0,173,0,6,0,0,0,237,0,255,0,75,0,59,0,213,0,70,0,172,0,0,0,189,0,0,0,116,0,182,0,140,0,21,0,0,0,53,0,0,0,164,0,139,0,45,0,180,0,35,0,0,0,19,0,179,0,150,0,237,0,111,0,8,0,58,0,153,0,21,0,219,0,208,0,66,0,144,0,151,0,0,0,114,0,158,0,16,0,45,0,0,0,80,0,86,0,47,0,66,0,126,0,8,0,22,0,0,0,18,0,0,0,0,0,0,0,65,0,125,0,182,0,174,0,138,0,75,0,219,0,111,0,99,0,35,0,0,0,6,0,93,0,149,0,220,0,114,0,0,0,95,0,19,0,78,0,189,0,88,0,49,0,230,0,0,0,157,0,106,0,253,0,173,0,198,0,0,0,66,0,33,0,197,0,110,0,0,0,0,0,205,0,0,0,31,0,132,0,71,0,95,0,190,0,68,0,112,0,254,0,27,0,16,0,20,0,0,0,21,0,0,0,5,0,244,0,96,0,62,0,66,0,0,0,247,0,50,0,0,0,213,0,164,0,0,0,95,0,7,0,188,0,154,0,69,0,0,0,96,0,166,0,0,0,46,0,86,0,204,0,0,0,254,0,191,0,0,0,232,0,215,0,252,0,122,0,79,0,82,0,171,0,6,0,127,0,0,0,0,0,156,0,0,0,84,0,236,0,0,0,102,0,54,0,9,0,176,0,49,0,48,0,206,0,0,0,132,0,0,0,250,0,63,0,158,0,65,0,0,0,76,0,0,0,205,0,69,0,130,0,0,0,166,0,220,0,207,0,244,0,248,0,244,0,68,0,214,0,255,0,0,0,188,0,48,0,41,0,0,0,0,0,166,0,159,0,108,0,125,0,0,0,68,0,234,0,132,0,47,0,224,0,191,0,209,0,248,0,78,0,108,0,154,0,4,0,177,0,135,0,243,0,0,0,0,0,140,0,70,0,0,0,63,0,0,0,53,0,155,0,18,0,0,0,163,0,109,0,0,0,47,0,0,0,65,0,95,0,53,0,40,0,254,0,21,0,105,0,86,0,250,0,137,0,22,0,0,0,11,0,253,0,37,0,149,0,142,0,252,0,0,0,20,0,0,0,0,0,0,0,0,0,61,0,242,0,162,0,30,0,90,0,84,0,0,0,137,0,90,0,131,0,176,0,248,0,127,0,15,0,0,0,160,0,254,0,0,0,0,0,0,0,19,0,36,0,197,0,0,0,200,0,176,0,0,0,0,0,44,0,23,0,9,0,89,0,0,0,200,0,79,0,78,0,65,0,141,0,90,0,0,0,9,0,0,0,179,0,178,0,29,0,152,0,191,0,179,0,0,0,202,0,145,0,156,0,242,0,160,0,2,0,82,0,0,0,0,0,183,0,161,0,164,0,0,0,153,0,219,0,0,0,160,0,179,0,169,0,220,0,0,0,142,0,94,0,248,0,23,0,160,0,62,0,108,0,64,0,226,0,0,0,243,0,10,0,15,0,0,0,179,0,36,0,0,0,174,0,21,0,191,0,53,0,95,0);
signal scenario_full  : scenario_type := (43,31,69,31,26,31,144,31,159,31,46,31,240,31,240,30,223,31,171,31,127,31,91,31,246,31,201,31,220,31,64,31,64,30,26,31,21,31,21,30,121,31,102,31,227,31,227,30,42,31,10,31,19,31,50,31,234,31,136,31,40,31,152,31,137,31,49,31,49,30,101,31,217,31,217,30,77,31,182,31,182,30,143,31,207,31,121,31,26,31,99,31,243,31,79,31,103,31,156,31,156,30,216,31,216,30,27,31,6,31,253,31,84,31,84,30,120,31,185,31,87,31,87,30,13,31,167,31,167,30,206,31,183,31,241,31,222,31,193,31,230,31,18,31,38,31,102,31,220,31,109,31,7,31,51,31,110,31,210,31,245,31,245,30,74,31,74,30,196,31,196,30,168,31,168,30,68,31,37,31,37,30,81,31,193,31,146,31,112,31,189,31,60,31,189,31,239,31,33,31,226,31,226,30,13,31,221,31,159,31,159,30,122,31,42,31,42,30,226,31,14,31,158,31,204,31,129,31,253,31,254,31,200,31,50,31,38,31,8,31,2,31,111,31,150,31,72,31,4,31,4,30,154,31,159,31,91,31,33,31,138,31,56,31,10,31,10,31,127,31,235,31,184,31,218,31,18,31,134,31,57,31,113,31,57,31,39,31,229,31,166,31,185,31,185,30,167,31,208,31,206,31,94,31,45,31,115,31,189,31,199,31,199,30,95,31,96,31,13,31,135,31,237,31,26,31,90,31,193,31,156,31,38,31,242,31,242,30,197,31,150,31,152,31,152,30,152,29,152,28,168,31,91,31,43,31,19,31,19,30,19,29,19,28,128,31,18,31,174,31,78,31,179,31,142,31,115,31,11,31,11,30,195,31,62,31,236,31,33,31,142,31,202,31,97,31,171,31,61,31,160,31,200,31,219,31,135,31,105,31,166,31,166,30,166,29,189,31,212,31,76,31,209,31,73,31,205,31,205,30,205,29,16,31,210,31,210,30,239,31,27,31,217,31,16,31,155,31,247,31,247,30,70,31,97,31,69,31,79,31,69,31,25,31,95,31,95,30,31,31,31,30,51,31,49,31,49,30,115,31,172,31,199,31,161,31,189,31,22,31,22,30,231,31,246,31,35,31,35,30,174,31,188,31,188,30,67,31,40,31,130,31,11,31,171,31,243,31,67,31,109,31,109,30,52,31,149,31,251,31,60,31,193,31,19,31,67,31,67,30,222,31,248,31,16,31,17,31,86,31,117,31,143,31,42,31,225,31,231,31,231,30,38,31,5,31,5,30,113,31,122,31,122,30,173,31,6,31,6,30,237,31,255,31,75,31,59,31,213,31,70,31,172,31,172,30,189,31,189,30,116,31,182,31,140,31,21,31,21,30,53,31,53,30,164,31,139,31,45,31,180,31,35,31,35,30,19,31,179,31,150,31,237,31,111,31,8,31,58,31,153,31,21,31,219,31,208,31,66,31,144,31,151,31,151,30,114,31,158,31,16,31,45,31,45,30,80,31,86,31,47,31,66,31,126,31,8,31,22,31,22,30,18,31,18,30,18,29,18,28,65,31,125,31,182,31,174,31,138,31,75,31,219,31,111,31,99,31,35,31,35,30,6,31,93,31,149,31,220,31,114,31,114,30,95,31,19,31,78,31,189,31,88,31,49,31,230,31,230,30,157,31,106,31,253,31,173,31,198,31,198,30,66,31,33,31,197,31,110,31,110,30,110,29,205,31,205,30,31,31,132,31,71,31,95,31,190,31,68,31,112,31,254,31,27,31,16,31,20,31,20,30,21,31,21,30,5,31,244,31,96,31,62,31,66,31,66,30,247,31,50,31,50,30,213,31,164,31,164,30,95,31,7,31,188,31,154,31,69,31,69,30,96,31,166,31,166,30,46,31,86,31,204,31,204,30,254,31,191,31,191,30,232,31,215,31,252,31,122,31,79,31,82,31,171,31,6,31,127,31,127,30,127,29,156,31,156,30,84,31,236,31,236,30,102,31,54,31,9,31,176,31,49,31,48,31,206,31,206,30,132,31,132,30,250,31,63,31,158,31,65,31,65,30,76,31,76,30,205,31,69,31,130,31,130,30,166,31,220,31,207,31,244,31,248,31,244,31,68,31,214,31,255,31,255,30,188,31,48,31,41,31,41,30,41,29,166,31,159,31,108,31,125,31,125,30,68,31,234,31,132,31,47,31,224,31,191,31,209,31,248,31,78,31,108,31,154,31,4,31,177,31,135,31,243,31,243,30,243,29,140,31,70,31,70,30,63,31,63,30,53,31,155,31,18,31,18,30,163,31,109,31,109,30,47,31,47,30,65,31,95,31,53,31,40,31,254,31,21,31,105,31,86,31,250,31,137,31,22,31,22,30,11,31,253,31,37,31,149,31,142,31,252,31,252,30,20,31,20,30,20,29,20,28,20,27,61,31,242,31,162,31,30,31,90,31,84,31,84,30,137,31,90,31,131,31,176,31,248,31,127,31,15,31,15,30,160,31,254,31,254,30,254,29,254,28,19,31,36,31,197,31,197,30,200,31,176,31,176,30,176,29,44,31,23,31,9,31,89,31,89,30,200,31,79,31,78,31,65,31,141,31,90,31,90,30,9,31,9,30,179,31,178,31,29,31,152,31,191,31,179,31,179,30,202,31,145,31,156,31,242,31,160,31,2,31,82,31,82,30,82,29,183,31,161,31,164,31,164,30,153,31,219,31,219,30,160,31,179,31,169,31,220,31,220,30,142,31,94,31,248,31,23,31,160,31,62,31,108,31,64,31,226,31,226,30,243,31,10,31,15,31,15,30,179,31,36,31,36,30,174,31,21,31,191,31,53,31,95,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
