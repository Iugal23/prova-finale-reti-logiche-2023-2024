-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 588;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (10,0,67,0,0,0,0,0,180,0,0,0,248,0,140,0,155,0,234,0,182,0,63,0,124,0,254,0,0,0,236,0,0,0,170,0,0,0,167,0,137,0,182,0,0,0,175,0,175,0,30,0,212,0,95,0,152,0,39,0,0,0,0,0,104,0,203,0,219,0,39,0,224,0,17,0,167,0,102,0,131,0,132,0,0,0,121,0,55,0,220,0,0,0,0,0,0,0,243,0,94,0,0,0,0,0,58,0,121,0,239,0,0,0,37,0,56,0,83,0,0,0,47,0,205,0,163,0,18,0,0,0,232,0,22,0,197,0,0,0,0,0,0,0,184,0,106,0,76,0,0,0,95,0,86,0,61,0,0,0,1,0,155,0,240,0,150,0,3,0,195,0,226,0,191,0,94,0,90,0,82,0,218,0,63,0,3,0,167,0,0,0,0,0,0,0,172,0,176,0,165,0,85,0,153,0,0,0,120,0,0,0,116,0,0,0,133,0,222,0,197,0,219,0,200,0,0,0,1,0,141,0,181,0,222,0,169,0,101,0,0,0,0,0,210,0,147,0,108,0,0,0,154,0,202,0,0,0,0,0,0,0,231,0,148,0,152,0,4,0,89,0,0,0,120,0,212,0,49,0,129,0,204,0,223,0,4,0,205,0,23,0,25,0,105,0,110,0,161,0,252,0,26,0,254,0,51,0,144,0,229,0,41,0,30,0,230,0,213,0,174,0,208,0,108,0,40,0,240,0,0,0,242,0,25,0,191,0,0,0,225,0,195,0,19,0,0,0,0,0,215,0,198,0,58,0,184,0,0,0,0,0,108,0,121,0,0,0,104,0,200,0,237,0,175,0,0,0,108,0,28,0,5,0,116,0,0,0,207,0,0,0,57,0,98,0,115,0,83,0,164,0,0,0,28,0,99,0,0,0,92,0,50,0,230,0,225,0,188,0,131,0,30,0,195,0,93,0,72,0,214,0,185,0,112,0,228,0,252,0,195,0,55,0,53,0,231,0,0,0,0,0,51,0,1,0,206,0,122,0,247,0,0,0,233,0,236,0,164,0,0,0,228,0,0,0,0,0,93,0,114,0,242,0,0,0,199,0,202,0,214,0,139,0,0,0,124,0,170,0,87,0,0,0,65,0,180,0,90,0,224,0,10,0,123,0,187,0,0,0,116,0,161,0,78,0,25,0,85,0,45,0,107,0,142,0,0,0,0,0,0,0,215,0,0,0,127,0,97,0,120,0,193,0,99,0,56,0,218,0,0,0,189,0,27,0,17,0,31,0,51,0,26,0,140,0,208,0,30,0,40,0,0,0,39,0,76,0,2,0,201,0,82,0,81,0,167,0,33,0,0,0,130,0,0,0,111,0,182,0,0,0,0,0,127,0,12,0,172,0,165,0,65,0,255,0,216,0,46,0,44,0,44,0,91,0,88,0,238,0,24,0,4,0,0,0,41,0,0,0,0,0,239,0,0,0,103,0,77,0,53,0,65,0,0,0,150,0,0,0,3,0,92,0,99,0,228,0,14,0,60,0,246,0,253,0,92,0,163,0,160,0,0,0,0,0,0,0,237,0,217,0,200,0,106,0,0,0,151,0,135,0,79,0,0,0,229,0,11,0,134,0,0,0,0,0,0,0,203,0,235,0,153,0,39,0,107,0,0,0,253,0,158,0,93,0,148,0,117,0,205,0,0,0,139,0,92,0,178,0,0,0,0,0,15,0,204,0,25,0,191,0,0,0,73,0,142,0,0,0,157,0,0,0,197,0,163,0,46,0,0,0,87,0,0,0,37,0,208,0,88,0,162,0,53,0,144,0,116,0,14,0,164,0,189,0,53,0,50,0,113,0,132,0,61,0,117,0,209,0,91,0,60,0,167,0,22,0,183,0,231,0,167,0,101,0,77,0,0,0,229,0,0,0,65,0,121,0,114,0,15,0,0,0,0,0,26,0,74,0,188,0,0,0,246,0,0,0,114,0,212,0,0,0,214,0,205,0,119,0,37,0,185,0,151,0,66,0,0,0,127,0,111,0,65,0,252,0,10,0,192,0,26,0,27,0,129,0,187,0,165,0,76,0,221,0,128,0,83,0,0,0,241,0,42,0,199,0,168,0,130,0,0,0,137,0,247,0,41,0,196,0,120,0,110,0,0,0,55,0,8,0,0,0,0,0,231,0,66,0,197,0,19,0,103,0,34,0,196,0,209,0,227,0,8,0,225,0,169,0,68,0,22,0,0,0,163,0,135,0,98,0,229,0,0,0,106,0,31,0,0,0,91,0,115,0,37,0,32,0,225,0,96,0,250,0,229,0,0,0,0,0,122,0,54,0,6,0,246,0,166,0,76,0,0,0,216,0,0,0,97,0,0,0,0,0,165,0,208,0,133,0,162,0,61,0,168,0,166,0,236,0,201,0,193,0,39,0,30,0,110,0,235,0,143,0,0,0,236,0,0,0,129,0,107,0,0,0,172,0,187,0,89,0,133,0,200,0,240,0,206,0,52,0,127,0,85,0,199,0,131,0,0,0,205,0,245,0,122,0,0,0,170,0,10,0,141,0,208,0,0,0,74,0,14,0,33,0,199,0,94,0,181,0,196,0,0,0,28,0,0,0,6,0,123,0,32,0,4,0,106,0,68,0,183,0);
signal scenario_full  : scenario_type := (10,31,67,31,67,30,67,29,180,31,180,30,248,31,140,31,155,31,234,31,182,31,63,31,124,31,254,31,254,30,236,31,236,30,170,31,170,30,167,31,137,31,182,31,182,30,175,31,175,31,30,31,212,31,95,31,152,31,39,31,39,30,39,29,104,31,203,31,219,31,39,31,224,31,17,31,167,31,102,31,131,31,132,31,132,30,121,31,55,31,220,31,220,30,220,29,220,28,243,31,94,31,94,30,94,29,58,31,121,31,239,31,239,30,37,31,56,31,83,31,83,30,47,31,205,31,163,31,18,31,18,30,232,31,22,31,197,31,197,30,197,29,197,28,184,31,106,31,76,31,76,30,95,31,86,31,61,31,61,30,1,31,155,31,240,31,150,31,3,31,195,31,226,31,191,31,94,31,90,31,82,31,218,31,63,31,3,31,167,31,167,30,167,29,167,28,172,31,176,31,165,31,85,31,153,31,153,30,120,31,120,30,116,31,116,30,133,31,222,31,197,31,219,31,200,31,200,30,1,31,141,31,181,31,222,31,169,31,101,31,101,30,101,29,210,31,147,31,108,31,108,30,154,31,202,31,202,30,202,29,202,28,231,31,148,31,152,31,4,31,89,31,89,30,120,31,212,31,49,31,129,31,204,31,223,31,4,31,205,31,23,31,25,31,105,31,110,31,161,31,252,31,26,31,254,31,51,31,144,31,229,31,41,31,30,31,230,31,213,31,174,31,208,31,108,31,40,31,240,31,240,30,242,31,25,31,191,31,191,30,225,31,195,31,19,31,19,30,19,29,215,31,198,31,58,31,184,31,184,30,184,29,108,31,121,31,121,30,104,31,200,31,237,31,175,31,175,30,108,31,28,31,5,31,116,31,116,30,207,31,207,30,57,31,98,31,115,31,83,31,164,31,164,30,28,31,99,31,99,30,92,31,50,31,230,31,225,31,188,31,131,31,30,31,195,31,93,31,72,31,214,31,185,31,112,31,228,31,252,31,195,31,55,31,53,31,231,31,231,30,231,29,51,31,1,31,206,31,122,31,247,31,247,30,233,31,236,31,164,31,164,30,228,31,228,30,228,29,93,31,114,31,242,31,242,30,199,31,202,31,214,31,139,31,139,30,124,31,170,31,87,31,87,30,65,31,180,31,90,31,224,31,10,31,123,31,187,31,187,30,116,31,161,31,78,31,25,31,85,31,45,31,107,31,142,31,142,30,142,29,142,28,215,31,215,30,127,31,97,31,120,31,193,31,99,31,56,31,218,31,218,30,189,31,27,31,17,31,31,31,51,31,26,31,140,31,208,31,30,31,40,31,40,30,39,31,76,31,2,31,201,31,82,31,81,31,167,31,33,31,33,30,130,31,130,30,111,31,182,31,182,30,182,29,127,31,12,31,172,31,165,31,65,31,255,31,216,31,46,31,44,31,44,31,91,31,88,31,238,31,24,31,4,31,4,30,41,31,41,30,41,29,239,31,239,30,103,31,77,31,53,31,65,31,65,30,150,31,150,30,3,31,92,31,99,31,228,31,14,31,60,31,246,31,253,31,92,31,163,31,160,31,160,30,160,29,160,28,237,31,217,31,200,31,106,31,106,30,151,31,135,31,79,31,79,30,229,31,11,31,134,31,134,30,134,29,134,28,203,31,235,31,153,31,39,31,107,31,107,30,253,31,158,31,93,31,148,31,117,31,205,31,205,30,139,31,92,31,178,31,178,30,178,29,15,31,204,31,25,31,191,31,191,30,73,31,142,31,142,30,157,31,157,30,197,31,163,31,46,31,46,30,87,31,87,30,37,31,208,31,88,31,162,31,53,31,144,31,116,31,14,31,164,31,189,31,53,31,50,31,113,31,132,31,61,31,117,31,209,31,91,31,60,31,167,31,22,31,183,31,231,31,167,31,101,31,77,31,77,30,229,31,229,30,65,31,121,31,114,31,15,31,15,30,15,29,26,31,74,31,188,31,188,30,246,31,246,30,114,31,212,31,212,30,214,31,205,31,119,31,37,31,185,31,151,31,66,31,66,30,127,31,111,31,65,31,252,31,10,31,192,31,26,31,27,31,129,31,187,31,165,31,76,31,221,31,128,31,83,31,83,30,241,31,42,31,199,31,168,31,130,31,130,30,137,31,247,31,41,31,196,31,120,31,110,31,110,30,55,31,8,31,8,30,8,29,231,31,66,31,197,31,19,31,103,31,34,31,196,31,209,31,227,31,8,31,225,31,169,31,68,31,22,31,22,30,163,31,135,31,98,31,229,31,229,30,106,31,31,31,31,30,91,31,115,31,37,31,32,31,225,31,96,31,250,31,229,31,229,30,229,29,122,31,54,31,6,31,246,31,166,31,76,31,76,30,216,31,216,30,97,31,97,30,97,29,165,31,208,31,133,31,162,31,61,31,168,31,166,31,236,31,201,31,193,31,39,31,30,31,110,31,235,31,143,31,143,30,236,31,236,30,129,31,107,31,107,30,172,31,187,31,89,31,133,31,200,31,240,31,206,31,52,31,127,31,85,31,199,31,131,31,131,30,205,31,245,31,122,31,122,30,170,31,10,31,141,31,208,31,208,30,74,31,14,31,33,31,199,31,94,31,181,31,196,31,196,30,28,31,28,30,6,31,123,31,32,31,4,31,106,31,68,31,183,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
