-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 905;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,71,0,193,0,0,0,98,0,202,0,249,0,0,0,53,0,151,0,0,0,238,0,134,0,0,0,132,0,198,0,84,0,0,0,34,0,0,0,0,0,228,0,172,0,207,0,200,0,165,0,224,0,60,0,59,0,52,0,180,0,150,0,93,0,0,0,246,0,176,0,15,0,180,0,221,0,138,0,189,0,0,0,114,0,69,0,0,0,0,0,51,0,181,0,92,0,211,0,182,0,0,0,131,0,166,0,24,0,0,0,0,0,44,0,0,0,77,0,69,0,0,0,225,0,157,0,21,0,32,0,0,0,23,0,172,0,176,0,0,0,103,0,8,0,0,0,93,0,0,0,9,0,0,0,169,0,46,0,0,0,39,0,20,0,153,0,180,0,201,0,171,0,229,0,22,0,0,0,76,0,141,0,237,0,112,0,6,0,0,0,84,0,0,0,0,0,22,0,21,0,51,0,70,0,106,0,0,0,0,0,106,0,61,0,103,0,8,0,82,0,209,0,101,0,29,0,142,0,48,0,68,0,126,0,104,0,97,0,179,0,0,0,185,0,165,0,243,0,196,0,124,0,0,0,173,0,101,0,150,0,225,0,239,0,159,0,125,0,175,0,0,0,0,0,17,0,41,0,148,0,42,0,0,0,0,0,169,0,184,0,38,0,0,0,140,0,190,0,31,0,249,0,204,0,2,0,227,0,156,0,232,0,0,0,0,0,218,0,91,0,105,0,170,0,171,0,182,0,163,0,0,0,223,0,183,0,245,0,80,0,176,0,189,0,46,0,225,0,0,0,206,0,204,0,60,0,223,0,13,0,22,0,203,0,124,0,185,0,75,0,62,0,47,0,21,0,186,0,212,0,36,0,13,0,165,0,75,0,68,0,217,0,213,0,153,0,198,0,12,0,0,0,85,0,33,0,135,0,116,0,190,0,81,0,153,0,201,0,235,0,28,0,211,0,0,0,0,0,67,0,8,0,3,0,44,0,201,0,119,0,198,0,0,0,170,0,185,0,151,0,223,0,197,0,18,0,14,0,0,0,0,0,10,0,0,0,37,0,158,0,195,0,203,0,20,0,157,0,118,0,0,0,127,0,154,0,72,0,154,0,174,0,75,0,253,0,178,0,0,0,220,0,63,0,226,0,130,0,166,0,0,0,19,0,18,0,0,0,177,0,161,0,58,0,142,0,177,0,0,0,72,0,114,0,40,0,187,0,0,0,219,0,62,0,113,0,209,0,0,0,12,0,244,0,199,0,139,0,240,0,0,0,155,0,83,0,81,0,47,0,43,0,180,0,236,0,28,0,47,0,153,0,22,0,62,0,1,0,179,0,98,0,172,0,0,0,57,0,68,0,136,0,1,0,25,0,79,0,194,0,198,0,24,0,0,0,156,0,150,0,89,0,181,0,199,0,132,0,105,0,0,0,0,0,61,0,208,0,97,0,198,0,151,0,229,0,115,0,76,0,171,0,123,0,161,0,238,0,5,0,195,0,172,0,45,0,0,0,104,0,157,0,61,0,60,0,14,0,14,0,45,0,230,0,238,0,231,0,159,0,39,0,53,0,0,0,92,0,61,0,178,0,159,0,254,0,105,0,0,0,0,0,160,0,45,0,141,0,221,0,0,0,0,0,135,0,107,0,30,0,5,0,111,0,196,0,0,0,9,0,125,0,201,0,101,0,0,0,220,0,141,0,225,0,0,0,159,0,136,0,44,0,6,0,201,0,252,0,139,0,17,0,172,0,115,0,0,0,113,0,70,0,7,0,252,0,25,0,90,0,70,0,0,0,0,0,0,0,0,0,100,0,232,0,18,0,235,0,190,0,169,0,0,0,226,0,17,0,0,0,120,0,253,0,0,0,0,0,228,0,157,0,158,0,0,0,55,0,232,0,0,0,188,0,136,0,91,0,250,0,53,0,175,0,123,0,123,0,78,0,105,0,196,0,209,0,232,0,217,0,0,0,36,0,220,0,57,0,175,0,12,0,89,0,0,0,0,0,45,0,109,0,125,0,73,0,0,0,217,0,56,0,0,0,128,0,0,0,168,0,0,0,0,0,193,0,207,0,138,0,0,0,172,0,36,0,214,0,0,0,184,0,149,0,246,0,229,0,8,0,43,0,224,0,195,0,64,0,172,0,162,0,114,0,157,0,8,0,97,0,174,0,185,0,162,0,177,0,74,0,195,0,163,0,115,0,160,0,138,0,197,0,253,0,0,0,62,0,210,0,126,0,214,0,43,0,34,0,204,0,197,0,225,0,166,0,124,0,192,0,4,0,118,0,242,0,31,0,226,0,242,0,0,0,198,0,0,0,53,0,25,0,173,0,177,0,0,0,198,0,45,0,164,0,142,0,0,0,21,0,153,0,47,0,0,0,210,0,132,0,195,0,0,0,74,0,97,0,154,0,65,0,186,0,66,0,183,0,0,0,100,0,0,0,207,0,0,0,88,0,166,0,48,0,56,0,107,0,73,0,0,0,195,0,0,0,0,0,154,0,231,0,83,0,147,0,157,0,42,0,252,0,0,0,32,0,13,0,221,0,160,0,0,0,0,0,0,0,56,0,13,0,108,0,103,0,0,0,3,0,243,0,95,0,0,0,0,0,225,0,143,0,173,0,47,0,183,0,105,0,0,0,133,0,19,0,128,0,7,0,89,0,0,0,247,0,73,0,0,0,232,0,153,0,239,0,85,0,92,0,181,0,103,0,145,0,37,0,17,0,214,0,175,0,127,0,193,0,5,0,24,0,0,0,76,0,182,0,10,0,235,0,41,0,175,0,0,0,0,0,150,0,3,0,139,0,154,0,159,0,38,0,102,0,116,0,201,0,0,0,128,0,0,0,92,0,27,0,97,0,205,0,0,0,163,0,49,0,183,0,110,0,0,0,252,0,0,0,75,0,124,0,208,0,0,0,39,0,0,0,141,0,121,0,166,0,23,0,184,0,13,0,163,0,171,0,162,0,192,0,18,0,74,0,33,0,123,0,122,0,47,0,28,0,19,0,8,0,240,0,39,0,87,0,34,0,251,0,34,0,26,0,86,0,228,0,9,0,0,0,1,0,238,0,129,0,155,0,110,0,0,0,124,0,0,0,45,0,122,0,178,0,45,0,32,0,103,0,84,0,10,0,94,0,73,0,78,0,159,0,227,0,127,0,71,0,0,0,21,0,191,0,110,0,187,0,182,0,139,0,214,0,183,0,0,0,126,0,25,0,18,0,190,0,165,0,22,0,233,0,57,0,66,0,79,0,94,0,6,0,231,0,172,0,160,0,0,0,55,0,245,0,223,0,73,0,18,0,16,0,247,0,15,0,232,0,240,0,123,0,22,0,35,0,207,0,248,0,169,0,0,0,225,0,148,0,0,0,97,0,0,0,111,0,19,0,0,0,62,0,231,0,20,0,176,0,220,0,24,0,136,0,241,0,0,0,212,0,40,0,0,0,39,0,178,0,0,0,0,0,204,0,88,0,246,0,249,0,96,0,72,0,208,0,44,0,64,0,161,0,142,0,222,0,189,0,165,0,100,0,119,0,51,0,0,0,71,0,0,0,129,0,209,0,16,0,152,0,31,0,53,0,154,0,0,0,124,0,110,0,0,0,196,0,249,0,20,0,116,0,175,0,181,0,0,0,156,0,217,0,188,0,74,0,187,0,7,0,116,0,193,0,0,0,128,0,70,0,254,0,136,0,112,0,230,0,124,0,0,0,227,0,0,0,196,0,203,0,86,0,129,0,86,0,235,0,39,0,244,0,207,0,0,0,0,0,96,0,131,0,107,0,254,0,0,0,248,0,0,0,8,0,113,0,228,0,0,0,96,0,138,0,0,0,42,0,6,0,28,0,0,0,108,0,80,0,0,0,0,0,215,0,69,0,3,0,196,0,194,0,73,0,3,0,242,0,0,0,62,0,41,0,107,0,238,0,250,0,21,0,52,0,18,0,222,0,73,0,96,0,0,0,108,0,0,0,149,0,95,0,149,0,121,0,23,0,114,0,39,0,106,0,0,0,130,0,219,0,198,0,179,0,0,0,80,0,97,0,198,0,249,0,0,0,214,0,33,0);
signal scenario_full  : scenario_type := (214,31,71,31,193,31,193,30,98,31,202,31,249,31,249,30,53,31,151,31,151,30,238,31,134,31,134,30,132,31,198,31,84,31,84,30,34,31,34,30,34,29,228,31,172,31,207,31,200,31,165,31,224,31,60,31,59,31,52,31,180,31,150,31,93,31,93,30,246,31,176,31,15,31,180,31,221,31,138,31,189,31,189,30,114,31,69,31,69,30,69,29,51,31,181,31,92,31,211,31,182,31,182,30,131,31,166,31,24,31,24,30,24,29,44,31,44,30,77,31,69,31,69,30,225,31,157,31,21,31,32,31,32,30,23,31,172,31,176,31,176,30,103,31,8,31,8,30,93,31,93,30,9,31,9,30,169,31,46,31,46,30,39,31,20,31,153,31,180,31,201,31,171,31,229,31,22,31,22,30,76,31,141,31,237,31,112,31,6,31,6,30,84,31,84,30,84,29,22,31,21,31,51,31,70,31,106,31,106,30,106,29,106,31,61,31,103,31,8,31,82,31,209,31,101,31,29,31,142,31,48,31,68,31,126,31,104,31,97,31,179,31,179,30,185,31,165,31,243,31,196,31,124,31,124,30,173,31,101,31,150,31,225,31,239,31,159,31,125,31,175,31,175,30,175,29,17,31,41,31,148,31,42,31,42,30,42,29,169,31,184,31,38,31,38,30,140,31,190,31,31,31,249,31,204,31,2,31,227,31,156,31,232,31,232,30,232,29,218,31,91,31,105,31,170,31,171,31,182,31,163,31,163,30,223,31,183,31,245,31,80,31,176,31,189,31,46,31,225,31,225,30,206,31,204,31,60,31,223,31,13,31,22,31,203,31,124,31,185,31,75,31,62,31,47,31,21,31,186,31,212,31,36,31,13,31,165,31,75,31,68,31,217,31,213,31,153,31,198,31,12,31,12,30,85,31,33,31,135,31,116,31,190,31,81,31,153,31,201,31,235,31,28,31,211,31,211,30,211,29,67,31,8,31,3,31,44,31,201,31,119,31,198,31,198,30,170,31,185,31,151,31,223,31,197,31,18,31,14,31,14,30,14,29,10,31,10,30,37,31,158,31,195,31,203,31,20,31,157,31,118,31,118,30,127,31,154,31,72,31,154,31,174,31,75,31,253,31,178,31,178,30,220,31,63,31,226,31,130,31,166,31,166,30,19,31,18,31,18,30,177,31,161,31,58,31,142,31,177,31,177,30,72,31,114,31,40,31,187,31,187,30,219,31,62,31,113,31,209,31,209,30,12,31,244,31,199,31,139,31,240,31,240,30,155,31,83,31,81,31,47,31,43,31,180,31,236,31,28,31,47,31,153,31,22,31,62,31,1,31,179,31,98,31,172,31,172,30,57,31,68,31,136,31,1,31,25,31,79,31,194,31,198,31,24,31,24,30,156,31,150,31,89,31,181,31,199,31,132,31,105,31,105,30,105,29,61,31,208,31,97,31,198,31,151,31,229,31,115,31,76,31,171,31,123,31,161,31,238,31,5,31,195,31,172,31,45,31,45,30,104,31,157,31,61,31,60,31,14,31,14,31,45,31,230,31,238,31,231,31,159,31,39,31,53,31,53,30,92,31,61,31,178,31,159,31,254,31,105,31,105,30,105,29,160,31,45,31,141,31,221,31,221,30,221,29,135,31,107,31,30,31,5,31,111,31,196,31,196,30,9,31,125,31,201,31,101,31,101,30,220,31,141,31,225,31,225,30,159,31,136,31,44,31,6,31,201,31,252,31,139,31,17,31,172,31,115,31,115,30,113,31,70,31,7,31,252,31,25,31,90,31,70,31,70,30,70,29,70,28,70,27,100,31,232,31,18,31,235,31,190,31,169,31,169,30,226,31,17,31,17,30,120,31,253,31,253,30,253,29,228,31,157,31,158,31,158,30,55,31,232,31,232,30,188,31,136,31,91,31,250,31,53,31,175,31,123,31,123,31,78,31,105,31,196,31,209,31,232,31,217,31,217,30,36,31,220,31,57,31,175,31,12,31,89,31,89,30,89,29,45,31,109,31,125,31,73,31,73,30,217,31,56,31,56,30,128,31,128,30,168,31,168,30,168,29,193,31,207,31,138,31,138,30,172,31,36,31,214,31,214,30,184,31,149,31,246,31,229,31,8,31,43,31,224,31,195,31,64,31,172,31,162,31,114,31,157,31,8,31,97,31,174,31,185,31,162,31,177,31,74,31,195,31,163,31,115,31,160,31,138,31,197,31,253,31,253,30,62,31,210,31,126,31,214,31,43,31,34,31,204,31,197,31,225,31,166,31,124,31,192,31,4,31,118,31,242,31,31,31,226,31,242,31,242,30,198,31,198,30,53,31,25,31,173,31,177,31,177,30,198,31,45,31,164,31,142,31,142,30,21,31,153,31,47,31,47,30,210,31,132,31,195,31,195,30,74,31,97,31,154,31,65,31,186,31,66,31,183,31,183,30,100,31,100,30,207,31,207,30,88,31,166,31,48,31,56,31,107,31,73,31,73,30,195,31,195,30,195,29,154,31,231,31,83,31,147,31,157,31,42,31,252,31,252,30,32,31,13,31,221,31,160,31,160,30,160,29,160,28,56,31,13,31,108,31,103,31,103,30,3,31,243,31,95,31,95,30,95,29,225,31,143,31,173,31,47,31,183,31,105,31,105,30,133,31,19,31,128,31,7,31,89,31,89,30,247,31,73,31,73,30,232,31,153,31,239,31,85,31,92,31,181,31,103,31,145,31,37,31,17,31,214,31,175,31,127,31,193,31,5,31,24,31,24,30,76,31,182,31,10,31,235,31,41,31,175,31,175,30,175,29,150,31,3,31,139,31,154,31,159,31,38,31,102,31,116,31,201,31,201,30,128,31,128,30,92,31,27,31,97,31,205,31,205,30,163,31,49,31,183,31,110,31,110,30,252,31,252,30,75,31,124,31,208,31,208,30,39,31,39,30,141,31,121,31,166,31,23,31,184,31,13,31,163,31,171,31,162,31,192,31,18,31,74,31,33,31,123,31,122,31,47,31,28,31,19,31,8,31,240,31,39,31,87,31,34,31,251,31,34,31,26,31,86,31,228,31,9,31,9,30,1,31,238,31,129,31,155,31,110,31,110,30,124,31,124,30,45,31,122,31,178,31,45,31,32,31,103,31,84,31,10,31,94,31,73,31,78,31,159,31,227,31,127,31,71,31,71,30,21,31,191,31,110,31,187,31,182,31,139,31,214,31,183,31,183,30,126,31,25,31,18,31,190,31,165,31,22,31,233,31,57,31,66,31,79,31,94,31,6,31,231,31,172,31,160,31,160,30,55,31,245,31,223,31,73,31,18,31,16,31,247,31,15,31,232,31,240,31,123,31,22,31,35,31,207,31,248,31,169,31,169,30,225,31,148,31,148,30,97,31,97,30,111,31,19,31,19,30,62,31,231,31,20,31,176,31,220,31,24,31,136,31,241,31,241,30,212,31,40,31,40,30,39,31,178,31,178,30,178,29,204,31,88,31,246,31,249,31,96,31,72,31,208,31,44,31,64,31,161,31,142,31,222,31,189,31,165,31,100,31,119,31,51,31,51,30,71,31,71,30,129,31,209,31,16,31,152,31,31,31,53,31,154,31,154,30,124,31,110,31,110,30,196,31,249,31,20,31,116,31,175,31,181,31,181,30,156,31,217,31,188,31,74,31,187,31,7,31,116,31,193,31,193,30,128,31,70,31,254,31,136,31,112,31,230,31,124,31,124,30,227,31,227,30,196,31,203,31,86,31,129,31,86,31,235,31,39,31,244,31,207,31,207,30,207,29,96,31,131,31,107,31,254,31,254,30,248,31,248,30,8,31,113,31,228,31,228,30,96,31,138,31,138,30,42,31,6,31,28,31,28,30,108,31,80,31,80,30,80,29,215,31,69,31,3,31,196,31,194,31,73,31,3,31,242,31,242,30,62,31,41,31,107,31,238,31,250,31,21,31,52,31,18,31,222,31,73,31,96,31,96,30,108,31,108,30,149,31,95,31,149,31,121,31,23,31,114,31,39,31,106,31,106,30,130,31,219,31,198,31,179,31,179,30,80,31,97,31,198,31,249,31,249,30,214,31,33,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
