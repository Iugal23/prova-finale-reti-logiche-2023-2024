-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 360;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,0,0,227,0,0,0,222,0,107,0,0,0,214,0,161,0,78,0,4,0,112,0,0,0,104,0,0,0,156,0,0,0,0,0,0,0,237,0,15,0,96,0,0,0,168,0,0,0,254,0,197,0,54,0,110,0,7,0,229,0,29,0,138,0,0,0,153,0,67,0,186,0,0,0,0,0,0,0,111,0,199,0,60,0,0,0,94,0,15,0,219,0,222,0,39,0,142,0,150,0,1,0,122,0,42,0,33,0,175,0,213,0,0,0,44,0,136,0,144,0,151,0,170,0,160,0,169,0,243,0,51,0,230,0,95,0,142,0,48,0,138,0,175,0,230,0,75,0,0,0,200,0,0,0,0,0,88,0,213,0,234,0,69,0,0,0,96,0,189,0,125,0,0,0,0,0,104,0,0,0,23,0,243,0,100,0,82,0,85,0,68,0,62,0,152,0,121,0,95,0,0,0,154,0,115,0,173,0,85,0,125,0,0,0,249,0,212,0,154,0,0,0,0,0,0,0,221,0,36,0,0,0,26,0,81,0,161,0,62,0,16,0,217,0,233,0,0,0,0,0,0,0,51,0,140,0,0,0,170,0,30,0,222,0,161,0,252,0,0,0,0,0,0,0,172,0,167,0,0,0,88,0,0,0,144,0,229,0,77,0,221,0,177,0,194,0,27,0,185,0,204,0,198,0,245,0,99,0,12,0,70,0,107,0,47,0,162,0,17,0,3,0,230,0,19,0,183,0,132,0,0,0,71,0,0,0,182,0,46,0,166,0,191,0,87,0,182,0,19,0,218,0,122,0,34,0,71,0,220,0,36,0,93,0,47,0,3,0,116,0,20,0,0,0,183,0,191,0,0,0,211,0,197,0,57,0,41,0,218,0,7,0,0,0,0,0,112,0,194,0,0,0,249,0,0,0,214,0,255,0,242,0,0,0,183,0,32,0,0,0,158,0,76,0,185,0,0,0,127,0,0,0,0,0,234,0,0,0,0,0,0,0,0,0,172,0,2,0,1,0,240,0,235,0,171,0,0,0,40,0,125,0,0,0,155,0,184,0,19,0,120,0,132,0,13,0,0,0,99,0,221,0,168,0,39,0,99,0,0,0,23,0,119,0,0,0,247,0,0,0,117,0,189,0,125,0,138,0,197,0,0,0,57,0,217,0,0,0,130,0,64,0,234,0,18,0,227,0,0,0,187,0,217,0,45,0,150,0,148,0,0,0,0,0,102,0,187,0,0,0,153,0,212,0,30,0,196,0,205,0,0,0,255,0,98,0,0,0,163,0,99,0,123,0,100,0,170,0,0,0,164,0,254,0,0,0,113,0,243,0,224,0,192,0,0,0,155,0,0,0,0,0,8,0,161,0,185,0,232,0,225,0,51,0,0,0,40,0,234,0,251,0,54,0,12,0,85,0,99,0,0,0,38,0,17,0,114,0,0,0,111,0,148,0,75,0,4,0,20,0,76,0,0,0,160,0,116,0,81,0,0,0,87,0,80,0,0,0,166,0,77,0,150,0,171,0,106,0,93,0,66,0,0,0,150,0,0,0,151,0,107,0,0,0,212,0,142,0,0,0,190,0,121,0,129,0,145,0,178,0,254,0,223,0,0,0,63,0);
signal scenario_full  : scenario_type := (133,31,133,30,227,31,227,30,222,31,107,31,107,30,214,31,161,31,78,31,4,31,112,31,112,30,104,31,104,30,156,31,156,30,156,29,156,28,237,31,15,31,96,31,96,30,168,31,168,30,254,31,197,31,54,31,110,31,7,31,229,31,29,31,138,31,138,30,153,31,67,31,186,31,186,30,186,29,186,28,111,31,199,31,60,31,60,30,94,31,15,31,219,31,222,31,39,31,142,31,150,31,1,31,122,31,42,31,33,31,175,31,213,31,213,30,44,31,136,31,144,31,151,31,170,31,160,31,169,31,243,31,51,31,230,31,95,31,142,31,48,31,138,31,175,31,230,31,75,31,75,30,200,31,200,30,200,29,88,31,213,31,234,31,69,31,69,30,96,31,189,31,125,31,125,30,125,29,104,31,104,30,23,31,243,31,100,31,82,31,85,31,68,31,62,31,152,31,121,31,95,31,95,30,154,31,115,31,173,31,85,31,125,31,125,30,249,31,212,31,154,31,154,30,154,29,154,28,221,31,36,31,36,30,26,31,81,31,161,31,62,31,16,31,217,31,233,31,233,30,233,29,233,28,51,31,140,31,140,30,170,31,30,31,222,31,161,31,252,31,252,30,252,29,252,28,172,31,167,31,167,30,88,31,88,30,144,31,229,31,77,31,221,31,177,31,194,31,27,31,185,31,204,31,198,31,245,31,99,31,12,31,70,31,107,31,47,31,162,31,17,31,3,31,230,31,19,31,183,31,132,31,132,30,71,31,71,30,182,31,46,31,166,31,191,31,87,31,182,31,19,31,218,31,122,31,34,31,71,31,220,31,36,31,93,31,47,31,3,31,116,31,20,31,20,30,183,31,191,31,191,30,211,31,197,31,57,31,41,31,218,31,7,31,7,30,7,29,112,31,194,31,194,30,249,31,249,30,214,31,255,31,242,31,242,30,183,31,32,31,32,30,158,31,76,31,185,31,185,30,127,31,127,30,127,29,234,31,234,30,234,29,234,28,234,27,172,31,2,31,1,31,240,31,235,31,171,31,171,30,40,31,125,31,125,30,155,31,184,31,19,31,120,31,132,31,13,31,13,30,99,31,221,31,168,31,39,31,99,31,99,30,23,31,119,31,119,30,247,31,247,30,117,31,189,31,125,31,138,31,197,31,197,30,57,31,217,31,217,30,130,31,64,31,234,31,18,31,227,31,227,30,187,31,217,31,45,31,150,31,148,31,148,30,148,29,102,31,187,31,187,30,153,31,212,31,30,31,196,31,205,31,205,30,255,31,98,31,98,30,163,31,99,31,123,31,100,31,170,31,170,30,164,31,254,31,254,30,113,31,243,31,224,31,192,31,192,30,155,31,155,30,155,29,8,31,161,31,185,31,232,31,225,31,51,31,51,30,40,31,234,31,251,31,54,31,12,31,85,31,99,31,99,30,38,31,17,31,114,31,114,30,111,31,148,31,75,31,4,31,20,31,76,31,76,30,160,31,116,31,81,31,81,30,87,31,80,31,80,30,166,31,77,31,150,31,171,31,106,31,93,31,66,31,66,30,150,31,150,30,151,31,107,31,107,30,212,31,142,31,142,30,190,31,121,31,129,31,145,31,178,31,254,31,223,31,223,30,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
