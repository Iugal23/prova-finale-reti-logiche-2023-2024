-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 776;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,32,0,0,0,238,0,117,0,0,0,177,0,48,0,109,0,0,0,178,0,136,0,160,0,109,0,187,0,154,0,204,0,200,0,0,0,94,0,176,0,139,0,95,0,0,0,89,0,141,0,100,0,211,0,155,0,193,0,18,0,134,0,193,0,0,0,95,0,0,0,83,0,57,0,91,0,72,0,120,0,218,0,245,0,16,0,176,0,75,0,161,0,0,0,55,0,89,0,160,0,112,0,248,0,117,0,0,0,87,0,207,0,171,0,54,0,55,0,217,0,160,0,0,0,38,0,0,0,8,0,22,0,17,0,0,0,139,0,14,0,20,0,183,0,212,0,152,0,0,0,157,0,71,0,85,0,0,0,124,0,5,0,192,0,154,0,31,0,196,0,184,0,58,0,31,0,18,0,0,0,92,0,228,0,91,0,85,0,0,0,0,0,57,0,0,0,19,0,102,0,57,0,161,0,103,0,118,0,117,0,97,0,235,0,124,0,185,0,0,0,117,0,249,0,87,0,230,0,70,0,41,0,190,0,118,0,24,0,0,0,222,0,188,0,0,0,26,0,57,0,253,0,156,0,13,0,62,0,118,0,65,0,218,0,81,0,82,0,246,0,15,0,65,0,22,0,14,0,0,0,61,0,0,0,0,0,223,0,0,0,0,0,253,0,114,0,166,0,0,0,230,0,0,0,0,0,104,0,204,0,47,0,0,0,129,0,158,0,0,0,246,0,205,0,244,0,0,0,0,0,194,0,32,0,90,0,0,0,147,0,37,0,133,0,37,0,212,0,230,0,69,0,255,0,40,0,138,0,11,0,47,0,0,0,0,0,206,0,50,0,252,0,26,0,0,0,64,0,0,0,190,0,141,0,177,0,122,0,238,0,136,0,0,0,182,0,171,0,247,0,219,0,225,0,164,0,92,0,0,0,201,0,217,0,210,0,149,0,0,0,215,0,0,0,230,0,184,0,17,0,6,0,55,0,0,0,7,0,184,0,14,0,0,0,23,0,156,0,148,0,20,0,52,0,55,0,140,0,82,0,21,0,123,0,101,0,144,0,217,0,0,0,0,0,237,0,86,0,59,0,56,0,204,0,235,0,8,0,59,0,152,0,245,0,211,0,46,0,0,0,0,0,13,0,194,0,87,0,111,0,137,0,28,0,196,0,0,0,199,0,0,0,206,0,0,0,82,0,81,0,0,0,77,0,167,0,206,0,218,0,246,0,38,0,131,0,211,0,0,0,0,0,97,0,0,0,4,0,215,0,0,0,155,0,0,0,191,0,172,0,74,0,147,0,0,0,0,0,153,0,170,0,155,0,0,0,17,0,0,0,161,0,185,0,72,0,0,0,221,0,174,0,221,0,201,0,84,0,221,0,94,0,0,0,26,0,0,0,98,0,166,0,253,0,135,0,13,0,238,0,51,0,0,0,138,0,210,0,35,0,120,0,126,0,126,0,11,0,225,0,160,0,248,0,115,0,110,0,0,0,6,0,223,0,249,0,254,0,223,0,199,0,110,0,253,0,228,0,194,0,191,0,213,0,233,0,0,0,152,0,127,0,0,0,146,0,243,0,0,0,32,0,178,0,0,0,100,0,0,0,0,0,57,0,62,0,78,0,207,0,78,0,130,0,210,0,239,0,120,0,202,0,0,0,167,0,174,0,0,0,168,0,35,0,173,0,172,0,85,0,0,0,171,0,214,0,0,0,211,0,196,0,126,0,92,0,208,0,22,0,236,0,155,0,191,0,0,0,209,0,0,0,21,0,10,0,0,0,114,0,238,0,165,0,236,0,90,0,0,0,0,0,184,0,203,0,186,0,212,0,9,0,0,0,213,0,147,0,148,0,153,0,155,0,99,0,9,0,253,0,11,0,233,0,0,0,166,0,86,0,48,0,132,0,252,0,244,0,230,0,0,0,0,0,104,0,79,0,218,0,141,0,0,0,241,0,31,0,214,0,171,0,0,0,66,0,111,0,205,0,214,0,0,0,87,0,0,0,117,0,132,0,54,0,0,0,0,0,163,0,123,0,0,0,202,0,0,0,0,0,0,0,116,0,214,0,243,0,28,0,0,0,150,0,60,0,151,0,194,0,204,0,233,0,32,0,58,0,0,0,216,0,241,0,182,0,2,0,234,0,0,0,0,0,0,0,7,0,127,0,0,0,253,0,91,0,42,0,248,0,0,0,163,0,0,0,205,0,16,0,235,0,136,0,0,0,128,0,83,0,122,0,171,0,143,0,205,0,0,0,99,0,150,0,0,0,196,0,20,0,0,0,23,0,87,0,57,0,74,0,197,0,253,0,49,0,236,0,198,0,40,0,77,0,0,0,88,0,184,0,0,0,20,0,117,0,94,0,48,0,146,0,23,0,23,0,0,0,19,0,10,0,101,0,63,0,33,0,180,0,48,0,135,0,85,0,0,0,0,0,131,0,245,0,123,0,253,0,41,0,112,0,0,0,187,0,0,0,125,0,71,0,204,0,161,0,84,0,110,0,111,0,0,0,212,0,223,0,238,0,53,0,232,0,192,0,142,0,76,0,220,0,0,0,54,0,42,0,226,0,0,0,71,0,243,0,25,0,102,0,17,0,87,0,3,0,0,0,0,0,106,0,52,0,160,0,53,0,199,0,215,0,31,0,191,0,34,0,0,0,57,0,234,0,87,0,190,0,0,0,0,0,120,0,136,0,171,0,160,0,0,0,73,0,114,0,10,0,99,0,142,0,23,0,0,0,113,0,0,0,0,0,18,0,124,0,76,0,13,0,146,0,254,0,158,0,200,0,252,0,137,0,193,0,203,0,60,0,66,0,161,0,201,0,220,0,195,0,141,0,218,0,66,0,54,0,99,0,229,0,227,0,90,0,11,0,234,0,53,0,31,0,175,0,224,0,185,0,0,0,169,0,171,0,16,0,192,0,249,0,29,0,216,0,101,0,131,0,161,0,214,0,119,0,129,0,105,0,109,0,121,0,113,0,152,0,218,0,0,0,91,0,29,0,29,0,59,0,52,0,91,0,157,0,170,0,226,0,96,0,167,0,0,0,0,0,4,0,0,0,221,0,222,0,42,0,33,0,230,0,226,0,67,0,66,0,171,0,0,0,43,0,99,0,61,0,0,0,0,0,8,0,138,0,195,0,61,0,0,0,209,0,60,0,37,0,194,0,117,0,191,0,116,0,95,0,40,0,247,0,153,0,0,0,139,0,184,0,0,0,0,0,105,0,168,0,92,0,126,0,0,0,99,0,56,0,84,0,0,0,216,0,0,0,23,0,50,0,195,0,41,0,25,0,0,0,144,0,211,0,156,0,10,0,173,0,116,0,183,0,77,0,181,0,174,0,0,0,0,0,9,0,14,0,0,0,0,0,224,0,0,0,159,0,9,0,0,0,203,0,0,0,46,0,182,0,45,0,120,0,90,0,138,0,162,0,31,0,71,0,51,0,7,0,0,0,243,0,226,0,225,0,0,0,167,0,6,0,159,0);
signal scenario_full  : scenario_type := (9,31,32,31,32,30,238,31,117,31,117,30,177,31,48,31,109,31,109,30,178,31,136,31,160,31,109,31,187,31,154,31,204,31,200,31,200,30,94,31,176,31,139,31,95,31,95,30,89,31,141,31,100,31,211,31,155,31,193,31,18,31,134,31,193,31,193,30,95,31,95,30,83,31,57,31,91,31,72,31,120,31,218,31,245,31,16,31,176,31,75,31,161,31,161,30,55,31,89,31,160,31,112,31,248,31,117,31,117,30,87,31,207,31,171,31,54,31,55,31,217,31,160,31,160,30,38,31,38,30,8,31,22,31,17,31,17,30,139,31,14,31,20,31,183,31,212,31,152,31,152,30,157,31,71,31,85,31,85,30,124,31,5,31,192,31,154,31,31,31,196,31,184,31,58,31,31,31,18,31,18,30,92,31,228,31,91,31,85,31,85,30,85,29,57,31,57,30,19,31,102,31,57,31,161,31,103,31,118,31,117,31,97,31,235,31,124,31,185,31,185,30,117,31,249,31,87,31,230,31,70,31,41,31,190,31,118,31,24,31,24,30,222,31,188,31,188,30,26,31,57,31,253,31,156,31,13,31,62,31,118,31,65,31,218,31,81,31,82,31,246,31,15,31,65,31,22,31,14,31,14,30,61,31,61,30,61,29,223,31,223,30,223,29,253,31,114,31,166,31,166,30,230,31,230,30,230,29,104,31,204,31,47,31,47,30,129,31,158,31,158,30,246,31,205,31,244,31,244,30,244,29,194,31,32,31,90,31,90,30,147,31,37,31,133,31,37,31,212,31,230,31,69,31,255,31,40,31,138,31,11,31,47,31,47,30,47,29,206,31,50,31,252,31,26,31,26,30,64,31,64,30,190,31,141,31,177,31,122,31,238,31,136,31,136,30,182,31,171,31,247,31,219,31,225,31,164,31,92,31,92,30,201,31,217,31,210,31,149,31,149,30,215,31,215,30,230,31,184,31,17,31,6,31,55,31,55,30,7,31,184,31,14,31,14,30,23,31,156,31,148,31,20,31,52,31,55,31,140,31,82,31,21,31,123,31,101,31,144,31,217,31,217,30,217,29,237,31,86,31,59,31,56,31,204,31,235,31,8,31,59,31,152,31,245,31,211,31,46,31,46,30,46,29,13,31,194,31,87,31,111,31,137,31,28,31,196,31,196,30,199,31,199,30,206,31,206,30,82,31,81,31,81,30,77,31,167,31,206,31,218,31,246,31,38,31,131,31,211,31,211,30,211,29,97,31,97,30,4,31,215,31,215,30,155,31,155,30,191,31,172,31,74,31,147,31,147,30,147,29,153,31,170,31,155,31,155,30,17,31,17,30,161,31,185,31,72,31,72,30,221,31,174,31,221,31,201,31,84,31,221,31,94,31,94,30,26,31,26,30,98,31,166,31,253,31,135,31,13,31,238,31,51,31,51,30,138,31,210,31,35,31,120,31,126,31,126,31,11,31,225,31,160,31,248,31,115,31,110,31,110,30,6,31,223,31,249,31,254,31,223,31,199,31,110,31,253,31,228,31,194,31,191,31,213,31,233,31,233,30,152,31,127,31,127,30,146,31,243,31,243,30,32,31,178,31,178,30,100,31,100,30,100,29,57,31,62,31,78,31,207,31,78,31,130,31,210,31,239,31,120,31,202,31,202,30,167,31,174,31,174,30,168,31,35,31,173,31,172,31,85,31,85,30,171,31,214,31,214,30,211,31,196,31,126,31,92,31,208,31,22,31,236,31,155,31,191,31,191,30,209,31,209,30,21,31,10,31,10,30,114,31,238,31,165,31,236,31,90,31,90,30,90,29,184,31,203,31,186,31,212,31,9,31,9,30,213,31,147,31,148,31,153,31,155,31,99,31,9,31,253,31,11,31,233,31,233,30,166,31,86,31,48,31,132,31,252,31,244,31,230,31,230,30,230,29,104,31,79,31,218,31,141,31,141,30,241,31,31,31,214,31,171,31,171,30,66,31,111,31,205,31,214,31,214,30,87,31,87,30,117,31,132,31,54,31,54,30,54,29,163,31,123,31,123,30,202,31,202,30,202,29,202,28,116,31,214,31,243,31,28,31,28,30,150,31,60,31,151,31,194,31,204,31,233,31,32,31,58,31,58,30,216,31,241,31,182,31,2,31,234,31,234,30,234,29,234,28,7,31,127,31,127,30,253,31,91,31,42,31,248,31,248,30,163,31,163,30,205,31,16,31,235,31,136,31,136,30,128,31,83,31,122,31,171,31,143,31,205,31,205,30,99,31,150,31,150,30,196,31,20,31,20,30,23,31,87,31,57,31,74,31,197,31,253,31,49,31,236,31,198,31,40,31,77,31,77,30,88,31,184,31,184,30,20,31,117,31,94,31,48,31,146,31,23,31,23,31,23,30,19,31,10,31,101,31,63,31,33,31,180,31,48,31,135,31,85,31,85,30,85,29,131,31,245,31,123,31,253,31,41,31,112,31,112,30,187,31,187,30,125,31,71,31,204,31,161,31,84,31,110,31,111,31,111,30,212,31,223,31,238,31,53,31,232,31,192,31,142,31,76,31,220,31,220,30,54,31,42,31,226,31,226,30,71,31,243,31,25,31,102,31,17,31,87,31,3,31,3,30,3,29,106,31,52,31,160,31,53,31,199,31,215,31,31,31,191,31,34,31,34,30,57,31,234,31,87,31,190,31,190,30,190,29,120,31,136,31,171,31,160,31,160,30,73,31,114,31,10,31,99,31,142,31,23,31,23,30,113,31,113,30,113,29,18,31,124,31,76,31,13,31,146,31,254,31,158,31,200,31,252,31,137,31,193,31,203,31,60,31,66,31,161,31,201,31,220,31,195,31,141,31,218,31,66,31,54,31,99,31,229,31,227,31,90,31,11,31,234,31,53,31,31,31,175,31,224,31,185,31,185,30,169,31,171,31,16,31,192,31,249,31,29,31,216,31,101,31,131,31,161,31,214,31,119,31,129,31,105,31,109,31,121,31,113,31,152,31,218,31,218,30,91,31,29,31,29,31,59,31,52,31,91,31,157,31,170,31,226,31,96,31,167,31,167,30,167,29,4,31,4,30,221,31,222,31,42,31,33,31,230,31,226,31,67,31,66,31,171,31,171,30,43,31,99,31,61,31,61,30,61,29,8,31,138,31,195,31,61,31,61,30,209,31,60,31,37,31,194,31,117,31,191,31,116,31,95,31,40,31,247,31,153,31,153,30,139,31,184,31,184,30,184,29,105,31,168,31,92,31,126,31,126,30,99,31,56,31,84,31,84,30,216,31,216,30,23,31,50,31,195,31,41,31,25,31,25,30,144,31,211,31,156,31,10,31,173,31,116,31,183,31,77,31,181,31,174,31,174,30,174,29,9,31,14,31,14,30,14,29,224,31,224,30,159,31,9,31,9,30,203,31,203,30,46,31,182,31,45,31,120,31,90,31,138,31,162,31,31,31,71,31,51,31,7,31,7,30,243,31,226,31,225,31,225,30,167,31,6,31,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
