-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 902;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (74,0,143,0,65,0,0,0,102,0,212,0,0,0,73,0,0,0,17,0,18,0,197,0,71,0,0,0,147,0,89,0,0,0,129,0,51,0,231,0,162,0,0,0,0,0,29,0,122,0,212,0,74,0,30,0,0,0,229,0,0,0,128,0,0,0,0,0,124,0,0,0,110,0,68,0,0,0,190,0,73,0,169,0,31,0,228,0,28,0,228,0,141,0,216,0,15,0,122,0,131,0,206,0,67,0,126,0,91,0,130,0,42,0,193,0,121,0,0,0,252,0,42,0,145,0,0,0,133,0,241,0,60,0,100,0,229,0,0,0,4,0,254,0,52,0,84,0,222,0,59,0,12,0,0,0,95,0,149,0,193,0,49,0,22,0,112,0,37,0,8,0,55,0,118,0,90,0,75,0,152,0,0,0,11,0,182,0,246,0,240,0,60,0,31,0,228,0,155,0,23,0,158,0,214,0,49,0,0,0,157,0,0,0,100,0,0,0,213,0,3,0,241,0,35,0,161,0,155,0,196,0,213,0,39,0,59,0,0,0,58,0,43,0,9,0,199,0,126,0,221,0,33,0,103,0,148,0,169,0,0,0,0,0,165,0,40,0,201,0,4,0,107,0,233,0,244,0,137,0,231,0,0,0,57,0,0,0,185,0,130,0,60,0,22,0,20,0,159,0,0,0,218,0,99,0,0,0,0,0,153,0,55,0,196,0,109,0,0,0,0,0,0,0,40,0,178,0,131,0,254,0,100,0,39,0,0,0,60,0,200,0,139,0,190,0,0,0,36,0,13,0,73,0,116,0,42,0,0,0,0,0,6,0,126,0,92,0,61,0,248,0,150,0,93,0,0,0,136,0,61,0,21,0,103,0,216,0,50,0,0,0,0,0,66,0,207,0,72,0,231,0,0,0,0,0,0,0,115,0,18,0,32,0,194,0,0,0,128,0,0,0,248,0,154,0,0,0,15,0,204,0,165,0,193,0,181,0,169,0,175,0,54,0,248,0,115,0,239,0,240,0,56,0,52,0,97,0,0,0,124,0,97,0,0,0,4,0,0,0,122,0,32,0,167,0,0,0,234,0,0,0,110,0,171,0,57,0,0,0,0,0,138,0,172,0,97,0,85,0,194,0,48,0,16,0,178,0,76,0,12,0,136,0,3,0,195,0,4,0,0,0,173,0,51,0,0,0,0,0,162,0,145,0,246,0,188,0,106,0,234,0,194,0,238,0,10,0,129,0,0,0,0,0,82,0,234,0,114,0,53,0,91,0,0,0,25,0,139,0,121,0,219,0,225,0,114,0,29,0,96,0,66,0,134,0,0,0,182,0,14,0,211,0,76,0,51,0,21,0,174,0,134,0,13,0,12,0,38,0,8,0,0,0,54,0,187,0,150,0,0,0,237,0,173,0,210,0,0,0,65,0,156,0,58,0,0,0,221,0,32,0,188,0,0,0,226,0,172,0,163,0,188,0,0,0,199,0,7,0,188,0,195,0,9,0,99,0,22,0,65,0,73,0,13,0,0,0,243,0,246,0,10,0,197,0,0,0,95,0,94,0,167,0,0,0,152,0,86,0,0,0,50,0,0,0,70,0,255,0,73,0,226,0,212,0,0,0,216,0,0,0,87,0,0,0,0,0,0,0,8,0,0,0,250,0,11,0,33,0,173,0,153,0,0,0,133,0,99,0,9,0,186,0,104,0,0,0,85,0,126,0,210,0,52,0,212,0,77,0,14,0,111,0,0,0,192,0,121,0,0,0,170,0,154,0,0,0,12,0,29,0,46,0,218,0,85,0,88,0,135,0,0,0,0,0,89,0,35,0,95,0,182,0,189,0,76,0,0,0,0,0,2,0,78,0,0,0,0,0,0,0,142,0,0,0,180,0,183,0,0,0,55,0,129,0,176,0,47,0,220,0,0,0,181,0,109,0,228,0,174,0,0,0,72,0,214,0,154,0,178,0,0,0,0,0,57,0,85,0,0,0,72,0,172,0,0,0,26,0,0,0,248,0,173,0,253,0,165,0,118,0,79,0,168,0,108,0,192,0,0,0,0,0,138,0,165,0,76,0,63,0,134,0,188,0,128,0,99,0,27,0,157,0,0,0,0,0,43,0,137,0,0,0,194,0,108,0,0,0,49,0,70,0,142,0,0,0,132,0,53,0,75,0,0,0,102,0,141,0,247,0,64,0,0,0,205,0,217,0,188,0,116,0,106,0,0,0,30,0,0,0,11,0,204,0,80,0,159,0,26,0,85,0,162,0,64,0,0,0,96,0,75,0,0,0,216,0,153,0,0,0,216,0,0,0,248,0,31,0,49,0,0,0,43,0,229,0,231,0,220,0,196,0,0,0,0,0,0,0,55,0,221,0,139,0,83,0,0,0,0,0,126,0,224,0,218,0,125,0,153,0,191,0,153,0,125,0,235,0,166,0,124,0,13,0,99,0,62,0,131,0,96,0,210,0,177,0,16,0,153,0,42,0,66,0,0,0,184,0,132,0,184,0,0,0,244,0,37,0,214,0,232,0,122,0,40,0,0,0,57,0,127,0,224,0,121,0,129,0,5,0,133,0,101,0,184,0,47,0,69,0,246,0,205,0,0,0,0,0,118,0,122,0,208,0,0,0,191,0,235,0,5,0,209,0,130,0,219,0,0,0,0,0,202,0,148,0,0,0,76,0,111,0,19,0,0,0,0,0,108,0,136,0,202,0,163,0,131,0,152,0,0,0,94,0,30,0,0,0,0,0,0,0,37,0,22,0,0,0,40,0,244,0,0,0,50,0,223,0,45,0,39,0,0,0,106,0,164,0,168,0,146,0,115,0,52,0,0,0,118,0,78,0,28,0,149,0,12,0,160,0,177,0,195,0,0,0,142,0,142,0,227,0,168,0,140,0,0,0,2,0,0,0,0,0,78,0,28,0,177,0,252,0,221,0,229,0,116,0,94,0,100,0,229,0,54,0,18,0,0,0,233,0,142,0,161,0,89,0,125,0,83,0,56,0,36,0,112,0,190,0,238,0,0,0,240,0,110,0,245,0,225,0,57,0,0,0,97,0,23,0,0,0,53,0,123,0,113,0,0,0,40,0,25,0,241,0,135,0,60,0,237,0,1,0,215,0,248,0,235,0,0,0,251,0,251,0,198,0,205,0,80,0,59,0,237,0,0,0,149,0,0,0,0,0,16,0,104,0,159,0,62,0,85,0,96,0,0,0,166,0,110,0,0,0,25,0,59,0,0,0,148,0,203,0,145,0,138,0,68,0,177,0,113,0,0,0,164,0,2,0,0,0,30,0,185,0,169,0,72,0,55,0,0,0,66,0,230,0,56,0,113,0,0,0,213,0,191,0,0,0,239,0,161,0,0,0,0,0,201,0,252,0,238,0,190,0,91,0,80,0,29,0,227,0,117,0,0,0,53,0,101,0,13,0,170,0,0,0,233,0,0,0,184,0,89,0,209,0,138,0,152,0,133,0,232,0,0,0,212,0,14,0,136,0,206,0,0,0,84,0,0,0,1,0,61,0,53,0,22,0,0,0,90,0,157,0,0,0,0,0,182,0,78,0,103,0,97,0,0,0,142,0,66,0,39,0,56,0,66,0,46,0,0,0,50,0,0,0,229,0,115,0,214,0,208,0,213,0,237,0,224,0,227,0,186,0,190,0,76,0,108,0,0,0,13,0,0,0,110,0,210,0,244,0,252,0,129,0,110,0,144,0,184,0,0,0,29,0,0,0,0,0,58,0,200,0,106,0,208,0,192,0,187,0,167,0,10,0,74,0,0,0,56,0,76,0,146,0,184,0,0,0,75,0,50,0,215,0,0,0,197,0,102,0,52,0,127,0,65,0,0,0,126,0,0,0,238,0,172,0,38,0,175,0,209,0,0,0,0,0,142,0,0,0,18,0,244,0,179,0,108,0,0,0,231,0,158,0,0,0,5,0,141,0,216,0,163,0,195,0,154,0,0,0,87,0,137,0,0,0,13,0,0,0,32,0,194,0,81,0,70,0,226,0,137,0,130,0,22,0,0,0,148,0,138,0,79,0,104,0,152,0);
signal scenario_full  : scenario_type := (74,31,143,31,65,31,65,30,102,31,212,31,212,30,73,31,73,30,17,31,18,31,197,31,71,31,71,30,147,31,89,31,89,30,129,31,51,31,231,31,162,31,162,30,162,29,29,31,122,31,212,31,74,31,30,31,30,30,229,31,229,30,128,31,128,30,128,29,124,31,124,30,110,31,68,31,68,30,190,31,73,31,169,31,31,31,228,31,28,31,228,31,141,31,216,31,15,31,122,31,131,31,206,31,67,31,126,31,91,31,130,31,42,31,193,31,121,31,121,30,252,31,42,31,145,31,145,30,133,31,241,31,60,31,100,31,229,31,229,30,4,31,254,31,52,31,84,31,222,31,59,31,12,31,12,30,95,31,149,31,193,31,49,31,22,31,112,31,37,31,8,31,55,31,118,31,90,31,75,31,152,31,152,30,11,31,182,31,246,31,240,31,60,31,31,31,228,31,155,31,23,31,158,31,214,31,49,31,49,30,157,31,157,30,100,31,100,30,213,31,3,31,241,31,35,31,161,31,155,31,196,31,213,31,39,31,59,31,59,30,58,31,43,31,9,31,199,31,126,31,221,31,33,31,103,31,148,31,169,31,169,30,169,29,165,31,40,31,201,31,4,31,107,31,233,31,244,31,137,31,231,31,231,30,57,31,57,30,185,31,130,31,60,31,22,31,20,31,159,31,159,30,218,31,99,31,99,30,99,29,153,31,55,31,196,31,109,31,109,30,109,29,109,28,40,31,178,31,131,31,254,31,100,31,39,31,39,30,60,31,200,31,139,31,190,31,190,30,36,31,13,31,73,31,116,31,42,31,42,30,42,29,6,31,126,31,92,31,61,31,248,31,150,31,93,31,93,30,136,31,61,31,21,31,103,31,216,31,50,31,50,30,50,29,66,31,207,31,72,31,231,31,231,30,231,29,231,28,115,31,18,31,32,31,194,31,194,30,128,31,128,30,248,31,154,31,154,30,15,31,204,31,165,31,193,31,181,31,169,31,175,31,54,31,248,31,115,31,239,31,240,31,56,31,52,31,97,31,97,30,124,31,97,31,97,30,4,31,4,30,122,31,32,31,167,31,167,30,234,31,234,30,110,31,171,31,57,31,57,30,57,29,138,31,172,31,97,31,85,31,194,31,48,31,16,31,178,31,76,31,12,31,136,31,3,31,195,31,4,31,4,30,173,31,51,31,51,30,51,29,162,31,145,31,246,31,188,31,106,31,234,31,194,31,238,31,10,31,129,31,129,30,129,29,82,31,234,31,114,31,53,31,91,31,91,30,25,31,139,31,121,31,219,31,225,31,114,31,29,31,96,31,66,31,134,31,134,30,182,31,14,31,211,31,76,31,51,31,21,31,174,31,134,31,13,31,12,31,38,31,8,31,8,30,54,31,187,31,150,31,150,30,237,31,173,31,210,31,210,30,65,31,156,31,58,31,58,30,221,31,32,31,188,31,188,30,226,31,172,31,163,31,188,31,188,30,199,31,7,31,188,31,195,31,9,31,99,31,22,31,65,31,73,31,13,31,13,30,243,31,246,31,10,31,197,31,197,30,95,31,94,31,167,31,167,30,152,31,86,31,86,30,50,31,50,30,70,31,255,31,73,31,226,31,212,31,212,30,216,31,216,30,87,31,87,30,87,29,87,28,8,31,8,30,250,31,11,31,33,31,173,31,153,31,153,30,133,31,99,31,9,31,186,31,104,31,104,30,85,31,126,31,210,31,52,31,212,31,77,31,14,31,111,31,111,30,192,31,121,31,121,30,170,31,154,31,154,30,12,31,29,31,46,31,218,31,85,31,88,31,135,31,135,30,135,29,89,31,35,31,95,31,182,31,189,31,76,31,76,30,76,29,2,31,78,31,78,30,78,29,78,28,142,31,142,30,180,31,183,31,183,30,55,31,129,31,176,31,47,31,220,31,220,30,181,31,109,31,228,31,174,31,174,30,72,31,214,31,154,31,178,31,178,30,178,29,57,31,85,31,85,30,72,31,172,31,172,30,26,31,26,30,248,31,173,31,253,31,165,31,118,31,79,31,168,31,108,31,192,31,192,30,192,29,138,31,165,31,76,31,63,31,134,31,188,31,128,31,99,31,27,31,157,31,157,30,157,29,43,31,137,31,137,30,194,31,108,31,108,30,49,31,70,31,142,31,142,30,132,31,53,31,75,31,75,30,102,31,141,31,247,31,64,31,64,30,205,31,217,31,188,31,116,31,106,31,106,30,30,31,30,30,11,31,204,31,80,31,159,31,26,31,85,31,162,31,64,31,64,30,96,31,75,31,75,30,216,31,153,31,153,30,216,31,216,30,248,31,31,31,49,31,49,30,43,31,229,31,231,31,220,31,196,31,196,30,196,29,196,28,55,31,221,31,139,31,83,31,83,30,83,29,126,31,224,31,218,31,125,31,153,31,191,31,153,31,125,31,235,31,166,31,124,31,13,31,99,31,62,31,131,31,96,31,210,31,177,31,16,31,153,31,42,31,66,31,66,30,184,31,132,31,184,31,184,30,244,31,37,31,214,31,232,31,122,31,40,31,40,30,57,31,127,31,224,31,121,31,129,31,5,31,133,31,101,31,184,31,47,31,69,31,246,31,205,31,205,30,205,29,118,31,122,31,208,31,208,30,191,31,235,31,5,31,209,31,130,31,219,31,219,30,219,29,202,31,148,31,148,30,76,31,111,31,19,31,19,30,19,29,108,31,136,31,202,31,163,31,131,31,152,31,152,30,94,31,30,31,30,30,30,29,30,28,37,31,22,31,22,30,40,31,244,31,244,30,50,31,223,31,45,31,39,31,39,30,106,31,164,31,168,31,146,31,115,31,52,31,52,30,118,31,78,31,28,31,149,31,12,31,160,31,177,31,195,31,195,30,142,31,142,31,227,31,168,31,140,31,140,30,2,31,2,30,2,29,78,31,28,31,177,31,252,31,221,31,229,31,116,31,94,31,100,31,229,31,54,31,18,31,18,30,233,31,142,31,161,31,89,31,125,31,83,31,56,31,36,31,112,31,190,31,238,31,238,30,240,31,110,31,245,31,225,31,57,31,57,30,97,31,23,31,23,30,53,31,123,31,113,31,113,30,40,31,25,31,241,31,135,31,60,31,237,31,1,31,215,31,248,31,235,31,235,30,251,31,251,31,198,31,205,31,80,31,59,31,237,31,237,30,149,31,149,30,149,29,16,31,104,31,159,31,62,31,85,31,96,31,96,30,166,31,110,31,110,30,25,31,59,31,59,30,148,31,203,31,145,31,138,31,68,31,177,31,113,31,113,30,164,31,2,31,2,30,30,31,185,31,169,31,72,31,55,31,55,30,66,31,230,31,56,31,113,31,113,30,213,31,191,31,191,30,239,31,161,31,161,30,161,29,201,31,252,31,238,31,190,31,91,31,80,31,29,31,227,31,117,31,117,30,53,31,101,31,13,31,170,31,170,30,233,31,233,30,184,31,89,31,209,31,138,31,152,31,133,31,232,31,232,30,212,31,14,31,136,31,206,31,206,30,84,31,84,30,1,31,61,31,53,31,22,31,22,30,90,31,157,31,157,30,157,29,182,31,78,31,103,31,97,31,97,30,142,31,66,31,39,31,56,31,66,31,46,31,46,30,50,31,50,30,229,31,115,31,214,31,208,31,213,31,237,31,224,31,227,31,186,31,190,31,76,31,108,31,108,30,13,31,13,30,110,31,210,31,244,31,252,31,129,31,110,31,144,31,184,31,184,30,29,31,29,30,29,29,58,31,200,31,106,31,208,31,192,31,187,31,167,31,10,31,74,31,74,30,56,31,76,31,146,31,184,31,184,30,75,31,50,31,215,31,215,30,197,31,102,31,52,31,127,31,65,31,65,30,126,31,126,30,238,31,172,31,38,31,175,31,209,31,209,30,209,29,142,31,142,30,18,31,244,31,179,31,108,31,108,30,231,31,158,31,158,30,5,31,141,31,216,31,163,31,195,31,154,31,154,30,87,31,137,31,137,30,13,31,13,30,32,31,194,31,81,31,70,31,226,31,137,31,130,31,22,31,22,30,148,31,138,31,79,31,104,31,152,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
