-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_487 is
end project_tb_487;

architecture project_tb_arch_487 of project_tb_487 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 873;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,147,0,177,0,171,0,0,0,112,0,0,0,0,0,165,0,129,0,200,0,41,0,41,0,128,0,2,0,213,0,141,0,239,0,153,0,150,0,0,0,241,0,55,0,211,0,205,0,0,0,222,0,172,0,68,0,7,0,0,0,0,0,0,0,0,0,145,0,46,0,228,0,0,0,205,0,0,0,53,0,0,0,208,0,148,0,0,0,94,0,128,0,94,0,182,0,117,0,2,0,133,0,126,0,244,0,0,0,10,0,173,0,15,0,16,0,0,0,87,0,192,0,176,0,187,0,28,0,28,0,0,0,214,0,32,0,172,0,157,0,141,0,0,0,114,0,136,0,245,0,0,0,48,0,40,0,226,0,8,0,0,0,108,0,123,0,41,0,23,0,169,0,221,0,41,0,66,0,211,0,0,0,73,0,0,0,83,0,0,0,183,0,205,0,0,0,0,0,129,0,0,0,212,0,138,0,0,0,129,0,35,0,214,0,81,0,173,0,0,0,39,0,227,0,60,0,36,0,241,0,120,0,96,0,43,0,0,0,52,0,0,0,220,0,167,0,84,0,214,0,44,0,253,0,132,0,99,0,243,0,0,0,0,0,180,0,70,0,102,0,180,0,7,0,113,0,110,0,0,0,198,0,86,0,105,0,50,0,0,0,0,0,132,0,49,0,111,0,147,0,137,0,150,0,0,0,0,0,37,0,250,0,76,0,98,0,168,0,172,0,193,0,187,0,24,0,40,0,157,0,14,0,171,0,199,0,50,0,81,0,42,0,33,0,132,0,0,0,0,0,131,0,198,0,121,0,0,0,102,0,0,0,243,0,0,0,128,0,101,0,0,0,0,0,0,0,45,0,147,0,105,0,17,0,0,0,42,0,245,0,5,0,0,0,0,0,152,0,90,0,194,0,0,0,0,0,6,0,0,0,201,0,78,0,87,0,0,0,86,0,76,0,132,0,249,0,113,0,38,0,70,0,0,0,83,0,97,0,0,0,0,0,22,0,60,0,76,0,0,0,36,0,212,0,227,0,24,0,70,0,210,0,35,0,155,0,80,0,13,0,76,0,0,0,130,0,0,0,27,0,244,0,0,0,0,0,20,0,0,0,0,0,138,0,0,0,0,0,0,0,134,0,78,0,239,0,64,0,0,0,22,0,42,0,191,0,55,0,0,0,0,0,208,0,224,0,124,0,0,0,205,0,213,0,0,0,107,0,51,0,49,0,24,0,129,0,75,0,19,0,145,0,0,0,242,0,194,0,142,0,213,0,176,0,232,0,16,0,47,0,172,0,245,0,108,0,232,0,241,0,0,0,135,0,95,0,39,0,96,0,182,0,0,0,0,0,0,0,117,0,227,0,0,0,17,0,0,0,2,0,191,0,232,0,33,0,101,0,61,0,205,0,6,0,146,0,115,0,141,0,135,0,7,0,0,0,86,0,34,0,77,0,199,0,148,0,225,0,232,0,121,0,57,0,82,0,55,0,34,0,0,0,0,0,209,0,90,0,169,0,22,0,93,0,60,0,160,0,29,0,22,0,69,0,107,0,0,0,0,0,214,0,46,0,7,0,245,0,141,0,199,0,5,0,218,0,184,0,60,0,252,0,199,0,29,0,247,0,102,0,23,0,114,0,150,0,251,0,0,0,172,0,79,0,168,0,198,0,29,0,124,0,130,0,204,0,0,0,62,0,84,0,146,0,191,0,128,0,2,0,102,0,0,0,2,0,227,0,118,0,0,0,131,0,0,0,140,0,194,0,218,0,128,0,242,0,1,0,168,0,64,0,17,0,57,0,146,0,73,0,0,0,106,0,57,0,0,0,222,0,251,0,242,0,0,0,123,0,228,0,143,0,128,0,99,0,24,0,255,0,33,0,183,0,244,0,109,0,16,0,90,0,120,0,46,0,215,0,211,0,60,0,172,0,189,0,0,0,220,0,104,0,85,0,11,0,0,0,0,0,21,0,77,0,217,0,199,0,49,0,199,0,67,0,0,0,184,0,43,0,0,0,93,0,199,0,209,0,83,0,215,0,212,0,0,0,142,0,84,0,121,0,0,0,120,0,153,0,29,0,144,0,5,0,0,0,35,0,52,0,0,0,89,0,0,0,0,0,225,0,240,0,19,0,167,0,254,0,199,0,51,0,55,0,171,0,195,0,0,0,0,0,177,0,7,0,0,0,113,0,57,0,85,0,0,0,43,0,0,0,148,0,43,0,22,0,176,0,18,0,134,0,60,0,116,0,117,0,0,0,224,0,0,0,226,0,91,0,51,0,134,0,218,0,150,0,124,0,92,0,209,0,214,0,101,0,56,0,208,0,255,0,238,0,210,0,252,0,150,0,89,0,0,0,0,0,98,0,198,0,239,0,142,0,0,0,24,0,47,0,205,0,43,0,0,0,169,0,232,0,158,0,84,0,218,0,153,0,37,0,38,0,247,0,242,0,163,0,0,0,167,0,79,0,200,0,185,0,236,0,172,0,9,0,0,0,0,0,139,0,74,0,190,0,8,0,155,0,105,0,125,0,114,0,0,0,235,0,125,0,164,0,96,0,169,0,0,0,128,0,148,0,146,0,0,0,0,0,223,0,0,0,76,0,0,0,53,0,3,0,215,0,216,0,183,0,121,0,49,0,150,0,62,0,225,0,16,0,27,0,0,0,33,0,0,0,1,0,86,0,46,0,0,0,64,0,91,0,151,0,0,0,82,0,30,0,117,0,186,0,101,0,87,0,0,0,161,0,170,0,140,0,17,0,146,0,62,0,130,0,22,0,117,0,128,0,59,0,0,0,150,0,95,0,185,0,182,0,0,0,125,0,177,0,173,0,85,0,60,0,133,0,167,0,0,0,138,0,140,0,160,0,152,0,208,0,136,0,53,0,28,0,196,0,0,0,93,0,46,0,71,0,0,0,62,0,126,0,223,0,224,0,23,0,203,0,145,0,63,0,251,0,243,0,9,0,188,0,146,0,63,0,197,0,209,0,102,0,0,0,205,0,0,0,91,0,143,0,64,0,199,0,212,0,183,0,48,0,68,0,219,0,45,0,0,0,41,0,0,0,174,0,137,0,3,0,0,0,92,0,0,0,3,0,213,0,185,0,152,0,253,0,0,0,243,0,32,0,58,0,184,0,69,0,77,0,0,0,0,0,74,0,11,0,156,0,0,0,181,0,97,0,120,0,0,0,185,0,193,0,77,0,29,0,28,0,163,0,83,0,228,0,87,0,0,0,41,0,72,0,77,0,0,0,107,0,169,0,0,0,138,0,34,0,1,0,24,0,60,0,57,0,55,0,108,0,27,0,73,0,188,0,234,0,54,0,32,0,0,0,0,0,3,0,0,0,122,0,84,0,217,0,226,0,91,0,80,0,193,0,219,0,69,0,77,0,102,0,222,0,189,0,194,0,236,0,227,0,117,0,219,0,0,0,250,0,82,0,182,0,228,0,188,0,109,0,0,0,247,0,231,0,47,0,75,0,182,0,92,0,244,0,31,0,139,0,206,0,249,0,0,0,233,0,28,0,0,0,46,0,8,0,166,0,0,0,73,0,12,0,221,0,90,0,0,0,252,0,80,0,110,0,190,0,166,0,0,0,123,0,0,0,105,0,28,0,0,0,63,0,31,0,201,0,176,0,235,0,252,0,132,0,217,0,87,0,0,0,3,0,198,0,0,0,0,0,187,0,231,0,0,0,250,0,187,0,206,0,31,0,0,0,0,0,0,0,0,0,0,0,85,0,107,0,200,0,0,0,43,0,77,0,61,0,124,0,63,0,0,0,0,0,231,0,0,0,145,0,0,0,27,0,181,0,194,0,121,0,0,0,108,0,87,0,169,0,141,0,187,0,32,0,128,0,15,0,249,0,242,0,0,0,123,0,122,0,31,0,0,0,128,0,113,0,178,0,200,0,160,0,5,0,185,0);
signal scenario_full  : scenario_type := (0,0,147,31,177,31,171,31,171,30,112,31,112,30,112,29,165,31,129,31,200,31,41,31,41,31,128,31,2,31,213,31,141,31,239,31,153,31,150,31,150,30,241,31,55,31,211,31,205,31,205,30,222,31,172,31,68,31,7,31,7,30,7,29,7,28,7,27,145,31,46,31,228,31,228,30,205,31,205,30,53,31,53,30,208,31,148,31,148,30,94,31,128,31,94,31,182,31,117,31,2,31,133,31,126,31,244,31,244,30,10,31,173,31,15,31,16,31,16,30,87,31,192,31,176,31,187,31,28,31,28,31,28,30,214,31,32,31,172,31,157,31,141,31,141,30,114,31,136,31,245,31,245,30,48,31,40,31,226,31,8,31,8,30,108,31,123,31,41,31,23,31,169,31,221,31,41,31,66,31,211,31,211,30,73,31,73,30,83,31,83,30,183,31,205,31,205,30,205,29,129,31,129,30,212,31,138,31,138,30,129,31,35,31,214,31,81,31,173,31,173,30,39,31,227,31,60,31,36,31,241,31,120,31,96,31,43,31,43,30,52,31,52,30,220,31,167,31,84,31,214,31,44,31,253,31,132,31,99,31,243,31,243,30,243,29,180,31,70,31,102,31,180,31,7,31,113,31,110,31,110,30,198,31,86,31,105,31,50,31,50,30,50,29,132,31,49,31,111,31,147,31,137,31,150,31,150,30,150,29,37,31,250,31,76,31,98,31,168,31,172,31,193,31,187,31,24,31,40,31,157,31,14,31,171,31,199,31,50,31,81,31,42,31,33,31,132,31,132,30,132,29,131,31,198,31,121,31,121,30,102,31,102,30,243,31,243,30,128,31,101,31,101,30,101,29,101,28,45,31,147,31,105,31,17,31,17,30,42,31,245,31,5,31,5,30,5,29,152,31,90,31,194,31,194,30,194,29,6,31,6,30,201,31,78,31,87,31,87,30,86,31,76,31,132,31,249,31,113,31,38,31,70,31,70,30,83,31,97,31,97,30,97,29,22,31,60,31,76,31,76,30,36,31,212,31,227,31,24,31,70,31,210,31,35,31,155,31,80,31,13,31,76,31,76,30,130,31,130,30,27,31,244,31,244,30,244,29,20,31,20,30,20,29,138,31,138,30,138,29,138,28,134,31,78,31,239,31,64,31,64,30,22,31,42,31,191,31,55,31,55,30,55,29,208,31,224,31,124,31,124,30,205,31,213,31,213,30,107,31,51,31,49,31,24,31,129,31,75,31,19,31,145,31,145,30,242,31,194,31,142,31,213,31,176,31,232,31,16,31,47,31,172,31,245,31,108,31,232,31,241,31,241,30,135,31,95,31,39,31,96,31,182,31,182,30,182,29,182,28,117,31,227,31,227,30,17,31,17,30,2,31,191,31,232,31,33,31,101,31,61,31,205,31,6,31,146,31,115,31,141,31,135,31,7,31,7,30,86,31,34,31,77,31,199,31,148,31,225,31,232,31,121,31,57,31,82,31,55,31,34,31,34,30,34,29,209,31,90,31,169,31,22,31,93,31,60,31,160,31,29,31,22,31,69,31,107,31,107,30,107,29,214,31,46,31,7,31,245,31,141,31,199,31,5,31,218,31,184,31,60,31,252,31,199,31,29,31,247,31,102,31,23,31,114,31,150,31,251,31,251,30,172,31,79,31,168,31,198,31,29,31,124,31,130,31,204,31,204,30,62,31,84,31,146,31,191,31,128,31,2,31,102,31,102,30,2,31,227,31,118,31,118,30,131,31,131,30,140,31,194,31,218,31,128,31,242,31,1,31,168,31,64,31,17,31,57,31,146,31,73,31,73,30,106,31,57,31,57,30,222,31,251,31,242,31,242,30,123,31,228,31,143,31,128,31,99,31,24,31,255,31,33,31,183,31,244,31,109,31,16,31,90,31,120,31,46,31,215,31,211,31,60,31,172,31,189,31,189,30,220,31,104,31,85,31,11,31,11,30,11,29,21,31,77,31,217,31,199,31,49,31,199,31,67,31,67,30,184,31,43,31,43,30,93,31,199,31,209,31,83,31,215,31,212,31,212,30,142,31,84,31,121,31,121,30,120,31,153,31,29,31,144,31,5,31,5,30,35,31,52,31,52,30,89,31,89,30,89,29,225,31,240,31,19,31,167,31,254,31,199,31,51,31,55,31,171,31,195,31,195,30,195,29,177,31,7,31,7,30,113,31,57,31,85,31,85,30,43,31,43,30,148,31,43,31,22,31,176,31,18,31,134,31,60,31,116,31,117,31,117,30,224,31,224,30,226,31,91,31,51,31,134,31,218,31,150,31,124,31,92,31,209,31,214,31,101,31,56,31,208,31,255,31,238,31,210,31,252,31,150,31,89,31,89,30,89,29,98,31,198,31,239,31,142,31,142,30,24,31,47,31,205,31,43,31,43,30,169,31,232,31,158,31,84,31,218,31,153,31,37,31,38,31,247,31,242,31,163,31,163,30,167,31,79,31,200,31,185,31,236,31,172,31,9,31,9,30,9,29,139,31,74,31,190,31,8,31,155,31,105,31,125,31,114,31,114,30,235,31,125,31,164,31,96,31,169,31,169,30,128,31,148,31,146,31,146,30,146,29,223,31,223,30,76,31,76,30,53,31,3,31,215,31,216,31,183,31,121,31,49,31,150,31,62,31,225,31,16,31,27,31,27,30,33,31,33,30,1,31,86,31,46,31,46,30,64,31,91,31,151,31,151,30,82,31,30,31,117,31,186,31,101,31,87,31,87,30,161,31,170,31,140,31,17,31,146,31,62,31,130,31,22,31,117,31,128,31,59,31,59,30,150,31,95,31,185,31,182,31,182,30,125,31,177,31,173,31,85,31,60,31,133,31,167,31,167,30,138,31,140,31,160,31,152,31,208,31,136,31,53,31,28,31,196,31,196,30,93,31,46,31,71,31,71,30,62,31,126,31,223,31,224,31,23,31,203,31,145,31,63,31,251,31,243,31,9,31,188,31,146,31,63,31,197,31,209,31,102,31,102,30,205,31,205,30,91,31,143,31,64,31,199,31,212,31,183,31,48,31,68,31,219,31,45,31,45,30,41,31,41,30,174,31,137,31,3,31,3,30,92,31,92,30,3,31,213,31,185,31,152,31,253,31,253,30,243,31,32,31,58,31,184,31,69,31,77,31,77,30,77,29,74,31,11,31,156,31,156,30,181,31,97,31,120,31,120,30,185,31,193,31,77,31,29,31,28,31,163,31,83,31,228,31,87,31,87,30,41,31,72,31,77,31,77,30,107,31,169,31,169,30,138,31,34,31,1,31,24,31,60,31,57,31,55,31,108,31,27,31,73,31,188,31,234,31,54,31,32,31,32,30,32,29,3,31,3,30,122,31,84,31,217,31,226,31,91,31,80,31,193,31,219,31,69,31,77,31,102,31,222,31,189,31,194,31,236,31,227,31,117,31,219,31,219,30,250,31,82,31,182,31,228,31,188,31,109,31,109,30,247,31,231,31,47,31,75,31,182,31,92,31,244,31,31,31,139,31,206,31,249,31,249,30,233,31,28,31,28,30,46,31,8,31,166,31,166,30,73,31,12,31,221,31,90,31,90,30,252,31,80,31,110,31,190,31,166,31,166,30,123,31,123,30,105,31,28,31,28,30,63,31,31,31,201,31,176,31,235,31,252,31,132,31,217,31,87,31,87,30,3,31,198,31,198,30,198,29,187,31,231,31,231,30,250,31,187,31,206,31,31,31,31,30,31,29,31,28,31,27,31,26,85,31,107,31,200,31,200,30,43,31,77,31,61,31,124,31,63,31,63,30,63,29,231,31,231,30,145,31,145,30,27,31,181,31,194,31,121,31,121,30,108,31,87,31,169,31,141,31,187,31,32,31,128,31,15,31,249,31,242,31,242,30,123,31,122,31,31,31,31,30,128,31,113,31,178,31,200,31,160,31,5,31,185,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
