-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 273;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (178,0,0,0,59,0,220,0,0,0,0,0,216,0,104,0,167,0,250,0,0,0,20,0,105,0,133,0,0,0,190,0,18,0,152,0,155,0,90,0,24,0,249,0,164,0,90,0,171,0,224,0,156,0,142,0,0,0,227,0,95,0,187,0,244,0,195,0,0,0,125,0,254,0,81,0,92,0,14,0,222,0,4,0,9,0,97,0,15,0,76,0,54,0,190,0,42,0,175,0,187,0,121,0,184,0,76,0,130,0,146,0,207,0,194,0,147,0,59,0,190,0,188,0,255,0,0,0,232,0,57,0,201,0,125,0,197,0,78,0,168,0,188,0,0,0,209,0,36,0,84,0,124,0,0,0,0,0,145,0,150,0,226,0,175,0,41,0,139,0,133,0,141,0,82,0,0,0,0,0,16,0,159,0,154,0,0,0,188,0,0,0,67,0,136,0,0,0,229,0,225,0,38,0,0,0,85,0,188,0,144,0,120,0,32,0,162,0,94,0,150,0,169,0,65,0,235,0,234,0,183,0,0,0,0,0,158,0,94,0,0,0,41,0,0,0,0,0,100,0,175,0,143,0,226,0,55,0,115,0,190,0,19,0,254,0,55,0,201,0,53,0,129,0,96,0,196,0,77,0,177,0,66,0,129,0,69,0,111,0,0,0,132,0,0,0,216,0,202,0,204,0,174,0,124,0,251,0,101,0,130,0,68,0,163,0,0,0,189,0,0,0,94,0,0,0,193,0,217,0,155,0,32,0,12,0,117,0,0,0,21,0,148,0,38,0,165,0,90,0,250,0,91,0,60,0,79,0,132,0,76,0,49,0,184,0,38,0,215,0,143,0,33,0,70,0,72,0,81,0,216,0,219,0,0,0,93,0,0,0,0,0,222,0,231,0,170,0,0,0,19,0,162,0,57,0,179,0,167,0,133,0,0,0,145,0,170,0,252,0,55,0,14,0,37,0,112,0,29,0,121,0,32,0,158,0,186,0,210,0,118,0,139,0,217,0,83,0,0,0,19,0,0,0,84,0,67,0,0,0,0,0,10,0,50,0,97,0,144,0,168,0,56,0,91,0,23,0,151,0,79,0,108,0,250,0,68,0,207,0,0,0,50,0,42,0,78,0,232,0,82,0,169,0,53,0,103,0,195,0,125,0,156,0,160,0,67,0,152,0,5,0,133,0,0,0,226,0,11,0,85,0,0,0,0,0,157,0,86,0,232,0,0,0,0,0);
signal scenario_full  : scenario_type := (178,31,178,30,59,31,220,31,220,30,220,29,216,31,104,31,167,31,250,31,250,30,20,31,105,31,133,31,133,30,190,31,18,31,152,31,155,31,90,31,24,31,249,31,164,31,90,31,171,31,224,31,156,31,142,31,142,30,227,31,95,31,187,31,244,31,195,31,195,30,125,31,254,31,81,31,92,31,14,31,222,31,4,31,9,31,97,31,15,31,76,31,54,31,190,31,42,31,175,31,187,31,121,31,184,31,76,31,130,31,146,31,207,31,194,31,147,31,59,31,190,31,188,31,255,31,255,30,232,31,57,31,201,31,125,31,197,31,78,31,168,31,188,31,188,30,209,31,36,31,84,31,124,31,124,30,124,29,145,31,150,31,226,31,175,31,41,31,139,31,133,31,141,31,82,31,82,30,82,29,16,31,159,31,154,31,154,30,188,31,188,30,67,31,136,31,136,30,229,31,225,31,38,31,38,30,85,31,188,31,144,31,120,31,32,31,162,31,94,31,150,31,169,31,65,31,235,31,234,31,183,31,183,30,183,29,158,31,94,31,94,30,41,31,41,30,41,29,100,31,175,31,143,31,226,31,55,31,115,31,190,31,19,31,254,31,55,31,201,31,53,31,129,31,96,31,196,31,77,31,177,31,66,31,129,31,69,31,111,31,111,30,132,31,132,30,216,31,202,31,204,31,174,31,124,31,251,31,101,31,130,31,68,31,163,31,163,30,189,31,189,30,94,31,94,30,193,31,217,31,155,31,32,31,12,31,117,31,117,30,21,31,148,31,38,31,165,31,90,31,250,31,91,31,60,31,79,31,132,31,76,31,49,31,184,31,38,31,215,31,143,31,33,31,70,31,72,31,81,31,216,31,219,31,219,30,93,31,93,30,93,29,222,31,231,31,170,31,170,30,19,31,162,31,57,31,179,31,167,31,133,31,133,30,145,31,170,31,252,31,55,31,14,31,37,31,112,31,29,31,121,31,32,31,158,31,186,31,210,31,118,31,139,31,217,31,83,31,83,30,19,31,19,30,84,31,67,31,67,30,67,29,10,31,50,31,97,31,144,31,168,31,56,31,91,31,23,31,151,31,79,31,108,31,250,31,68,31,207,31,207,30,50,31,42,31,78,31,232,31,82,31,169,31,53,31,103,31,195,31,125,31,156,31,160,31,67,31,152,31,5,31,133,31,133,30,226,31,11,31,85,31,85,30,85,29,157,31,86,31,232,31,232,30,232,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
