-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 317;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,92,0,151,0,129,0,255,0,139,0,39,0,0,0,0,0,172,0,182,0,220,0,138,0,66,0,135,0,184,0,139,0,22,0,0,0,10,0,56,0,211,0,243,0,180,0,25,0,124,0,218,0,245,0,34,0,138,0,108,0,97,0,0,0,59,0,0,0,242,0,0,0,165,0,23,0,5,0,104,0,207,0,178,0,152,0,26,0,92,0,7,0,230,0,105,0,25,0,128,0,147,0,206,0,73,0,0,0,137,0,0,0,190,0,0,0,170,0,0,0,4,0,140,0,71,0,146,0,31,0,0,0,42,0,163,0,192,0,121,0,207,0,197,0,68,0,77,0,222,0,1,0,0,0,89,0,231,0,252,0,82,0,75,0,204,0,157,0,0,0,59,0,9,0,0,0,0,0,0,0,44,0,8,0,1,0,167,0,32,0,215,0,4,0,0,0,97,0,0,0,0,0,0,0,254,0,114,0,0,0,52,0,10,0,197,0,202,0,0,0,182,0,0,0,239,0,233,0,0,0,0,0,0,0,137,0,0,0,86,0,138,0,0,0,22,0,243,0,133,0,169,0,250,0,127,0,235,0,197,0,52,0,71,0,189,0,0,0,0,0,151,0,75,0,153,0,31,0,0,0,66,0,0,0,165,0,38,0,0,0,90,0,249,0,72,0,100,0,84,0,208,0,0,0,0,0,172,0,7,0,18,0,155,0,0,0,195,0,198,0,50,0,28,0,85,0,239,0,247,0,162,0,145,0,0,0,0,0,0,0,122,0,125,0,133,0,0,0,98,0,166,0,0,0,0,0,120,0,236,0,169,0,248,0,79,0,168,0,0,0,0,0,126,0,120,0,14,0,65,0,165,0,196,0,0,0,229,0,233,0,90,0,165,0,73,0,191,0,0,0,17,0,104,0,233,0,0,0,189,0,137,0,0,0,190,0,88,0,231,0,0,0,0,0,0,0,79,0,145,0,0,0,26,0,0,0,244,0,50,0,27,0,4,0,42,0,0,0,57,0,120,0,0,0,35,0,0,0,28,0,218,0,137,0,225,0,0,0,212,0,77,0,48,0,30,0,154,0,0,0,121,0,226,0,0,0,2,0,80,0,185,0,191,0,0,0,28,0,38,0,195,0,51,0,205,0,45,0,147,0,204,0,36,0,218,0,83,0,194,0,172,0,253,0,72,0,237,0,58,0,0,0,45,0,66,0,20,0,57,0,225,0,0,0,154,0,182,0,42,0,136,0,235,0,0,0,127,0,171,0,179,0,0,0,0,0,182,0,26,0,78,0,208,0,0,0,119,0,179,0,29,0,203,0,246,0,187,0,169,0,131,0,9,0,46,0,88,0,101,0,255,0,135,0,159,0,32,0,225,0,32,0,0,0,237,0,169,0,0,0,248,0,97,0,168,0,198,0,239,0,96,0);
signal scenario_full  : scenario_type := (40,31,92,31,151,31,129,31,255,31,139,31,39,31,39,30,39,29,172,31,182,31,220,31,138,31,66,31,135,31,184,31,139,31,22,31,22,30,10,31,56,31,211,31,243,31,180,31,25,31,124,31,218,31,245,31,34,31,138,31,108,31,97,31,97,30,59,31,59,30,242,31,242,30,165,31,23,31,5,31,104,31,207,31,178,31,152,31,26,31,92,31,7,31,230,31,105,31,25,31,128,31,147,31,206,31,73,31,73,30,137,31,137,30,190,31,190,30,170,31,170,30,4,31,140,31,71,31,146,31,31,31,31,30,42,31,163,31,192,31,121,31,207,31,197,31,68,31,77,31,222,31,1,31,1,30,89,31,231,31,252,31,82,31,75,31,204,31,157,31,157,30,59,31,9,31,9,30,9,29,9,28,44,31,8,31,1,31,167,31,32,31,215,31,4,31,4,30,97,31,97,30,97,29,97,28,254,31,114,31,114,30,52,31,10,31,197,31,202,31,202,30,182,31,182,30,239,31,233,31,233,30,233,29,233,28,137,31,137,30,86,31,138,31,138,30,22,31,243,31,133,31,169,31,250,31,127,31,235,31,197,31,52,31,71,31,189,31,189,30,189,29,151,31,75,31,153,31,31,31,31,30,66,31,66,30,165,31,38,31,38,30,90,31,249,31,72,31,100,31,84,31,208,31,208,30,208,29,172,31,7,31,18,31,155,31,155,30,195,31,198,31,50,31,28,31,85,31,239,31,247,31,162,31,145,31,145,30,145,29,145,28,122,31,125,31,133,31,133,30,98,31,166,31,166,30,166,29,120,31,236,31,169,31,248,31,79,31,168,31,168,30,168,29,126,31,120,31,14,31,65,31,165,31,196,31,196,30,229,31,233,31,90,31,165,31,73,31,191,31,191,30,17,31,104,31,233,31,233,30,189,31,137,31,137,30,190,31,88,31,231,31,231,30,231,29,231,28,79,31,145,31,145,30,26,31,26,30,244,31,50,31,27,31,4,31,42,31,42,30,57,31,120,31,120,30,35,31,35,30,28,31,218,31,137,31,225,31,225,30,212,31,77,31,48,31,30,31,154,31,154,30,121,31,226,31,226,30,2,31,80,31,185,31,191,31,191,30,28,31,38,31,195,31,51,31,205,31,45,31,147,31,204,31,36,31,218,31,83,31,194,31,172,31,253,31,72,31,237,31,58,31,58,30,45,31,66,31,20,31,57,31,225,31,225,30,154,31,182,31,42,31,136,31,235,31,235,30,127,31,171,31,179,31,179,30,179,29,182,31,26,31,78,31,208,31,208,30,119,31,179,31,29,31,203,31,246,31,187,31,169,31,131,31,9,31,46,31,88,31,101,31,255,31,135,31,159,31,32,31,225,31,32,31,32,30,237,31,169,31,169,30,248,31,97,31,168,31,198,31,239,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
