-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_717 is
end project_tb_717;

architecture project_tb_arch_717 of project_tb_717 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 950;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,204,0,0,0,115,0,230,0,191,0,186,0,121,0,89,0,28,0,6,0,24,0,0,0,109,0,74,0,95,0,161,0,198,0,0,0,158,0,79,0,90,0,0,0,0,0,207,0,210,0,0,0,20,0,242,0,28,0,254,0,0,0,179,0,103,0,84,0,133,0,113,0,16,0,77,0,155,0,206,0,0,0,5,0,60,0,0,0,241,0,122,0,0,0,0,0,21,0,168,0,235,0,0,0,209,0,65,0,0,0,188,0,4,0,24,0,209,0,75,0,0,0,16,0,24,0,189,0,0,0,122,0,167,0,0,0,47,0,16,0,0,0,0,0,126,0,31,0,20,0,30,0,93,0,48,0,254,0,252,0,0,0,0,0,0,0,170,0,0,0,0,0,219,0,248,0,65,0,79,0,133,0,165,0,61,0,249,0,5,0,116,0,201,0,188,0,179,0,0,0,90,0,238,0,0,0,248,0,140,0,254,0,24,0,130,0,54,0,111,0,196,0,160,0,69,0,72,0,74,0,158,0,83,0,58,0,106,0,0,0,184,0,52,0,128,0,214,0,251,0,4,0,14,0,184,0,104,0,231,0,0,0,0,0,46,0,0,0,150,0,197,0,165,0,0,0,34,0,219,0,59,0,34,0,106,0,73,0,0,0,191,0,16,0,189,0,0,0,32,0,178,0,232,0,10,0,39,0,152,0,40,0,95,0,150,0,0,0,0,0,173,0,109,0,198,0,195,0,151,0,142,0,224,0,142,0,111,0,130,0,207,0,13,0,48,0,0,0,137,0,123,0,131,0,143,0,91,0,176,0,169,0,84,0,209,0,129,0,123,0,0,0,189,0,0,0,0,0,134,0,197,0,93,0,0,0,171,0,89,0,130,0,167,0,141,0,101,0,153,0,124,0,244,0,119,0,0,0,117,0,0,0,0,0,46,0,243,0,153,0,135,0,77,0,0,0,0,0,0,0,98,0,116,0,114,0,0,0,19,0,119,0,0,0,0,0,145,0,0,0,182,0,91,0,4,0,0,0,0,0,247,0,223,0,85,0,65,0,54,0,0,0,206,0,57,0,106,0,241,0,0,0,217,0,144,0,2,0,0,0,229,0,156,0,12,0,0,0,106,0,34,0,157,0,23,0,0,0,144,0,18,0,0,0,188,0,79,0,0,0,254,0,146,0,0,0,244,0,121,0,52,0,175,0,198,0,164,0,0,0,244,0,152,0,49,0,109,0,149,0,130,0,154,0,0,0,226,0,184,0,0,0,188,0,0,0,0,0,0,0,0,0,0,0,207,0,147,0,135,0,0,0,0,0,23,0,103,0,148,0,174,0,0,0,0,0,98,0,30,0,11,0,188,0,135,0,0,0,27,0,209,0,58,0,214,0,0,0,114,0,57,0,5,0,117,0,110,0,0,0,71,0,225,0,145,0,239,0,225,0,101,0,240,0,232,0,192,0,128,0,199,0,121,0,0,0,124,0,171,0,12,0,6,0,94,0,126,0,0,0,172,0,138,0,35,0,246,0,45,0,88,0,0,0,113,0,10,0,210,0,123,0,90,0,44,0,123,0,221,0,222,0,200,0,142,0,122,0,16,0,129,0,15,0,93,0,93,0,0,0,108,0,171,0,200,0,0,0,0,0,66,0,164,0,53,0,164,0,25,0,51,0,0,0,135,0,97,0,114,0,0,0,86,0,210,0,228,0,216,0,37,0,171,0,121,0,198,0,19,0,240,0,241,0,111,0,0,0,169,0,191,0,43,0,218,0,207,0,0,0,250,0,0,0,108,0,192,0,172,0,0,0,36,0,149,0,95,0,230,0,0,0,216,0,91,0,0,0,70,0,64,0,2,0,144,0,198,0,37,0,0,0,127,0,96,0,105,0,206,0,218,0,0,0,92,0,0,0,199,0,188,0,205,0,44,0,55,0,0,0,150,0,9,0,130,0,0,0,168,0,24,0,99,0,0,0,251,0,0,0,106,0,126,0,168,0,34,0,130,0,100,0,227,0,214,0,188,0,219,0,0,0,227,0,95,0,18,0,237,0,131,0,153,0,79,0,225,0,89,0,23,0,109,0,224,0,123,0,101,0,0,0,179,0,248,0,0,0,0,0,184,0,137,0,88,0,105,0,37,0,59,0,0,0,35,0,205,0,0,0,0,0,253,0,0,0,141,0,159,0,177,0,185,0,254,0,0,0,234,0,0,0,55,0,0,0,0,0,0,0,251,0,0,0,216,0,149,0,0,0,220,0,251,0,0,0,235,0,16,0,151,0,228,0,0,0,110,0,207,0,27,0,54,0,14,0,49,0,0,0,0,0,128,0,0,0,135,0,253,0,3,0,109,0,108,0,43,0,197,0,225,0,0,0,0,0,239,0,202,0,209,0,9,0,227,0,99,0,152,0,45,0,28,0,64,0,253,0,0,0,134,0,141,0,104,0,184,0,108,0,134,0,142,0,85,0,0,0,53,0,189,0,0,0,155,0,0,0,0,0,105,0,243,0,207,0,242,0,237,0,27,0,160,0,190,0,150,0,72,0,0,0,217,0,125,0,0,0,27,0,251,0,150,0,67,0,148,0,0,0,83,0,45,0,0,0,8,0,0,0,0,0,173,0,109,0,190,0,0,0,15,0,213,0,159,0,234,0,64,0,138,0,199,0,0,0,0,0,186,0,0,0,176,0,198,0,37,0,0,0,248,0,0,0,135,0,136,0,0,0,221,0,91,0,23,0,68,0,13,0,184,0,200,0,184,0,45,0,94,0,111,0,186,0,188,0,150,0,107,0,21,0,149,0,119,0,191,0,133,0,221,0,53,0,48,0,214,0,58,0,0,0,160,0,0,0,0,0,253,0,247,0,159,0,129,0,0,0,47,0,0,0,157,0,200,0,155,0,0,0,82,0,239,0,173,0,135,0,0,0,114,0,33,0,32,0,235,0,108,0,78,0,98,0,200,0,96,0,225,0,179,0,84,0,0,0,147,0,15,0,233,0,177,0,0,0,133,0,103,0,155,0,15,0,246,0,0,0,148,0,148,0,134,0,189,0,187,0,76,0,217,0,131,0,0,0,0,0,119,0,152,0,138,0,105,0,0,0,0,0,202,0,191,0,0,0,108,0,190,0,192,0,122,0,244,0,0,0,32,0,0,0,17,0,0,0,186,0,208,0,207,0,112,0,179,0,178,0,108,0,98,0,0,0,0,0,72,0,46,0,116,0,68,0,117,0,74,0,10,0,56,0,66,0,0,0,55,0,65,0,19,0,250,0,132,0,34,0,0,0,0,0,64,0,55,0,113,0,103,0,230,0,255,0,133,0,207,0,99,0,243,0,0,0,59,0,107,0,0,0,0,0,0,0,105,0,218,0,68,0,0,0,123,0,198,0,18,0,2,0,0,0,232,0,202,0,12,0,240,0,173,0,159,0,75,0,205,0,0,0,0,0,0,0,217,0,211,0,199,0,58,0,121,0,3,0,42,0,199,0,0,0,0,0,0,0,13,0,35,0,138,0,7,0,113,0,225,0,0,0,226,0,170,0,186,0,144,0,0,0,46,0,168,0,164,0,78,0,123,0,0,0,140,0,240,0,184,0,0,0,0,0,31,0,0,0,156,0,214,0,159,0,51,0,162,0,97,0,63,0,0,0,149,0,0,0,204,0,6,0,246,0,191,0,254,0,142,0,212,0,0,0,207,0,0,0,25,0,187,0,186,0,207,0,16,0,201,0,0,0,90,0,9,0,167,0,174,0,64,0,188,0,5,0,0,0,0,0,170,0,0,0,0,0,245,0,57,0,168,0,95,0,0,0,141,0,154,0,0,0,62,0,229,0,199,0,96,0,190,0,142,0,57,0,33,0,15,0,0,0,0,0,252,0,89,0,221,0,91,0,87,0,9,0,250,0,229,0,0,0,176,0,50,0,237,0,47,0,178,0,23,0,41,0,198,0,90,0,155,0,0,0,43,0,142,0,0,0,40,0,56,0,41,0,0,0,248,0,97,0,29,0,25,0,231,0,187,0,156,0,69,0,254,0,0,0,108,0,253,0,0,0,0,0,2,0,87,0,0,0,193,0,219,0,1,0,128,0,98,0,240,0,0,0,28,0,39,0,0,0,54,0,25,0,0,0,194,0,106,0,188,0,40,0,79,0,191,0,117,0,2,0,235,0,80,0,230,0,16,0,1,0,0,0,255,0,0,0,161,0,72,0,0,0,104,0,122,0,230,0,175,0,125,0,5,0,239,0,18,0,231,0,237,0,175,0,0,0);
signal scenario_full  : scenario_type := (0,0,204,31,204,30,115,31,230,31,191,31,186,31,121,31,89,31,28,31,6,31,24,31,24,30,109,31,74,31,95,31,161,31,198,31,198,30,158,31,79,31,90,31,90,30,90,29,207,31,210,31,210,30,20,31,242,31,28,31,254,31,254,30,179,31,103,31,84,31,133,31,113,31,16,31,77,31,155,31,206,31,206,30,5,31,60,31,60,30,241,31,122,31,122,30,122,29,21,31,168,31,235,31,235,30,209,31,65,31,65,30,188,31,4,31,24,31,209,31,75,31,75,30,16,31,24,31,189,31,189,30,122,31,167,31,167,30,47,31,16,31,16,30,16,29,126,31,31,31,20,31,30,31,93,31,48,31,254,31,252,31,252,30,252,29,252,28,170,31,170,30,170,29,219,31,248,31,65,31,79,31,133,31,165,31,61,31,249,31,5,31,116,31,201,31,188,31,179,31,179,30,90,31,238,31,238,30,248,31,140,31,254,31,24,31,130,31,54,31,111,31,196,31,160,31,69,31,72,31,74,31,158,31,83,31,58,31,106,31,106,30,184,31,52,31,128,31,214,31,251,31,4,31,14,31,184,31,104,31,231,31,231,30,231,29,46,31,46,30,150,31,197,31,165,31,165,30,34,31,219,31,59,31,34,31,106,31,73,31,73,30,191,31,16,31,189,31,189,30,32,31,178,31,232,31,10,31,39,31,152,31,40,31,95,31,150,31,150,30,150,29,173,31,109,31,198,31,195,31,151,31,142,31,224,31,142,31,111,31,130,31,207,31,13,31,48,31,48,30,137,31,123,31,131,31,143,31,91,31,176,31,169,31,84,31,209,31,129,31,123,31,123,30,189,31,189,30,189,29,134,31,197,31,93,31,93,30,171,31,89,31,130,31,167,31,141,31,101,31,153,31,124,31,244,31,119,31,119,30,117,31,117,30,117,29,46,31,243,31,153,31,135,31,77,31,77,30,77,29,77,28,98,31,116,31,114,31,114,30,19,31,119,31,119,30,119,29,145,31,145,30,182,31,91,31,4,31,4,30,4,29,247,31,223,31,85,31,65,31,54,31,54,30,206,31,57,31,106,31,241,31,241,30,217,31,144,31,2,31,2,30,229,31,156,31,12,31,12,30,106,31,34,31,157,31,23,31,23,30,144,31,18,31,18,30,188,31,79,31,79,30,254,31,146,31,146,30,244,31,121,31,52,31,175,31,198,31,164,31,164,30,244,31,152,31,49,31,109,31,149,31,130,31,154,31,154,30,226,31,184,31,184,30,188,31,188,30,188,29,188,28,188,27,188,26,207,31,147,31,135,31,135,30,135,29,23,31,103,31,148,31,174,31,174,30,174,29,98,31,30,31,11,31,188,31,135,31,135,30,27,31,209,31,58,31,214,31,214,30,114,31,57,31,5,31,117,31,110,31,110,30,71,31,225,31,145,31,239,31,225,31,101,31,240,31,232,31,192,31,128,31,199,31,121,31,121,30,124,31,171,31,12,31,6,31,94,31,126,31,126,30,172,31,138,31,35,31,246,31,45,31,88,31,88,30,113,31,10,31,210,31,123,31,90,31,44,31,123,31,221,31,222,31,200,31,142,31,122,31,16,31,129,31,15,31,93,31,93,31,93,30,108,31,171,31,200,31,200,30,200,29,66,31,164,31,53,31,164,31,25,31,51,31,51,30,135,31,97,31,114,31,114,30,86,31,210,31,228,31,216,31,37,31,171,31,121,31,198,31,19,31,240,31,241,31,111,31,111,30,169,31,191,31,43,31,218,31,207,31,207,30,250,31,250,30,108,31,192,31,172,31,172,30,36,31,149,31,95,31,230,31,230,30,216,31,91,31,91,30,70,31,64,31,2,31,144,31,198,31,37,31,37,30,127,31,96,31,105,31,206,31,218,31,218,30,92,31,92,30,199,31,188,31,205,31,44,31,55,31,55,30,150,31,9,31,130,31,130,30,168,31,24,31,99,31,99,30,251,31,251,30,106,31,126,31,168,31,34,31,130,31,100,31,227,31,214,31,188,31,219,31,219,30,227,31,95,31,18,31,237,31,131,31,153,31,79,31,225,31,89,31,23,31,109,31,224,31,123,31,101,31,101,30,179,31,248,31,248,30,248,29,184,31,137,31,88,31,105,31,37,31,59,31,59,30,35,31,205,31,205,30,205,29,253,31,253,30,141,31,159,31,177,31,185,31,254,31,254,30,234,31,234,30,55,31,55,30,55,29,55,28,251,31,251,30,216,31,149,31,149,30,220,31,251,31,251,30,235,31,16,31,151,31,228,31,228,30,110,31,207,31,27,31,54,31,14,31,49,31,49,30,49,29,128,31,128,30,135,31,253,31,3,31,109,31,108,31,43,31,197,31,225,31,225,30,225,29,239,31,202,31,209,31,9,31,227,31,99,31,152,31,45,31,28,31,64,31,253,31,253,30,134,31,141,31,104,31,184,31,108,31,134,31,142,31,85,31,85,30,53,31,189,31,189,30,155,31,155,30,155,29,105,31,243,31,207,31,242,31,237,31,27,31,160,31,190,31,150,31,72,31,72,30,217,31,125,31,125,30,27,31,251,31,150,31,67,31,148,31,148,30,83,31,45,31,45,30,8,31,8,30,8,29,173,31,109,31,190,31,190,30,15,31,213,31,159,31,234,31,64,31,138,31,199,31,199,30,199,29,186,31,186,30,176,31,198,31,37,31,37,30,248,31,248,30,135,31,136,31,136,30,221,31,91,31,23,31,68,31,13,31,184,31,200,31,184,31,45,31,94,31,111,31,186,31,188,31,150,31,107,31,21,31,149,31,119,31,191,31,133,31,221,31,53,31,48,31,214,31,58,31,58,30,160,31,160,30,160,29,253,31,247,31,159,31,129,31,129,30,47,31,47,30,157,31,200,31,155,31,155,30,82,31,239,31,173,31,135,31,135,30,114,31,33,31,32,31,235,31,108,31,78,31,98,31,200,31,96,31,225,31,179,31,84,31,84,30,147,31,15,31,233,31,177,31,177,30,133,31,103,31,155,31,15,31,246,31,246,30,148,31,148,31,134,31,189,31,187,31,76,31,217,31,131,31,131,30,131,29,119,31,152,31,138,31,105,31,105,30,105,29,202,31,191,31,191,30,108,31,190,31,192,31,122,31,244,31,244,30,32,31,32,30,17,31,17,30,186,31,208,31,207,31,112,31,179,31,178,31,108,31,98,31,98,30,98,29,72,31,46,31,116,31,68,31,117,31,74,31,10,31,56,31,66,31,66,30,55,31,65,31,19,31,250,31,132,31,34,31,34,30,34,29,64,31,55,31,113,31,103,31,230,31,255,31,133,31,207,31,99,31,243,31,243,30,59,31,107,31,107,30,107,29,107,28,105,31,218,31,68,31,68,30,123,31,198,31,18,31,2,31,2,30,232,31,202,31,12,31,240,31,173,31,159,31,75,31,205,31,205,30,205,29,205,28,217,31,211,31,199,31,58,31,121,31,3,31,42,31,199,31,199,30,199,29,199,28,13,31,35,31,138,31,7,31,113,31,225,31,225,30,226,31,170,31,186,31,144,31,144,30,46,31,168,31,164,31,78,31,123,31,123,30,140,31,240,31,184,31,184,30,184,29,31,31,31,30,156,31,214,31,159,31,51,31,162,31,97,31,63,31,63,30,149,31,149,30,204,31,6,31,246,31,191,31,254,31,142,31,212,31,212,30,207,31,207,30,25,31,187,31,186,31,207,31,16,31,201,31,201,30,90,31,9,31,167,31,174,31,64,31,188,31,5,31,5,30,5,29,170,31,170,30,170,29,245,31,57,31,168,31,95,31,95,30,141,31,154,31,154,30,62,31,229,31,199,31,96,31,190,31,142,31,57,31,33,31,15,31,15,30,15,29,252,31,89,31,221,31,91,31,87,31,9,31,250,31,229,31,229,30,176,31,50,31,237,31,47,31,178,31,23,31,41,31,198,31,90,31,155,31,155,30,43,31,142,31,142,30,40,31,56,31,41,31,41,30,248,31,97,31,29,31,25,31,231,31,187,31,156,31,69,31,254,31,254,30,108,31,253,31,253,30,253,29,2,31,87,31,87,30,193,31,219,31,1,31,128,31,98,31,240,31,240,30,28,31,39,31,39,30,54,31,25,31,25,30,194,31,106,31,188,31,40,31,79,31,191,31,117,31,2,31,235,31,80,31,230,31,16,31,1,31,1,30,255,31,255,30,161,31,72,31,72,30,104,31,122,31,230,31,175,31,125,31,5,31,239,31,18,31,231,31,237,31,175,31,175,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
