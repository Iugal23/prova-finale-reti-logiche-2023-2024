-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_385 is
end project_tb_385;

architecture project_tb_arch_385 of project_tb_385 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 233;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,242,0,169,0,153,0,0,0,124,0,203,0,175,0,176,0,161,0,200,0,0,0,42,0,11,0,229,0,88,0,151,0,9,0,0,0,87,0,10,0,0,0,131,0,177,0,0,0,142,0,14,0,255,0,0,0,0,0,177,0,180,0,0,0,79,0,0,0,152,0,109,0,127,0,69,0,0,0,0,0,156,0,185,0,0,0,113,0,247,0,0,0,146,0,0,0,163,0,0,0,95,0,71,0,251,0,0,0,152,0,203,0,0,0,227,0,182,0,221,0,0,0,0,0,252,0,51,0,39,0,0,0,94,0,169,0,197,0,116,0,46,0,140,0,0,0,40,0,147,0,103,0,87,0,125,0,121,0,68,0,145,0,0,0,102,0,177,0,0,0,24,0,0,0,235,0,61,0,90,0,0,0,0,0,185,0,144,0,251,0,138,0,255,0,23,0,224,0,112,0,47,0,140,0,144,0,84,0,60,0,178,0,51,0,18,0,0,0,206,0,0,0,0,0,143,0,75,0,22,0,105,0,7,0,130,0,206,0,142,0,63,0,254,0,0,0,94,0,164,0,108,0,93,0,0,0,0,0,169,0,164,0,45,0,229,0,3,0,123,0,216,0,73,0,5,0,54,0,149,0,0,0,29,0,92,0,194,0,236,0,9,0,105,0,137,0,14,0,59,0,32,0,197,0,41,0,0,0,119,0,36,0,49,0,96,0,0,0,209,0,31,0,28,0,169,0,249,0,0,0,12,0,182,0,169,0,0,0,99,0,0,0,210,0,234,0,94,0,77,0,93,0,0,0,51,0,0,0,172,0,234,0,120,0,0,0,16,0,108,0,253,0,39,0,182,0,68,0,182,0,178,0,0,0,127,0,211,0,69,0,0,0,42,0,107,0,0,0,87,0,99,0,0,0,239,0,141,0,138,0,167,0,158,0,84,0,0,0,125,0,0,0,25,0,172,0,150,0,27,0,176,0,128,0,42,0,50,0,105,0,208,0,0,0,0,0,51,0,122,0,0,0,60,0,33,0,65,0,188,0,243,0,125,0);
signal scenario_full  : scenario_type := (49,31,242,31,169,31,153,31,153,30,124,31,203,31,175,31,176,31,161,31,200,31,200,30,42,31,11,31,229,31,88,31,151,31,9,31,9,30,87,31,10,31,10,30,131,31,177,31,177,30,142,31,14,31,255,31,255,30,255,29,177,31,180,31,180,30,79,31,79,30,152,31,109,31,127,31,69,31,69,30,69,29,156,31,185,31,185,30,113,31,247,31,247,30,146,31,146,30,163,31,163,30,95,31,71,31,251,31,251,30,152,31,203,31,203,30,227,31,182,31,221,31,221,30,221,29,252,31,51,31,39,31,39,30,94,31,169,31,197,31,116,31,46,31,140,31,140,30,40,31,147,31,103,31,87,31,125,31,121,31,68,31,145,31,145,30,102,31,177,31,177,30,24,31,24,30,235,31,61,31,90,31,90,30,90,29,185,31,144,31,251,31,138,31,255,31,23,31,224,31,112,31,47,31,140,31,144,31,84,31,60,31,178,31,51,31,18,31,18,30,206,31,206,30,206,29,143,31,75,31,22,31,105,31,7,31,130,31,206,31,142,31,63,31,254,31,254,30,94,31,164,31,108,31,93,31,93,30,93,29,169,31,164,31,45,31,229,31,3,31,123,31,216,31,73,31,5,31,54,31,149,31,149,30,29,31,92,31,194,31,236,31,9,31,105,31,137,31,14,31,59,31,32,31,197,31,41,31,41,30,119,31,36,31,49,31,96,31,96,30,209,31,31,31,28,31,169,31,249,31,249,30,12,31,182,31,169,31,169,30,99,31,99,30,210,31,234,31,94,31,77,31,93,31,93,30,51,31,51,30,172,31,234,31,120,31,120,30,16,31,108,31,253,31,39,31,182,31,68,31,182,31,178,31,178,30,127,31,211,31,69,31,69,30,42,31,107,31,107,30,87,31,99,31,99,30,239,31,141,31,138,31,167,31,158,31,84,31,84,30,125,31,125,30,25,31,172,31,150,31,27,31,176,31,128,31,42,31,50,31,105,31,208,31,208,30,208,29,51,31,122,31,122,30,60,31,33,31,65,31,188,31,243,31,125,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
