-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 199;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,4,0,23,0,16,0,89,0,0,0,12,0,171,0,214,0,113,0,0,0,151,0,0,0,0,0,49,0,85,0,189,0,41,0,5,0,166,0,224,0,152,0,206,0,247,0,228,0,0,0,191,0,67,0,0,0,2,0,115,0,16,0,85,0,179,0,187,0,181,0,145,0,168,0,68,0,12,0,87,0,0,0,242,0,0,0,0,0,7,0,20,0,0,0,25,0,136,0,114,0,238,0,73,0,0,0,0,0,232,0,54,0,23,0,150,0,76,0,9,0,15,0,103,0,219,0,152,0,0,0,253,0,165,0,0,0,84,0,61,0,0,0,0,0,48,0,0,0,75,0,192,0,196,0,110,0,194,0,58,0,244,0,0,0,38,0,213,0,0,0,163,0,189,0,32,0,110,0,0,0,20,0,10,0,150,0,0,0,99,0,61,0,160,0,199,0,254,0,178,0,126,0,243,0,120,0,26,0,0,0,87,0,29,0,163,0,4,0,43,0,37,0,108,0,227,0,153,0,27,0,75,0,0,0,150,0,201,0,75,0,0,0,14,0,36,0,106,0,0,0,0,0,87,0,0,0,176,0,252,0,236,0,120,0,113,0,228,0,231,0,0,0,131,0,154,0,227,0,106,0,0,0,206,0,49,0,168,0,101,0,15,0,52,0,115,0,239,0,0,0,115,0,0,0,185,0,0,0,200,0,66,0,0,0,0,0,52,0,235,0,0,0,201,0,139,0,2,0,85,0,125,0,0,0,105,0,246,0,211,0,41,0,0,0,194,0,83,0,5,0,224,0,119,0,113,0,154,0,145,0,64,0,108,0,251,0,191,0,194,0,106,0,158,0,67,0,58,0,0,0,57,0,103,0,211,0,147,0,248,0,0,0,250,0,164,0);
signal scenario_full  : scenario_type := (0,0,4,31,23,31,16,31,89,31,89,30,12,31,171,31,214,31,113,31,113,30,151,31,151,30,151,29,49,31,85,31,189,31,41,31,5,31,166,31,224,31,152,31,206,31,247,31,228,31,228,30,191,31,67,31,67,30,2,31,115,31,16,31,85,31,179,31,187,31,181,31,145,31,168,31,68,31,12,31,87,31,87,30,242,31,242,30,242,29,7,31,20,31,20,30,25,31,136,31,114,31,238,31,73,31,73,30,73,29,232,31,54,31,23,31,150,31,76,31,9,31,15,31,103,31,219,31,152,31,152,30,253,31,165,31,165,30,84,31,61,31,61,30,61,29,48,31,48,30,75,31,192,31,196,31,110,31,194,31,58,31,244,31,244,30,38,31,213,31,213,30,163,31,189,31,32,31,110,31,110,30,20,31,10,31,150,31,150,30,99,31,61,31,160,31,199,31,254,31,178,31,126,31,243,31,120,31,26,31,26,30,87,31,29,31,163,31,4,31,43,31,37,31,108,31,227,31,153,31,27,31,75,31,75,30,150,31,201,31,75,31,75,30,14,31,36,31,106,31,106,30,106,29,87,31,87,30,176,31,252,31,236,31,120,31,113,31,228,31,231,31,231,30,131,31,154,31,227,31,106,31,106,30,206,31,49,31,168,31,101,31,15,31,52,31,115,31,239,31,239,30,115,31,115,30,185,31,185,30,200,31,66,31,66,30,66,29,52,31,235,31,235,30,201,31,139,31,2,31,85,31,125,31,125,30,105,31,246,31,211,31,41,31,41,30,194,31,83,31,5,31,224,31,119,31,113,31,154,31,145,31,64,31,108,31,251,31,191,31,194,31,106,31,158,31,67,31,58,31,58,30,57,31,103,31,211,31,147,31,248,31,248,30,250,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
