-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_338 is
end project_tb_338;

architecture project_tb_arch_338 of project_tb_338 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 658;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,234,0,118,0,0,0,0,0,167,0,114,0,108,0,33,0,182,0,0,0,104,0,168,0,0,0,178,0,37,0,33,0,163,0,0,0,0,0,177,0,209,0,120,0,121,0,31,0,88,0,200,0,0,0,13,0,235,0,0,0,81,0,0,0,63,0,222,0,43,0,20,0,139,0,119,0,150,0,0,0,0,0,97,0,0,0,0,0,164,0,56,0,0,0,29,0,0,0,180,0,106,0,81,0,146,0,0,0,138,0,0,0,207,0,3,0,67,0,8,0,233,0,175,0,144,0,204,0,28,0,0,0,51,0,0,0,163,0,24,0,0,0,0,0,30,0,55,0,149,0,98,0,14,0,0,0,18,0,21,0,47,0,160,0,89,0,18,0,160,0,0,0,175,0,228,0,243,0,184,0,238,0,241,0,0,0,82,0,36,0,11,0,136,0,0,0,193,0,132,0,0,0,98,0,207,0,63,0,253,0,99,0,89,0,5,0,214,0,208,0,36,0,51,0,229,0,0,0,0,0,0,0,65,0,69,0,55,0,87,0,101,0,0,0,0,0,139,0,6,0,0,0,0,0,0,0,201,0,32,0,0,0,121,0,247,0,0,0,44,0,4,0,191,0,212,0,186,0,116,0,99,0,189,0,5,0,0,0,33,0,84,0,120,0,0,0,191,0,204,0,145,0,128,0,133,0,203,0,228,0,61,0,92,0,82,0,2,0,164,0,0,0,159,0,84,0,180,0,170,0,150,0,61,0,124,0,249,0,48,0,49,0,0,0,75,0,171,0,0,0,43,0,0,0,172,0,214,0,160,0,11,0,144,0,76,0,0,0,192,0,235,0,6,0,69,0,63,0,231,0,232,0,35,0,248,0,0,0,0,0,167,0,40,0,112,0,220,0,82,0,70,0,112,0,39,0,80,0,143,0,92,0,239,0,212,0,112,0,42,0,212,0,91,0,236,0,95,0,251,0,14,0,0,0,64,0,142,0,0,0,151,0,68,0,83,0,129,0,0,0,201,0,39,0,136,0,0,0,3,0,18,0,210,0,174,0,176,0,53,0,104,0,159,0,47,0,136,0,135,0,46,0,186,0,101,0,25,0,44,0,139,0,0,0,123,0,77,0,201,0,206,0,45,0,0,0,27,0,0,0,248,0,118,0,7,0,103,0,14,0,0,0,67,0,57,0,21,0,149,0,107,0,123,0,7,0,0,0,0,0,8,0,136,0,52,0,38,0,80,0,153,0,7,0,22,0,0,0,68,0,0,0,120,0,85,0,225,0,74,0,144,0,92,0,238,0,36,0,224,0,49,0,239,0,88,0,49,0,184,0,90,0,243,0,222,0,112,0,94,0,223,0,91,0,55,0,183,0,164,0,189,0,182,0,0,0,31,0,180,0,158,0,137,0,170,0,127,0,20,0,59,0,0,0,0,0,178,0,0,0,0,0,0,0,201,0,196,0,0,0,122,0,166,0,133,0,211,0,0,0,236,0,119,0,97,0,0,0,197,0,152,0,251,0,0,0,205,0,0,0,0,0,0,0,84,0,223,0,179,0,132,0,138,0,115,0,128,0,196,0,0,0,0,0,171,0,0,0,193,0,0,0,47,0,240,0,58,0,0,0,185,0,0,0,62,0,165,0,157,0,85,0,21,0,115,0,28,0,65,0,0,0,125,0,0,0,113,0,53,0,143,0,119,0,116,0,163,0,0,0,171,0,0,0,250,0,86,0,189,0,240,0,24,0,141,0,0,0,223,0,159,0,136,0,0,0,90,0,238,0,0,0,240,0,0,0,18,0,230,0,0,0,177,0,85,0,56,0,226,0,76,0,43,0,167,0,192,0,0,0,15,0,0,0,0,0,230,0,2,0,125,0,0,0,230,0,0,0,176,0,16,0,80,0,42,0,0,0,129,0,113,0,46,0,93,0,49,0,217,0,0,0,93,0,235,0,83,0,241,0,0,0,0,0,154,0,203,0,7,0,248,0,157,0,125,0,8,0,23,0,154,0,30,0,0,0,93,0,182,0,6,0,236,0,0,0,118,0,83,0,166,0,37,0,0,0,151,0,170,0,12,0,241,0,130,0,39,0,155,0,93,0,0,0,246,0,197,0,194,0,116,0,43,0,113,0,250,0,76,0,53,0,67,0,209,0,229,0,238,0,221,0,129,0,226,0,79,0,0,0,183,0,0,0,252,0,193,0,41,0,195,0,220,0,214,0,207,0,112,0,166,0,190,0,246,0,50,0,253,0,51,0,47,0,5,0,30,0,49,0,89,0,197,0,228,0,181,0,0,0,226,0,0,0,156,0,186,0,0,0,138,0,15,0,205,0,96,0,39,0,33,0,160,0,17,0,0,0,71,0,251,0,0,0,58,0,211,0,231,0,249,0,194,0,252,0,159,0,65,0,0,0,247,0,176,0,152,0,142,0,0,0,126,0,50,0,142,0,109,0,199,0,0,0,0,0,189,0,0,0,91,0,186,0,239,0,109,0,0,0,0,0,79,0,0,0,117,0,76,0,88,0,0,0,9,0,0,0,228,0,177,0,235,0,116,0,224,0,67,0,114,0,199,0,84,0,18,0,56,0,32,0,0,0,0,0,210,0,218,0,102,0,0,0,0,0,106,0,102,0,0,0,0,0,201,0,0,0,210,0,115,0,47,0,48,0,245,0,236,0,0,0,0,0,0,0,82,0,228,0,180,0,129,0,0,0,243,0,159,0,0,0,94,0,206,0,0,0,0,0,207,0,56,0,0,0,78,0,191,0,225,0,170,0,213,0,98,0,61,0,114,0,93,0,237,0,248,0,0,0,95,0,21,0,148,0,126,0,8,0,203,0,241,0,174,0,147,0,201,0,87,0,77,0,164,0,4,0,0,0,146,0,120,0,66,0,47,0,0,0,25,0,49,0,137,0,168,0,0,0,22,0,0,0,0,0,80,0,1,0,188,0,25,0);
signal scenario_full  : scenario_type := (0,0,234,31,118,31,118,30,118,29,167,31,114,31,108,31,33,31,182,31,182,30,104,31,168,31,168,30,178,31,37,31,33,31,163,31,163,30,163,29,177,31,209,31,120,31,121,31,31,31,88,31,200,31,200,30,13,31,235,31,235,30,81,31,81,30,63,31,222,31,43,31,20,31,139,31,119,31,150,31,150,30,150,29,97,31,97,30,97,29,164,31,56,31,56,30,29,31,29,30,180,31,106,31,81,31,146,31,146,30,138,31,138,30,207,31,3,31,67,31,8,31,233,31,175,31,144,31,204,31,28,31,28,30,51,31,51,30,163,31,24,31,24,30,24,29,30,31,55,31,149,31,98,31,14,31,14,30,18,31,21,31,47,31,160,31,89,31,18,31,160,31,160,30,175,31,228,31,243,31,184,31,238,31,241,31,241,30,82,31,36,31,11,31,136,31,136,30,193,31,132,31,132,30,98,31,207,31,63,31,253,31,99,31,89,31,5,31,214,31,208,31,36,31,51,31,229,31,229,30,229,29,229,28,65,31,69,31,55,31,87,31,101,31,101,30,101,29,139,31,6,31,6,30,6,29,6,28,201,31,32,31,32,30,121,31,247,31,247,30,44,31,4,31,191,31,212,31,186,31,116,31,99,31,189,31,5,31,5,30,33,31,84,31,120,31,120,30,191,31,204,31,145,31,128,31,133,31,203,31,228,31,61,31,92,31,82,31,2,31,164,31,164,30,159,31,84,31,180,31,170,31,150,31,61,31,124,31,249,31,48,31,49,31,49,30,75,31,171,31,171,30,43,31,43,30,172,31,214,31,160,31,11,31,144,31,76,31,76,30,192,31,235,31,6,31,69,31,63,31,231,31,232,31,35,31,248,31,248,30,248,29,167,31,40,31,112,31,220,31,82,31,70,31,112,31,39,31,80,31,143,31,92,31,239,31,212,31,112,31,42,31,212,31,91,31,236,31,95,31,251,31,14,31,14,30,64,31,142,31,142,30,151,31,68,31,83,31,129,31,129,30,201,31,39,31,136,31,136,30,3,31,18,31,210,31,174,31,176,31,53,31,104,31,159,31,47,31,136,31,135,31,46,31,186,31,101,31,25,31,44,31,139,31,139,30,123,31,77,31,201,31,206,31,45,31,45,30,27,31,27,30,248,31,118,31,7,31,103,31,14,31,14,30,67,31,57,31,21,31,149,31,107,31,123,31,7,31,7,30,7,29,8,31,136,31,52,31,38,31,80,31,153,31,7,31,22,31,22,30,68,31,68,30,120,31,85,31,225,31,74,31,144,31,92,31,238,31,36,31,224,31,49,31,239,31,88,31,49,31,184,31,90,31,243,31,222,31,112,31,94,31,223,31,91,31,55,31,183,31,164,31,189,31,182,31,182,30,31,31,180,31,158,31,137,31,170,31,127,31,20,31,59,31,59,30,59,29,178,31,178,30,178,29,178,28,201,31,196,31,196,30,122,31,166,31,133,31,211,31,211,30,236,31,119,31,97,31,97,30,197,31,152,31,251,31,251,30,205,31,205,30,205,29,205,28,84,31,223,31,179,31,132,31,138,31,115,31,128,31,196,31,196,30,196,29,171,31,171,30,193,31,193,30,47,31,240,31,58,31,58,30,185,31,185,30,62,31,165,31,157,31,85,31,21,31,115,31,28,31,65,31,65,30,125,31,125,30,113,31,53,31,143,31,119,31,116,31,163,31,163,30,171,31,171,30,250,31,86,31,189,31,240,31,24,31,141,31,141,30,223,31,159,31,136,31,136,30,90,31,238,31,238,30,240,31,240,30,18,31,230,31,230,30,177,31,85,31,56,31,226,31,76,31,43,31,167,31,192,31,192,30,15,31,15,30,15,29,230,31,2,31,125,31,125,30,230,31,230,30,176,31,16,31,80,31,42,31,42,30,129,31,113,31,46,31,93,31,49,31,217,31,217,30,93,31,235,31,83,31,241,31,241,30,241,29,154,31,203,31,7,31,248,31,157,31,125,31,8,31,23,31,154,31,30,31,30,30,93,31,182,31,6,31,236,31,236,30,118,31,83,31,166,31,37,31,37,30,151,31,170,31,12,31,241,31,130,31,39,31,155,31,93,31,93,30,246,31,197,31,194,31,116,31,43,31,113,31,250,31,76,31,53,31,67,31,209,31,229,31,238,31,221,31,129,31,226,31,79,31,79,30,183,31,183,30,252,31,193,31,41,31,195,31,220,31,214,31,207,31,112,31,166,31,190,31,246,31,50,31,253,31,51,31,47,31,5,31,30,31,49,31,89,31,197,31,228,31,181,31,181,30,226,31,226,30,156,31,186,31,186,30,138,31,15,31,205,31,96,31,39,31,33,31,160,31,17,31,17,30,71,31,251,31,251,30,58,31,211,31,231,31,249,31,194,31,252,31,159,31,65,31,65,30,247,31,176,31,152,31,142,31,142,30,126,31,50,31,142,31,109,31,199,31,199,30,199,29,189,31,189,30,91,31,186,31,239,31,109,31,109,30,109,29,79,31,79,30,117,31,76,31,88,31,88,30,9,31,9,30,228,31,177,31,235,31,116,31,224,31,67,31,114,31,199,31,84,31,18,31,56,31,32,31,32,30,32,29,210,31,218,31,102,31,102,30,102,29,106,31,102,31,102,30,102,29,201,31,201,30,210,31,115,31,47,31,48,31,245,31,236,31,236,30,236,29,236,28,82,31,228,31,180,31,129,31,129,30,243,31,159,31,159,30,94,31,206,31,206,30,206,29,207,31,56,31,56,30,78,31,191,31,225,31,170,31,213,31,98,31,61,31,114,31,93,31,237,31,248,31,248,30,95,31,21,31,148,31,126,31,8,31,203,31,241,31,174,31,147,31,201,31,87,31,77,31,164,31,4,31,4,30,146,31,120,31,66,31,47,31,47,30,25,31,49,31,137,31,168,31,168,30,22,31,22,30,22,29,80,31,1,31,188,31,25,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
