-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 782;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,6,0,253,0,202,0,182,0,0,0,0,0,119,0,39,0,199,0,136,0,12,0,0,0,179,0,208,0,0,0,69,0,3,0,119,0,186,0,0,0,0,0,0,0,129,0,205,0,27,0,35,0,125,0,80,0,235,0,181,0,0,0,249,0,248,0,149,0,0,0,150,0,201,0,170,0,12,0,247,0,195,0,131,0,203,0,31,0,0,0,14,0,213,0,174,0,234,0,92,0,244,0,176,0,129,0,110,0,133,0,0,0,104,0,0,0,165,0,199,0,12,0,182,0,127,0,146,0,203,0,52,0,0,0,0,0,113,0,0,0,59,0,78,0,53,0,132,0,173,0,0,0,172,0,158,0,86,0,57,0,170,0,145,0,227,0,13,0,215,0,131,0,206,0,100,0,167,0,116,0,0,0,178,0,92,0,200,0,149,0,124,0,0,0,107,0,0,0,148,0,254,0,206,0,178,0,220,0,64,0,196,0,209,0,26,0,111,0,0,0,230,0,245,0,224,0,61,0,247,0,151,0,250,0,0,0,0,0,4,0,198,0,56,0,139,0,147,0,0,0,0,0,187,0,156,0,107,0,0,0,236,0,83,0,0,0,83,0,0,0,110,0,0,0,94,0,241,0,179,0,211,0,22,0,67,0,27,0,254,0,90,0,57,0,144,0,132,0,21,0,163,0,0,0,3,0,46,0,243,0,110,0,0,0,71,0,87,0,0,0,196,0,228,0,68,0,0,0,97,0,32,0,120,0,81,0,12,0,66,0,0,0,0,0,202,0,0,0,0,0,104,0,61,0,152,0,0,0,122,0,161,0,105,0,137,0,236,0,0,0,176,0,0,0,70,0,211,0,0,0,0,0,241,0,222,0,218,0,161,0,250,0,0,0,150,0,186,0,0,0,0,0,30,0,86,0,0,0,19,0,199,0,67,0,0,0,105,0,170,0,66,0,0,0,45,0,11,0,112,0,147,0,120,0,125,0,88,0,0,0,151,0,248,0,0,0,169,0,0,0,89,0,0,0,237,0,34,0,22,0,226,0,0,0,0,0,0,0,75,0,98,0,226,0,187,0,18,0,40,0,0,0,107,0,153,0,195,0,188,0,175,0,36,0,20,0,129,0,41,0,134,0,0,0,0,0,94,0,0,0,142,0,127,0,152,0,22,0,39,0,124,0,224,0,250,0,0,0,7,0,120,0,109,0,0,0,13,0,116,0,104,0,0,0,0,0,25,0,196,0,57,0,66,0,0,0,13,0,196,0,184,0,0,0,240,0,53,0,0,0,79,0,250,0,97,0,44,0,130,0,188,0,181,0,86,0,185,0,119,0,242,0,70,0,0,0,202,0,167,0,214,0,164,0,49,0,0,0,180,0,56,0,9,0,0,0,206,0,225,0,196,0,154,0,0,0,247,0,178,0,35,0,112,0,163,0,69,0,73,0,0,0,237,0,108,0,104,0,38,0,172,0,0,0,61,0,211,0,122,0,0,0,122,0,64,0,43,0,220,0,0,0,229,0,0,0,97,0,134,0,245,0,171,0,29,0,29,0,116,0,0,0,123,0,0,0,108,0,14,0,0,0,40,0,164,0,62,0,128,0,57,0,229,0,0,0,200,0,177,0,72,0,200,0,217,0,0,0,173,0,0,0,144,0,5,0,76,0,0,0,59,0,103,0,209,0,0,0,177,0,240,0,173,0,46,0,238,0,172,0,23,0,238,0,51,0,79,0,97,0,0,0,0,0,43,0,137,0,0,0,48,0,185,0,94,0,82,0,37,0,65,0,61,0,120,0,255,0,123,0,102,0,250,0,252,0,0,0,154,0,205,0,159,0,109,0,182,0,221,0,244,0,239,0,5,0,0,0,176,0,231,0,137,0,0,0,113,0,147,0,172,0,48,0,246,0,121,0,147,0,0,0,120,0,60,0,233,0,243,0,0,0,0,0,0,0,138,0,0,0,27,0,0,0,205,0,0,0,167,0,0,0,252,0,69,0,51,0,0,0,0,0,248,0,0,0,0,0,103,0,173,0,175,0,17,0,136,0,0,0,40,0,119,0,0,0,0,0,0,0,0,0,0,0,250,0,0,0,245,0,0,0,233,0,151,0,22,0,0,0,203,0,0,0,172,0,106,0,0,0,168,0,92,0,147,0,129,0,5,0,138,0,180,0,177,0,0,0,103,0,143,0,3,0,18,0,131,0,35,0,21,0,208,0,119,0,216,0,220,0,0,0,56,0,187,0,0,0,167,0,183,0,235,0,131,0,0,0,0,0,173,0,255,0,135,0,0,0,225,0,0,0,21,0,0,0,14,0,0,0,0,0,134,0,204,0,86,0,77,0,0,0,25,0,4,0,0,0,205,0,141,0,8,0,223,0,0,0,0,0,0,0,0,0,57,0,0,0,247,0,31,0,49,0,0,0,127,0,118,0,80,0,129,0,103,0,20,0,3,0,172,0,0,0,0,0,97,0,99,0,126,0,166,0,0,0,49,0,251,0,42,0,179,0,217,0,138,0,0,0,207,0,174,0,71,0,17,0,133,0,203,0,0,0,153,0,74,0,0,0,10,0,137,0,186,0,3,0,60,0,37,0,239,0,60,0,0,0,14,0,73,0,27,0,100,0,44,0,41,0,0,0,241,0,0,0,58,0,0,0,174,0,68,0,43,0,50,0,217,0,46,0,233,0,124,0,23,0,0,0,71,0,85,0,0,0,191,0,115,0,138,0,0,0,0,0,217,0,44,0,87,0,0,0,5,0,212,0,86,0,6,0,198,0,195,0,230,0,0,0,0,0,181,0,181,0,151,0,27,0,130,0,0,0,214,0,27,0,70,0,122,0,22,0,0,0,0,0,157,0,0,0,50,0,154,0,152,0,29,0,0,0,3,0,159,0,0,0,252,0,40,0,109,0,82,0,115,0,56,0,120,0,188,0,54,0,123,0,101,0,0,0,139,0,43,0,193,0,203,0,234,0,89,0,226,0,0,0,203,0,15,0,0,0,0,0,0,0,0,0,176,0,243,0,0,0,229,0,95,0,0,0,184,0,0,0,98,0,8,0,107,0,56,0,90,0,0,0,173,0,98,0,238,0,0,0,87,0,0,0,28,0,0,0,8,0,0,0,247,0,205,0,91,0,53,0,30,0,92,0,141,0,0,0,0,0,7,0,1,0,70,0,202,0,158,0,182,0,133,0,112,0,0,0,60,0,0,0,43,0,154,0,149,0,231,0,41,0,223,0,13,0,0,0,0,0,0,0,254,0,231,0,0,0,13,0,139,0,189,0,117,0,47,0,158,0,167,0,117,0,34,0,66,0,0,0,214,0,143,0,148,0,14,0,69,0,149,0,143,0,206,0,99,0,130,0,0,0,0,0,0,0,166,0,231,0,64,0,233,0,0,0,34,0,253,0,179,0,150,0,105,0,0,0,61,0,0,0,0,0,0,0,0,0,0,0,121,0,133,0,208,0,27,0,0,0,90,0,165,0,164,0,23,0,13,0,153,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,6,31,253,31,202,31,182,31,182,30,182,29,119,31,39,31,199,31,136,31,12,31,12,30,179,31,208,31,208,30,69,31,3,31,119,31,186,31,186,30,186,29,186,28,129,31,205,31,27,31,35,31,125,31,80,31,235,31,181,31,181,30,249,31,248,31,149,31,149,30,150,31,201,31,170,31,12,31,247,31,195,31,131,31,203,31,31,31,31,30,14,31,213,31,174,31,234,31,92,31,244,31,176,31,129,31,110,31,133,31,133,30,104,31,104,30,165,31,199,31,12,31,182,31,127,31,146,31,203,31,52,31,52,30,52,29,113,31,113,30,59,31,78,31,53,31,132,31,173,31,173,30,172,31,158,31,86,31,57,31,170,31,145,31,227,31,13,31,215,31,131,31,206,31,100,31,167,31,116,31,116,30,178,31,92,31,200,31,149,31,124,31,124,30,107,31,107,30,148,31,254,31,206,31,178,31,220,31,64,31,196,31,209,31,26,31,111,31,111,30,230,31,245,31,224,31,61,31,247,31,151,31,250,31,250,30,250,29,4,31,198,31,56,31,139,31,147,31,147,30,147,29,187,31,156,31,107,31,107,30,236,31,83,31,83,30,83,31,83,30,110,31,110,30,94,31,241,31,179,31,211,31,22,31,67,31,27,31,254,31,90,31,57,31,144,31,132,31,21,31,163,31,163,30,3,31,46,31,243,31,110,31,110,30,71,31,87,31,87,30,196,31,228,31,68,31,68,30,97,31,32,31,120,31,81,31,12,31,66,31,66,30,66,29,202,31,202,30,202,29,104,31,61,31,152,31,152,30,122,31,161,31,105,31,137,31,236,31,236,30,176,31,176,30,70,31,211,31,211,30,211,29,241,31,222,31,218,31,161,31,250,31,250,30,150,31,186,31,186,30,186,29,30,31,86,31,86,30,19,31,199,31,67,31,67,30,105,31,170,31,66,31,66,30,45,31,11,31,112,31,147,31,120,31,125,31,88,31,88,30,151,31,248,31,248,30,169,31,169,30,89,31,89,30,237,31,34,31,22,31,226,31,226,30,226,29,226,28,75,31,98,31,226,31,187,31,18,31,40,31,40,30,107,31,153,31,195,31,188,31,175,31,36,31,20,31,129,31,41,31,134,31,134,30,134,29,94,31,94,30,142,31,127,31,152,31,22,31,39,31,124,31,224,31,250,31,250,30,7,31,120,31,109,31,109,30,13,31,116,31,104,31,104,30,104,29,25,31,196,31,57,31,66,31,66,30,13,31,196,31,184,31,184,30,240,31,53,31,53,30,79,31,250,31,97,31,44,31,130,31,188,31,181,31,86,31,185,31,119,31,242,31,70,31,70,30,202,31,167,31,214,31,164,31,49,31,49,30,180,31,56,31,9,31,9,30,206,31,225,31,196,31,154,31,154,30,247,31,178,31,35,31,112,31,163,31,69,31,73,31,73,30,237,31,108,31,104,31,38,31,172,31,172,30,61,31,211,31,122,31,122,30,122,31,64,31,43,31,220,31,220,30,229,31,229,30,97,31,134,31,245,31,171,31,29,31,29,31,116,31,116,30,123,31,123,30,108,31,14,31,14,30,40,31,164,31,62,31,128,31,57,31,229,31,229,30,200,31,177,31,72,31,200,31,217,31,217,30,173,31,173,30,144,31,5,31,76,31,76,30,59,31,103,31,209,31,209,30,177,31,240,31,173,31,46,31,238,31,172,31,23,31,238,31,51,31,79,31,97,31,97,30,97,29,43,31,137,31,137,30,48,31,185,31,94,31,82,31,37,31,65,31,61,31,120,31,255,31,123,31,102,31,250,31,252,31,252,30,154,31,205,31,159,31,109,31,182,31,221,31,244,31,239,31,5,31,5,30,176,31,231,31,137,31,137,30,113,31,147,31,172,31,48,31,246,31,121,31,147,31,147,30,120,31,60,31,233,31,243,31,243,30,243,29,243,28,138,31,138,30,27,31,27,30,205,31,205,30,167,31,167,30,252,31,69,31,51,31,51,30,51,29,248,31,248,30,248,29,103,31,173,31,175,31,17,31,136,31,136,30,40,31,119,31,119,30,119,29,119,28,119,27,119,26,250,31,250,30,245,31,245,30,233,31,151,31,22,31,22,30,203,31,203,30,172,31,106,31,106,30,168,31,92,31,147,31,129,31,5,31,138,31,180,31,177,31,177,30,103,31,143,31,3,31,18,31,131,31,35,31,21,31,208,31,119,31,216,31,220,31,220,30,56,31,187,31,187,30,167,31,183,31,235,31,131,31,131,30,131,29,173,31,255,31,135,31,135,30,225,31,225,30,21,31,21,30,14,31,14,30,14,29,134,31,204,31,86,31,77,31,77,30,25,31,4,31,4,30,205,31,141,31,8,31,223,31,223,30,223,29,223,28,223,27,57,31,57,30,247,31,31,31,49,31,49,30,127,31,118,31,80,31,129,31,103,31,20,31,3,31,172,31,172,30,172,29,97,31,99,31,126,31,166,31,166,30,49,31,251,31,42,31,179,31,217,31,138,31,138,30,207,31,174,31,71,31,17,31,133,31,203,31,203,30,153,31,74,31,74,30,10,31,137,31,186,31,3,31,60,31,37,31,239,31,60,31,60,30,14,31,73,31,27,31,100,31,44,31,41,31,41,30,241,31,241,30,58,31,58,30,174,31,68,31,43,31,50,31,217,31,46,31,233,31,124,31,23,31,23,30,71,31,85,31,85,30,191,31,115,31,138,31,138,30,138,29,217,31,44,31,87,31,87,30,5,31,212,31,86,31,6,31,198,31,195,31,230,31,230,30,230,29,181,31,181,31,151,31,27,31,130,31,130,30,214,31,27,31,70,31,122,31,22,31,22,30,22,29,157,31,157,30,50,31,154,31,152,31,29,31,29,30,3,31,159,31,159,30,252,31,40,31,109,31,82,31,115,31,56,31,120,31,188,31,54,31,123,31,101,31,101,30,139,31,43,31,193,31,203,31,234,31,89,31,226,31,226,30,203,31,15,31,15,30,15,29,15,28,15,27,176,31,243,31,243,30,229,31,95,31,95,30,184,31,184,30,98,31,8,31,107,31,56,31,90,31,90,30,173,31,98,31,238,31,238,30,87,31,87,30,28,31,28,30,8,31,8,30,247,31,205,31,91,31,53,31,30,31,92,31,141,31,141,30,141,29,7,31,1,31,70,31,202,31,158,31,182,31,133,31,112,31,112,30,60,31,60,30,43,31,154,31,149,31,231,31,41,31,223,31,13,31,13,30,13,29,13,28,254,31,231,31,231,30,13,31,139,31,189,31,117,31,47,31,158,31,167,31,117,31,34,31,66,31,66,30,214,31,143,31,148,31,14,31,69,31,149,31,143,31,206,31,99,31,130,31,130,30,130,29,130,28,166,31,231,31,64,31,233,31,233,30,34,31,253,31,179,31,150,31,105,31,105,30,61,31,61,30,61,29,61,28,61,27,61,26,121,31,133,31,208,31,27,31,27,30,90,31,165,31,164,31,23,31,13,31,153,31,153,30,153,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
