-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_36 is
end project_tb_36;

architecture project_tb_arch_36 of project_tb_36 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,20,0,72,0,0,0,0,0,226,0,74,0,25,0,121,0,101,0,190,0,0,0,243,0,0,0,0,0,29,0,0,0,132,0,117,0,246,0,171,0,0,0,207,0,58,0,0,0,95,0,136,0,136,0,13,0,137,0,28,0,132,0,246,0,185,0,1,0,185,0,171,0,0,0,136,0,48,0,250,0,195,0,0,0,0,0,62,0,175,0,244,0,235,0,240,0,96,0,122,0,110,0,0,0,66,0,37,0,0,0,69,0,6,0,0,0,118,0,0,0,26,0,66,0,0,0,179,0,187,0,71,0,16,0,25,0,133,0,0,0,65,0,72,0,95,0,158,0,0,0,52,0,190,0,252,0,177,0,186,0,170,0,240,0,106,0,0,0,215,0,167,0,45,0,0,0,8,0,3,0,56,0,116,0,0,0,0,0,11,0,30,0,70,0,86,0,212,0,138,0,180,0,253,0,71,0,159,0,59,0,130,0,85,0,0,0,232,0,170,0,146,0,36,0,84,0,0,0,26,0,112,0,165,0,244,0,0,0,127,0,216,0,0,0,216,0,106,0,39,0,104,0,201,0,166,0,229,0,0,0,36,0,216,0,56,0,0,0,0,0,0,0,108,0,208,0,180,0,127,0,0,0,13,0,20,0,201,0,188,0,0,0,97,0,65,0,182,0,0,0,52,0,27,0,222,0,61,0,0,0,0,0,0,0,161,0,1,0,129,0,100,0,250,0,142,0,0,0,120,0,20,0,63,0,217,0,99,0,165,0,227,0,163,0,183,0,113,0,0,0,227,0,79,0,35,0,35,0,122,0,140,0,0,0,178,0,0,0,127,0,42,0,0,0,197,0,253,0,56,0,194,0,121,0,215,0,113,0,51,0,66,0,41,0,209,0,167,0,0,0,39,0,243,0,14,0,0,0,0,0,251,0,100,0,180,0,213,0,0,0,141,0,177,0,255,0,0,0,0,0,253,0,13,0,142,0,198,0,230,0,0,0,103,0,252,0,109,0,175,0,204,0,68,0,174,0,68,0,0,0,0,0,39,0,0,0,175,0,211,0,4,0,0,0,0,0,237,0,133,0,13,0,154,0,87,0,29,0,0,0,234,0,182,0,0,0,210,0,131,0,52,0,215,0,156,0,251,0,73,0,0,0,151,0,0,0,131,0,64,0,170,0,68,0,198,0,171,0,142,0,20,0,157,0,201,0,72,0,40,0,222,0,197,0,42,0,210,0,165,0,148,0,120,0,248,0,116,0,75,0,0,0,243,0,218,0,159,0,0,0,191,0,0,0,217,0,15,0,142,0,167,0,127,0,253,0,199,0,78,0,61,0,71,0,0,0,0,0,17,0,83,0,136,0,132,0,109,0,129,0,0,0,130,0,140,0,176,0,92,0,0,0,29,0,82,0,252,0,248,0,203,0,0,0,214,0,189,0,9,0,9,0,35,0,146,0,53,0,217,0,255,0,128,0,97,0,172,0,174,0,0,0,6,0,158,0,25,0,220,0,0,0,40,0,144,0,0,0,7,0,1,0,120,0,0,0,126,0,111,0,142,0,0,0,30,0,35,0,84,0,9,0,148,0,222,0,43,0,13,0,28,0,139,0,27,0,152,0,8,0,81,0,0,0,161,0,23,0,0,0,44,0,136,0,0,0,0,0,0,0,0,0,173,0,136,0,93,0,234,0,0,0,216,0,9,0,151,0,244,0,81,0,0,0,254,0,156,0,209,0,150,0,150,0,193,0,237,0,17,0,0,0,33,0,0,0,0,0,42,0,151,0,61,0,39,0,52,0,187,0,84,0,137,0,201,0,0,0,92,0,116,0,0,0,0,0,173,0,0,0,254,0,0,0,155,0,153,0,86,0,16,0,76,0,65,0,114,0,121,0,124,0,124,0,0,0,196,0,179,0,66,0,248,0,141,0,235,0,0,0,53,0,144,0,177,0,213,0,129,0,205,0,177,0,0,0,233,0,16,0,106,0,198,0,42,0,221,0,61,0,153,0,32,0,149,0,66,0,81,0,0,0,130,0,203,0,0,0,27,0,228,0,157,0,235,0,186,0,219,0,21,0,135,0,73,0,63,0,209,0,127,0,0,0,15,0,255,0,250,0,0,0,242,0,0,0,48,0,100,0,53,0,131,0,105,0,221,0,0,0,162,0,81,0,233,0,158,0,227,0,240,0,200,0,184,0,131,0,130,0,63,0,58,0,0,0,0,0,118,0,0,0,209,0,0,0,122,0,0,0,219,0,242,0,107,0,117,0,254,0,5,0,138,0,18,0,0,0,52,0,151,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,114,0,0,0,204,0,49,0,72,0,220,0,0,0,0,0,55,0,100,0,224,0,90,0,0,0,253,0,40,0,167,0,183,0,0,0,103,0,180,0,163,0,0,0,0,0,139,0,137,0,143,0,156,0,178,0,195,0,169,0,143,0,239,0,225,0,69,0,34,0,211,0,50,0,229,0,250,0,0,0,172,0,0,0,250,0,0,0,19,0,23,0,179,0,144,0,29,0,129,0,0,0,18,0,29,0,0,0,148,0,0,0,64,0,147,0,169,0,0,0,171,0,149,0,158,0,124,0,51,0,0,0,250,0,119,0,109,0,54,0,230,0,0,0,57,0,205,0,107,0,0,0,61,0,205,0,35,0,248,0,166,0,179,0,72,0,108,0,101,0,41,0,215,0,0,0,224,0,200,0,40,0,156,0,72,0,98,0,116,0,176,0,126,0,78,0,0,0,28,0,53,0,171,0,86,0,0,0,124,0,8,0,43,0,0,0,150,0,118,0,132,0,104,0,140,0,53,0,40,0,0,0,227,0,0,0,191,0,240,0,0,0,147,0,186,0,214,0,115,0,134,0);
signal scenario_full  : scenario_type := (0,0,0,0,20,31,72,31,72,30,72,29,226,31,74,31,25,31,121,31,101,31,190,31,190,30,243,31,243,30,243,29,29,31,29,30,132,31,117,31,246,31,171,31,171,30,207,31,58,31,58,30,95,31,136,31,136,31,13,31,137,31,28,31,132,31,246,31,185,31,1,31,185,31,171,31,171,30,136,31,48,31,250,31,195,31,195,30,195,29,62,31,175,31,244,31,235,31,240,31,96,31,122,31,110,31,110,30,66,31,37,31,37,30,69,31,6,31,6,30,118,31,118,30,26,31,66,31,66,30,179,31,187,31,71,31,16,31,25,31,133,31,133,30,65,31,72,31,95,31,158,31,158,30,52,31,190,31,252,31,177,31,186,31,170,31,240,31,106,31,106,30,215,31,167,31,45,31,45,30,8,31,3,31,56,31,116,31,116,30,116,29,11,31,30,31,70,31,86,31,212,31,138,31,180,31,253,31,71,31,159,31,59,31,130,31,85,31,85,30,232,31,170,31,146,31,36,31,84,31,84,30,26,31,112,31,165,31,244,31,244,30,127,31,216,31,216,30,216,31,106,31,39,31,104,31,201,31,166,31,229,31,229,30,36,31,216,31,56,31,56,30,56,29,56,28,108,31,208,31,180,31,127,31,127,30,13,31,20,31,201,31,188,31,188,30,97,31,65,31,182,31,182,30,52,31,27,31,222,31,61,31,61,30,61,29,61,28,161,31,1,31,129,31,100,31,250,31,142,31,142,30,120,31,20,31,63,31,217,31,99,31,165,31,227,31,163,31,183,31,113,31,113,30,227,31,79,31,35,31,35,31,122,31,140,31,140,30,178,31,178,30,127,31,42,31,42,30,197,31,253,31,56,31,194,31,121,31,215,31,113,31,51,31,66,31,41,31,209,31,167,31,167,30,39,31,243,31,14,31,14,30,14,29,251,31,100,31,180,31,213,31,213,30,141,31,177,31,255,31,255,30,255,29,253,31,13,31,142,31,198,31,230,31,230,30,103,31,252,31,109,31,175,31,204,31,68,31,174,31,68,31,68,30,68,29,39,31,39,30,175,31,211,31,4,31,4,30,4,29,237,31,133,31,13,31,154,31,87,31,29,31,29,30,234,31,182,31,182,30,210,31,131,31,52,31,215,31,156,31,251,31,73,31,73,30,151,31,151,30,131,31,64,31,170,31,68,31,198,31,171,31,142,31,20,31,157,31,201,31,72,31,40,31,222,31,197,31,42,31,210,31,165,31,148,31,120,31,248,31,116,31,75,31,75,30,243,31,218,31,159,31,159,30,191,31,191,30,217,31,15,31,142,31,167,31,127,31,253,31,199,31,78,31,61,31,71,31,71,30,71,29,17,31,83,31,136,31,132,31,109,31,129,31,129,30,130,31,140,31,176,31,92,31,92,30,29,31,82,31,252,31,248,31,203,31,203,30,214,31,189,31,9,31,9,31,35,31,146,31,53,31,217,31,255,31,128,31,97,31,172,31,174,31,174,30,6,31,158,31,25,31,220,31,220,30,40,31,144,31,144,30,7,31,1,31,120,31,120,30,126,31,111,31,142,31,142,30,30,31,35,31,84,31,9,31,148,31,222,31,43,31,13,31,28,31,139,31,27,31,152,31,8,31,81,31,81,30,161,31,23,31,23,30,44,31,136,31,136,30,136,29,136,28,136,27,173,31,136,31,93,31,234,31,234,30,216,31,9,31,151,31,244,31,81,31,81,30,254,31,156,31,209,31,150,31,150,31,193,31,237,31,17,31,17,30,33,31,33,30,33,29,42,31,151,31,61,31,39,31,52,31,187,31,84,31,137,31,201,31,201,30,92,31,116,31,116,30,116,29,173,31,173,30,254,31,254,30,155,31,153,31,86,31,16,31,76,31,65,31,114,31,121,31,124,31,124,31,124,30,196,31,179,31,66,31,248,31,141,31,235,31,235,30,53,31,144,31,177,31,213,31,129,31,205,31,177,31,177,30,233,31,16,31,106,31,198,31,42,31,221,31,61,31,153,31,32,31,149,31,66,31,81,31,81,30,130,31,203,31,203,30,27,31,228,31,157,31,235,31,186,31,219,31,21,31,135,31,73,31,63,31,209,31,127,31,127,30,15,31,255,31,250,31,250,30,242,31,242,30,48,31,100,31,53,31,131,31,105,31,221,31,221,30,162,31,81,31,233,31,158,31,227,31,240,31,200,31,184,31,131,31,130,31,63,31,58,31,58,30,58,29,118,31,118,30,209,31,209,30,122,31,122,30,219,31,242,31,107,31,117,31,254,31,5,31,138,31,18,31,18,30,52,31,151,31,151,30,151,29,151,28,151,27,151,26,151,25,151,24,114,31,114,30,204,31,49,31,72,31,220,31,220,30,220,29,55,31,100,31,224,31,90,31,90,30,253,31,40,31,167,31,183,31,183,30,103,31,180,31,163,31,163,30,163,29,139,31,137,31,143,31,156,31,178,31,195,31,169,31,143,31,239,31,225,31,69,31,34,31,211,31,50,31,229,31,250,31,250,30,172,31,172,30,250,31,250,30,19,31,23,31,179,31,144,31,29,31,129,31,129,30,18,31,29,31,29,30,148,31,148,30,64,31,147,31,169,31,169,30,171,31,149,31,158,31,124,31,51,31,51,30,250,31,119,31,109,31,54,31,230,31,230,30,57,31,205,31,107,31,107,30,61,31,205,31,35,31,248,31,166,31,179,31,72,31,108,31,101,31,41,31,215,31,215,30,224,31,200,31,40,31,156,31,72,31,98,31,116,31,176,31,126,31,78,31,78,30,28,31,53,31,171,31,86,31,86,30,124,31,8,31,43,31,43,30,150,31,118,31,132,31,104,31,140,31,53,31,40,31,40,30,227,31,227,30,191,31,240,31,240,30,147,31,186,31,214,31,115,31,134,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
