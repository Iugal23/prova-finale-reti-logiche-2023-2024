-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_685 is
end project_tb_685;

architecture project_tb_arch_685 of project_tb_685 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 379;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,177,0,232,0,156,0,198,0,242,0,0,0,35,0,138,0,224,0,117,0,125,0,214,0,20,0,85,0,33,0,11,0,72,0,199,0,134,0,38,0,139,0,18,0,44,0,81,0,157,0,0,0,0,0,0,0,59,0,0,0,70,0,34,0,115,0,10,0,0,0,108,0,69,0,49,0,12,0,0,0,0,0,0,0,114,0,3,0,163,0,0,0,55,0,188,0,102,0,115,0,170,0,136,0,243,0,207,0,74,0,244,0,135,0,90,0,204,0,0,0,0,0,202,0,200,0,191,0,212,0,96,0,169,0,0,0,107,0,150,0,157,0,0,0,190,0,31,0,0,0,0,0,48,0,0,0,2,0,62,0,7,0,0,0,0,0,32,0,210,0,15,0,0,0,0,0,14,0,0,0,133,0,91,0,235,0,65,0,46,0,88,0,235,0,163,0,217,0,0,0,0,0,0,0,130,0,0,0,46,0,235,0,9,0,150,0,67,0,0,0,229,0,0,0,0,0,96,0,136,0,100,0,42,0,30,0,217,0,34,0,214,0,56,0,251,0,0,0,139,0,242,0,0,0,143,0,191,0,0,0,76,0,0,0,0,0,234,0,25,0,87,0,250,0,0,0,109,0,112,0,80,0,167,0,0,0,0,0,148,0,158,0,0,0,103,0,152,0,209,0,170,0,200,0,8,0,86,0,72,0,47,0,0,0,0,0,128,0,52,0,186,0,69,0,150,0,0,0,59,0,30,0,166,0,213,0,0,0,141,0,75,0,129,0,0,0,0,0,251,0,0,0,118,0,127,0,0,0,234,0,205,0,24,0,0,0,135,0,2,0,137,0,155,0,136,0,180,0,150,0,0,0,219,0,92,0,131,0,75,0,235,0,158,0,202,0,179,0,227,0,39,0,0,0,0,0,21,0,70,0,183,0,75,0,37,0,140,0,135,0,116,0,115,0,243,0,141,0,41,0,0,0,96,0,41,0,0,0,7,0,239,0,69,0,184,0,49,0,103,0,179,0,27,0,163,0,195,0,55,0,91,0,0,0,112,0,88,0,0,0,229,0,84,0,0,0,0,0,209,0,0,0,140,0,117,0,113,0,173,0,164,0,125,0,121,0,226,0,24,0,175,0,125,0,0,0,22,0,248,0,212,0,31,0,54,0,108,0,220,0,0,0,46,0,52,0,124,0,10,0,0,0,19,0,0,0,54,0,35,0,164,0,0,0,247,0,0,0,172,0,67,0,58,0,230,0,248,0,57,0,0,0,0,0,145,0,119,0,0,0,249,0,0,0,250,0,181,0,220,0,195,0,86,0,50,0,240,0,75,0,32,0,107,0,102,0,173,0,102,0,70,0,0,0,71,0,10,0,137,0,56,0,240,0,0,0,160,0,0,0,124,0,0,0,134,0,49,0,123,0,25,0,0,0,208,0,162,0,188,0,234,0,0,0,72,0,247,0,46,0,187,0,130,0,0,0,39,0,0,0,40,0,59,0,0,0,106,0,103,0,29,0,91,0,0,0,245,0,213,0,253,0,119,0,0,0,73,0,0,0,109,0,120,0,110,0,43,0,79,0,0,0,90,0,5,0,17,0,162,0,0,0,186,0,243,0,207,0,60,0,77,0,0,0,89,0,137,0,97,0,41,0,126,0,199,0,252,0,198,0,227,0,222,0,193,0,0,0,0,0,0,0,138,0,93,0);
signal scenario_full  : scenario_type := (214,31,177,31,232,31,156,31,198,31,242,31,242,30,35,31,138,31,224,31,117,31,125,31,214,31,20,31,85,31,33,31,11,31,72,31,199,31,134,31,38,31,139,31,18,31,44,31,81,31,157,31,157,30,157,29,157,28,59,31,59,30,70,31,34,31,115,31,10,31,10,30,108,31,69,31,49,31,12,31,12,30,12,29,12,28,114,31,3,31,163,31,163,30,55,31,188,31,102,31,115,31,170,31,136,31,243,31,207,31,74,31,244,31,135,31,90,31,204,31,204,30,204,29,202,31,200,31,191,31,212,31,96,31,169,31,169,30,107,31,150,31,157,31,157,30,190,31,31,31,31,30,31,29,48,31,48,30,2,31,62,31,7,31,7,30,7,29,32,31,210,31,15,31,15,30,15,29,14,31,14,30,133,31,91,31,235,31,65,31,46,31,88,31,235,31,163,31,217,31,217,30,217,29,217,28,130,31,130,30,46,31,235,31,9,31,150,31,67,31,67,30,229,31,229,30,229,29,96,31,136,31,100,31,42,31,30,31,217,31,34,31,214,31,56,31,251,31,251,30,139,31,242,31,242,30,143,31,191,31,191,30,76,31,76,30,76,29,234,31,25,31,87,31,250,31,250,30,109,31,112,31,80,31,167,31,167,30,167,29,148,31,158,31,158,30,103,31,152,31,209,31,170,31,200,31,8,31,86,31,72,31,47,31,47,30,47,29,128,31,52,31,186,31,69,31,150,31,150,30,59,31,30,31,166,31,213,31,213,30,141,31,75,31,129,31,129,30,129,29,251,31,251,30,118,31,127,31,127,30,234,31,205,31,24,31,24,30,135,31,2,31,137,31,155,31,136,31,180,31,150,31,150,30,219,31,92,31,131,31,75,31,235,31,158,31,202,31,179,31,227,31,39,31,39,30,39,29,21,31,70,31,183,31,75,31,37,31,140,31,135,31,116,31,115,31,243,31,141,31,41,31,41,30,96,31,41,31,41,30,7,31,239,31,69,31,184,31,49,31,103,31,179,31,27,31,163,31,195,31,55,31,91,31,91,30,112,31,88,31,88,30,229,31,84,31,84,30,84,29,209,31,209,30,140,31,117,31,113,31,173,31,164,31,125,31,121,31,226,31,24,31,175,31,125,31,125,30,22,31,248,31,212,31,31,31,54,31,108,31,220,31,220,30,46,31,52,31,124,31,10,31,10,30,19,31,19,30,54,31,35,31,164,31,164,30,247,31,247,30,172,31,67,31,58,31,230,31,248,31,57,31,57,30,57,29,145,31,119,31,119,30,249,31,249,30,250,31,181,31,220,31,195,31,86,31,50,31,240,31,75,31,32,31,107,31,102,31,173,31,102,31,70,31,70,30,71,31,10,31,137,31,56,31,240,31,240,30,160,31,160,30,124,31,124,30,134,31,49,31,123,31,25,31,25,30,208,31,162,31,188,31,234,31,234,30,72,31,247,31,46,31,187,31,130,31,130,30,39,31,39,30,40,31,59,31,59,30,106,31,103,31,29,31,91,31,91,30,245,31,213,31,253,31,119,31,119,30,73,31,73,30,109,31,120,31,110,31,43,31,79,31,79,30,90,31,5,31,17,31,162,31,162,30,186,31,243,31,207,31,60,31,77,31,77,30,89,31,137,31,97,31,41,31,126,31,199,31,252,31,198,31,227,31,222,31,193,31,193,30,193,29,193,28,138,31,93,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
