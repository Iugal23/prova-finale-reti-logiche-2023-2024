-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_936 is
end project_tb_936;

architecture project_tb_arch_936 of project_tb_936 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 709;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (78,0,0,0,184,0,197,0,104,0,224,0,222,0,75,0,194,0,194,0,0,0,118,0,142,0,0,0,125,0,0,0,143,0,177,0,0,0,60,0,32,0,200,0,147,0,103,0,145,0,23,0,105,0,203,0,196,0,0,0,105,0,0,0,141,0,75,0,158,0,0,0,182,0,61,0,9,0,82,0,72,0,126,0,0,0,169,0,103,0,69,0,212,0,0,0,0,0,147,0,51,0,171,0,133,0,226,0,0,0,46,0,65,0,116,0,132,0,0,0,50,0,11,0,0,0,179,0,254,0,243,0,0,0,210,0,183,0,29,0,117,0,233,0,141,0,42,0,0,0,0,0,10,0,110,0,124,0,0,0,51,0,205,0,149,0,126,0,189,0,230,0,190,0,176,0,44,0,169,0,93,0,105,0,163,0,113,0,125,0,0,0,125,0,0,0,82,0,55,0,0,0,174,0,61,0,0,0,0,0,97,0,95,0,65,0,140,0,80,0,31,0,35,0,0,0,213,0,107,0,0,0,175,0,158,0,251,0,152,0,137,0,62,0,151,0,46,0,8,0,30,0,157,0,47,0,247,0,0,0,136,0,133,0,1,0,144,0,0,0,24,0,0,0,255,0,78,0,0,0,209,0,101,0,69,0,136,0,34,0,66,0,0,0,0,0,131,0,196,0,139,0,181,0,113,0,191,0,46,0,108,0,92,0,101,0,34,0,242,0,6,0,232,0,75,0,205,0,0,0,63,0,112,0,89,0,17,0,0,0,0,0,227,0,0,0,0,0,0,0,0,0,211,0,97,0,100,0,15,0,26,0,4,0,74,0,186,0,141,0,196,0,0,0,19,0,185,0,104,0,0,0,199,0,110,0,48,0,136,0,246,0,66,0,96,0,203,0,201,0,0,0,18,0,58,0,102,0,222,0,0,0,246,0,137,0,246,0,218,0,45,0,167,0,0,0,0,0,0,0,106,0,123,0,60,0,164,0,0,0,58,0,83,0,98,0,148,0,0,0,0,0,27,0,129,0,237,0,19,0,205,0,0,0,120,0,180,0,143,0,153,0,247,0,141,0,0,0,109,0,40,0,42,0,11,0,0,0,0,0,240,0,173,0,189,0,66,0,20,0,0,0,0,0,163,0,172,0,204,0,0,0,251,0,69,0,132,0,237,0,245,0,80,0,123,0,247,0,0,0,252,0,98,0,182,0,170,0,0,0,248,0,218,0,216,0,126,0,96,0,117,0,116,0,239,0,200,0,204,0,35,0,131,0,232,0,169,0,161,0,0,0,0,0,50,0,27,0,195,0,153,0,0,0,44,0,36,0,0,0,0,0,215,0,179,0,15,0,0,0,98,0,87,0,119,0,0,0,134,0,252,0,156,0,159,0,0,0,167,0,45,0,175,0,62,0,215,0,210,0,113,0,61,0,83,0,4,0,17,0,23,0,15,0,130,0,237,0,88,0,251,0,0,0,19,0,231,0,133,0,120,0,105,0,0,0,56,0,101,0,164,0,128,0,141,0,0,0,170,0,13,0,249,0,95,0,113,0,57,0,29,0,53,0,224,0,47,0,35,0,224,0,170,0,77,0,149,0,203,0,0,0,53,0,233,0,64,0,143,0,21,0,32,0,0,0,70,0,72,0,203,0,113,0,0,0,140,0,142,0,0,0,0,0,96,0,217,0,0,0,0,0,75,0,105,0,199,0,51,0,83,0,0,0,126,0,202,0,182,0,80,0,79,0,95,0,118,0,131,0,239,0,42,0,44,0,0,0,236,0,170,0,199,0,152,0,237,0,0,0,191,0,111,0,83,0,14,0,222,0,35,0,60,0,113,0,89,0,21,0,50,0,0,0,157,0,184,0,225,0,0,0,233,0,217,0,107,0,53,0,255,0,96,0,39,0,0,0,143,0,19,0,44,0,10,0,228,0,0,0,0,0,3,0,36,0,0,0,0,0,34,0,138,0,95,0,74,0,243,0,0,0,0,0,149,0,59,0,97,0,28,0,0,0,30,0,0,0,0,0,255,0,0,0,30,0,0,0,120,0,121,0,209,0,60,0,228,0,193,0,87,0,41,0,46,0,190,0,34,0,0,0,172,0,160,0,0,0,212,0,196,0,164,0,25,0,52,0,158,0,37,0,247,0,170,0,0,0,163,0,144,0,0,0,169,0,234,0,162,0,231,0,169,0,209,0,61,0,174,0,209,0,53,0,192,0,0,0,108,0,0,0,0,0,252,0,0,0,0,0,113,0,32,0,207,0,79,0,231,0,0,0,0,0,180,0,60,0,68,0,68,0,253,0,20,0,112,0,3,0,0,0,12,0,0,0,129,0,214,0,2,0,93,0,65,0,75,0,0,0,0,0,157,0,167,0,91,0,0,0,202,0,7,0,0,0,0,0,83,0,0,0,142,0,214,0,0,0,11,0,0,0,0,0,254,0,51,0,0,0,20,0,232,0,48,0,0,0,57,0,0,0,217,0,27,0,143,0,22,0,229,0,70,0,109,0,138,0,60,0,205,0,183,0,233,0,191,0,210,0,0,0,0,0,141,0,129,0,231,0,24,0,10,0,117,0,128,0,0,0,31,0,8,0,192,0,189,0,87,0,140,0,143,0,20,0,136,0,210,0,0,0,153,0,34,0,1,0,226,0,74,0,35,0,197,0,6,0,47,0,0,0,100,0,174,0,23,0,76,0,52,0,103,0,61,0,123,0,230,0,42,0,95,0,0,0,130,0,0,0,19,0,111,0,0,0,133,0,0,0,69,0,101,0,34,0,173,0,0,0,209,0,243,0,205,0,165,0,8,0,0,0,0,0,100,0,92,0,33,0,172,0,0,0,0,0,125,0,46,0,137,0,0,0,111,0,198,0,0,0,203,0,206,0,0,0,60,0,224,0,253,0,245,0,196,0,0,0,0,0,250,0,226,0,34,0,235,0,230,0,0,0,0,0,118,0,83,0,51,0,243,0,57,0,0,0,43,0,30,0,183,0,0,0,35,0,69,0,157,0,146,0,164,0,163,0,198,0,138,0,116,0,208,0,124,0,48,0,129,0,187,0,234,0,0,0,0,0,74,0,215,0,228,0,241,0,0,0,197,0,254,0,0,0,176,0,0,0,251,0,173,0,191,0,0,0,0,0,0,0,184,0,0,0,0,0,88,0,53,0,33,0,234,0,33,0,83,0);
signal scenario_full  : scenario_type := (78,31,78,30,184,31,197,31,104,31,224,31,222,31,75,31,194,31,194,31,194,30,118,31,142,31,142,30,125,31,125,30,143,31,177,31,177,30,60,31,32,31,200,31,147,31,103,31,145,31,23,31,105,31,203,31,196,31,196,30,105,31,105,30,141,31,75,31,158,31,158,30,182,31,61,31,9,31,82,31,72,31,126,31,126,30,169,31,103,31,69,31,212,31,212,30,212,29,147,31,51,31,171,31,133,31,226,31,226,30,46,31,65,31,116,31,132,31,132,30,50,31,11,31,11,30,179,31,254,31,243,31,243,30,210,31,183,31,29,31,117,31,233,31,141,31,42,31,42,30,42,29,10,31,110,31,124,31,124,30,51,31,205,31,149,31,126,31,189,31,230,31,190,31,176,31,44,31,169,31,93,31,105,31,163,31,113,31,125,31,125,30,125,31,125,30,82,31,55,31,55,30,174,31,61,31,61,30,61,29,97,31,95,31,65,31,140,31,80,31,31,31,35,31,35,30,213,31,107,31,107,30,175,31,158,31,251,31,152,31,137,31,62,31,151,31,46,31,8,31,30,31,157,31,47,31,247,31,247,30,136,31,133,31,1,31,144,31,144,30,24,31,24,30,255,31,78,31,78,30,209,31,101,31,69,31,136,31,34,31,66,31,66,30,66,29,131,31,196,31,139,31,181,31,113,31,191,31,46,31,108,31,92,31,101,31,34,31,242,31,6,31,232,31,75,31,205,31,205,30,63,31,112,31,89,31,17,31,17,30,17,29,227,31,227,30,227,29,227,28,227,27,211,31,97,31,100,31,15,31,26,31,4,31,74,31,186,31,141,31,196,31,196,30,19,31,185,31,104,31,104,30,199,31,110,31,48,31,136,31,246,31,66,31,96,31,203,31,201,31,201,30,18,31,58,31,102,31,222,31,222,30,246,31,137,31,246,31,218,31,45,31,167,31,167,30,167,29,167,28,106,31,123,31,60,31,164,31,164,30,58,31,83,31,98,31,148,31,148,30,148,29,27,31,129,31,237,31,19,31,205,31,205,30,120,31,180,31,143,31,153,31,247,31,141,31,141,30,109,31,40,31,42,31,11,31,11,30,11,29,240,31,173,31,189,31,66,31,20,31,20,30,20,29,163,31,172,31,204,31,204,30,251,31,69,31,132,31,237,31,245,31,80,31,123,31,247,31,247,30,252,31,98,31,182,31,170,31,170,30,248,31,218,31,216,31,126,31,96,31,117,31,116,31,239,31,200,31,204,31,35,31,131,31,232,31,169,31,161,31,161,30,161,29,50,31,27,31,195,31,153,31,153,30,44,31,36,31,36,30,36,29,215,31,179,31,15,31,15,30,98,31,87,31,119,31,119,30,134,31,252,31,156,31,159,31,159,30,167,31,45,31,175,31,62,31,215,31,210,31,113,31,61,31,83,31,4,31,17,31,23,31,15,31,130,31,237,31,88,31,251,31,251,30,19,31,231,31,133,31,120,31,105,31,105,30,56,31,101,31,164,31,128,31,141,31,141,30,170,31,13,31,249,31,95,31,113,31,57,31,29,31,53,31,224,31,47,31,35,31,224,31,170,31,77,31,149,31,203,31,203,30,53,31,233,31,64,31,143,31,21,31,32,31,32,30,70,31,72,31,203,31,113,31,113,30,140,31,142,31,142,30,142,29,96,31,217,31,217,30,217,29,75,31,105,31,199,31,51,31,83,31,83,30,126,31,202,31,182,31,80,31,79,31,95,31,118,31,131,31,239,31,42,31,44,31,44,30,236,31,170,31,199,31,152,31,237,31,237,30,191,31,111,31,83,31,14,31,222,31,35,31,60,31,113,31,89,31,21,31,50,31,50,30,157,31,184,31,225,31,225,30,233,31,217,31,107,31,53,31,255,31,96,31,39,31,39,30,143,31,19,31,44,31,10,31,228,31,228,30,228,29,3,31,36,31,36,30,36,29,34,31,138,31,95,31,74,31,243,31,243,30,243,29,149,31,59,31,97,31,28,31,28,30,30,31,30,30,30,29,255,31,255,30,30,31,30,30,120,31,121,31,209,31,60,31,228,31,193,31,87,31,41,31,46,31,190,31,34,31,34,30,172,31,160,31,160,30,212,31,196,31,164,31,25,31,52,31,158,31,37,31,247,31,170,31,170,30,163,31,144,31,144,30,169,31,234,31,162,31,231,31,169,31,209,31,61,31,174,31,209,31,53,31,192,31,192,30,108,31,108,30,108,29,252,31,252,30,252,29,113,31,32,31,207,31,79,31,231,31,231,30,231,29,180,31,60,31,68,31,68,31,253,31,20,31,112,31,3,31,3,30,12,31,12,30,129,31,214,31,2,31,93,31,65,31,75,31,75,30,75,29,157,31,167,31,91,31,91,30,202,31,7,31,7,30,7,29,83,31,83,30,142,31,214,31,214,30,11,31,11,30,11,29,254,31,51,31,51,30,20,31,232,31,48,31,48,30,57,31,57,30,217,31,27,31,143,31,22,31,229,31,70,31,109,31,138,31,60,31,205,31,183,31,233,31,191,31,210,31,210,30,210,29,141,31,129,31,231,31,24,31,10,31,117,31,128,31,128,30,31,31,8,31,192,31,189,31,87,31,140,31,143,31,20,31,136,31,210,31,210,30,153,31,34,31,1,31,226,31,74,31,35,31,197,31,6,31,47,31,47,30,100,31,174,31,23,31,76,31,52,31,103,31,61,31,123,31,230,31,42,31,95,31,95,30,130,31,130,30,19,31,111,31,111,30,133,31,133,30,69,31,101,31,34,31,173,31,173,30,209,31,243,31,205,31,165,31,8,31,8,30,8,29,100,31,92,31,33,31,172,31,172,30,172,29,125,31,46,31,137,31,137,30,111,31,198,31,198,30,203,31,206,31,206,30,60,31,224,31,253,31,245,31,196,31,196,30,196,29,250,31,226,31,34,31,235,31,230,31,230,30,230,29,118,31,83,31,51,31,243,31,57,31,57,30,43,31,30,31,183,31,183,30,35,31,69,31,157,31,146,31,164,31,163,31,198,31,138,31,116,31,208,31,124,31,48,31,129,31,187,31,234,31,234,30,234,29,74,31,215,31,228,31,241,31,241,30,197,31,254,31,254,30,176,31,176,30,251,31,173,31,191,31,191,30,191,29,191,28,184,31,184,30,184,29,88,31,53,31,33,31,234,31,33,31,83,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
