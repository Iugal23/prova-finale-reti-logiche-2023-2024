-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 986;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (187,0,167,0,234,0,0,0,0,0,0,0,55,0,0,0,148,0,117,0,248,0,67,0,169,0,0,0,0,0,19,0,66,0,0,0,0,0,55,0,211,0,225,0,235,0,110,0,219,0,0,0,123,0,5,0,172,0,170,0,143,0,189,0,34,0,100,0,58,0,24,0,170,0,5,0,0,0,59,0,0,0,183,0,177,0,122,0,0,0,172,0,0,0,0,0,51,0,0,0,149,0,187,0,21,0,172,0,10,0,231,0,45,0,237,0,192,0,188,0,196,0,113,0,157,0,187,0,140,0,0,0,184,0,214,0,108,0,0,0,57,0,186,0,167,0,97,0,40,0,0,0,13,0,30,0,96,0,71,0,224,0,148,0,149,0,47,0,122,0,179,0,55,0,175,0,137,0,0,0,99,0,94,0,235,0,94,0,0,0,73,0,49,0,247,0,0,0,137,0,133,0,0,0,156,0,0,0,227,0,193,0,0,0,119,0,248,0,10,0,214,0,213,0,134,0,135,0,154,0,0,0,23,0,226,0,80,0,0,0,44,0,38,0,166,0,49,0,188,0,47,0,160,0,0,0,17,0,185,0,52,0,147,0,117,0,133,0,166,0,124,0,113,0,216,0,33,0,203,0,58,0,217,0,0,0,233,0,252,0,40,0,192,0,168,0,0,0,114,0,0,0,0,0,48,0,0,0,0,0,82,0,0,0,149,0,83,0,167,0,212,0,160,0,155,0,0,0,36,0,201,0,53,0,0,0,152,0,37,0,169,0,93,0,241,0,253,0,101,0,162,0,162,0,65,0,84,0,0,0,0,0,54,0,145,0,234,0,136,0,152,0,35,0,45,0,171,0,40,0,0,0,216,0,0,0,206,0,164,0,83,0,200,0,0,0,0,0,0,0,44,0,80,0,194,0,170,0,220,0,118,0,248,0,92,0,245,0,47,0,141,0,72,0,0,0,224,0,111,0,0,0,0,0,70,0,0,0,189,0,110,0,224,0,162,0,244,0,91,0,154,0,0,0,185,0,18,0,10,0,0,0,15,0,213,0,31,0,0,0,183,0,0,0,138,0,36,0,216,0,29,0,150,0,0,0,132,0,78,0,0,0,211,0,141,0,53,0,0,0,201,0,0,0,170,0,16,0,162,0,0,0,127,0,0,0,109,0,165,0,247,0,37,0,0,0,162,0,0,0,91,0,0,0,0,0,181,0,73,0,63,0,225,0,207,0,166,0,241,0,201,0,110,0,254,0,110,0,186,0,111,0,0,0,199,0,4,0,104,0,186,0,109,0,83,0,0,0,159,0,228,0,0,0,187,0,154,0,253,0,172,0,0,0,144,0,131,0,251,0,55,0,123,0,196,0,71,0,0,0,85,0,207,0,60,0,253,0,236,0,41,0,0,0,117,0,149,0,162,0,149,0,108,0,131,0,49,0,30,0,0,0,235,0,72,0,0,0,248,0,20,0,25,0,80,0,82,0,0,0,157,0,186,0,49,0,71,0,0,0,33,0,118,0,145,0,127,0,211,0,219,0,0,0,37,0,251,0,14,0,137,0,223,0,0,0,96,0,0,0,155,0,219,0,0,0,96,0,0,0,206,0,44,0,62,0,100,0,68,0,180,0,0,0,91,0,182,0,53,0,14,0,227,0,143,0,208,0,139,0,192,0,184,0,202,0,5,0,253,0,171,0,197,0,186,0,209,0,9,0,163,0,29,0,31,0,100,0,9,0,215,0,44,0,57,0,0,0,85,0,14,0,0,0,83,0,0,0,139,0,156,0,80,0,0,0,0,0,190,0,46,0,210,0,216,0,36,0,0,0,172,0,0,0,0,0,76,0,238,0,134,0,161,0,130,0,0,0,222,0,176,0,0,0,199,0,67,0,0,0,0,0,164,0,80,0,27,0,170,0,191,0,80,0,13,0,143,0,13,0,19,0,7,0,247,0,36,0,123,0,125,0,32,0,79,0,0,0,107,0,0,0,140,0,57,0,0,0,232,0,17,0,153,0,34,0,218,0,162,0,94,0,140,0,195,0,242,0,95,0,51,0,142,0,20,0,35,0,0,0,58,0,253,0,139,0,143,0,247,0,0,0,26,0,35,0,103,0,86,0,0,0,0,0,23,0,7,0,159,0,177,0,113,0,166,0,0,0,0,0,10,0,20,0,200,0,117,0,157,0,0,0,143,0,91,0,0,0,31,0,130,0,222,0,18,0,44,0,6,0,0,0,159,0,0,0,42,0,0,0,224,0,0,0,0,0,20,0,182,0,101,0,0,0,84,0,52,0,130,0,200,0,0,0,66,0,91,0,14,0,92,0,31,0,129,0,171,0,79,0,0,0,216,0,0,0,170,0,78,0,241,0,0,0,49,0,0,0,0,0,167,0,100,0,148,0,0,0,198,0,0,0,133,0,254,0,140,0,93,0,116,0,107,0,94,0,21,0,117,0,0,0,73,0,157,0,0,0,40,0,206,0,19,0,35,0,0,0,211,0,187,0,65,0,138,0,66,0,65,0,0,0,40,0,240,0,196,0,233,0,44,0,126,0,0,0,0,0,0,0,211,0,99,0,186,0,39,0,27,0,0,0,0,0,111,0,0,0,241,0,118,0,37,0,175,0,43,0,247,0,89,0,147,0,19,0,198,0,0,0,0,0,208,0,134,0,0,0,63,0,62,0,135,0,0,0,45,0,192,0,0,0,0,0,175,0,0,0,17,0,245,0,230,0,37,0,0,0,68,0,162,0,0,0,0,0,18,0,151,0,232,0,0,0,0,0,0,0,173,0,174,0,197,0,16,0,177,0,207,0,21,0,0,0,191,0,0,0,4,0,238,0,77,0,194,0,0,0,127,0,7,0,215,0,81,0,201,0,196,0,90,0,105,0,58,0,165,0,0,0,0,0,115,0,223,0,139,0,163,0,43,0,128,0,65,0,44,0,94,0,85,0,170,0,159,0,0,0,57,0,27,0,119,0,0,0,93,0,58,0,0,0,0,0,205,0,250,0,155,0,177,0,115,0,28,0,122,0,192,0,200,0,218,0,255,0,224,0,56,0,220,0,0,0,118,0,246,0,237,0,108,0,0,0,135,0,181,0,226,0,0,0,0,0,0,0,185,0,0,0,74,0,0,0,33,0,135,0,168,0,0,0,134,0,210,0,166,0,52,0,234,0,32,0,0,0,246,0,202,0,193,0,175,0,136,0,0,0,0,0,88,0,0,0,4,0,50,0,0,0,115,0,30,0,218,0,179,0,0,0,176,0,174,0,99,0,191,0,153,0,118,0,233,0,146,0,9,0,6,0,91,0,12,0,47,0,0,0,114,0,115,0,232,0,163,0,133,0,0,0,0,0,179,0,0,0,37,0,173,0,113,0,143,0,199,0,169,0,237,0,74,0,167,0,12,0,238,0,203,0,232,0,219,0,169,0,174,0,0,0,0,0,73,0,244,0,0,0,0,0,0,0,0,0,110,0,0,0,0,0,31,0,212,0,0,0,41,0,156,0,228,0,236,0,0,0,100,0,175,0,0,0,134,0,100,0,155,0,63,0,0,0,0,0,114,0,226,0,78,0,174,0,83,0,7,0,111,0,0,0,219,0,0,0,183,0,63,0,125,0,0,0,89,0,10,0,191,0,49,0,230,0,136,0,85,0,105,0,174,0,0,0,0,0,90,0,0,0,11,0,205,0,0,0,123,0,200,0,186,0,63,0,12,0,125,0,0,0,0,0,94,0,0,0,223,0,0,0,131,0,12,0,20,0,126,0,41,0,106,0,80,0,60,0,73,0,48,0,202,0,104,0,212,0,5,0,0,0,107,0,129,0,161,0,0,0,218,0,102,0,224,0,198,0,134,0,19,0,251,0,146,0,34,0,160,0,77,0,32,0,204,0,123,0,0,0,0,0,0,0,155,0,118,0,109,0,49,0,203,0,247,0,98,0,26,0,0,0,7,0,254,0,210,0,154,0,0,0,2,0,10,0,182,0,26,0,202,0,195,0,0,0,165,0,169,0,101,0,96,0,40,0,124,0,0,0,193,0,36,0,75,0,0,0,0,0,119,0,134,0,0,0,217,0,204,0,43,0,162,0,115,0,90,0,18,0,97,0,93,0,59,0,149,0,234,0,120,0,72,0,0,0,0,0,73,0,144,0,9,0,185,0,8,0,35,0,150,0,194,0,146,0,93,0,56,0,113,0,15,0,218,0,38,0,56,0,0,0,126,0,156,0,0,0,0,0,224,0,36,0,122,0,110,0,75,0,23,0,205,0,169,0,225,0,66,0,102,0,0,0,202,0,186,0,60,0,134,0,33,0,0,0,184,0,183,0,229,0,225,0,242,0,209,0,158,0,24,0,60,0,0,0,169,0,0,0,0,0,91,0,0,0,0,0,93,0,138,0,0,0,215,0,75,0,0,0,66,0,0,0,242,0);
signal scenario_full  : scenario_type := (187,31,167,31,234,31,234,30,234,29,234,28,55,31,55,30,148,31,117,31,248,31,67,31,169,31,169,30,169,29,19,31,66,31,66,30,66,29,55,31,211,31,225,31,235,31,110,31,219,31,219,30,123,31,5,31,172,31,170,31,143,31,189,31,34,31,100,31,58,31,24,31,170,31,5,31,5,30,59,31,59,30,183,31,177,31,122,31,122,30,172,31,172,30,172,29,51,31,51,30,149,31,187,31,21,31,172,31,10,31,231,31,45,31,237,31,192,31,188,31,196,31,113,31,157,31,187,31,140,31,140,30,184,31,214,31,108,31,108,30,57,31,186,31,167,31,97,31,40,31,40,30,13,31,30,31,96,31,71,31,224,31,148,31,149,31,47,31,122,31,179,31,55,31,175,31,137,31,137,30,99,31,94,31,235,31,94,31,94,30,73,31,49,31,247,31,247,30,137,31,133,31,133,30,156,31,156,30,227,31,193,31,193,30,119,31,248,31,10,31,214,31,213,31,134,31,135,31,154,31,154,30,23,31,226,31,80,31,80,30,44,31,38,31,166,31,49,31,188,31,47,31,160,31,160,30,17,31,185,31,52,31,147,31,117,31,133,31,166,31,124,31,113,31,216,31,33,31,203,31,58,31,217,31,217,30,233,31,252,31,40,31,192,31,168,31,168,30,114,31,114,30,114,29,48,31,48,30,48,29,82,31,82,30,149,31,83,31,167,31,212,31,160,31,155,31,155,30,36,31,201,31,53,31,53,30,152,31,37,31,169,31,93,31,241,31,253,31,101,31,162,31,162,31,65,31,84,31,84,30,84,29,54,31,145,31,234,31,136,31,152,31,35,31,45,31,171,31,40,31,40,30,216,31,216,30,206,31,164,31,83,31,200,31,200,30,200,29,200,28,44,31,80,31,194,31,170,31,220,31,118,31,248,31,92,31,245,31,47,31,141,31,72,31,72,30,224,31,111,31,111,30,111,29,70,31,70,30,189,31,110,31,224,31,162,31,244,31,91,31,154,31,154,30,185,31,18,31,10,31,10,30,15,31,213,31,31,31,31,30,183,31,183,30,138,31,36,31,216,31,29,31,150,31,150,30,132,31,78,31,78,30,211,31,141,31,53,31,53,30,201,31,201,30,170,31,16,31,162,31,162,30,127,31,127,30,109,31,165,31,247,31,37,31,37,30,162,31,162,30,91,31,91,30,91,29,181,31,73,31,63,31,225,31,207,31,166,31,241,31,201,31,110,31,254,31,110,31,186,31,111,31,111,30,199,31,4,31,104,31,186,31,109,31,83,31,83,30,159,31,228,31,228,30,187,31,154,31,253,31,172,31,172,30,144,31,131,31,251,31,55,31,123,31,196,31,71,31,71,30,85,31,207,31,60,31,253,31,236,31,41,31,41,30,117,31,149,31,162,31,149,31,108,31,131,31,49,31,30,31,30,30,235,31,72,31,72,30,248,31,20,31,25,31,80,31,82,31,82,30,157,31,186,31,49,31,71,31,71,30,33,31,118,31,145,31,127,31,211,31,219,31,219,30,37,31,251,31,14,31,137,31,223,31,223,30,96,31,96,30,155,31,219,31,219,30,96,31,96,30,206,31,44,31,62,31,100,31,68,31,180,31,180,30,91,31,182,31,53,31,14,31,227,31,143,31,208,31,139,31,192,31,184,31,202,31,5,31,253,31,171,31,197,31,186,31,209,31,9,31,163,31,29,31,31,31,100,31,9,31,215,31,44,31,57,31,57,30,85,31,14,31,14,30,83,31,83,30,139,31,156,31,80,31,80,30,80,29,190,31,46,31,210,31,216,31,36,31,36,30,172,31,172,30,172,29,76,31,238,31,134,31,161,31,130,31,130,30,222,31,176,31,176,30,199,31,67,31,67,30,67,29,164,31,80,31,27,31,170,31,191,31,80,31,13,31,143,31,13,31,19,31,7,31,247,31,36,31,123,31,125,31,32,31,79,31,79,30,107,31,107,30,140,31,57,31,57,30,232,31,17,31,153,31,34,31,218,31,162,31,94,31,140,31,195,31,242,31,95,31,51,31,142,31,20,31,35,31,35,30,58,31,253,31,139,31,143,31,247,31,247,30,26,31,35,31,103,31,86,31,86,30,86,29,23,31,7,31,159,31,177,31,113,31,166,31,166,30,166,29,10,31,20,31,200,31,117,31,157,31,157,30,143,31,91,31,91,30,31,31,130,31,222,31,18,31,44,31,6,31,6,30,159,31,159,30,42,31,42,30,224,31,224,30,224,29,20,31,182,31,101,31,101,30,84,31,52,31,130,31,200,31,200,30,66,31,91,31,14,31,92,31,31,31,129,31,171,31,79,31,79,30,216,31,216,30,170,31,78,31,241,31,241,30,49,31,49,30,49,29,167,31,100,31,148,31,148,30,198,31,198,30,133,31,254,31,140,31,93,31,116,31,107,31,94,31,21,31,117,31,117,30,73,31,157,31,157,30,40,31,206,31,19,31,35,31,35,30,211,31,187,31,65,31,138,31,66,31,65,31,65,30,40,31,240,31,196,31,233,31,44,31,126,31,126,30,126,29,126,28,211,31,99,31,186,31,39,31,27,31,27,30,27,29,111,31,111,30,241,31,118,31,37,31,175,31,43,31,247,31,89,31,147,31,19,31,198,31,198,30,198,29,208,31,134,31,134,30,63,31,62,31,135,31,135,30,45,31,192,31,192,30,192,29,175,31,175,30,17,31,245,31,230,31,37,31,37,30,68,31,162,31,162,30,162,29,18,31,151,31,232,31,232,30,232,29,232,28,173,31,174,31,197,31,16,31,177,31,207,31,21,31,21,30,191,31,191,30,4,31,238,31,77,31,194,31,194,30,127,31,7,31,215,31,81,31,201,31,196,31,90,31,105,31,58,31,165,31,165,30,165,29,115,31,223,31,139,31,163,31,43,31,128,31,65,31,44,31,94,31,85,31,170,31,159,31,159,30,57,31,27,31,119,31,119,30,93,31,58,31,58,30,58,29,205,31,250,31,155,31,177,31,115,31,28,31,122,31,192,31,200,31,218,31,255,31,224,31,56,31,220,31,220,30,118,31,246,31,237,31,108,31,108,30,135,31,181,31,226,31,226,30,226,29,226,28,185,31,185,30,74,31,74,30,33,31,135,31,168,31,168,30,134,31,210,31,166,31,52,31,234,31,32,31,32,30,246,31,202,31,193,31,175,31,136,31,136,30,136,29,88,31,88,30,4,31,50,31,50,30,115,31,30,31,218,31,179,31,179,30,176,31,174,31,99,31,191,31,153,31,118,31,233,31,146,31,9,31,6,31,91,31,12,31,47,31,47,30,114,31,115,31,232,31,163,31,133,31,133,30,133,29,179,31,179,30,37,31,173,31,113,31,143,31,199,31,169,31,237,31,74,31,167,31,12,31,238,31,203,31,232,31,219,31,169,31,174,31,174,30,174,29,73,31,244,31,244,30,244,29,244,28,244,27,110,31,110,30,110,29,31,31,212,31,212,30,41,31,156,31,228,31,236,31,236,30,100,31,175,31,175,30,134,31,100,31,155,31,63,31,63,30,63,29,114,31,226,31,78,31,174,31,83,31,7,31,111,31,111,30,219,31,219,30,183,31,63,31,125,31,125,30,89,31,10,31,191,31,49,31,230,31,136,31,85,31,105,31,174,31,174,30,174,29,90,31,90,30,11,31,205,31,205,30,123,31,200,31,186,31,63,31,12,31,125,31,125,30,125,29,94,31,94,30,223,31,223,30,131,31,12,31,20,31,126,31,41,31,106,31,80,31,60,31,73,31,48,31,202,31,104,31,212,31,5,31,5,30,107,31,129,31,161,31,161,30,218,31,102,31,224,31,198,31,134,31,19,31,251,31,146,31,34,31,160,31,77,31,32,31,204,31,123,31,123,30,123,29,123,28,155,31,118,31,109,31,49,31,203,31,247,31,98,31,26,31,26,30,7,31,254,31,210,31,154,31,154,30,2,31,10,31,182,31,26,31,202,31,195,31,195,30,165,31,169,31,101,31,96,31,40,31,124,31,124,30,193,31,36,31,75,31,75,30,75,29,119,31,134,31,134,30,217,31,204,31,43,31,162,31,115,31,90,31,18,31,97,31,93,31,59,31,149,31,234,31,120,31,72,31,72,30,72,29,73,31,144,31,9,31,185,31,8,31,35,31,150,31,194,31,146,31,93,31,56,31,113,31,15,31,218,31,38,31,56,31,56,30,126,31,156,31,156,30,156,29,224,31,36,31,122,31,110,31,75,31,23,31,205,31,169,31,225,31,66,31,102,31,102,30,202,31,186,31,60,31,134,31,33,31,33,30,184,31,183,31,229,31,225,31,242,31,209,31,158,31,24,31,60,31,60,30,169,31,169,30,169,29,91,31,91,30,91,29,93,31,138,31,138,30,215,31,75,31,75,30,66,31,66,30,242,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
