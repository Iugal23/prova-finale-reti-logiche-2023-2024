-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 635;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (228,0,51,0,149,0,167,0,49,0,102,0,0,0,252,0,0,0,68,0,161,0,105,0,247,0,0,0,216,0,248,0,231,0,30,0,0,0,19,0,0,0,240,0,0,0,227,0,240,0,0,0,78,0,224,0,29,0,56,0,10,0,231,0,0,0,77,0,72,0,149,0,216,0,49,0,20,0,185,0,140,0,47,0,86,0,67,0,0,0,0,0,171,0,131,0,141,0,0,0,7,0,0,0,239,0,170,0,61,0,124,0,11,0,0,0,145,0,136,0,230,0,39,0,124,0,0,0,36,0,234,0,211,0,113,0,0,0,147,0,254,0,87,0,111,0,59,0,0,0,143,0,95,0,10,0,57,0,100,0,40,0,75,0,128,0,133,0,0,0,36,0,15,0,19,0,165,0,151,0,222,0,62,0,0,0,144,0,0,0,0,0,0,0,112,0,95,0,0,0,0,0,173,0,0,0,38,0,250,0,16,0,17,0,233,0,198,0,73,0,178,0,219,0,58,0,251,0,243,0,142,0,178,0,0,0,219,0,21,0,255,0,220,0,75,0,0,0,250,0,209,0,0,0,178,0,171,0,215,0,79,0,0,0,0,0,4,0,181,0,204,0,33,0,0,0,95,0,160,0,251,0,38,0,0,0,233,0,2,0,41,0,112,0,0,0,42,0,221,0,0,0,95,0,0,0,107,0,218,0,0,0,152,0,77,0,98,0,142,0,140,0,19,0,84,0,0,0,167,0,248,0,0,0,79,0,0,0,110,0,2,0,0,0,0,0,253,0,130,0,0,0,44,0,0,0,94,0,219,0,95,0,0,0,127,0,106,0,83,0,104,0,62,0,205,0,244,0,35,0,0,0,111,0,100,0,152,0,190,0,84,0,80,0,199,0,200,0,18,0,94,0,153,0,31,0,233,0,0,0,0,0,0,0,221,0,100,0,223,0,9,0,0,0,104,0,55,0,162,0,208,0,40,0,186,0,84,0,144,0,221,0,70,0,0,0,122,0,0,0,51,0,142,0,230,0,0,0,92,0,0,0,13,0,198,0,116,0,0,0,0,0,0,0,183,0,77,0,48,0,149,0,25,0,33,0,106,0,67,0,253,0,0,0,175,0,0,0,98,0,246,0,250,0,244,0,170,0,161,0,103,0,102,0,214,0,163,0,182,0,0,0,134,0,20,0,160,0,212,0,0,0,0,0,159,0,0,0,0,0,222,0,217,0,0,0,114,0,0,0,100,0,0,0,0,0,238,0,239,0,232,0,165,0,0,0,0,0,0,0,245,0,111,0,211,0,6,0,84,0,62,0,159,0,183,0,129,0,13,0,142,0,232,0,49,0,0,0,16,0,44,0,240,0,204,0,214,0,0,0,42,0,133,0,223,0,166,0,236,0,117,0,28,0,9,0,0,0,0,0,0,0,0,0,208,0,130,0,207,0,160,0,190,0,42,0,176,0,161,0,239,0,28,0,0,0,106,0,141,0,161,0,40,0,0,0,242,0,119,0,101,0,166,0,126,0,204,0,3,0,182,0,155,0,60,0,154,0,110,0,0,0,0,0,0,0,160,0,78,0,251,0,0,0,141,0,0,0,84,0,200,0,0,0,243,0,184,0,8,0,4,0,164,0,17,0,242,0,53,0,0,0,16,0,138,0,120,0,80,0,245,0,0,0,197,0,53,0,172,0,155,0,126,0,161,0,150,0,246,0,43,0,52,0,124,0,0,0,154,0,104,0,48,0,214,0,0,0,0,0,64,0,0,0,106,0,249,0,100,0,247,0,199,0,26,0,0,0,126,0,136,0,210,0,59,0,0,0,97,0,15,0,160,0,196,0,0,0,42,0,110,0,0,0,165,0,21,0,195,0,0,0,175,0,188,0,243,0,1,0,138,0,29,0,195,0,0,0,144,0,79,0,127,0,39,0,190,0,132,0,52,0,0,0,33,0,96,0,22,0,246,0,1,0,139,0,128,0,113,0,75,0,95,0,0,0,220,0,0,0,0,0,177,0,0,0,100,0,184,0,0,0,0,0,36,0,21,0,42,0,106,0,5,0,35,0,99,0,0,0,77,0,237,0,171,0,76,0,85,0,0,0,0,0,42,0,0,0,0,0,36,0,0,0,133,0,166,0,0,0,76,0,30,0,153,0,230,0,131,0,39,0,0,0,190,0,67,0,102,0,71,0,0,0,225,0,244,0,0,0,17,0,0,0,0,0,103,0,0,0,172,0,151,0,75,0,0,0,235,0,235,0,0,0,22,0,253,0,0,0,85,0,226,0,0,0,70,0,217,0,1,0,174,0,242,0,0,0,0,0,0,0,2,0,0,0,0,0,124,0,176,0,255,0,204,0,99,0,0,0,135,0,126,0,123,0,230,0,224,0,154,0,141,0,73,0,131,0,239,0,0,0,32,0,93,0,251,0,72,0,101,0,80,0,0,0,100,0,177,0,0,0,36,0,57,0,232,0,0,0,254,0,130,0,0,0,28,0,34,0,114,0,197,0,213,0,223,0,142,0,205,0,0,0,54,0,195,0,50,0,117,0,88,0,0,0,139,0,0,0,0,0,47,0,0,0,109,0,0,0,0,0,0,0,113,0,52,0,159,0,41,0,0,0,0,0,33,0,0,0,37,0,62,0,142,0,0,0,0,0,231,0,144,0,96,0,213,0,247,0,179,0,127,0,89,0,0,0,16,0,0,0,241,0,89,0,193,0,68,0,154,0,56,0,44,0,82,0,109,0,125,0,147,0,233,0,0,0,169,0,0,0,78,0,119,0,207,0,0,0,129,0,18,0,145,0,243,0,131,0,218,0,144,0,0,0,155,0,0,0,115,0,0,0,128,0,0,0,76,0);
signal scenario_full  : scenario_type := (228,31,51,31,149,31,167,31,49,31,102,31,102,30,252,31,252,30,68,31,161,31,105,31,247,31,247,30,216,31,248,31,231,31,30,31,30,30,19,31,19,30,240,31,240,30,227,31,240,31,240,30,78,31,224,31,29,31,56,31,10,31,231,31,231,30,77,31,72,31,149,31,216,31,49,31,20,31,185,31,140,31,47,31,86,31,67,31,67,30,67,29,171,31,131,31,141,31,141,30,7,31,7,30,239,31,170,31,61,31,124,31,11,31,11,30,145,31,136,31,230,31,39,31,124,31,124,30,36,31,234,31,211,31,113,31,113,30,147,31,254,31,87,31,111,31,59,31,59,30,143,31,95,31,10,31,57,31,100,31,40,31,75,31,128,31,133,31,133,30,36,31,15,31,19,31,165,31,151,31,222,31,62,31,62,30,144,31,144,30,144,29,144,28,112,31,95,31,95,30,95,29,173,31,173,30,38,31,250,31,16,31,17,31,233,31,198,31,73,31,178,31,219,31,58,31,251,31,243,31,142,31,178,31,178,30,219,31,21,31,255,31,220,31,75,31,75,30,250,31,209,31,209,30,178,31,171,31,215,31,79,31,79,30,79,29,4,31,181,31,204,31,33,31,33,30,95,31,160,31,251,31,38,31,38,30,233,31,2,31,41,31,112,31,112,30,42,31,221,31,221,30,95,31,95,30,107,31,218,31,218,30,152,31,77,31,98,31,142,31,140,31,19,31,84,31,84,30,167,31,248,31,248,30,79,31,79,30,110,31,2,31,2,30,2,29,253,31,130,31,130,30,44,31,44,30,94,31,219,31,95,31,95,30,127,31,106,31,83,31,104,31,62,31,205,31,244,31,35,31,35,30,111,31,100,31,152,31,190,31,84,31,80,31,199,31,200,31,18,31,94,31,153,31,31,31,233,31,233,30,233,29,233,28,221,31,100,31,223,31,9,31,9,30,104,31,55,31,162,31,208,31,40,31,186,31,84,31,144,31,221,31,70,31,70,30,122,31,122,30,51,31,142,31,230,31,230,30,92,31,92,30,13,31,198,31,116,31,116,30,116,29,116,28,183,31,77,31,48,31,149,31,25,31,33,31,106,31,67,31,253,31,253,30,175,31,175,30,98,31,246,31,250,31,244,31,170,31,161,31,103,31,102,31,214,31,163,31,182,31,182,30,134,31,20,31,160,31,212,31,212,30,212,29,159,31,159,30,159,29,222,31,217,31,217,30,114,31,114,30,100,31,100,30,100,29,238,31,239,31,232,31,165,31,165,30,165,29,165,28,245,31,111,31,211,31,6,31,84,31,62,31,159,31,183,31,129,31,13,31,142,31,232,31,49,31,49,30,16,31,44,31,240,31,204,31,214,31,214,30,42,31,133,31,223,31,166,31,236,31,117,31,28,31,9,31,9,30,9,29,9,28,9,27,208,31,130,31,207,31,160,31,190,31,42,31,176,31,161,31,239,31,28,31,28,30,106,31,141,31,161,31,40,31,40,30,242,31,119,31,101,31,166,31,126,31,204,31,3,31,182,31,155,31,60,31,154,31,110,31,110,30,110,29,110,28,160,31,78,31,251,31,251,30,141,31,141,30,84,31,200,31,200,30,243,31,184,31,8,31,4,31,164,31,17,31,242,31,53,31,53,30,16,31,138,31,120,31,80,31,245,31,245,30,197,31,53,31,172,31,155,31,126,31,161,31,150,31,246,31,43,31,52,31,124,31,124,30,154,31,104,31,48,31,214,31,214,30,214,29,64,31,64,30,106,31,249,31,100,31,247,31,199,31,26,31,26,30,126,31,136,31,210,31,59,31,59,30,97,31,15,31,160,31,196,31,196,30,42,31,110,31,110,30,165,31,21,31,195,31,195,30,175,31,188,31,243,31,1,31,138,31,29,31,195,31,195,30,144,31,79,31,127,31,39,31,190,31,132,31,52,31,52,30,33,31,96,31,22,31,246,31,1,31,139,31,128,31,113,31,75,31,95,31,95,30,220,31,220,30,220,29,177,31,177,30,100,31,184,31,184,30,184,29,36,31,21,31,42,31,106,31,5,31,35,31,99,31,99,30,77,31,237,31,171,31,76,31,85,31,85,30,85,29,42,31,42,30,42,29,36,31,36,30,133,31,166,31,166,30,76,31,30,31,153,31,230,31,131,31,39,31,39,30,190,31,67,31,102,31,71,31,71,30,225,31,244,31,244,30,17,31,17,30,17,29,103,31,103,30,172,31,151,31,75,31,75,30,235,31,235,31,235,30,22,31,253,31,253,30,85,31,226,31,226,30,70,31,217,31,1,31,174,31,242,31,242,30,242,29,242,28,2,31,2,30,2,29,124,31,176,31,255,31,204,31,99,31,99,30,135,31,126,31,123,31,230,31,224,31,154,31,141,31,73,31,131,31,239,31,239,30,32,31,93,31,251,31,72,31,101,31,80,31,80,30,100,31,177,31,177,30,36,31,57,31,232,31,232,30,254,31,130,31,130,30,28,31,34,31,114,31,197,31,213,31,223,31,142,31,205,31,205,30,54,31,195,31,50,31,117,31,88,31,88,30,139,31,139,30,139,29,47,31,47,30,109,31,109,30,109,29,109,28,113,31,52,31,159,31,41,31,41,30,41,29,33,31,33,30,37,31,62,31,142,31,142,30,142,29,231,31,144,31,96,31,213,31,247,31,179,31,127,31,89,31,89,30,16,31,16,30,241,31,89,31,193,31,68,31,154,31,56,31,44,31,82,31,109,31,125,31,147,31,233,31,233,30,169,31,169,30,78,31,119,31,207,31,207,30,129,31,18,31,145,31,243,31,131,31,218,31,144,31,144,30,155,31,155,30,115,31,115,30,128,31,128,30,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
