-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_63 is
end project_tb_63;

architecture project_tb_arch_63 of project_tb_63 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 694;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,125,0,243,0,0,0,125,0,197,0,238,0,230,0,0,0,85,0,109,0,80,0,74,0,0,0,176,0,64,0,144,0,55,0,31,0,90,0,63,0,133,0,0,0,229,0,8,0,0,0,0,0,0,0,0,0,139,0,103,0,0,0,0,0,135,0,218,0,143,0,190,0,34,0,24,0,0,0,13,0,212,0,0,0,177,0,11,0,137,0,0,0,244,0,223,0,7,0,53,0,163,0,21,0,161,0,128,0,57,0,0,0,0,0,31,0,180,0,0,0,15,0,101,0,247,0,65,0,59,0,131,0,53,0,48,0,124,0,237,0,235,0,160,0,10,0,26,0,0,0,0,0,58,0,57,0,0,0,0,0,91,0,225,0,103,0,62,0,0,0,110,0,242,0,0,0,182,0,127,0,97,0,151,0,254,0,82,0,251,0,162,0,177,0,172,0,29,0,0,0,171,0,151,0,40,0,128,0,116,0,0,0,74,0,48,0,96,0,64,0,85,0,0,0,111,0,196,0,138,0,249,0,250,0,87,0,65,0,209,0,194,0,0,0,116,0,0,0,250,0,219,0,115,0,125,0,44,0,70,0,160,0,10,0,82,0,113,0,198,0,94,0,241,0,164,0,231,0,155,0,152,0,184,0,107,0,0,0,91,0,0,0,0,0,218,0,50,0,0,0,36,0,47,0,110,0,0,0,217,0,15,0,54,0,230,0,221,0,200,0,117,0,0,0,26,0,0,0,0,0,93,0,92,0,38,0,179,0,222,0,103,0,216,0,210,0,107,0,86,0,20,0,9,0,231,0,4,0,59,0,207,0,62,0,194,0,175,0,95,0,212,0,0,0,136,0,214,0,0,0,127,0,0,0,49,0,215,0,0,0,0,0,19,0,230,0,158,0,0,0,218,0,25,0,179,0,190,0,69,0,49,0,129,0,26,0,228,0,169,0,0,0,74,0,134,0,166,0,111,0,131,0,69,0,74,0,218,0,0,0,0,0,96,0,118,0,3,0,215,0,33,0,0,0,0,0,0,0,243,0,239,0,0,0,220,0,15,0,116,0,102,0,0,0,0,0,242,0,218,0,30,0,187,0,193,0,0,0,79,0,1,0,7,0,2,0,0,0,1,0,137,0,76,0,221,0,55,0,238,0,98,0,0,0,238,0,55,0,6,0,252,0,0,0,23,0,114,0,224,0,241,0,0,0,91,0,0,0,133,0,0,0,140,0,240,0,189,0,0,0,174,0,0,0,190,0,244,0,0,0,89,0,169,0,0,0,0,0,127,0,180,0,165,0,189,0,211,0,80,0,32,0,248,0,19,0,0,0,179,0,32,0,120,0,0,0,177,0,32,0,11,0,98,0,136,0,50,0,0,0,0,0,215,0,0,0,173,0,99,0,254,0,52,0,208,0,0,0,75,0,76,0,60,0,190,0,172,0,92,0,104,0,120,0,76,0,76,0,166,0,226,0,149,0,177,0,136,0,124,0,60,0,210,0,82,0,236,0,191,0,0,0,250,0,139,0,60,0,0,0,154,0,236,0,84,0,0,0,64,0,181,0,94,0,163,0,227,0,105,0,151,0,71,0,142,0,104,0,212,0,0,0,0,0,218,0,37,0,32,0,191,0,230,0,0,0,233,0,249,0,122,0,54,0,2,0,0,0,34,0,82,0,63,0,23,0,215,0,0,0,56,0,0,0,100,0,0,0,247,0,148,0,0,0,0,0,164,0,147,0,53,0,88,0,177,0,151,0,194,0,21,0,163,0,140,0,211,0,244,0,0,0,0,0,220,0,0,0,0,0,75,0,0,0,116,0,50,0,103,0,59,0,0,0,22,0,19,0,253,0,13,0,197,0,42,0,0,0,0,0,172,0,37,0,127,0,235,0,216,0,233,0,223,0,113,0,0,0,43,0,187,0,207,0,159,0,90,0,0,0,94,0,176,0,162,0,190,0,0,0,178,0,49,0,0,0,77,0,198,0,111,0,216,0,20,0,59,0,83,0,2,0,0,0,149,0,0,0,244,0,144,0,0,0,0,0,0,0,44,0,24,0,200,0,68,0,248,0,80,0,72,0,204,0,105,0,206,0,173,0,0,0,118,0,130,0,54,0,34,0,55,0,251,0,0,0,113,0,127,0,15,0,0,0,200,0,0,0,129,0,75,0,0,0,239,0,0,0,15,0,0,0,207,0,240,0,189,0,185,0,254,0,16,0,131,0,0,0,194,0,157,0,15,0,188,0,4,0,173,0,111,0,122,0,118,0,0,0,51,0,195,0,0,0,145,0,2,0,204,0,0,0,32,0,120,0,227,0,19,0,0,0,0,0,189,0,148,0,105,0,27,0,151,0,94,0,126,0,50,0,97,0,98,0,191,0,0,0,217,0,19,0,92,0,158,0,73,0,0,0,135,0,0,0,115,0,0,0,0,0,111,0,0,0,233,0,248,0,132,0,228,0,186,0,0,0,0,0,88,0,58,0,9,0,199,0,18,0,0,0,72,0,13,0,239,0,238,0,222,0,0,0,232,0,122,0,190,0,163,0,0,0,236,0,123,0,185,0,229,0,0,0,131,0,131,0,191,0,0,0,242,0,0,0,138,0,249,0,252,0,230,0,48,0,120,0,240,0,61,0,37,0,169,0,233,0,0,0,90,0,91,0,97,0,57,0,160,0,95,0,254,0,30,0,36,0,248,0,0,0,173,0,38,0,50,0,229,0,170,0,86,0,52,0,0,0,159,0,134,0,30,0,149,0,160,0,164,0,108,0,86,0,110,0,143,0,0,0,0,0,229,0,250,0,111,0,11,0,32,0,207,0,36,0,208,0,236,0,83,0,52,0,0,0,167,0,216,0,66,0,89,0,176,0,202,0,50,0,238,0,0,0,159,0,201,0,0,0,234,0,88,0,145,0,94,0,26,0,130,0,110,0,161,0,68,0,114,0,208,0,133,0,255,0,25,0,0,0,86,0,103,0,195,0,0,0,105,0,0,0,0,0,107,0,108,0,196,0,248,0,0,0,0,0,219,0,205,0,253,0,20,0,0,0,0,0,84,0,19,0,196,0,15,0,114,0,91,0,85,0,0,0,41,0,183,0,0,0,68,0,41,0,208,0,30,0);
signal scenario_full  : scenario_type := (0,0,125,31,243,31,243,30,125,31,197,31,238,31,230,31,230,30,85,31,109,31,80,31,74,31,74,30,176,31,64,31,144,31,55,31,31,31,90,31,63,31,133,31,133,30,229,31,8,31,8,30,8,29,8,28,8,27,139,31,103,31,103,30,103,29,135,31,218,31,143,31,190,31,34,31,24,31,24,30,13,31,212,31,212,30,177,31,11,31,137,31,137,30,244,31,223,31,7,31,53,31,163,31,21,31,161,31,128,31,57,31,57,30,57,29,31,31,180,31,180,30,15,31,101,31,247,31,65,31,59,31,131,31,53,31,48,31,124,31,237,31,235,31,160,31,10,31,26,31,26,30,26,29,58,31,57,31,57,30,57,29,91,31,225,31,103,31,62,31,62,30,110,31,242,31,242,30,182,31,127,31,97,31,151,31,254,31,82,31,251,31,162,31,177,31,172,31,29,31,29,30,171,31,151,31,40,31,128,31,116,31,116,30,74,31,48,31,96,31,64,31,85,31,85,30,111,31,196,31,138,31,249,31,250,31,87,31,65,31,209,31,194,31,194,30,116,31,116,30,250,31,219,31,115,31,125,31,44,31,70,31,160,31,10,31,82,31,113,31,198,31,94,31,241,31,164,31,231,31,155,31,152,31,184,31,107,31,107,30,91,31,91,30,91,29,218,31,50,31,50,30,36,31,47,31,110,31,110,30,217,31,15,31,54,31,230,31,221,31,200,31,117,31,117,30,26,31,26,30,26,29,93,31,92,31,38,31,179,31,222,31,103,31,216,31,210,31,107,31,86,31,20,31,9,31,231,31,4,31,59,31,207,31,62,31,194,31,175,31,95,31,212,31,212,30,136,31,214,31,214,30,127,31,127,30,49,31,215,31,215,30,215,29,19,31,230,31,158,31,158,30,218,31,25,31,179,31,190,31,69,31,49,31,129,31,26,31,228,31,169,31,169,30,74,31,134,31,166,31,111,31,131,31,69,31,74,31,218,31,218,30,218,29,96,31,118,31,3,31,215,31,33,31,33,30,33,29,33,28,243,31,239,31,239,30,220,31,15,31,116,31,102,31,102,30,102,29,242,31,218,31,30,31,187,31,193,31,193,30,79,31,1,31,7,31,2,31,2,30,1,31,137,31,76,31,221,31,55,31,238,31,98,31,98,30,238,31,55,31,6,31,252,31,252,30,23,31,114,31,224,31,241,31,241,30,91,31,91,30,133,31,133,30,140,31,240,31,189,31,189,30,174,31,174,30,190,31,244,31,244,30,89,31,169,31,169,30,169,29,127,31,180,31,165,31,189,31,211,31,80,31,32,31,248,31,19,31,19,30,179,31,32,31,120,31,120,30,177,31,32,31,11,31,98,31,136,31,50,31,50,30,50,29,215,31,215,30,173,31,99,31,254,31,52,31,208,31,208,30,75,31,76,31,60,31,190,31,172,31,92,31,104,31,120,31,76,31,76,31,166,31,226,31,149,31,177,31,136,31,124,31,60,31,210,31,82,31,236,31,191,31,191,30,250,31,139,31,60,31,60,30,154,31,236,31,84,31,84,30,64,31,181,31,94,31,163,31,227,31,105,31,151,31,71,31,142,31,104,31,212,31,212,30,212,29,218,31,37,31,32,31,191,31,230,31,230,30,233,31,249,31,122,31,54,31,2,31,2,30,34,31,82,31,63,31,23,31,215,31,215,30,56,31,56,30,100,31,100,30,247,31,148,31,148,30,148,29,164,31,147,31,53,31,88,31,177,31,151,31,194,31,21,31,163,31,140,31,211,31,244,31,244,30,244,29,220,31,220,30,220,29,75,31,75,30,116,31,50,31,103,31,59,31,59,30,22,31,19,31,253,31,13,31,197,31,42,31,42,30,42,29,172,31,37,31,127,31,235,31,216,31,233,31,223,31,113,31,113,30,43,31,187,31,207,31,159,31,90,31,90,30,94,31,176,31,162,31,190,31,190,30,178,31,49,31,49,30,77,31,198,31,111,31,216,31,20,31,59,31,83,31,2,31,2,30,149,31,149,30,244,31,144,31,144,30,144,29,144,28,44,31,24,31,200,31,68,31,248,31,80,31,72,31,204,31,105,31,206,31,173,31,173,30,118,31,130,31,54,31,34,31,55,31,251,31,251,30,113,31,127,31,15,31,15,30,200,31,200,30,129,31,75,31,75,30,239,31,239,30,15,31,15,30,207,31,240,31,189,31,185,31,254,31,16,31,131,31,131,30,194,31,157,31,15,31,188,31,4,31,173,31,111,31,122,31,118,31,118,30,51,31,195,31,195,30,145,31,2,31,204,31,204,30,32,31,120,31,227,31,19,31,19,30,19,29,189,31,148,31,105,31,27,31,151,31,94,31,126,31,50,31,97,31,98,31,191,31,191,30,217,31,19,31,92,31,158,31,73,31,73,30,135,31,135,30,115,31,115,30,115,29,111,31,111,30,233,31,248,31,132,31,228,31,186,31,186,30,186,29,88,31,58,31,9,31,199,31,18,31,18,30,72,31,13,31,239,31,238,31,222,31,222,30,232,31,122,31,190,31,163,31,163,30,236,31,123,31,185,31,229,31,229,30,131,31,131,31,191,31,191,30,242,31,242,30,138,31,249,31,252,31,230,31,48,31,120,31,240,31,61,31,37,31,169,31,233,31,233,30,90,31,91,31,97,31,57,31,160,31,95,31,254,31,30,31,36,31,248,31,248,30,173,31,38,31,50,31,229,31,170,31,86,31,52,31,52,30,159,31,134,31,30,31,149,31,160,31,164,31,108,31,86,31,110,31,143,31,143,30,143,29,229,31,250,31,111,31,11,31,32,31,207,31,36,31,208,31,236,31,83,31,52,31,52,30,167,31,216,31,66,31,89,31,176,31,202,31,50,31,238,31,238,30,159,31,201,31,201,30,234,31,88,31,145,31,94,31,26,31,130,31,110,31,161,31,68,31,114,31,208,31,133,31,255,31,25,31,25,30,86,31,103,31,195,31,195,30,105,31,105,30,105,29,107,31,108,31,196,31,248,31,248,30,248,29,219,31,205,31,253,31,20,31,20,30,20,29,84,31,19,31,196,31,15,31,114,31,91,31,85,31,85,30,41,31,183,31,183,30,68,31,41,31,208,31,30,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
