-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1019;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (243,0,0,0,58,0,0,0,78,0,113,0,51,0,91,0,39,0,125,0,252,0,72,0,138,0,50,0,0,0,225,0,0,0,175,0,0,0,206,0,75,0,45,0,87,0,0,0,0,0,1,0,77,0,170,0,185,0,115,0,11,0,48,0,0,0,111,0,225,0,209,0,166,0,237,0,221,0,96,0,31,0,149,0,0,0,12,0,244,0,101,0,226,0,93,0,191,0,253,0,247,0,9,0,7,0,133,0,0,0,21,0,0,0,216,0,141,0,165,0,10,0,80,0,130,0,0,0,199,0,62,0,47,0,69,0,0,0,197,0,0,0,74,0,0,0,0,0,0,0,0,0,65,0,191,0,222,0,198,0,0,0,53,0,0,0,0,0,243,0,245,0,233,0,225,0,13,0,0,0,6,0,123,0,49,0,125,0,229,0,0,0,46,0,0,0,10,0,201,0,0,0,97,0,177,0,46,0,0,0,254,0,138,0,82,0,169,0,0,0,152,0,104,0,83,0,55,0,0,0,176,0,0,0,202,0,203,0,0,0,240,0,96,0,7,0,3,0,8,0,0,0,0,0,6,0,34,0,57,0,0,0,1,0,0,0,249,0,134,0,0,0,168,0,223,0,187,0,0,0,21,0,29,0,17,0,76,0,246,0,1,0,111,0,0,0,7,0,148,0,26,0,0,0,0,0,36,0,62,0,16,0,0,0,41,0,179,0,0,0,0,0,165,0,207,0,0,0,94,0,189,0,182,0,126,0,145,0,84,0,11,0,175,0,193,0,125,0,0,0,93,0,102,0,26,0,152,0,0,0,99,0,124,0,255,0,59,0,153,0,235,0,149,0,52,0,225,0,0,0,132,0,0,0,55,0,110,0,209,0,167,0,25,0,19,0,163,0,175,0,91,0,0,0,0,0,228,0,37,0,0,0,0,0,102,0,198,0,36,0,185,0,0,0,174,0,205,0,214,0,0,0,183,0,229,0,211,0,136,0,0,0,133,0,173,0,0,0,142,0,174,0,109,0,83,0,130,0,0,0,249,0,26,0,61,0,18,0,0,0,71,0,14,0,0,0,163,0,250,0,2,0,0,0,0,0,0,0,118,0,188,0,182,0,194,0,21,0,153,0,0,0,48,0,140,0,247,0,154,0,0,0,18,0,20,0,30,0,55,0,0,0,8,0,0,0,171,0,0,0,17,0,57,0,245,0,0,0,230,0,158,0,162,0,164,0,92,0,123,0,239,0,136,0,73,0,120,0,80,0,165,0,0,0,11,0,210,0,23,0,0,0,118,0,251,0,108,0,0,0,42,0,29,0,11,0,41,0,243,0,196,0,0,0,224,0,212,0,0,0,242,0,132,0,7,0,149,0,193,0,0,0,3,0,252,0,168,0,74,0,0,0,176,0,236,0,9,0,111,0,188,0,0,0,109,0,154,0,200,0,37,0,230,0,19,0,105,0,0,0,177,0,248,0,13,0,39,0,0,0,113,0,88,0,117,0,0,0,45,0,160,0,118,0,88,0,53,0,104,0,0,0,0,0,0,0,144,0,76,0,89,0,252,0,242,0,210,0,82,0,0,0,0,0,176,0,0,0,0,0,0,0,51,0,0,0,118,0,251,0,0,0,81,0,0,0,157,0,251,0,85,0,216,0,0,0,245,0,71,0,0,0,0,0,0,0,40,0,185,0,16,0,187,0,0,0,51,0,157,0,153,0,165,0,60,0,107,0,0,0,199,0,55,0,198,0,96,0,163,0,0,0,3,0,0,0,47,0,150,0,235,0,237,0,0,0,124,0,78,0,163,0,245,0,65,0,208,0,159,0,222,0,175,0,86,0,88,0,125,0,167,0,121,0,206,0,0,0,193,0,1,0,61,0,48,0,182,0,229,0,242,0,236,0,0,0,163,0,0,0,251,0,98,0,36,0,250,0,191,0,76,0,0,0,17,0,62,0,75,0,0,0,18,0,179,0,251,0,36,0,0,0,100,0,142,0,161,0,247,0,59,0,39,0,206,0,0,0,114,0,0,0,0,0,0,0,209,0,14,0,0,0,142,0,61,0,201,0,107,0,0,0,255,0,204,0,70,0,247,0,141,0,50,0,247,0,161,0,102,0,0,0,26,0,0,0,61,0,238,0,163,0,35,0,78,0,130,0,240,0,0,0,0,0,113,0,98,0,10,0,27,0,108,0,61,0,247,0,0,0,43,0,146,0,147,0,0,0,250,0,154,0,0,0,196,0,0,0,141,0,92,0,0,0,0,0,249,0,16,0,242,0,109,0,186,0,222,0,0,0,167,0,48,0,60,0,10,0,68,0,120,0,136,0,0,0,0,0,163,0,0,0,58,0,211,0,162,0,106,0,0,0,0,0,17,0,199,0,113,0,192,0,190,0,236,0,104,0,162,0,0,0,0,0,38,0,153,0,43,0,99,0,216,0,183,0,108,0,186,0,109,0,219,0,61,0,231,0,22,0,111,0,214,0,145,0,126,0,60,0,15,0,200,0,0,0,193,0,46,0,18,0,79,0,11,0,0,0,0,0,23,0,0,0,113,0,245,0,0,0,37,0,223,0,0,0,143,0,163,0,138,0,0,0,164,0,51,0,157,0,26,0,128,0,172,0,167,0,0,0,113,0,184,0,146,0,190,0,46,0,150,0,81,0,139,0,0,0,229,0,0,0,243,0,241,0,77,0,0,0,0,0,207,0,114,0,0,0,0,0,89,0,67,0,24,0,40,0,0,0,117,0,205,0,131,0,0,0,109,0,183,0,166,0,68,0,0,0,67,0,40,0,115,0,119,0,52,0,92,0,6,0,244,0,221,0,180,0,255,0,217,0,0,0,0,0,157,0,0,0,34,0,46,0,138,0,67,0,91,0,240,0,237,0,112,0,205,0,175,0,238,0,175,0,186,0,165,0,70,0,154,0,11,0,213,0,0,0,74,0,2,0,253,0,177,0,178,0,163,0,114,0,166,0,0,0,0,0,36,0,236,0,246,0,46,0,143,0,0,0,21,0,252,0,221,0,8,0,145,0,0,0,211,0,53,0,0,0,222,0,0,0,1,0,228,0,237,0,38,0,119,0,0,0,187,0,231,0,0,0,186,0,154,0,254,0,64,0,132,0,155,0,172,0,76,0,0,0,219,0,160,0,221,0,252,0,248,0,0,0,2,0,66,0,0,0,0,0,98,0,34,0,157,0,0,0,46,0,0,0,168,0,111,0,38,0,169,0,0,0,211,0,223,0,223,0,0,0,69,0,47,0,126,0,203,0,144,0,73,0,4,0,229,0,116,0,230,0,86,0,0,0,203,0,102,0,37,0,0,0,233,0,134,0,49,0,246,0,105,0,156,0,0,0,51,0,0,0,108,0,100,0,0,0,137,0,15,0,208,0,95,0,117,0,252,0,0,0,0,0,0,0,187,0,110,0,106,0,59,0,72,0,50,0,162,0,68,0,70,0,255,0,205,0,163,0,0,0,220,0,0,0,113,0,255,0,173,0,0,0,97,0,175,0,35,0,138,0,0,0,42,0,229,0,0,0,55,0,52,0,33,0,59,0,101,0,182,0,10,0,55,0,0,0,213,0,0,0,179,0,0,0,0,0,225,0,36,0,169,0,146,0,98,0,105,0,115,0,26,0,14,0,164,0,44,0,137,0,55,0,95,0,59,0,210,0,160,0,4,0,16,0,63,0,227,0,28,0,168,0,30,0,0,0,43,0,58,0,202,0,97,0,0,0,112,0,218,0,239,0,137,0,5,0,69,0,0,0,0,0,252,0,117,0,193,0,172,0,0,0,183,0,90,0,152,0,9,0,30,0,217,0,111,0,0,0,43,0,155,0,53,0,139,0,0,0,161,0,33,0,95,0,0,0,160,0,33,0,120,0,145,0,133,0,21,0,0,0,191,0,81,0,0,0,202,0,126,0,0,0,83,0,22,0,117,0,77,0,249,0,71,0,0,0,0,0,127,0,151,0,241,0,131,0,123,0,217,0,86,0,125,0,0,0,226,0,65,0,232,0,131,0,195,0,0,0,0,0,101,0,167,0,246,0,22,0,121,0,88,0,75,0,0,0,0,0,23,0,172,0,59,0,64,0,17,0,174,0,92,0,0,0,54,0,244,0,219,0,0,0,174,0,90,0,212,0,0,0,229,0,141,0,89,0,239,0,194,0,195,0,152,0,0,0,121,0,176,0,122,0,98,0,169,0,0,0,221,0,28,0,127,0,0,0,186,0,0,0,224,0,221,0,185,0,199,0,134,0,0,0,182,0,49,0,132,0,0,0,0,0,0,0,182,0,48,0,57,0,62,0,170,0,87,0,0,0,0,0,39,0,87,0,0,0,0,0,32,0,129,0,238,0,182,0,229,0,52,0,81,0,0,0,155,0,103,0,2,0,0,0,2,0,29,0,0,0,75,0,222,0,0,0,131,0,30,0,87,0,226,0,218,0,66,0,0,0,79,0,208,0,17,0,95,0,0,0,35,0,0,0,219,0,54,0,81,0,225,0,46,0,28,0,0,0,0,0,32,0,159,0,19,0,115,0,18,0,234,0,0,0,57,0,23,0,0,0,222,0);
signal scenario_full  : scenario_type := (243,31,243,30,58,31,58,30,78,31,113,31,51,31,91,31,39,31,125,31,252,31,72,31,138,31,50,31,50,30,225,31,225,30,175,31,175,30,206,31,75,31,45,31,87,31,87,30,87,29,1,31,77,31,170,31,185,31,115,31,11,31,48,31,48,30,111,31,225,31,209,31,166,31,237,31,221,31,96,31,31,31,149,31,149,30,12,31,244,31,101,31,226,31,93,31,191,31,253,31,247,31,9,31,7,31,133,31,133,30,21,31,21,30,216,31,141,31,165,31,10,31,80,31,130,31,130,30,199,31,62,31,47,31,69,31,69,30,197,31,197,30,74,31,74,30,74,29,74,28,74,27,65,31,191,31,222,31,198,31,198,30,53,31,53,30,53,29,243,31,245,31,233,31,225,31,13,31,13,30,6,31,123,31,49,31,125,31,229,31,229,30,46,31,46,30,10,31,201,31,201,30,97,31,177,31,46,31,46,30,254,31,138,31,82,31,169,31,169,30,152,31,104,31,83,31,55,31,55,30,176,31,176,30,202,31,203,31,203,30,240,31,96,31,7,31,3,31,8,31,8,30,8,29,6,31,34,31,57,31,57,30,1,31,1,30,249,31,134,31,134,30,168,31,223,31,187,31,187,30,21,31,29,31,17,31,76,31,246,31,1,31,111,31,111,30,7,31,148,31,26,31,26,30,26,29,36,31,62,31,16,31,16,30,41,31,179,31,179,30,179,29,165,31,207,31,207,30,94,31,189,31,182,31,126,31,145,31,84,31,11,31,175,31,193,31,125,31,125,30,93,31,102,31,26,31,152,31,152,30,99,31,124,31,255,31,59,31,153,31,235,31,149,31,52,31,225,31,225,30,132,31,132,30,55,31,110,31,209,31,167,31,25,31,19,31,163,31,175,31,91,31,91,30,91,29,228,31,37,31,37,30,37,29,102,31,198,31,36,31,185,31,185,30,174,31,205,31,214,31,214,30,183,31,229,31,211,31,136,31,136,30,133,31,173,31,173,30,142,31,174,31,109,31,83,31,130,31,130,30,249,31,26,31,61,31,18,31,18,30,71,31,14,31,14,30,163,31,250,31,2,31,2,30,2,29,2,28,118,31,188,31,182,31,194,31,21,31,153,31,153,30,48,31,140,31,247,31,154,31,154,30,18,31,20,31,30,31,55,31,55,30,8,31,8,30,171,31,171,30,17,31,57,31,245,31,245,30,230,31,158,31,162,31,164,31,92,31,123,31,239,31,136,31,73,31,120,31,80,31,165,31,165,30,11,31,210,31,23,31,23,30,118,31,251,31,108,31,108,30,42,31,29,31,11,31,41,31,243,31,196,31,196,30,224,31,212,31,212,30,242,31,132,31,7,31,149,31,193,31,193,30,3,31,252,31,168,31,74,31,74,30,176,31,236,31,9,31,111,31,188,31,188,30,109,31,154,31,200,31,37,31,230,31,19,31,105,31,105,30,177,31,248,31,13,31,39,31,39,30,113,31,88,31,117,31,117,30,45,31,160,31,118,31,88,31,53,31,104,31,104,30,104,29,104,28,144,31,76,31,89,31,252,31,242,31,210,31,82,31,82,30,82,29,176,31,176,30,176,29,176,28,51,31,51,30,118,31,251,31,251,30,81,31,81,30,157,31,251,31,85,31,216,31,216,30,245,31,71,31,71,30,71,29,71,28,40,31,185,31,16,31,187,31,187,30,51,31,157,31,153,31,165,31,60,31,107,31,107,30,199,31,55,31,198,31,96,31,163,31,163,30,3,31,3,30,47,31,150,31,235,31,237,31,237,30,124,31,78,31,163,31,245,31,65,31,208,31,159,31,222,31,175,31,86,31,88,31,125,31,167,31,121,31,206,31,206,30,193,31,1,31,61,31,48,31,182,31,229,31,242,31,236,31,236,30,163,31,163,30,251,31,98,31,36,31,250,31,191,31,76,31,76,30,17,31,62,31,75,31,75,30,18,31,179,31,251,31,36,31,36,30,100,31,142,31,161,31,247,31,59,31,39,31,206,31,206,30,114,31,114,30,114,29,114,28,209,31,14,31,14,30,142,31,61,31,201,31,107,31,107,30,255,31,204,31,70,31,247,31,141,31,50,31,247,31,161,31,102,31,102,30,26,31,26,30,61,31,238,31,163,31,35,31,78,31,130,31,240,31,240,30,240,29,113,31,98,31,10,31,27,31,108,31,61,31,247,31,247,30,43,31,146,31,147,31,147,30,250,31,154,31,154,30,196,31,196,30,141,31,92,31,92,30,92,29,249,31,16,31,242,31,109,31,186,31,222,31,222,30,167,31,48,31,60,31,10,31,68,31,120,31,136,31,136,30,136,29,163,31,163,30,58,31,211,31,162,31,106,31,106,30,106,29,17,31,199,31,113,31,192,31,190,31,236,31,104,31,162,31,162,30,162,29,38,31,153,31,43,31,99,31,216,31,183,31,108,31,186,31,109,31,219,31,61,31,231,31,22,31,111,31,214,31,145,31,126,31,60,31,15,31,200,31,200,30,193,31,46,31,18,31,79,31,11,31,11,30,11,29,23,31,23,30,113,31,245,31,245,30,37,31,223,31,223,30,143,31,163,31,138,31,138,30,164,31,51,31,157,31,26,31,128,31,172,31,167,31,167,30,113,31,184,31,146,31,190,31,46,31,150,31,81,31,139,31,139,30,229,31,229,30,243,31,241,31,77,31,77,30,77,29,207,31,114,31,114,30,114,29,89,31,67,31,24,31,40,31,40,30,117,31,205,31,131,31,131,30,109,31,183,31,166,31,68,31,68,30,67,31,40,31,115,31,119,31,52,31,92,31,6,31,244,31,221,31,180,31,255,31,217,31,217,30,217,29,157,31,157,30,34,31,46,31,138,31,67,31,91,31,240,31,237,31,112,31,205,31,175,31,238,31,175,31,186,31,165,31,70,31,154,31,11,31,213,31,213,30,74,31,2,31,253,31,177,31,178,31,163,31,114,31,166,31,166,30,166,29,36,31,236,31,246,31,46,31,143,31,143,30,21,31,252,31,221,31,8,31,145,31,145,30,211,31,53,31,53,30,222,31,222,30,1,31,228,31,237,31,38,31,119,31,119,30,187,31,231,31,231,30,186,31,154,31,254,31,64,31,132,31,155,31,172,31,76,31,76,30,219,31,160,31,221,31,252,31,248,31,248,30,2,31,66,31,66,30,66,29,98,31,34,31,157,31,157,30,46,31,46,30,168,31,111,31,38,31,169,31,169,30,211,31,223,31,223,31,223,30,69,31,47,31,126,31,203,31,144,31,73,31,4,31,229,31,116,31,230,31,86,31,86,30,203,31,102,31,37,31,37,30,233,31,134,31,49,31,246,31,105,31,156,31,156,30,51,31,51,30,108,31,100,31,100,30,137,31,15,31,208,31,95,31,117,31,252,31,252,30,252,29,252,28,187,31,110,31,106,31,59,31,72,31,50,31,162,31,68,31,70,31,255,31,205,31,163,31,163,30,220,31,220,30,113,31,255,31,173,31,173,30,97,31,175,31,35,31,138,31,138,30,42,31,229,31,229,30,55,31,52,31,33,31,59,31,101,31,182,31,10,31,55,31,55,30,213,31,213,30,179,31,179,30,179,29,225,31,36,31,169,31,146,31,98,31,105,31,115,31,26,31,14,31,164,31,44,31,137,31,55,31,95,31,59,31,210,31,160,31,4,31,16,31,63,31,227,31,28,31,168,31,30,31,30,30,43,31,58,31,202,31,97,31,97,30,112,31,218,31,239,31,137,31,5,31,69,31,69,30,69,29,252,31,117,31,193,31,172,31,172,30,183,31,90,31,152,31,9,31,30,31,217,31,111,31,111,30,43,31,155,31,53,31,139,31,139,30,161,31,33,31,95,31,95,30,160,31,33,31,120,31,145,31,133,31,21,31,21,30,191,31,81,31,81,30,202,31,126,31,126,30,83,31,22,31,117,31,77,31,249,31,71,31,71,30,71,29,127,31,151,31,241,31,131,31,123,31,217,31,86,31,125,31,125,30,226,31,65,31,232,31,131,31,195,31,195,30,195,29,101,31,167,31,246,31,22,31,121,31,88,31,75,31,75,30,75,29,23,31,172,31,59,31,64,31,17,31,174,31,92,31,92,30,54,31,244,31,219,31,219,30,174,31,90,31,212,31,212,30,229,31,141,31,89,31,239,31,194,31,195,31,152,31,152,30,121,31,176,31,122,31,98,31,169,31,169,30,221,31,28,31,127,31,127,30,186,31,186,30,224,31,221,31,185,31,199,31,134,31,134,30,182,31,49,31,132,31,132,30,132,29,132,28,182,31,48,31,57,31,62,31,170,31,87,31,87,30,87,29,39,31,87,31,87,30,87,29,32,31,129,31,238,31,182,31,229,31,52,31,81,31,81,30,155,31,103,31,2,31,2,30,2,31,29,31,29,30,75,31,222,31,222,30,131,31,30,31,87,31,226,31,218,31,66,31,66,30,79,31,208,31,17,31,95,31,95,30,35,31,35,30,219,31,54,31,81,31,225,31,46,31,28,31,28,30,28,29,32,31,159,31,19,31,115,31,18,31,234,31,234,30,57,31,23,31,23,30,222,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
