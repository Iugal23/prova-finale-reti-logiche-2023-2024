-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,6,0,67,0,42,0,119,0,170,0,227,0,132,0,175,0,0,0,126,0,88,0,0,0,169,0,0,0,73,0,252,0,108,0,255,0,57,0,111,0,51,0,67,0,162,0,94,0,10,0,137,0,167,0,66,0,0,0,241,0,174,0,0,0,91,0,47,0,0,0,197,0,138,0,15,0,0,0,62,0,164,0,221,0,0,0,18,0,168,0,226,0,40,0,181,0,86,0,40,0,249,0,235,0,24,0,0,0,234,0,37,0,154,0,0,0,69,0,104,0,55,0,54,0,242,0,40,0,50,0,150,0,151,0,219,0,117,0,136,0,0,0,212,0,0,0,19,0,101,0,168,0,16,0,27,0,155,0,77,0,116,0,220,0,232,0,51,0,0,0,0,0,136,0,146,0,143,0,190,0,219,0,29,0,193,0,58,0,19,0,0,0,91,0,175,0,82,0,40,0,74,0,139,0,36,0,129,0,33,0,182,0,213,0,90,0,107,0,0,0,183,0,29,0,136,0,179,0,240,0,0,0,23,0,0,0,75,0,0,0,38,0,162,0,20,0,0,0,23,0,213,0,0,0,0,0,176,0,97,0,176,0,163,0,238,0,168,0,79,0,31,0,136,0,174,0,0,0,0,0,0,0,5,0,127,0,160,0,0,0,219,0,112,0,0,0,125,0,224,0,223,0,129,0,218,0,98,0,54,0,149,0,0,0,78,0,38,0,0,0,98,0,147,0,117,0,172,0,239,0,60,0,130,0,0,0,15,0,3,0,0,0,240,0,226,0,191,0,57,0,76,0,227,0,213,0,0,0,42,0,106,0,170,0,0,0,115,0,188,0,152,0,10,0,204,0,0,0,6,0,0,0,66,0,199,0,0,0,7,0,0,0,0,0,0,0,241,0,216,0,0,0,47,0,251,0,201,0,144,0,254,0,145,0,0,0,32,0,0,0,19,0,139,0,0,0,158,0,0,0,6,0,132,0,250,0,0,0,4,0,233,0,97,0,242,0,29,0,233,0,21,0,0,0,112,0,122,0,28,0,99,0,0,0,249,0,198,0,152,0,134,0,46,0,205,0,0,0,72,0,68,0,0,0,130,0,125,0,178,0,58,0,108,0,147,0,155,0,220,0,170,0,0,0,0,0,119,0,222,0,71,0,211,0,0,0,143,0,123,0,172,0,78,0,150,0,0,0,46,0,5,0,17,0,118,0,136,0,0,0,203,0,105,0,0,0,62,0,153,0,29,0,1,0,0,0,0,0,2,0,241,0,176,0,73,0,98,0,155,0,148,0,166,0,107,0,150,0,175,0,250,0,159,0,112,0,176,0,173,0,44,0,0,0,103,0,189,0,0,0,0,0,247,0,232,0,0,0,0,0,251,0,75,0,88,0,115,0,35,0,226,0,76,0,144,0,210,0,0,0,118,0,36,0,0,0,217,0,0,0,223,0,28,0,118,0,114,0,122,0,208,0,10,0,218,0,109,0,66,0,27,0,0,0,85,0,0,0,167,0,0,0,223,0,0,0,60,0,235,0,170,0,185,0,139,0,105,0,0,0,80,0,0,0,64,0,66,0,47,0,190,0,125,0,119,0,0,0,65,0,172,0,51,0,82,0,136,0,0,0,59,0,13,0,0,0,75,0,17,0,0,0,0,0,242,0,231,0,0,0,0,0,132,0,104,0,194,0,26,0,240,0,188,0,222,0,188,0,31,0,185,0,249,0,0,0,192,0,178,0,84,0,0,0,88,0,134,0,71,0,178,0,191,0,18,0,184,0,0,0,198,0,0,0,8,0,211,0,43,0,6,0,126,0,165,0,45,0,1,0,206,0,0,0,43,0,14,0,65,0,83,0,140,0,0,0,22,0,155,0,234,0,205,0,33,0,40,0,26,0,209,0,0,0,74,0,80,0,0,0,234,0,161,0,0,0,155,0,144,0,20,0,136,0,0,0,57,0,57,0,238,0,195,0,214,0,99,0,139,0,167,0,169,0,214,0,0,0,173,0,247,0,156,0,96,0,244,0,105,0,151,0,0,0,47,0,218,0,143,0,247,0,93,0,24,0,0,0,29,0,228,0,168,0,0,0,0,0,243,0,0,0,172,0,78,0,53,0,75,0,0,0,62,0,0,0,224,0,176,0,73,0,57,0,90,0,103,0,241,0,55,0,113,0,0,0,188,0,0,0,36,0,244,0,98,0,56,0,122,0,3,0,0,0,244,0,250,0,140,0,39,0,173,0,0,0,0,0,205,0,0,0,0,0,229,0,0,0,0,0,98,0,11,0,215,0,0,0,0,0,9,0,90,0,0,0,77,0,120,0,5,0,183,0,0,0,92,0,0,0,4,0,148,0,23,0,191,0,44,0,185,0,225,0,102,0,202,0,0,0,117,0,243,0,69,0,60,0,91,0,0,0,29,0,197,0,0,0,33,0,211,0,96,0,178,0,106,0,195,0,117,0,0,0,141,0,157,0,238,0,0,0,181,0,0,0,0,0,19,0,22,0,0,0,47,0,119,0,0,0,0,0,0,0,51,0,116,0,47,0,139,0,78,0,134,0,0,0,83,0,118,0,40,0,2,0,170,0,0,0,74,0,102,0,222,0,184,0,81,0,19,0,0,0,255,0,216,0,162,0,0,0,0,0,36,0,239,0,78,0,251,0,81,0,83,0,127,0,29,0,232,0,225,0,130,0,128,0,68,0,173,0,0,0,254,0,0,0,63,0,19,0,198,0,0,0,104,0,243,0,147,0,158,0,0,0,76,0,15,0,94,0,98,0,197,0,93,0,8,0,64,0,128,0,98,0,0,0,109,0,196,0,142,0,104,0,10,0,184,0,30,0,130,0,91,0,128,0,52,0,94,0,36,0,137,0,218,0,0,0,47,0,0,0,18,0,132,0,0,0,0,0,36,0,0,0,28,0,213,0,136,0,235,0,0,0,250,0,165,0,0,0,248,0,0,0,113,0,0,0,235,0,42,0,251,0,236,0,65,0,0,0,6,0,51,0,53,0,0,0,249,0,189,0,102,0,43,0,185,0,0,0,181,0,246,0,45,0,252,0,33,0,125,0,36,0,34,0,212,0,114,0,190,0,91,0,229,0,15,0,30,0,0,0,65,0,19,0,157,0,191,0,217,0,0,0,242,0,43,0,159,0,167,0,14,0,0,0,106,0,0,0,251,0,85,0,220,0,92,0,214,0,1,0,210,0,0,0,63,0,62,0,244,0,65,0,180,0,124,0,160,0,169,0,74,0,219,0,1,0,156,0,85,0,148,0,113,0,169,0,212,0,252,0,109,0,0,0,138,0,125,0,194,0,155,0,8,0,29,0,27,0,185,0,253,0,0,0,226,0,138,0,47,0,122,0,47,0,186,0,6,0,141,0,0,0,40,0,165,0,188,0,103,0,224,0,81,0,63,0,168,0,83,0,140,0,224,0,0,0,33,0,239,0,102,0,0,0,9,0,46,0,83,0,225,0,148,0,137,0,165,0,0,0,0,0,213,0,0,0,241,0,17,0,0,0,220,0,0,0,70,0,0,0,25,0,119,0,0,0,117,0,43,0,179,0,0,0,53,0,194,0,0,0,163,0,116,0,13,0,0,0,252,0,71,0,0,0,36,0,205,0,223,0,235,0,149,0,220,0,3,0,69,0,175,0,0,0,49,0,232,0,213,0,0,0,14,0,228,0,28,0,164,0,167,0,35,0,8,0,13,0,0,0,0,0,169,0,1,0,250,0,34,0,0,0,0,0,0,0,251,0,235,0,241,0,0,0,49,0,151,0,114,0,0,0,98,0,131,0,0,0,99,0,89,0,127,0,113,0,1,0,0,0,36,0,0,0,94,0,237,0,157,0,0,0,151,0,135,0,73,0,0,0,213,0,148,0,140,0,7,0,173,0,41,0,188,0,188,0,255,0,0,0,65,0,127,0,172,0,61,0,157,0,0,0,0,0,99,0,72,0,100,0,15,0,193,0,0,0,140,0,225,0,248,0,227,0,80,0,0,0,195,0,106,0,0,0,246,0,91,0,62,0,58,0,0,0,144,0,14,0,0,0,106,0,83,0,80,0,212,0,223,0,76,0,21,0,25,0,197,0,74,0,0,0,247,0,97,0,91,0,118,0,173,0,238,0,153,0,36,0,91,0,103,0,0,0,99,0,131,0,142,0,97,0,60,0,0,0,10,0,11,0,67,0,67,0,240,0,106,0,14,0,151,0,160,0,18,0,219,0,251,0,82,0,0,0,0,0,130,0,228,0,0,0,94,0,173,0,107,0,102,0,0,0,0,0,235,0,68,0,0,0,246,0,0,0,109,0,0,0,46,0,197,0,202,0,0,0,120,0,155,0,238,0,0,0,219,0,30,0,0,0,169,0,0,0);
signal scenario_full  : scenario_type := (0,0,6,31,67,31,42,31,119,31,170,31,227,31,132,31,175,31,175,30,126,31,88,31,88,30,169,31,169,30,73,31,252,31,108,31,255,31,57,31,111,31,51,31,67,31,162,31,94,31,10,31,137,31,167,31,66,31,66,30,241,31,174,31,174,30,91,31,47,31,47,30,197,31,138,31,15,31,15,30,62,31,164,31,221,31,221,30,18,31,168,31,226,31,40,31,181,31,86,31,40,31,249,31,235,31,24,31,24,30,234,31,37,31,154,31,154,30,69,31,104,31,55,31,54,31,242,31,40,31,50,31,150,31,151,31,219,31,117,31,136,31,136,30,212,31,212,30,19,31,101,31,168,31,16,31,27,31,155,31,77,31,116,31,220,31,232,31,51,31,51,30,51,29,136,31,146,31,143,31,190,31,219,31,29,31,193,31,58,31,19,31,19,30,91,31,175,31,82,31,40,31,74,31,139,31,36,31,129,31,33,31,182,31,213,31,90,31,107,31,107,30,183,31,29,31,136,31,179,31,240,31,240,30,23,31,23,30,75,31,75,30,38,31,162,31,20,31,20,30,23,31,213,31,213,30,213,29,176,31,97,31,176,31,163,31,238,31,168,31,79,31,31,31,136,31,174,31,174,30,174,29,174,28,5,31,127,31,160,31,160,30,219,31,112,31,112,30,125,31,224,31,223,31,129,31,218,31,98,31,54,31,149,31,149,30,78,31,38,31,38,30,98,31,147,31,117,31,172,31,239,31,60,31,130,31,130,30,15,31,3,31,3,30,240,31,226,31,191,31,57,31,76,31,227,31,213,31,213,30,42,31,106,31,170,31,170,30,115,31,188,31,152,31,10,31,204,31,204,30,6,31,6,30,66,31,199,31,199,30,7,31,7,30,7,29,7,28,241,31,216,31,216,30,47,31,251,31,201,31,144,31,254,31,145,31,145,30,32,31,32,30,19,31,139,31,139,30,158,31,158,30,6,31,132,31,250,31,250,30,4,31,233,31,97,31,242,31,29,31,233,31,21,31,21,30,112,31,122,31,28,31,99,31,99,30,249,31,198,31,152,31,134,31,46,31,205,31,205,30,72,31,68,31,68,30,130,31,125,31,178,31,58,31,108,31,147,31,155,31,220,31,170,31,170,30,170,29,119,31,222,31,71,31,211,31,211,30,143,31,123,31,172,31,78,31,150,31,150,30,46,31,5,31,17,31,118,31,136,31,136,30,203,31,105,31,105,30,62,31,153,31,29,31,1,31,1,30,1,29,2,31,241,31,176,31,73,31,98,31,155,31,148,31,166,31,107,31,150,31,175,31,250,31,159,31,112,31,176,31,173,31,44,31,44,30,103,31,189,31,189,30,189,29,247,31,232,31,232,30,232,29,251,31,75,31,88,31,115,31,35,31,226,31,76,31,144,31,210,31,210,30,118,31,36,31,36,30,217,31,217,30,223,31,28,31,118,31,114,31,122,31,208,31,10,31,218,31,109,31,66,31,27,31,27,30,85,31,85,30,167,31,167,30,223,31,223,30,60,31,235,31,170,31,185,31,139,31,105,31,105,30,80,31,80,30,64,31,66,31,47,31,190,31,125,31,119,31,119,30,65,31,172,31,51,31,82,31,136,31,136,30,59,31,13,31,13,30,75,31,17,31,17,30,17,29,242,31,231,31,231,30,231,29,132,31,104,31,194,31,26,31,240,31,188,31,222,31,188,31,31,31,185,31,249,31,249,30,192,31,178,31,84,31,84,30,88,31,134,31,71,31,178,31,191,31,18,31,184,31,184,30,198,31,198,30,8,31,211,31,43,31,6,31,126,31,165,31,45,31,1,31,206,31,206,30,43,31,14,31,65,31,83,31,140,31,140,30,22,31,155,31,234,31,205,31,33,31,40,31,26,31,209,31,209,30,74,31,80,31,80,30,234,31,161,31,161,30,155,31,144,31,20,31,136,31,136,30,57,31,57,31,238,31,195,31,214,31,99,31,139,31,167,31,169,31,214,31,214,30,173,31,247,31,156,31,96,31,244,31,105,31,151,31,151,30,47,31,218,31,143,31,247,31,93,31,24,31,24,30,29,31,228,31,168,31,168,30,168,29,243,31,243,30,172,31,78,31,53,31,75,31,75,30,62,31,62,30,224,31,176,31,73,31,57,31,90,31,103,31,241,31,55,31,113,31,113,30,188,31,188,30,36,31,244,31,98,31,56,31,122,31,3,31,3,30,244,31,250,31,140,31,39,31,173,31,173,30,173,29,205,31,205,30,205,29,229,31,229,30,229,29,98,31,11,31,215,31,215,30,215,29,9,31,90,31,90,30,77,31,120,31,5,31,183,31,183,30,92,31,92,30,4,31,148,31,23,31,191,31,44,31,185,31,225,31,102,31,202,31,202,30,117,31,243,31,69,31,60,31,91,31,91,30,29,31,197,31,197,30,33,31,211,31,96,31,178,31,106,31,195,31,117,31,117,30,141,31,157,31,238,31,238,30,181,31,181,30,181,29,19,31,22,31,22,30,47,31,119,31,119,30,119,29,119,28,51,31,116,31,47,31,139,31,78,31,134,31,134,30,83,31,118,31,40,31,2,31,170,31,170,30,74,31,102,31,222,31,184,31,81,31,19,31,19,30,255,31,216,31,162,31,162,30,162,29,36,31,239,31,78,31,251,31,81,31,83,31,127,31,29,31,232,31,225,31,130,31,128,31,68,31,173,31,173,30,254,31,254,30,63,31,19,31,198,31,198,30,104,31,243,31,147,31,158,31,158,30,76,31,15,31,94,31,98,31,197,31,93,31,8,31,64,31,128,31,98,31,98,30,109,31,196,31,142,31,104,31,10,31,184,31,30,31,130,31,91,31,128,31,52,31,94,31,36,31,137,31,218,31,218,30,47,31,47,30,18,31,132,31,132,30,132,29,36,31,36,30,28,31,213,31,136,31,235,31,235,30,250,31,165,31,165,30,248,31,248,30,113,31,113,30,235,31,42,31,251,31,236,31,65,31,65,30,6,31,51,31,53,31,53,30,249,31,189,31,102,31,43,31,185,31,185,30,181,31,246,31,45,31,252,31,33,31,125,31,36,31,34,31,212,31,114,31,190,31,91,31,229,31,15,31,30,31,30,30,65,31,19,31,157,31,191,31,217,31,217,30,242,31,43,31,159,31,167,31,14,31,14,30,106,31,106,30,251,31,85,31,220,31,92,31,214,31,1,31,210,31,210,30,63,31,62,31,244,31,65,31,180,31,124,31,160,31,169,31,74,31,219,31,1,31,156,31,85,31,148,31,113,31,169,31,212,31,252,31,109,31,109,30,138,31,125,31,194,31,155,31,8,31,29,31,27,31,185,31,253,31,253,30,226,31,138,31,47,31,122,31,47,31,186,31,6,31,141,31,141,30,40,31,165,31,188,31,103,31,224,31,81,31,63,31,168,31,83,31,140,31,224,31,224,30,33,31,239,31,102,31,102,30,9,31,46,31,83,31,225,31,148,31,137,31,165,31,165,30,165,29,213,31,213,30,241,31,17,31,17,30,220,31,220,30,70,31,70,30,25,31,119,31,119,30,117,31,43,31,179,31,179,30,53,31,194,31,194,30,163,31,116,31,13,31,13,30,252,31,71,31,71,30,36,31,205,31,223,31,235,31,149,31,220,31,3,31,69,31,175,31,175,30,49,31,232,31,213,31,213,30,14,31,228,31,28,31,164,31,167,31,35,31,8,31,13,31,13,30,13,29,169,31,1,31,250,31,34,31,34,30,34,29,34,28,251,31,235,31,241,31,241,30,49,31,151,31,114,31,114,30,98,31,131,31,131,30,99,31,89,31,127,31,113,31,1,31,1,30,36,31,36,30,94,31,237,31,157,31,157,30,151,31,135,31,73,31,73,30,213,31,148,31,140,31,7,31,173,31,41,31,188,31,188,31,255,31,255,30,65,31,127,31,172,31,61,31,157,31,157,30,157,29,99,31,72,31,100,31,15,31,193,31,193,30,140,31,225,31,248,31,227,31,80,31,80,30,195,31,106,31,106,30,246,31,91,31,62,31,58,31,58,30,144,31,14,31,14,30,106,31,83,31,80,31,212,31,223,31,76,31,21,31,25,31,197,31,74,31,74,30,247,31,97,31,91,31,118,31,173,31,238,31,153,31,36,31,91,31,103,31,103,30,99,31,131,31,142,31,97,31,60,31,60,30,10,31,11,31,67,31,67,31,240,31,106,31,14,31,151,31,160,31,18,31,219,31,251,31,82,31,82,30,82,29,130,31,228,31,228,30,94,31,173,31,107,31,102,31,102,30,102,29,235,31,68,31,68,30,246,31,246,30,109,31,109,30,46,31,197,31,202,31,202,30,120,31,155,31,238,31,238,30,219,31,30,31,30,30,169,31,169,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
