-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 160;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,231,0,72,0,16,0,0,0,60,0,58,0,0,0,0,0,228,0,35,0,43,0,237,0,202,0,129,0,223,0,0,0,234,0,130,0,105,0,250,0,241,0,12,0,244,0,7,0,0,0,0,0,30,0,71,0,189,0,48,0,83,0,126,0,28,0,199,0,148,0,184,0,59,0,59,0,187,0,77,0,184,0,242,0,49,0,0,0,0,0,153,0,159,0,157,0,188,0,0,0,0,0,124,0,175,0,88,0,150,0,111,0,66,0,190,0,0,0,113,0,152,0,103,0,198,0,224,0,49,0,0,0,175,0,216,0,223,0,53,0,174,0,0,0,74,0,125,0,74,0,0,0,97,0,203,0,213,0,0,0,214,0,0,0,123,0,166,0,98,0,133,0,110,0,195,0,0,0,126,0,137,0,215,0,87,0,200,0,7,0,54,0,88,0,142,0,0,0,172,0,94,0,194,0,0,0,176,0,0,0,93,0,0,0,216,0,0,0,65,0,35,0,0,0,0,0,234,0,211,0,0,0,22,0,0,0,235,0,47,0,0,0,43,0,46,0,62,0,173,0,218,0,85,0,222,0,0,0,0,0,237,0,248,0,112,0,163,0,14,0,236,0,147,0,22,0,160,0,106,0,71,0,54,0,254,0,231,0,77,0,173,0,91,0,206,0,202,0,215,0,0,0,210,0,176,0,222,0,136,0,223,0,161,0,0,0,220,0);
signal scenario_full  : scenario_type := (0,0,231,31,72,31,16,31,16,30,60,31,58,31,58,30,58,29,228,31,35,31,43,31,237,31,202,31,129,31,223,31,223,30,234,31,130,31,105,31,250,31,241,31,12,31,244,31,7,31,7,30,7,29,30,31,71,31,189,31,48,31,83,31,126,31,28,31,199,31,148,31,184,31,59,31,59,31,187,31,77,31,184,31,242,31,49,31,49,30,49,29,153,31,159,31,157,31,188,31,188,30,188,29,124,31,175,31,88,31,150,31,111,31,66,31,190,31,190,30,113,31,152,31,103,31,198,31,224,31,49,31,49,30,175,31,216,31,223,31,53,31,174,31,174,30,74,31,125,31,74,31,74,30,97,31,203,31,213,31,213,30,214,31,214,30,123,31,166,31,98,31,133,31,110,31,195,31,195,30,126,31,137,31,215,31,87,31,200,31,7,31,54,31,88,31,142,31,142,30,172,31,94,31,194,31,194,30,176,31,176,30,93,31,93,30,216,31,216,30,65,31,35,31,35,30,35,29,234,31,211,31,211,30,22,31,22,30,235,31,47,31,47,30,43,31,46,31,62,31,173,31,218,31,85,31,222,31,222,30,222,29,237,31,248,31,112,31,163,31,14,31,236,31,147,31,22,31,160,31,106,31,71,31,54,31,254,31,231,31,77,31,173,31,91,31,206,31,202,31,215,31,215,30,210,31,176,31,222,31,136,31,223,31,161,31,161,30,220,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
