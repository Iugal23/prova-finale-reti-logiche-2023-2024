-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_147 is
end project_tb_147;

architecture project_tb_arch_147 of project_tb_147 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 573;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,165,0,56,0,64,0,95,0,226,0,237,0,44,0,173,0,0,0,220,0,128,0,126,0,0,0,255,0,152,0,215,0,0,0,203,0,76,0,153,0,139,0,59,0,161,0,246,0,35,0,0,0,0,0,192,0,0,0,148,0,246,0,0,0,137,0,21,0,144,0,0,0,47,0,86,0,0,0,184,0,116,0,8,0,228,0,180,0,198,0,154,0,0,0,16,0,0,0,118,0,240,0,64,0,0,0,212,0,194,0,164,0,82,0,0,0,204,0,236,0,138,0,231,0,0,0,83,0,135,0,86,0,76,0,6,0,83,0,203,0,202,0,37,0,200,0,137,0,0,0,52,0,209,0,177,0,0,0,0,0,29,0,140,0,117,0,69,0,0,0,0,0,7,0,86,0,0,0,35,0,146,0,0,0,177,0,140,0,151,0,249,0,41,0,237,0,0,0,127,0,21,0,106,0,0,0,175,0,99,0,4,0,186,0,74,0,205,0,77,0,125,0,0,0,0,0,0,0,4,0,149,0,61,0,55,0,99,0,0,0,68,0,175,0,29,0,39,0,148,0,37,0,140,0,170,0,19,0,45,0,102,0,91,0,67,0,215,0,55,0,115,0,152,0,4,0,176,0,163,0,162,0,214,0,139,0,0,0,156,0,4,0,188,0,62,0,0,0,223,0,42,0,34,0,192,0,155,0,216,0,68,0,111,0,112,0,164,0,120,0,9,0,32,0,118,0,0,0,0,0,50,0,0,0,218,0,0,0,106,0,69,0,167,0,144,0,16,0,38,0,75,0,242,0,130,0,242,0,223,0,245,0,141,0,62,0,153,0,0,0,0,0,106,0,65,0,168,0,223,0,198,0,102,0,50,0,161,0,51,0,124,0,51,0,240,0,189,0,0,0,240,0,0,0,65,0,113,0,0,0,229,0,175,0,129,0,0,0,97,0,172,0,31,0,199,0,226,0,179,0,91,0,111,0,0,0,102,0,0,0,10,0,163,0,239,0,0,0,54,0,0,0,167,0,127,0,212,0,204,0,188,0,0,0,199,0,11,0,0,0,0,0,161,0,0,0,0,0,160,0,119,0,237,0,18,0,242,0,26,0,253,0,12,0,0,0,49,0,106,0,127,0,0,0,148,0,162,0,0,0,124,0,203,0,55,0,0,0,66,0,222,0,0,0,0,0,143,0,48,0,171,0,0,0,117,0,28,0,241,0,209,0,228,0,68,0,154,0,19,0,195,0,248,0,137,0,254,0,209,0,170,0,0,0,22,0,202,0,153,0,170,0,25,0,105,0,0,0,238,0,152,0,0,0,0,0,0,0,65,0,185,0,166,0,193,0,79,0,177,0,235,0,0,0,243,0,57,0,155,0,249,0,63,0,0,0,65,0,234,0,19,0,232,0,130,0,107,0,1,0,11,0,132,0,148,0,159,0,35,0,228,0,57,0,79,0,114,0,215,0,108,0,126,0,202,0,75,0,200,0,221,0,236,0,151,0,0,0,175,0,193,0,163,0,209,0,126,0,154,0,0,0,58,0,17,0,59,0,99,0,97,0,71,0,234,0,32,0,13,0,39,0,111,0,33,0,185,0,70,0,0,0,170,0,45,0,0,0,14,0,202,0,229,0,0,0,239,0,24,0,156,0,78,0,184,0,192,0,0,0,226,0,131,0,201,0,73,0,0,0,198,0,131,0,242,0,0,0,0,0,36,0,194,0,231,0,209,0,188,0,43,0,231,0,0,0,242,0,84,0,51,0,0,0,112,0,252,0,72,0,219,0,166,0,71,0,88,0,247,0,97,0,36,0,28,0,13,0,101,0,1,0,0,0,0,0,73,0,24,0,41,0,231,0,0,0,230,0,50,0,148,0,37,0,82,0,0,0,231,0,148,0,205,0,0,0,26,0,161,0,0,0,206,0,202,0,0,0,0,0,13,0,191,0,216,0,0,0,0,0,24,0,249,0,162,0,0,0,184,0,0,0,87,0,0,0,44,0,54,0,0,0,107,0,0,0,63,0,49,0,11,0,78,0,112,0,122,0,211,0,87,0,180,0,138,0,0,0,54,0,58,0,113,0,62,0,226,0,0,0,185,0,30,0,134,0,161,0,0,0,145,0,191,0,172,0,108,0,155,0,97,0,175,0,186,0,0,0,176,0,115,0,98,0,163,0,0,0,0,0,241,0,0,0,65,0,0,0,61,0,63,0,0,0,170,0,101,0,154,0,20,0,50,0,66,0,73,0,242,0,206,0,231,0,82,0,249,0,0,0,144,0,212,0,27,0,0,0,0,0,123,0,87,0,123,0,172,0,31,0,158,0,0,0,65,0,118,0,36,0,0,0,134,0,45,0,0,0,243,0,65,0,18,0,0,0,0,0,124,0,65,0,0,0,0,0,3,0,165,0,114,0,0,0,0,0,37,0,198,0,0,0,18,0,239,0,0,0,0,0,58,0,0,0,0,0,89,0,10,0,0,0,0,0,62,0,251,0,42,0,38,0,87,0,129,0,0,0,43,0,69,0,42,0,113,0,116,0,0,0,20,0,179,0,10,0,146,0,9,0,98,0,121,0);
signal scenario_full  : scenario_type := (0,0,165,31,56,31,64,31,95,31,226,31,237,31,44,31,173,31,173,30,220,31,128,31,126,31,126,30,255,31,152,31,215,31,215,30,203,31,76,31,153,31,139,31,59,31,161,31,246,31,35,31,35,30,35,29,192,31,192,30,148,31,246,31,246,30,137,31,21,31,144,31,144,30,47,31,86,31,86,30,184,31,116,31,8,31,228,31,180,31,198,31,154,31,154,30,16,31,16,30,118,31,240,31,64,31,64,30,212,31,194,31,164,31,82,31,82,30,204,31,236,31,138,31,231,31,231,30,83,31,135,31,86,31,76,31,6,31,83,31,203,31,202,31,37,31,200,31,137,31,137,30,52,31,209,31,177,31,177,30,177,29,29,31,140,31,117,31,69,31,69,30,69,29,7,31,86,31,86,30,35,31,146,31,146,30,177,31,140,31,151,31,249,31,41,31,237,31,237,30,127,31,21,31,106,31,106,30,175,31,99,31,4,31,186,31,74,31,205,31,77,31,125,31,125,30,125,29,125,28,4,31,149,31,61,31,55,31,99,31,99,30,68,31,175,31,29,31,39,31,148,31,37,31,140,31,170,31,19,31,45,31,102,31,91,31,67,31,215,31,55,31,115,31,152,31,4,31,176,31,163,31,162,31,214,31,139,31,139,30,156,31,4,31,188,31,62,31,62,30,223,31,42,31,34,31,192,31,155,31,216,31,68,31,111,31,112,31,164,31,120,31,9,31,32,31,118,31,118,30,118,29,50,31,50,30,218,31,218,30,106,31,69,31,167,31,144,31,16,31,38,31,75,31,242,31,130,31,242,31,223,31,245,31,141,31,62,31,153,31,153,30,153,29,106,31,65,31,168,31,223,31,198,31,102,31,50,31,161,31,51,31,124,31,51,31,240,31,189,31,189,30,240,31,240,30,65,31,113,31,113,30,229,31,175,31,129,31,129,30,97,31,172,31,31,31,199,31,226,31,179,31,91,31,111,31,111,30,102,31,102,30,10,31,163,31,239,31,239,30,54,31,54,30,167,31,127,31,212,31,204,31,188,31,188,30,199,31,11,31,11,30,11,29,161,31,161,30,161,29,160,31,119,31,237,31,18,31,242,31,26,31,253,31,12,31,12,30,49,31,106,31,127,31,127,30,148,31,162,31,162,30,124,31,203,31,55,31,55,30,66,31,222,31,222,30,222,29,143,31,48,31,171,31,171,30,117,31,28,31,241,31,209,31,228,31,68,31,154,31,19,31,195,31,248,31,137,31,254,31,209,31,170,31,170,30,22,31,202,31,153,31,170,31,25,31,105,31,105,30,238,31,152,31,152,30,152,29,152,28,65,31,185,31,166,31,193,31,79,31,177,31,235,31,235,30,243,31,57,31,155,31,249,31,63,31,63,30,65,31,234,31,19,31,232,31,130,31,107,31,1,31,11,31,132,31,148,31,159,31,35,31,228,31,57,31,79,31,114,31,215,31,108,31,126,31,202,31,75,31,200,31,221,31,236,31,151,31,151,30,175,31,193,31,163,31,209,31,126,31,154,31,154,30,58,31,17,31,59,31,99,31,97,31,71,31,234,31,32,31,13,31,39,31,111,31,33,31,185,31,70,31,70,30,170,31,45,31,45,30,14,31,202,31,229,31,229,30,239,31,24,31,156,31,78,31,184,31,192,31,192,30,226,31,131,31,201,31,73,31,73,30,198,31,131,31,242,31,242,30,242,29,36,31,194,31,231,31,209,31,188,31,43,31,231,31,231,30,242,31,84,31,51,31,51,30,112,31,252,31,72,31,219,31,166,31,71,31,88,31,247,31,97,31,36,31,28,31,13,31,101,31,1,31,1,30,1,29,73,31,24,31,41,31,231,31,231,30,230,31,50,31,148,31,37,31,82,31,82,30,231,31,148,31,205,31,205,30,26,31,161,31,161,30,206,31,202,31,202,30,202,29,13,31,191,31,216,31,216,30,216,29,24,31,249,31,162,31,162,30,184,31,184,30,87,31,87,30,44,31,54,31,54,30,107,31,107,30,63,31,49,31,11,31,78,31,112,31,122,31,211,31,87,31,180,31,138,31,138,30,54,31,58,31,113,31,62,31,226,31,226,30,185,31,30,31,134,31,161,31,161,30,145,31,191,31,172,31,108,31,155,31,97,31,175,31,186,31,186,30,176,31,115,31,98,31,163,31,163,30,163,29,241,31,241,30,65,31,65,30,61,31,63,31,63,30,170,31,101,31,154,31,20,31,50,31,66,31,73,31,242,31,206,31,231,31,82,31,249,31,249,30,144,31,212,31,27,31,27,30,27,29,123,31,87,31,123,31,172,31,31,31,158,31,158,30,65,31,118,31,36,31,36,30,134,31,45,31,45,30,243,31,65,31,18,31,18,30,18,29,124,31,65,31,65,30,65,29,3,31,165,31,114,31,114,30,114,29,37,31,198,31,198,30,18,31,239,31,239,30,239,29,58,31,58,30,58,29,89,31,10,31,10,30,10,29,62,31,251,31,42,31,38,31,87,31,129,31,129,30,43,31,69,31,42,31,113,31,116,31,116,30,20,31,179,31,10,31,146,31,9,31,98,31,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
