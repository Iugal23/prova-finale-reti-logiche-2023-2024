-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_595 is
end project_tb_595;

architecture project_tb_arch_595 of project_tb_595 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 464;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (15,0,224,0,98,0,5,0,0,0,86,0,160,0,37,0,0,0,173,0,96,0,0,0,0,0,231,0,100,0,0,0,16,0,251,0,103,0,101,0,0,0,0,0,73,0,0,0,183,0,54,0,17,0,81,0,153,0,179,0,70,0,164,0,125,0,236,0,68,0,245,0,123,0,126,0,100,0,218,0,115,0,0,0,245,0,198,0,0,0,190,0,244,0,30,0,243,0,160,0,133,0,0,0,7,0,58,0,221,0,51,0,66,0,191,0,179,0,0,0,0,0,212,0,0,0,0,0,51,0,43,0,21,0,161,0,31,0,97,0,93,0,0,0,234,0,42,0,0,0,215,0,240,0,71,0,0,0,0,0,2,0,66,0,0,0,0,0,22,0,168,0,168,0,0,0,0,0,137,0,229,0,134,0,0,0,0,0,109,0,0,0,0,0,178,0,0,0,228,0,111,0,0,0,107,0,251,0,15,0,102,0,169,0,0,0,230,0,14,0,0,0,86,0,137,0,67,0,108,0,248,0,245,0,119,0,133,0,243,0,152,0,175,0,149,0,0,0,0,0,92,0,87,0,213,0,255,0,237,0,244,0,207,0,140,0,128,0,143,0,38,0,0,0,24,0,108,0,0,0,0,0,0,0,83,0,215,0,0,0,105,0,176,0,152,0,0,0,41,0,116,0,78,0,100,0,0,0,53,0,71,0,224,0,225,0,0,0,168,0,0,0,209,0,208,0,196,0,0,0,89,0,145,0,231,0,19,0,78,0,0,0,5,0,0,0,201,0,64,0,171,0,9,0,10,0,46,0,104,0,157,0,188,0,162,0,195,0,0,0,152,0,196,0,122,0,31,0,17,0,0,0,174,0,237,0,177,0,11,0,128,0,29,0,223,0,111,0,216,0,0,0,126,0,234,0,154,0,165,0,63,0,240,0,97,0,138,0,240,0,0,0,121,0,253,0,76,0,0,0,185,0,127,0,44,0,228,0,11,0,230,0,0,0,64,0,53,0,204,0,203,0,88,0,207,0,0,0,19,0,45,0,110,0,28,0,96,0,0,0,0,0,223,0,0,0,179,0,209,0,0,0,213,0,186,0,243,0,237,0,71,0,67,0,0,0,178,0,73,0,176,0,134,0,244,0,180,0,68,0,42,0,237,0,138,0,16,0,0,0,234,0,127,0,111,0,160,0,150,0,187,0,165,0,0,0,45,0,14,0,0,0,0,0,84,0,92,0,78,0,208,0,118,0,132,0,96,0,227,0,88,0,93,0,115,0,223,0,208,0,200,0,249,0,96,0,219,0,57,0,102,0,110,0,247,0,0,0,190,0,126,0,118,0,197,0,38,0,63,0,4,0,82,0,32,0,155,0,163,0,0,0,88,0,156,0,215,0,97,0,224,0,144,0,149,0,116,0,0,0,205,0,83,0,247,0,212,0,119,0,191,0,39,0,201,0,128,0,171,0,23,0,168,0,171,0,38,0,180,0,102,0,206,0,215,0,2,0,156,0,210,0,29,0,162,0,205,0,54,0,46,0,212,0,0,0,55,0,52,0,203,0,44,0,201,0,246,0,119,0,0,0,3,0,7,0,0,0,74,0,184,0,0,0,202,0,253,0,183,0,0,0,75,0,75,0,0,0,0,0,248,0,147,0,79,0,0,0,165,0,252,0,186,0,0,0,88,0,129,0,177,0,0,0,247,0,56,0,23,0,204,0,180,0,0,0,18,0,106,0,173,0,65,0,129,0,32,0,0,0,92,0,36,0,0,0,225,0,66,0,0,0,84,0,0,0,174,0,82,0,172,0,109,0,0,0,205,0,179,0,0,0,42,0,0,0,196,0,66,0,0,0,0,0,0,0,123,0,58,0,0,0,254,0,0,0,0,0,102,0,245,0,204,0,205,0,239,0,79,0,0,0,210,0,89,0,0,0,4,0,180,0,254,0,62,0,107,0,180,0,199,0,0,0,46,0,223,0,187,0,115,0,0,0,108,0,228,0,74,0,28,0,61,0,95,0,0,0,129,0,0,0,0,0,111,0,229,0,92,0,114,0,116,0,75,0,0,0,130,0,62,0,75,0,59,0,149,0);
signal scenario_full  : scenario_type := (15,31,224,31,98,31,5,31,5,30,86,31,160,31,37,31,37,30,173,31,96,31,96,30,96,29,231,31,100,31,100,30,16,31,251,31,103,31,101,31,101,30,101,29,73,31,73,30,183,31,54,31,17,31,81,31,153,31,179,31,70,31,164,31,125,31,236,31,68,31,245,31,123,31,126,31,100,31,218,31,115,31,115,30,245,31,198,31,198,30,190,31,244,31,30,31,243,31,160,31,133,31,133,30,7,31,58,31,221,31,51,31,66,31,191,31,179,31,179,30,179,29,212,31,212,30,212,29,51,31,43,31,21,31,161,31,31,31,97,31,93,31,93,30,234,31,42,31,42,30,215,31,240,31,71,31,71,30,71,29,2,31,66,31,66,30,66,29,22,31,168,31,168,31,168,30,168,29,137,31,229,31,134,31,134,30,134,29,109,31,109,30,109,29,178,31,178,30,228,31,111,31,111,30,107,31,251,31,15,31,102,31,169,31,169,30,230,31,14,31,14,30,86,31,137,31,67,31,108,31,248,31,245,31,119,31,133,31,243,31,152,31,175,31,149,31,149,30,149,29,92,31,87,31,213,31,255,31,237,31,244,31,207,31,140,31,128,31,143,31,38,31,38,30,24,31,108,31,108,30,108,29,108,28,83,31,215,31,215,30,105,31,176,31,152,31,152,30,41,31,116,31,78,31,100,31,100,30,53,31,71,31,224,31,225,31,225,30,168,31,168,30,209,31,208,31,196,31,196,30,89,31,145,31,231,31,19,31,78,31,78,30,5,31,5,30,201,31,64,31,171,31,9,31,10,31,46,31,104,31,157,31,188,31,162,31,195,31,195,30,152,31,196,31,122,31,31,31,17,31,17,30,174,31,237,31,177,31,11,31,128,31,29,31,223,31,111,31,216,31,216,30,126,31,234,31,154,31,165,31,63,31,240,31,97,31,138,31,240,31,240,30,121,31,253,31,76,31,76,30,185,31,127,31,44,31,228,31,11,31,230,31,230,30,64,31,53,31,204,31,203,31,88,31,207,31,207,30,19,31,45,31,110,31,28,31,96,31,96,30,96,29,223,31,223,30,179,31,209,31,209,30,213,31,186,31,243,31,237,31,71,31,67,31,67,30,178,31,73,31,176,31,134,31,244,31,180,31,68,31,42,31,237,31,138,31,16,31,16,30,234,31,127,31,111,31,160,31,150,31,187,31,165,31,165,30,45,31,14,31,14,30,14,29,84,31,92,31,78,31,208,31,118,31,132,31,96,31,227,31,88,31,93,31,115,31,223,31,208,31,200,31,249,31,96,31,219,31,57,31,102,31,110,31,247,31,247,30,190,31,126,31,118,31,197,31,38,31,63,31,4,31,82,31,32,31,155,31,163,31,163,30,88,31,156,31,215,31,97,31,224,31,144,31,149,31,116,31,116,30,205,31,83,31,247,31,212,31,119,31,191,31,39,31,201,31,128,31,171,31,23,31,168,31,171,31,38,31,180,31,102,31,206,31,215,31,2,31,156,31,210,31,29,31,162,31,205,31,54,31,46,31,212,31,212,30,55,31,52,31,203,31,44,31,201,31,246,31,119,31,119,30,3,31,7,31,7,30,74,31,184,31,184,30,202,31,253,31,183,31,183,30,75,31,75,31,75,30,75,29,248,31,147,31,79,31,79,30,165,31,252,31,186,31,186,30,88,31,129,31,177,31,177,30,247,31,56,31,23,31,204,31,180,31,180,30,18,31,106,31,173,31,65,31,129,31,32,31,32,30,92,31,36,31,36,30,225,31,66,31,66,30,84,31,84,30,174,31,82,31,172,31,109,31,109,30,205,31,179,31,179,30,42,31,42,30,196,31,66,31,66,30,66,29,66,28,123,31,58,31,58,30,254,31,254,30,254,29,102,31,245,31,204,31,205,31,239,31,79,31,79,30,210,31,89,31,89,30,4,31,180,31,254,31,62,31,107,31,180,31,199,31,199,30,46,31,223,31,187,31,115,31,115,30,108,31,228,31,74,31,28,31,61,31,95,31,95,30,129,31,129,30,129,29,111,31,229,31,92,31,114,31,116,31,75,31,75,30,130,31,62,31,75,31,59,31,149,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
