-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 742;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (193,0,122,0,81,0,90,0,166,0,176,0,16,0,194,0,0,0,0,0,0,0,239,0,143,0,163,0,135,0,83,0,0,0,80,0,80,0,0,0,47,0,203,0,31,0,0,0,0,0,71,0,93,0,0,0,72,0,4,0,0,0,0,0,45,0,0,0,0,0,127,0,27,0,52,0,127,0,254,0,106,0,28,0,86,0,84,0,194,0,0,0,57,0,143,0,0,0,244,0,120,0,243,0,200,0,253,0,53,0,217,0,0,0,99,0,21,0,173,0,0,0,215,0,158,0,147,0,233,0,214,0,180,0,245,0,87,0,105,0,0,0,58,0,231,0,75,0,218,0,33,0,96,0,10,0,132,0,0,0,54,0,172,0,203,0,0,0,189,0,7,0,252,0,51,0,0,0,165,0,94,0,166,0,74,0,201,0,106,0,0,0,0,0,218,0,164,0,174,0,182,0,0,0,171,0,196,0,72,0,155,0,237,0,0,0,145,0,27,0,0,0,0,0,217,0,238,0,109,0,247,0,243,0,77,0,214,0,122,0,90,0,114,0,156,0,227,0,0,0,0,0,249,0,193,0,248,0,85,0,86,0,9,0,245,0,247,0,0,0,81,0,0,0,142,0,125,0,107,0,198,0,117,0,252,0,241,0,69,0,0,0,38,0,178,0,38,0,207,0,63,0,163,0,114,0,180,0,0,0,108,0,171,0,0,0,17,0,120,0,254,0,15,0,79,0,0,0,14,0,250,0,61,0,72,0,130,0,0,0,31,0,0,0,0,0,25,0,0,0,144,0,254,0,120,0,48,0,53,0,115,0,126,0,80,0,216,0,19,0,211,0,0,0,34,0,58,0,15,0,239,0,230,0,2,0,90,0,0,0,0,0,87,0,148,0,14,0,53,0,0,0,117,0,144,0,0,0,156,0,15,0,0,0,133,0,0,0,0,0,73,0,0,0,0,0,156,0,0,0,179,0,0,0,157,0,0,0,99,0,189,0,121,0,126,0,0,0,74,0,114,0,179,0,115,0,0,0,0,0,2,0,133,0,66,0,204,0,165,0,248,0,91,0,0,0,248,0,252,0,216,0,0,0,93,0,242,0,130,0,202,0,179,0,70,0,188,0,0,0,194,0,181,0,200,0,0,0,220,0,5,0,47,0,191,0,189,0,239,0,0,0,92,0,0,0,0,0,92,0,240,0,126,0,0,0,251,0,0,0,0,0,102,0,95,0,1,0,250,0,51,0,192,0,89,0,22,0,233,0,0,0,62,0,109,0,0,0,0,0,101,0,219,0,196,0,88,0,161,0,100,0,42,0,14,0,137,0,115,0,118,0,241,0,171,0,249,0,41,0,0,0,0,0,156,0,155,0,0,0,114,0,38,0,207,0,198,0,198,0,0,0,15,0,29,0,202,0,0,0,222,0,0,0,0,0,177,0,131,0,254,0,22,0,200,0,253,0,0,0,32,0,31,0,91,0,160,0,0,0,92,0,146,0,232,0,0,0,7,0,0,0,31,0,19,0,0,0,231,0,191,0,0,0,82,0,126,0,211,0,226,0,16,0,237,0,113,0,46,0,0,0,248,0,171,0,0,0,221,0,187,0,220,0,59,0,0,0,212,0,0,0,87,0,75,0,58,0,144,0,189,0,150,0,29,0,220,0,145,0,244,0,123,0,13,0,0,0,199,0,228,0,27,0,0,0,87,0,221,0,152,0,143,0,115,0,19,0,75,0,164,0,193,0,4,0,96,0,0,0,79,0,147,0,34,0,229,0,73,0,130,0,0,0,240,0,0,0,255,0,110,0,19,0,253,0,254,0,250,0,156,0,177,0,253,0,0,0,0,0,235,0,116,0,0,0,100,0,5,0,25,0,0,0,176,0,195,0,26,0,103,0,245,0,103,0,252,0,0,0,206,0,242,0,63,0,134,0,0,0,0,0,209,0,125,0,207,0,208,0,0,0,220,0,99,0,28,0,128,0,111,0,206,0,191,0,29,0,10,0,0,0,35,0,127,0,196,0,252,0,203,0,146,0,132,0,168,0,236,0,222,0,48,0,181,0,57,0,37,0,155,0,0,0,144,0,0,0,43,0,214,0,227,0,206,0,45,0,70,0,239,0,61,0,0,0,35,0,0,0,100,0,0,0,142,0,202,0,218,0,0,0,62,0,0,0,29,0,48,0,0,0,205,0,234,0,244,0,173,0,137,0,57,0,132,0,54,0,238,0,0,0,51,0,228,0,99,0,121,0,73,0,137,0,35,0,124,0,219,0,42,0,48,0,150,0,192,0,168,0,0,0,205,0,208,0,98,0,0,0,116,0,198,0,63,0,188,0,39,0,36,0,0,0,0,0,80,0,0,0,44,0,0,0,187,0,217,0,40,0,0,0,65,0,123,0,48,0,51,0,45,0,0,0,108,0,178,0,237,0,35,0,0,0,201,0,0,0,7,0,145,0,108,0,112,0,7,0,0,0,114,0,152,0,88,0,83,0,0,0,31,0,13,0,0,0,0,0,0,0,238,0,27,0,0,0,170,0,80,0,217,0,32,0,0,0,145,0,148,0,204,0,0,0,187,0,113,0,225,0,131,0,0,0,0,0,143,0,0,0,230,0,166,0,0,0,213,0,0,0,0,0,42,0,72,0,27,0,0,0,91,0,0,0,0,0,217,0,125,0,0,0,156,0,232,0,27,0,224,0,235,0,132,0,193,0,234,0,234,0,79,0,39,0,87,0,245,0,51,0,0,0,123,0,199,0,198,0,0,0,218,0,189,0,177,0,0,0,152,0,19,0,183,0,164,0,96,0,238,0,250,0,68,0,0,0,101,0,188,0,0,0,0,0,14,0,110,0,172,0,178,0,252,0,0,0,215,0,186,0,101,0,111,0,61,0,0,0,106,0,183,0,104,0,0,0,113,0,6,0,250,0,63,0,0,0,212,0,195,0,0,0,62,0,158,0,153,0,0,0,45,0,63,0,101,0,0,0,0,0,240,0,19,0,119,0,0,0,195,0,189,0,0,0,191,0,151,0,173,0,151,0,89,0,95,0,36,0,46,0,221,0,73,0,155,0,0,0,143,0,81,0,40,0,61,0,218,0,203,0,0,0,233,0,53,0,0,0,0,0,45,0,137,0,228,0,4,0,86,0,101,0,88,0,232,0,34,0,242,0,204,0,0,0,0,0,144,0,0,0,76,0,201,0,0,0,181,0,216,0,230,0,141,0,0,0,113,0,33,0,70,0,0,0,47,0,0,0,243,0,140,0,127,0,191,0,20,0,3,0,194,0,121,0,93,0,40,0,0,0,146,0,232,0,19,0,229,0,18,0,83,0,139,0);
signal scenario_full  : scenario_type := (193,31,122,31,81,31,90,31,166,31,176,31,16,31,194,31,194,30,194,29,194,28,239,31,143,31,163,31,135,31,83,31,83,30,80,31,80,31,80,30,47,31,203,31,31,31,31,30,31,29,71,31,93,31,93,30,72,31,4,31,4,30,4,29,45,31,45,30,45,29,127,31,27,31,52,31,127,31,254,31,106,31,28,31,86,31,84,31,194,31,194,30,57,31,143,31,143,30,244,31,120,31,243,31,200,31,253,31,53,31,217,31,217,30,99,31,21,31,173,31,173,30,215,31,158,31,147,31,233,31,214,31,180,31,245,31,87,31,105,31,105,30,58,31,231,31,75,31,218,31,33,31,96,31,10,31,132,31,132,30,54,31,172,31,203,31,203,30,189,31,7,31,252,31,51,31,51,30,165,31,94,31,166,31,74,31,201,31,106,31,106,30,106,29,218,31,164,31,174,31,182,31,182,30,171,31,196,31,72,31,155,31,237,31,237,30,145,31,27,31,27,30,27,29,217,31,238,31,109,31,247,31,243,31,77,31,214,31,122,31,90,31,114,31,156,31,227,31,227,30,227,29,249,31,193,31,248,31,85,31,86,31,9,31,245,31,247,31,247,30,81,31,81,30,142,31,125,31,107,31,198,31,117,31,252,31,241,31,69,31,69,30,38,31,178,31,38,31,207,31,63,31,163,31,114,31,180,31,180,30,108,31,171,31,171,30,17,31,120,31,254,31,15,31,79,31,79,30,14,31,250,31,61,31,72,31,130,31,130,30,31,31,31,30,31,29,25,31,25,30,144,31,254,31,120,31,48,31,53,31,115,31,126,31,80,31,216,31,19,31,211,31,211,30,34,31,58,31,15,31,239,31,230,31,2,31,90,31,90,30,90,29,87,31,148,31,14,31,53,31,53,30,117,31,144,31,144,30,156,31,15,31,15,30,133,31,133,30,133,29,73,31,73,30,73,29,156,31,156,30,179,31,179,30,157,31,157,30,99,31,189,31,121,31,126,31,126,30,74,31,114,31,179,31,115,31,115,30,115,29,2,31,133,31,66,31,204,31,165,31,248,31,91,31,91,30,248,31,252,31,216,31,216,30,93,31,242,31,130,31,202,31,179,31,70,31,188,31,188,30,194,31,181,31,200,31,200,30,220,31,5,31,47,31,191,31,189,31,239,31,239,30,92,31,92,30,92,29,92,31,240,31,126,31,126,30,251,31,251,30,251,29,102,31,95,31,1,31,250,31,51,31,192,31,89,31,22,31,233,31,233,30,62,31,109,31,109,30,109,29,101,31,219,31,196,31,88,31,161,31,100,31,42,31,14,31,137,31,115,31,118,31,241,31,171,31,249,31,41,31,41,30,41,29,156,31,155,31,155,30,114,31,38,31,207,31,198,31,198,31,198,30,15,31,29,31,202,31,202,30,222,31,222,30,222,29,177,31,131,31,254,31,22,31,200,31,253,31,253,30,32,31,31,31,91,31,160,31,160,30,92,31,146,31,232,31,232,30,7,31,7,30,31,31,19,31,19,30,231,31,191,31,191,30,82,31,126,31,211,31,226,31,16,31,237,31,113,31,46,31,46,30,248,31,171,31,171,30,221,31,187,31,220,31,59,31,59,30,212,31,212,30,87,31,75,31,58,31,144,31,189,31,150,31,29,31,220,31,145,31,244,31,123,31,13,31,13,30,199,31,228,31,27,31,27,30,87,31,221,31,152,31,143,31,115,31,19,31,75,31,164,31,193,31,4,31,96,31,96,30,79,31,147,31,34,31,229,31,73,31,130,31,130,30,240,31,240,30,255,31,110,31,19,31,253,31,254,31,250,31,156,31,177,31,253,31,253,30,253,29,235,31,116,31,116,30,100,31,5,31,25,31,25,30,176,31,195,31,26,31,103,31,245,31,103,31,252,31,252,30,206,31,242,31,63,31,134,31,134,30,134,29,209,31,125,31,207,31,208,31,208,30,220,31,99,31,28,31,128,31,111,31,206,31,191,31,29,31,10,31,10,30,35,31,127,31,196,31,252,31,203,31,146,31,132,31,168,31,236,31,222,31,48,31,181,31,57,31,37,31,155,31,155,30,144,31,144,30,43,31,214,31,227,31,206,31,45,31,70,31,239,31,61,31,61,30,35,31,35,30,100,31,100,30,142,31,202,31,218,31,218,30,62,31,62,30,29,31,48,31,48,30,205,31,234,31,244,31,173,31,137,31,57,31,132,31,54,31,238,31,238,30,51,31,228,31,99,31,121,31,73,31,137,31,35,31,124,31,219,31,42,31,48,31,150,31,192,31,168,31,168,30,205,31,208,31,98,31,98,30,116,31,198,31,63,31,188,31,39,31,36,31,36,30,36,29,80,31,80,30,44,31,44,30,187,31,217,31,40,31,40,30,65,31,123,31,48,31,51,31,45,31,45,30,108,31,178,31,237,31,35,31,35,30,201,31,201,30,7,31,145,31,108,31,112,31,7,31,7,30,114,31,152,31,88,31,83,31,83,30,31,31,13,31,13,30,13,29,13,28,238,31,27,31,27,30,170,31,80,31,217,31,32,31,32,30,145,31,148,31,204,31,204,30,187,31,113,31,225,31,131,31,131,30,131,29,143,31,143,30,230,31,166,31,166,30,213,31,213,30,213,29,42,31,72,31,27,31,27,30,91,31,91,30,91,29,217,31,125,31,125,30,156,31,232,31,27,31,224,31,235,31,132,31,193,31,234,31,234,31,79,31,39,31,87,31,245,31,51,31,51,30,123,31,199,31,198,31,198,30,218,31,189,31,177,31,177,30,152,31,19,31,183,31,164,31,96,31,238,31,250,31,68,31,68,30,101,31,188,31,188,30,188,29,14,31,110,31,172,31,178,31,252,31,252,30,215,31,186,31,101,31,111,31,61,31,61,30,106,31,183,31,104,31,104,30,113,31,6,31,250,31,63,31,63,30,212,31,195,31,195,30,62,31,158,31,153,31,153,30,45,31,63,31,101,31,101,30,101,29,240,31,19,31,119,31,119,30,195,31,189,31,189,30,191,31,151,31,173,31,151,31,89,31,95,31,36,31,46,31,221,31,73,31,155,31,155,30,143,31,81,31,40,31,61,31,218,31,203,31,203,30,233,31,53,31,53,30,53,29,45,31,137,31,228,31,4,31,86,31,101,31,88,31,232,31,34,31,242,31,204,31,204,30,204,29,144,31,144,30,76,31,201,31,201,30,181,31,216,31,230,31,141,31,141,30,113,31,33,31,70,31,70,30,47,31,47,30,243,31,140,31,127,31,191,31,20,31,3,31,194,31,121,31,93,31,40,31,40,30,146,31,232,31,19,31,229,31,18,31,83,31,139,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
