-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_438 is
end project_tb_438;

architecture project_tb_arch_438 of project_tb_438 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 845;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,173,0,0,0,0,0,90,0,51,0,52,0,0,0,0,0,150,0,168,0,0,0,65,0,136,0,0,0,236,0,83,0,0,0,0,0,0,0,186,0,0,0,11,0,170,0,146,0,9,0,75,0,0,0,160,0,215,0,192,0,100,0,0,0,0,0,0,0,9,0,81,0,0,0,0,0,100,0,4,0,199,0,35,0,220,0,32,0,150,0,75,0,208,0,0,0,0,0,160,0,0,0,142,0,0,0,0,0,46,0,0,0,228,0,43,0,134,0,27,0,58,0,90,0,0,0,0,0,0,0,91,0,201,0,76,0,0,0,0,0,110,0,96,0,97,0,0,0,0,0,0,0,0,0,20,0,163,0,29,0,6,0,30,0,176,0,153,0,15,0,170,0,4,0,122,0,8,0,55,0,22,0,255,0,0,0,0,0,0,0,40,0,0,0,0,0,0,0,246,0,0,0,181,0,252,0,128,0,124,0,99,0,253,0,57,0,62,0,72,0,161,0,8,0,212,0,0,0,60,0,148,0,58,0,196,0,202,0,219,0,0,0,0,0,253,0,0,0,0,0,0,0,0,0,0,0,131,0,124,0,85,0,22,0,211,0,215,0,0,0,123,0,49,0,0,0,72,0,186,0,137,0,0,0,104,0,203,0,230,0,0,0,9,0,146,0,179,0,0,0,170,0,143,0,187,0,128,0,94,0,39,0,92,0,220,0,0,0,11,0,203,0,145,0,188,0,240,0,37,0,31,0,32,0,186,0,60,0,175,0,182,0,35,0,0,0,142,0,59,0,112,0,74,0,241,0,21,0,156,0,215,0,223,0,72,0,239,0,140,0,138,0,74,0,234,0,213,0,118,0,150,0,26,0,51,0,62,0,51,0,206,0,0,0,123,0,0,0,181,0,125,0,0,0,37,0,88,0,43,0,84,0,21,0,0,0,104,0,85,0,0,0,47,0,40,0,0,0,118,0,232,0,95,0,139,0,83,0,175,0,104,0,191,0,170,0,184,0,186,0,204,0,118,0,217,0,186,0,0,0,111,0,25,0,126,0,213,0,0,0,50,0,239,0,134,0,29,0,63,0,170,0,36,0,0,0,139,0,138,0,30,0,0,0,0,0,138,0,0,0,76,0,0,0,0,0,17,0,201,0,209,0,122,0,34,0,107,0,146,0,180,0,0,0,134,0,63,0,7,0,231,0,68,0,53,0,151,0,138,0,96,0,19,0,103,0,66,0,36,0,160,0,163,0,0,0,28,0,246,0,163,0,85,0,0,0,0,0,8,0,62,0,102,0,204,0,36,0,191,0,164,0,11,0,84,0,147,0,91,0,36,0,108,0,0,0,0,0,0,0,63,0,116,0,189,0,0,0,14,0,166,0,207,0,107,0,229,0,79,0,110,0,99,0,98,0,0,0,99,0,0,0,62,0,62,0,0,0,186,0,179,0,0,0,216,0,180,0,228,0,115,0,10,0,0,0,228,0,240,0,116,0,20,0,0,0,185,0,163,0,145,0,175,0,176,0,9,0,0,0,107,0,236,0,254,0,0,0,0,0,208,0,178,0,223,0,0,0,89,0,41,0,29,0,86,0,134,0,0,0,55,0,184,0,191,0,52,0,0,0,5,0,64,0,195,0,52,0,92,0,169,0,0,0,189,0,0,0,207,0,167,0,18,0,187,0,48,0,0,0,145,0,74,0,43,0,187,0,0,0,243,0,83,0,51,0,14,0,0,0,243,0,7,0,37,0,194,0,226,0,8,0,0,0,90,0,157,0,98,0,0,0,216,0,25,0,57,0,234,0,237,0,211,0,0,0,47,0,154,0,0,0,78,0,175,0,58,0,239,0,201,0,221,0,0,0,34,0,201,0,147,0,107,0,151,0,30,0,0,0,244,0,203,0,14,0,71,0,179,0,0,0,0,0,195,0,182,0,0,0,175,0,0,0,215,0,30,0,21,0,217,0,248,0,0,0,213,0,0,0,14,0,0,0,42,0,116,0,211,0,0,0,239,0,61,0,164,0,68,0,106,0,0,0,27,0,135,0,119,0,0,0,0,0,0,0,0,0,238,0,35,0,0,0,155,0,214,0,83,0,169,0,238,0,220,0,107,0,77,0,0,0,85,0,0,0,140,0,170,0,0,0,51,0,0,0,152,0,29,0,119,0,217,0,148,0,0,0,177,0,0,0,0,0,229,0,184,0,143,0,120,0,0,0,226,0,35,0,0,0,18,0,247,0,235,0,246,0,0,0,141,0,74,0,0,0,18,0,184,0,0,0,102,0,119,0,167,0,157,0,0,0,167,0,229,0,141,0,169,0,0,0,25,0,61,0,209,0,205,0,0,0,192,0,0,0,0,0,0,0,174,0,236,0,45,0,136,0,0,0,149,0,177,0,229,0,237,0,134,0,53,0,219,0,126,0,131,0,0,0,117,0,120,0,0,0,105,0,123,0,177,0,53,0,8,0,116,0,203,0,117,0,19,0,118,0,0,0,202,0,93,0,241,0,26,0,0,0,248,0,36,0,0,0,0,0,0,0,159,0,180,0,203,0,0,0,244,0,0,0,37,0,110,0,0,0,104,0,179,0,222,0,0,0,67,0,184,0,182,0,0,0,151,0,105,0,3,0,228,0,56,0,230,0,146,0,7,0,253,0,142,0,0,0,117,0,0,0,226,0,0,0,0,0,30,0,115,0,24,0,154,0,201,0,190,0,63,0,124,0,234,0,240,0,132,0,92,0,194,0,163,0,78,0,0,0,34,0,60,0,80,0,43,0,7,0,10,0,69,0,39,0,184,0,0,0,111,0,144,0,84,0,28,0,251,0,0,0,216,0,251,0,6,0,0,0,111,0,205,0,0,0,0,0,135,0,152,0,0,0,191,0,234,0,255,0,0,0,146,0,119,0,42,0,0,0,97,0,14,0,130,0,177,0,166,0,49,0,32,0,0,0,38,0,213,0,232,0,69,0,45,0,0,0,244,0,141,0,59,0,124,0,74,0,0,0,215,0,15,0,148,0,154,0,45,0,48,0,165,0,130,0,165,0,191,0,15,0,249,0,219,0,5,0,77,0,151,0,0,0,186,0,0,0,126,0,24,0,0,0,46,0,230,0,127,0,3,0,26,0,41,0,64,0,163,0,0,0,201,0,161,0,252,0,162,0,66,0,47,0,248,0,0,0,99,0,41,0,57,0,242,0,0,0,233,0,238,0,145,0,194,0,71,0,85,0,59,0,111,0,0,0,254,0,115,0,77,0,226,0,138,0,46,0,156,0,188,0,101,0,203,0,0,0,121,0,0,0,136,0,126,0,139,0,33,0,39,0,115,0,0,0,68,0,86,0,159,0,210,0,13,0,153,0,180,0,25,0,31,0,210,0,66,0,254,0,68,0,0,0,168,0,82,0,182,0,0,0,19,0,168,0,0,0,0,0,100,0,124,0,224,0,187,0,0,0,0,0,128,0,0,0,182,0,0,0,204,0,241,0,231,0,98,0,79,0,217,0,0,0,158,0,123,0,241,0,53,0,28,0,210,0,120,0,219,0,149,0,196,0,0,0,0,0,252,0,198,0,84,0,119,0,55,0,0,0,78,0,178,0,192,0,85,0,180,0,236,0,3,0,0,0,0,0,79,0,0,0,210,0,31,0,7,0,73,0,196,0,0,0,95,0,139,0,130,0,130,0,167,0,100,0,0,0,210,0,214,0,166,0,196,0,101,0,18,0,139,0,116,0,158,0,79,0,238,0,26,0,190,0,104,0,0,0,59,0,12,0,69,0,0,0,103,0,137,0,228,0);
signal scenario_full  : scenario_type := (0,0,173,31,173,30,173,29,90,31,51,31,52,31,52,30,52,29,150,31,168,31,168,30,65,31,136,31,136,30,236,31,83,31,83,30,83,29,83,28,186,31,186,30,11,31,170,31,146,31,9,31,75,31,75,30,160,31,215,31,192,31,100,31,100,30,100,29,100,28,9,31,81,31,81,30,81,29,100,31,4,31,199,31,35,31,220,31,32,31,150,31,75,31,208,31,208,30,208,29,160,31,160,30,142,31,142,30,142,29,46,31,46,30,228,31,43,31,134,31,27,31,58,31,90,31,90,30,90,29,90,28,91,31,201,31,76,31,76,30,76,29,110,31,96,31,97,31,97,30,97,29,97,28,97,27,20,31,163,31,29,31,6,31,30,31,176,31,153,31,15,31,170,31,4,31,122,31,8,31,55,31,22,31,255,31,255,30,255,29,255,28,40,31,40,30,40,29,40,28,246,31,246,30,181,31,252,31,128,31,124,31,99,31,253,31,57,31,62,31,72,31,161,31,8,31,212,31,212,30,60,31,148,31,58,31,196,31,202,31,219,31,219,30,219,29,253,31,253,30,253,29,253,28,253,27,253,26,131,31,124,31,85,31,22,31,211,31,215,31,215,30,123,31,49,31,49,30,72,31,186,31,137,31,137,30,104,31,203,31,230,31,230,30,9,31,146,31,179,31,179,30,170,31,143,31,187,31,128,31,94,31,39,31,92,31,220,31,220,30,11,31,203,31,145,31,188,31,240,31,37,31,31,31,32,31,186,31,60,31,175,31,182,31,35,31,35,30,142,31,59,31,112,31,74,31,241,31,21,31,156,31,215,31,223,31,72,31,239,31,140,31,138,31,74,31,234,31,213,31,118,31,150,31,26,31,51,31,62,31,51,31,206,31,206,30,123,31,123,30,181,31,125,31,125,30,37,31,88,31,43,31,84,31,21,31,21,30,104,31,85,31,85,30,47,31,40,31,40,30,118,31,232,31,95,31,139,31,83,31,175,31,104,31,191,31,170,31,184,31,186,31,204,31,118,31,217,31,186,31,186,30,111,31,25,31,126,31,213,31,213,30,50,31,239,31,134,31,29,31,63,31,170,31,36,31,36,30,139,31,138,31,30,31,30,30,30,29,138,31,138,30,76,31,76,30,76,29,17,31,201,31,209,31,122,31,34,31,107,31,146,31,180,31,180,30,134,31,63,31,7,31,231,31,68,31,53,31,151,31,138,31,96,31,19,31,103,31,66,31,36,31,160,31,163,31,163,30,28,31,246,31,163,31,85,31,85,30,85,29,8,31,62,31,102,31,204,31,36,31,191,31,164,31,11,31,84,31,147,31,91,31,36,31,108,31,108,30,108,29,108,28,63,31,116,31,189,31,189,30,14,31,166,31,207,31,107,31,229,31,79,31,110,31,99,31,98,31,98,30,99,31,99,30,62,31,62,31,62,30,186,31,179,31,179,30,216,31,180,31,228,31,115,31,10,31,10,30,228,31,240,31,116,31,20,31,20,30,185,31,163,31,145,31,175,31,176,31,9,31,9,30,107,31,236,31,254,31,254,30,254,29,208,31,178,31,223,31,223,30,89,31,41,31,29,31,86,31,134,31,134,30,55,31,184,31,191,31,52,31,52,30,5,31,64,31,195,31,52,31,92,31,169,31,169,30,189,31,189,30,207,31,167,31,18,31,187,31,48,31,48,30,145,31,74,31,43,31,187,31,187,30,243,31,83,31,51,31,14,31,14,30,243,31,7,31,37,31,194,31,226,31,8,31,8,30,90,31,157,31,98,31,98,30,216,31,25,31,57,31,234,31,237,31,211,31,211,30,47,31,154,31,154,30,78,31,175,31,58,31,239,31,201,31,221,31,221,30,34,31,201,31,147,31,107,31,151,31,30,31,30,30,244,31,203,31,14,31,71,31,179,31,179,30,179,29,195,31,182,31,182,30,175,31,175,30,215,31,30,31,21,31,217,31,248,31,248,30,213,31,213,30,14,31,14,30,42,31,116,31,211,31,211,30,239,31,61,31,164,31,68,31,106,31,106,30,27,31,135,31,119,31,119,30,119,29,119,28,119,27,238,31,35,31,35,30,155,31,214,31,83,31,169,31,238,31,220,31,107,31,77,31,77,30,85,31,85,30,140,31,170,31,170,30,51,31,51,30,152,31,29,31,119,31,217,31,148,31,148,30,177,31,177,30,177,29,229,31,184,31,143,31,120,31,120,30,226,31,35,31,35,30,18,31,247,31,235,31,246,31,246,30,141,31,74,31,74,30,18,31,184,31,184,30,102,31,119,31,167,31,157,31,157,30,167,31,229,31,141,31,169,31,169,30,25,31,61,31,209,31,205,31,205,30,192,31,192,30,192,29,192,28,174,31,236,31,45,31,136,31,136,30,149,31,177,31,229,31,237,31,134,31,53,31,219,31,126,31,131,31,131,30,117,31,120,31,120,30,105,31,123,31,177,31,53,31,8,31,116,31,203,31,117,31,19,31,118,31,118,30,202,31,93,31,241,31,26,31,26,30,248,31,36,31,36,30,36,29,36,28,159,31,180,31,203,31,203,30,244,31,244,30,37,31,110,31,110,30,104,31,179,31,222,31,222,30,67,31,184,31,182,31,182,30,151,31,105,31,3,31,228,31,56,31,230,31,146,31,7,31,253,31,142,31,142,30,117,31,117,30,226,31,226,30,226,29,30,31,115,31,24,31,154,31,201,31,190,31,63,31,124,31,234,31,240,31,132,31,92,31,194,31,163,31,78,31,78,30,34,31,60,31,80,31,43,31,7,31,10,31,69,31,39,31,184,31,184,30,111,31,144,31,84,31,28,31,251,31,251,30,216,31,251,31,6,31,6,30,111,31,205,31,205,30,205,29,135,31,152,31,152,30,191,31,234,31,255,31,255,30,146,31,119,31,42,31,42,30,97,31,14,31,130,31,177,31,166,31,49,31,32,31,32,30,38,31,213,31,232,31,69,31,45,31,45,30,244,31,141,31,59,31,124,31,74,31,74,30,215,31,15,31,148,31,154,31,45,31,48,31,165,31,130,31,165,31,191,31,15,31,249,31,219,31,5,31,77,31,151,31,151,30,186,31,186,30,126,31,24,31,24,30,46,31,230,31,127,31,3,31,26,31,41,31,64,31,163,31,163,30,201,31,161,31,252,31,162,31,66,31,47,31,248,31,248,30,99,31,41,31,57,31,242,31,242,30,233,31,238,31,145,31,194,31,71,31,85,31,59,31,111,31,111,30,254,31,115,31,77,31,226,31,138,31,46,31,156,31,188,31,101,31,203,31,203,30,121,31,121,30,136,31,126,31,139,31,33,31,39,31,115,31,115,30,68,31,86,31,159,31,210,31,13,31,153,31,180,31,25,31,31,31,210,31,66,31,254,31,68,31,68,30,168,31,82,31,182,31,182,30,19,31,168,31,168,30,168,29,100,31,124,31,224,31,187,31,187,30,187,29,128,31,128,30,182,31,182,30,204,31,241,31,231,31,98,31,79,31,217,31,217,30,158,31,123,31,241,31,53,31,28,31,210,31,120,31,219,31,149,31,196,31,196,30,196,29,252,31,198,31,84,31,119,31,55,31,55,30,78,31,178,31,192,31,85,31,180,31,236,31,3,31,3,30,3,29,79,31,79,30,210,31,31,31,7,31,73,31,196,31,196,30,95,31,139,31,130,31,130,31,167,31,100,31,100,30,210,31,214,31,166,31,196,31,101,31,18,31,139,31,116,31,158,31,79,31,238,31,26,31,190,31,104,31,104,30,59,31,12,31,69,31,69,30,103,31,137,31,228,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
