-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_556 is
end project_tb_556;

architecture project_tb_arch_556 of project_tb_556 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 773;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (186,0,0,0,202,0,212,0,97,0,254,0,0,0,252,0,187,0,184,0,139,0,0,0,25,0,0,0,147,0,66,0,99,0,0,0,22,0,0,0,0,0,0,0,0,0,158,0,236,0,52,0,0,0,143,0,244,0,147,0,129,0,16,0,0,0,179,0,151,0,0,0,122,0,0,0,0,0,159,0,86,0,163,0,0,0,249,0,231,0,127,0,107,0,232,0,246,0,159,0,178,0,98,0,191,0,35,0,53,0,183,0,20,0,207,0,0,0,102,0,0,0,179,0,0,0,255,0,0,0,0,0,112,0,27,0,244,0,217,0,148,0,24,0,39,0,111,0,21,0,0,0,71,0,10,0,0,0,159,0,0,0,0,0,189,0,167,0,187,0,0,0,234,0,215,0,115,0,44,0,132,0,137,0,0,0,83,0,50,0,44,0,198,0,11,0,0,0,0,0,0,0,3,0,205,0,0,0,148,0,67,0,19,0,99,0,30,0,0,0,196,0,0,0,43,0,0,0,7,0,150,0,0,0,0,0,46,0,8,0,179,0,244,0,167,0,0,0,89,0,27,0,0,0,203,0,203,0,90,0,72,0,7,0,34,0,74,0,0,0,0,0,102,0,243,0,0,0,0,0,11,0,99,0,182,0,236,0,59,0,179,0,245,0,105,0,0,0,244,0,217,0,227,0,138,0,30,0,60,0,77,0,42,0,0,0,150,0,197,0,0,0,62,0,0,0,229,0,154,0,52,0,0,0,176,0,186,0,61,0,107,0,127,0,141,0,129,0,86,0,0,0,167,0,252,0,166,0,196,0,18,0,225,0,97,0,0,0,225,0,204,0,86,0,134,0,0,0,209,0,212,0,87,0,89,0,175,0,154,0,61,0,234,0,0,0,29,0,0,0,211,0,245,0,95,0,140,0,0,0,147,0,195,0,177,0,0,0,0,0,17,0,44,0,251,0,114,0,229,0,218,0,125,0,179,0,39,0,48,0,123,0,74,0,0,0,240,0,198,0,193,0,97,0,0,0,0,0,227,0,0,0,49,0,154,0,224,0,57,0,0,0,24,0,47,0,0,0,74,0,127,0,241,0,246,0,0,0,0,0,110,0,0,0,117,0,0,0,190,0,115,0,110,0,0,0,96,0,156,0,0,0,231,0,68,0,211,0,0,0,18,0,96,0,38,0,43,0,5,0,1,0,45,0,123,0,66,0,4,0,64,0,216,0,122,0,115,0,99,0,122,0,219,0,94,0,141,0,91,0,0,0,20,0,122,0,16,0,0,0,247,0,185,0,0,0,80,0,55,0,83,0,96,0,219,0,211,0,216,0,0,0,182,0,48,0,5,0,0,0,254,0,215,0,0,0,146,0,188,0,0,0,42,0,200,0,114,0,0,0,13,0,81,0,50,0,92,0,168,0,0,0,58,0,168,0,0,0,0,0,197,0,0,0,190,0,135,0,157,0,22,0,8,0,0,0,60,0,0,0,35,0,223,0,0,0,144,0,80,0,0,0,0,0,95,0,34,0,50,0,100,0,205,0,22,0,86,0,131,0,2,0,0,0,216,0,31,0,178,0,59,0,0,0,0,0,0,0,149,0,0,0,113,0,193,0,203,0,116,0,0,0,45,0,134,0,0,0,175,0,0,0,0,0,130,0,16,0,62,0,0,0,231,0,47,0,24,0,92,0,0,0,207,0,67,0,8,0,184,0,139,0,203,0,17,0,0,0,163,0,62,0,29,0,252,0,149,0,248,0,0,0,197,0,43,0,166,0,0,0,67,0,137,0,0,0,217,0,150,0,190,0,107,0,216,0,36,0,150,0,186,0,84,0,82,0,91,0,0,0,165,0,35,0,0,0,15,0,29,0,0,0,0,0,127,0,96,0,158,0,131,0,0,0,94,0,0,0,189,0,0,0,210,0,83,0,229,0,202,0,163,0,30,0,154,0,120,0,212,0,76,0,182,0,10,0,0,0,0,0,76,0,131,0,235,0,206,0,134,0,139,0,151,0,0,0,84,0,148,0,117,0,0,0,171,0,151,0,28,0,216,0,0,0,106,0,0,0,137,0,146,0,252,0,157,0,169,0,92,0,213,0,0,0,242,0,179,0,0,0,0,0,132,0,110,0,69,0,0,0,203,0,163,0,207,0,189,0,51,0,183,0,69,0,184,0,141,0,213,0,25,0,234,0,100,0,62,0,15,0,151,0,50,0,9,0,249,0,47,0,0,0,9,0,97,0,167,0,233,0,113,0,129,0,0,0,51,0,72,0,245,0,45,0,177,0,5,0,87,0,228,0,0,0,0,0,0,0,0,0,242,0,222,0,185,0,0,0,189,0,128,0,0,0,204,0,0,0,206,0,75,0,166,0,4,0,237,0,224,0,230,0,0,0,200,0,174,0,0,0,0,0,64,0,0,0,22,0,162,0,16,0,6,0,123,0,19,0,24,0,174,0,88,0,188,0,35,0,0,0,245,0,6,0,0,0,0,0,199,0,222,0,125,0,0,0,179,0,93,0,118,0,26,0,1,0,30,0,167,0,3,0,18,0,85,0,147,0,205,0,245,0,0,0,58,0,146,0,55,0,0,0,180,0,147,0,234,0,0,0,195,0,0,0,25,0,56,0,37,0,247,0,1,0,8,0,132,0,68,0,81,0,0,0,129,0,71,0,0,0,232,0,253,0,89,0,0,0,186,0,105,0,0,0,209,0,0,0,158,0,98,0,222,0,200,0,172,0,198,0,0,0,39,0,0,0,178,0,60,0,172,0,17,0,27,0,210,0,40,0,121,0,0,0,211,0,67,0,30,0,49,0,87,0,0,0,9,0,91,0,152,0,71,0,24,0,90,0,77,0,89,0,24,0,240,0,203,0,0,0,4,0,122,0,52,0,52,0,134,0,155,0,0,0,249,0,45,0,49,0,127,0,29,0,0,0,215,0,22,0,0,0,103,0,205,0,156,0,162,0,87,0,121,0,57,0,163,0,118,0,225,0,172,0,162,0,247,0,95,0,151,0,212,0,14,0,140,0,43,0,169,0,153,0,149,0,9,0,163,0,172,0,211,0,153,0,121,0,0,0,195,0,249,0,193,0,255,0,24,0,66,0,48,0,151,0,90,0,159,0,86,0,26,0,202,0,0,0,34,0,50,0,0,0,35,0,0,0,189,0,0,0,186,0,0,0,93,0,27,0,17,0,124,0,189,0,0,0,110,0,249,0,120,0,102,0,97,0,176,0,16,0,51,0,157,0,7,0,162,0,0,0,141,0,67,0,88,0,108,0,40,0,130,0,37,0,0,0,21,0,236,0,145,0,16,0,100,0,21,0,224,0,229,0,142,0,0,0,74,0,78,0,99,0,1,0,238,0,0,0,37,0,36,0,53,0,190,0,166,0,178,0,74,0,0,0,180,0,52,0,0,0,240,0,239,0,178,0,142,0,0,0,0,0,29,0,51,0,0,0,105,0,92,0,58,0);
signal scenario_full  : scenario_type := (186,31,186,30,202,31,212,31,97,31,254,31,254,30,252,31,187,31,184,31,139,31,139,30,25,31,25,30,147,31,66,31,99,31,99,30,22,31,22,30,22,29,22,28,22,27,158,31,236,31,52,31,52,30,143,31,244,31,147,31,129,31,16,31,16,30,179,31,151,31,151,30,122,31,122,30,122,29,159,31,86,31,163,31,163,30,249,31,231,31,127,31,107,31,232,31,246,31,159,31,178,31,98,31,191,31,35,31,53,31,183,31,20,31,207,31,207,30,102,31,102,30,179,31,179,30,255,31,255,30,255,29,112,31,27,31,244,31,217,31,148,31,24,31,39,31,111,31,21,31,21,30,71,31,10,31,10,30,159,31,159,30,159,29,189,31,167,31,187,31,187,30,234,31,215,31,115,31,44,31,132,31,137,31,137,30,83,31,50,31,44,31,198,31,11,31,11,30,11,29,11,28,3,31,205,31,205,30,148,31,67,31,19,31,99,31,30,31,30,30,196,31,196,30,43,31,43,30,7,31,150,31,150,30,150,29,46,31,8,31,179,31,244,31,167,31,167,30,89,31,27,31,27,30,203,31,203,31,90,31,72,31,7,31,34,31,74,31,74,30,74,29,102,31,243,31,243,30,243,29,11,31,99,31,182,31,236,31,59,31,179,31,245,31,105,31,105,30,244,31,217,31,227,31,138,31,30,31,60,31,77,31,42,31,42,30,150,31,197,31,197,30,62,31,62,30,229,31,154,31,52,31,52,30,176,31,186,31,61,31,107,31,127,31,141,31,129,31,86,31,86,30,167,31,252,31,166,31,196,31,18,31,225,31,97,31,97,30,225,31,204,31,86,31,134,31,134,30,209,31,212,31,87,31,89,31,175,31,154,31,61,31,234,31,234,30,29,31,29,30,211,31,245,31,95,31,140,31,140,30,147,31,195,31,177,31,177,30,177,29,17,31,44,31,251,31,114,31,229,31,218,31,125,31,179,31,39,31,48,31,123,31,74,31,74,30,240,31,198,31,193,31,97,31,97,30,97,29,227,31,227,30,49,31,154,31,224,31,57,31,57,30,24,31,47,31,47,30,74,31,127,31,241,31,246,31,246,30,246,29,110,31,110,30,117,31,117,30,190,31,115,31,110,31,110,30,96,31,156,31,156,30,231,31,68,31,211,31,211,30,18,31,96,31,38,31,43,31,5,31,1,31,45,31,123,31,66,31,4,31,64,31,216,31,122,31,115,31,99,31,122,31,219,31,94,31,141,31,91,31,91,30,20,31,122,31,16,31,16,30,247,31,185,31,185,30,80,31,55,31,83,31,96,31,219,31,211,31,216,31,216,30,182,31,48,31,5,31,5,30,254,31,215,31,215,30,146,31,188,31,188,30,42,31,200,31,114,31,114,30,13,31,81,31,50,31,92,31,168,31,168,30,58,31,168,31,168,30,168,29,197,31,197,30,190,31,135,31,157,31,22,31,8,31,8,30,60,31,60,30,35,31,223,31,223,30,144,31,80,31,80,30,80,29,95,31,34,31,50,31,100,31,205,31,22,31,86,31,131,31,2,31,2,30,216,31,31,31,178,31,59,31,59,30,59,29,59,28,149,31,149,30,113,31,193,31,203,31,116,31,116,30,45,31,134,31,134,30,175,31,175,30,175,29,130,31,16,31,62,31,62,30,231,31,47,31,24,31,92,31,92,30,207,31,67,31,8,31,184,31,139,31,203,31,17,31,17,30,163,31,62,31,29,31,252,31,149,31,248,31,248,30,197,31,43,31,166,31,166,30,67,31,137,31,137,30,217,31,150,31,190,31,107,31,216,31,36,31,150,31,186,31,84,31,82,31,91,31,91,30,165,31,35,31,35,30,15,31,29,31,29,30,29,29,127,31,96,31,158,31,131,31,131,30,94,31,94,30,189,31,189,30,210,31,83,31,229,31,202,31,163,31,30,31,154,31,120,31,212,31,76,31,182,31,10,31,10,30,10,29,76,31,131,31,235,31,206,31,134,31,139,31,151,31,151,30,84,31,148,31,117,31,117,30,171,31,151,31,28,31,216,31,216,30,106,31,106,30,137,31,146,31,252,31,157,31,169,31,92,31,213,31,213,30,242,31,179,31,179,30,179,29,132,31,110,31,69,31,69,30,203,31,163,31,207,31,189,31,51,31,183,31,69,31,184,31,141,31,213,31,25,31,234,31,100,31,62,31,15,31,151,31,50,31,9,31,249,31,47,31,47,30,9,31,97,31,167,31,233,31,113,31,129,31,129,30,51,31,72,31,245,31,45,31,177,31,5,31,87,31,228,31,228,30,228,29,228,28,228,27,242,31,222,31,185,31,185,30,189,31,128,31,128,30,204,31,204,30,206,31,75,31,166,31,4,31,237,31,224,31,230,31,230,30,200,31,174,31,174,30,174,29,64,31,64,30,22,31,162,31,16,31,6,31,123,31,19,31,24,31,174,31,88,31,188,31,35,31,35,30,245,31,6,31,6,30,6,29,199,31,222,31,125,31,125,30,179,31,93,31,118,31,26,31,1,31,30,31,167,31,3,31,18,31,85,31,147,31,205,31,245,31,245,30,58,31,146,31,55,31,55,30,180,31,147,31,234,31,234,30,195,31,195,30,25,31,56,31,37,31,247,31,1,31,8,31,132,31,68,31,81,31,81,30,129,31,71,31,71,30,232,31,253,31,89,31,89,30,186,31,105,31,105,30,209,31,209,30,158,31,98,31,222,31,200,31,172,31,198,31,198,30,39,31,39,30,178,31,60,31,172,31,17,31,27,31,210,31,40,31,121,31,121,30,211,31,67,31,30,31,49,31,87,31,87,30,9,31,91,31,152,31,71,31,24,31,90,31,77,31,89,31,24,31,240,31,203,31,203,30,4,31,122,31,52,31,52,31,134,31,155,31,155,30,249,31,45,31,49,31,127,31,29,31,29,30,215,31,22,31,22,30,103,31,205,31,156,31,162,31,87,31,121,31,57,31,163,31,118,31,225,31,172,31,162,31,247,31,95,31,151,31,212,31,14,31,140,31,43,31,169,31,153,31,149,31,9,31,163,31,172,31,211,31,153,31,121,31,121,30,195,31,249,31,193,31,255,31,24,31,66,31,48,31,151,31,90,31,159,31,86,31,26,31,202,31,202,30,34,31,50,31,50,30,35,31,35,30,189,31,189,30,186,31,186,30,93,31,27,31,17,31,124,31,189,31,189,30,110,31,249,31,120,31,102,31,97,31,176,31,16,31,51,31,157,31,7,31,162,31,162,30,141,31,67,31,88,31,108,31,40,31,130,31,37,31,37,30,21,31,236,31,145,31,16,31,100,31,21,31,224,31,229,31,142,31,142,30,74,31,78,31,99,31,1,31,238,31,238,30,37,31,36,31,53,31,190,31,166,31,178,31,74,31,74,30,180,31,52,31,52,30,240,31,239,31,178,31,142,31,142,30,142,29,29,31,51,31,51,30,105,31,92,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
