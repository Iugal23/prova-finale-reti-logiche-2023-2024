-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 759;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,30,0,252,0,30,0,232,0,165,0,11,0,205,0,0,0,118,0,0,0,0,0,226,0,0,0,0,0,0,0,0,0,0,0,10,0,0,0,120,0,0,0,108,0,19,0,0,0,19,0,207,0,98,0,102,0,208,0,65,0,199,0,0,0,60,0,152,0,224,0,108,0,214,0,0,0,103,0,115,0,0,0,0,0,138,0,6,0,35,0,50,0,0,0,209,0,83,0,63,0,66,0,251,0,50,0,204,0,132,0,68,0,166,0,141,0,128,0,161,0,0,0,33,0,0,0,0,0,244,0,162,0,58,0,80,0,0,0,48,0,62,0,229,0,77,0,125,0,10,0,124,0,142,0,138,0,236,0,150,0,0,0,0,0,209,0,94,0,53,0,244,0,0,0,73,0,142,0,219,0,0,0,80,0,23,0,117,0,49,0,72,0,255,0,242,0,202,0,91,0,154,0,118,0,25,0,156,0,90,0,2,0,22,0,175,0,73,0,113,0,77,0,214,0,0,0,225,0,166,0,26,0,0,0,117,0,0,0,204,0,9,0,69,0,23,0,224,0,194,0,185,0,235,0,141,0,251,0,229,0,7,0,59,0,164,0,235,0,149,0,235,0,0,0,0,0,0,0,0,0,112,0,234,0,93,0,0,0,58,0,0,0,129,0,100,0,109,0,159,0,0,0,247,0,197,0,0,0,107,0,143,0,135,0,33,0,209,0,98,0,248,0,143,0,55,0,0,0,210,0,162,0,0,0,243,0,222,0,116,0,110,0,47,0,0,0,107,0,93,0,182,0,151,0,108,0,115,0,0,0,0,0,10,0,211,0,94,0,0,0,0,0,3,0,48,0,145,0,202,0,143,0,48,0,46,0,227,0,62,0,59,0,0,0,0,0,0,0,117,0,0,0,118,0,137,0,4,0,250,0,42,0,135,0,238,0,91,0,142,0,0,0,137,0,203,0,105,0,164,0,0,0,35,0,0,0,190,0,141,0,248,0,81,0,226,0,218,0,4,0,249,0,128,0,134,0,34,0,27,0,17,0,0,0,208,0,75,0,11,0,92,0,164,0,162,0,0,0,0,0,0,0,77,0,114,0,61,0,0,0,56,0,171,0,114,0,148,0,163,0,248,0,39,0,152,0,89,0,0,0,22,0,0,0,52,0,169,0,3,0,0,0,0,0,8,0,225,0,196,0,10,0,0,0,224,0,138,0,167,0,20,0,0,0,63,0,199,0,141,0,207,0,196,0,50,0,49,0,5,0,115,0,217,0,219,0,151,0,0,0,178,0,84,0,0,0,195,0,92,0,208,0,211,0,54,0,0,0,129,0,123,0,97,0,141,0,0,0,74,0,146,0,237,0,0,0,0,0,211,0,102,0,240,0,136,0,63,0,116,0,0,0,0,0,253,0,0,0,90,0,76,0,16,0,35,0,199,0,0,0,0,0,49,0,34,0,128,0,212,0,119,0,0,0,199,0,82,0,0,0,20,0,178,0,83,0,152,0,33,0,35,0,199,0,67,0,36,0,240,0,252,0,0,0,25,0,100,0,0,0,211,0,28,0,27,0,227,0,84,0,0,0,233,0,1,0,0,0,0,0,212,0,124,0,64,0,125,0,248,0,32,0,38,0,27,0,0,0,31,0,94,0,0,0,0,0,16,0,25,0,0,0,0,0,0,0,0,0,0,0,215,0,53,0,7,0,0,0,0,0,206,0,54,0,0,0,64,0,85,0,0,0,111,0,218,0,23,0,167,0,0,0,118,0,217,0,0,0,196,0,0,0,0,0,111,0,180,0,31,0,241,0,213,0,22,0,113,0,211,0,128,0,20,0,205,0,161,0,58,0,0,0,146,0,233,0,110,0,254,0,43,0,2,0,204,0,226,0,51,0,33,0,142,0,40,0,44,0,123,0,0,0,47,0,212,0,0,0,80,0,0,0,69,0,37,0,189,0,0,0,74,0,10,0,203,0,83,0,128,0,169,0,0,0,185,0,0,0,4,0,28,0,108,0,157,0,50,0,179,0,175,0,99,0,88,0,11,0,91,0,0,0,214,0,109,0,151,0,72,0,213,0,232,0,221,0,226,0,21,0,133,0,9,0,106,0,146,0,243,0,138,0,0,0,199,0,28,0,114,0,0,0,0,0,0,0,0,0,0,0,81,0,138,0,102,0,86,0,8,0,28,0,34,0,186,0,38,0,146,0,79,0,121,0,0,0,155,0,157,0,0,0,30,0,0,0,0,0,139,0,87,0,179,0,117,0,0,0,0,0,232,0,120,0,54,0,0,0,62,0,216,0,251,0,215,0,0,0,0,0,64,0,237,0,189,0,255,0,25,0,87,0,163,0,114,0,91,0,0,0,35,0,2,0,0,0,121,0,172,0,0,0,117,0,0,0,185,0,11,0,53,0,130,0,253,0,62,0,183,0,0,0,179,0,128,0,0,0,249,0,207,0,42,0,14,0,0,0,1,0,57,0,214,0,78,0,98,0,0,0,134,0,94,0,53,0,80,0,0,0,0,0,163,0,193,0,13,0,0,0,179,0,131,0,223,0,28,0,95,0,251,0,164,0,0,0,152,0,139,0,14,0,0,0,215,0,63,0,0,0,220,0,0,0,0,0,129,0,73,0,102,0,172,0,36,0,141,0,225,0,244,0,252,0,206,0,42,0,58,0,120,0,72,0,219,0,163,0,52,0,0,0,235,0,56,0,0,0,56,0,0,0,0,0,134,0,189,0,105,0,56,0,218,0,180,0,4,0,249,0,185,0,240,0,0,0,226,0,95,0,46,0,38,0,129,0,0,0,149,0,0,0,186,0,134,0,0,0,145,0,88,0,231,0,184,0,216,0,0,0,4,0,0,0,0,0,59,0,48,0,45,0,169,0,198,0,123,0,0,0,0,0,0,0,197,0,204,0,225,0,159,0,205,0,0,0,252,0,187,0,127,0,83,0,110,0,231,0,168,0,242,0,212,0,229,0,0,0,68,0,91,0,0,0,136,0,132,0,0,0,121,0,23,0,250,0,0,0,164,0,188,0,0,0,164,0,0,0,0,0,121,0,133,0,51,0,177,0,185,0,1,0,113,0,153,0,225,0,30,0,162,0,166,0,0,0,0,0,244,0,128,0,2,0,58,0,0,0,207,0,172,0,0,0,12,0,237,0,64,0,0,0,76,0,212,0,105,0,88,0,73,0,244,0,59,0,9,0,122,0,73,0,74,0,24,0,52,0,58,0,118,0,0,0,139,0,0,0,232,0,138,0,218,0,157,0,107,0,191,0,119,0,64,0,0,0,0,0,211,0,133,0,92,0,177,0,0,0,163,0,100,0,0,0,135,0,69,0,117,0,53,0,141,0,114,0,138,0,0,0,71,0,116,0,29,0,22,0,0,0,12,0,209,0,11,0);
signal scenario_full  : scenario_type := (0,0,30,31,252,31,30,31,232,31,165,31,11,31,205,31,205,30,118,31,118,30,118,29,226,31,226,30,226,29,226,28,226,27,226,26,10,31,10,30,120,31,120,30,108,31,19,31,19,30,19,31,207,31,98,31,102,31,208,31,65,31,199,31,199,30,60,31,152,31,224,31,108,31,214,31,214,30,103,31,115,31,115,30,115,29,138,31,6,31,35,31,50,31,50,30,209,31,83,31,63,31,66,31,251,31,50,31,204,31,132,31,68,31,166,31,141,31,128,31,161,31,161,30,33,31,33,30,33,29,244,31,162,31,58,31,80,31,80,30,48,31,62,31,229,31,77,31,125,31,10,31,124,31,142,31,138,31,236,31,150,31,150,30,150,29,209,31,94,31,53,31,244,31,244,30,73,31,142,31,219,31,219,30,80,31,23,31,117,31,49,31,72,31,255,31,242,31,202,31,91,31,154,31,118,31,25,31,156,31,90,31,2,31,22,31,175,31,73,31,113,31,77,31,214,31,214,30,225,31,166,31,26,31,26,30,117,31,117,30,204,31,9,31,69,31,23,31,224,31,194,31,185,31,235,31,141,31,251,31,229,31,7,31,59,31,164,31,235,31,149,31,235,31,235,30,235,29,235,28,235,27,112,31,234,31,93,31,93,30,58,31,58,30,129,31,100,31,109,31,159,31,159,30,247,31,197,31,197,30,107,31,143,31,135,31,33,31,209,31,98,31,248,31,143,31,55,31,55,30,210,31,162,31,162,30,243,31,222,31,116,31,110,31,47,31,47,30,107,31,93,31,182,31,151,31,108,31,115,31,115,30,115,29,10,31,211,31,94,31,94,30,94,29,3,31,48,31,145,31,202,31,143,31,48,31,46,31,227,31,62,31,59,31,59,30,59,29,59,28,117,31,117,30,118,31,137,31,4,31,250,31,42,31,135,31,238,31,91,31,142,31,142,30,137,31,203,31,105,31,164,31,164,30,35,31,35,30,190,31,141,31,248,31,81,31,226,31,218,31,4,31,249,31,128,31,134,31,34,31,27,31,17,31,17,30,208,31,75,31,11,31,92,31,164,31,162,31,162,30,162,29,162,28,77,31,114,31,61,31,61,30,56,31,171,31,114,31,148,31,163,31,248,31,39,31,152,31,89,31,89,30,22,31,22,30,52,31,169,31,3,31,3,30,3,29,8,31,225,31,196,31,10,31,10,30,224,31,138,31,167,31,20,31,20,30,63,31,199,31,141,31,207,31,196,31,50,31,49,31,5,31,115,31,217,31,219,31,151,31,151,30,178,31,84,31,84,30,195,31,92,31,208,31,211,31,54,31,54,30,129,31,123,31,97,31,141,31,141,30,74,31,146,31,237,31,237,30,237,29,211,31,102,31,240,31,136,31,63,31,116,31,116,30,116,29,253,31,253,30,90,31,76,31,16,31,35,31,199,31,199,30,199,29,49,31,34,31,128,31,212,31,119,31,119,30,199,31,82,31,82,30,20,31,178,31,83,31,152,31,33,31,35,31,199,31,67,31,36,31,240,31,252,31,252,30,25,31,100,31,100,30,211,31,28,31,27,31,227,31,84,31,84,30,233,31,1,31,1,30,1,29,212,31,124,31,64,31,125,31,248,31,32,31,38,31,27,31,27,30,31,31,94,31,94,30,94,29,16,31,25,31,25,30,25,29,25,28,25,27,25,26,215,31,53,31,7,31,7,30,7,29,206,31,54,31,54,30,64,31,85,31,85,30,111,31,218,31,23,31,167,31,167,30,118,31,217,31,217,30,196,31,196,30,196,29,111,31,180,31,31,31,241,31,213,31,22,31,113,31,211,31,128,31,20,31,205,31,161,31,58,31,58,30,146,31,233,31,110,31,254,31,43,31,2,31,204,31,226,31,51,31,33,31,142,31,40,31,44,31,123,31,123,30,47,31,212,31,212,30,80,31,80,30,69,31,37,31,189,31,189,30,74,31,10,31,203,31,83,31,128,31,169,31,169,30,185,31,185,30,4,31,28,31,108,31,157,31,50,31,179,31,175,31,99,31,88,31,11,31,91,31,91,30,214,31,109,31,151,31,72,31,213,31,232,31,221,31,226,31,21,31,133,31,9,31,106,31,146,31,243,31,138,31,138,30,199,31,28,31,114,31,114,30,114,29,114,28,114,27,114,26,81,31,138,31,102,31,86,31,8,31,28,31,34,31,186,31,38,31,146,31,79,31,121,31,121,30,155,31,157,31,157,30,30,31,30,30,30,29,139,31,87,31,179,31,117,31,117,30,117,29,232,31,120,31,54,31,54,30,62,31,216,31,251,31,215,31,215,30,215,29,64,31,237,31,189,31,255,31,25,31,87,31,163,31,114,31,91,31,91,30,35,31,2,31,2,30,121,31,172,31,172,30,117,31,117,30,185,31,11,31,53,31,130,31,253,31,62,31,183,31,183,30,179,31,128,31,128,30,249,31,207,31,42,31,14,31,14,30,1,31,57,31,214,31,78,31,98,31,98,30,134,31,94,31,53,31,80,31,80,30,80,29,163,31,193,31,13,31,13,30,179,31,131,31,223,31,28,31,95,31,251,31,164,31,164,30,152,31,139,31,14,31,14,30,215,31,63,31,63,30,220,31,220,30,220,29,129,31,73,31,102,31,172,31,36,31,141,31,225,31,244,31,252,31,206,31,42,31,58,31,120,31,72,31,219,31,163,31,52,31,52,30,235,31,56,31,56,30,56,31,56,30,56,29,134,31,189,31,105,31,56,31,218,31,180,31,4,31,249,31,185,31,240,31,240,30,226,31,95,31,46,31,38,31,129,31,129,30,149,31,149,30,186,31,134,31,134,30,145,31,88,31,231,31,184,31,216,31,216,30,4,31,4,30,4,29,59,31,48,31,45,31,169,31,198,31,123,31,123,30,123,29,123,28,197,31,204,31,225,31,159,31,205,31,205,30,252,31,187,31,127,31,83,31,110,31,231,31,168,31,242,31,212,31,229,31,229,30,68,31,91,31,91,30,136,31,132,31,132,30,121,31,23,31,250,31,250,30,164,31,188,31,188,30,164,31,164,30,164,29,121,31,133,31,51,31,177,31,185,31,1,31,113,31,153,31,225,31,30,31,162,31,166,31,166,30,166,29,244,31,128,31,2,31,58,31,58,30,207,31,172,31,172,30,12,31,237,31,64,31,64,30,76,31,212,31,105,31,88,31,73,31,244,31,59,31,9,31,122,31,73,31,74,31,24,31,52,31,58,31,118,31,118,30,139,31,139,30,232,31,138,31,218,31,157,31,107,31,191,31,119,31,64,31,64,30,64,29,211,31,133,31,92,31,177,31,177,30,163,31,100,31,100,30,135,31,69,31,117,31,53,31,141,31,114,31,138,31,138,30,71,31,116,31,29,31,22,31,22,30,12,31,209,31,11,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
