-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_174 is
end project_tb_174;

architecture project_tb_arch_174 of project_tb_174 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 977;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (176,0,85,0,75,0,109,0,42,0,19,0,7,0,0,0,47,0,110,0,252,0,142,0,56,0,200,0,161,0,16,0,0,0,183,0,190,0,103,0,117,0,165,0,173,0,76,0,218,0,58,0,55,0,178,0,20,0,30,0,253,0,39,0,38,0,253,0,155,0,0,0,0,0,124,0,153,0,78,0,205,0,129,0,0,0,0,0,0,0,0,0,69,0,95,0,125,0,175,0,0,0,20,0,74,0,0,0,94,0,0,0,18,0,55,0,238,0,0,0,115,0,188,0,121,0,227,0,143,0,137,0,0,0,9,0,235,0,2,0,188,0,55,0,174,0,106,0,145,0,13,0,232,0,164,0,118,0,226,0,162,0,63,0,44,0,0,0,214,0,0,0,228,0,60,0,0,0,207,0,179,0,0,0,160,0,218,0,139,0,182,0,0,0,184,0,168,0,251,0,131,0,0,0,137,0,83,0,96,0,182,0,249,0,189,0,44,0,0,0,0,0,244,0,53,0,145,0,0,0,149,0,206,0,88,0,0,0,137,0,0,0,0,0,34,0,186,0,107,0,123,0,175,0,110,0,158,0,179,0,181,0,0,0,157,0,0,0,241,0,222,0,50,0,81,0,0,0,241,0,78,0,86,0,0,0,157,0,1,0,0,0,236,0,51,0,200,0,18,0,98,0,230,0,130,0,190,0,63,0,0,0,248,0,33,0,0,0,0,0,0,0,39,0,0,0,116,0,246,0,68,0,88,0,0,0,7,0,92,0,169,0,211,0,50,0,150,0,25,0,0,0,175,0,0,0,91,0,7,0,159,0,189,0,63,0,0,0,0,0,206,0,34,0,8,0,88,0,181,0,148,0,179,0,176,0,97,0,117,0,71,0,0,0,194,0,155,0,25,0,130,0,161,0,0,0,165,0,109,0,0,0,196,0,74,0,0,0,139,0,167,0,162,0,255,0,221,0,102,0,166,0,0,0,112,0,145,0,49,0,187,0,171,0,156,0,176,0,96,0,0,0,235,0,243,0,218,0,136,0,33,0,240,0,205,0,0,0,0,0,92,0,158,0,71,0,0,0,235,0,0,0,0,0,111,0,26,0,203,0,0,0,164,0,151,0,149,0,88,0,130,0,64,0,201,0,0,0,15,0,120,0,134,0,0,0,10,0,140,0,209,0,0,0,227,0,75,0,127,0,0,0,0,0,134,0,0,0,95,0,211,0,138,0,59,0,103,0,243,0,209,0,0,0,32,0,244,0,154,0,0,0,0,0,234,0,222,0,235,0,0,0,15,0,43,0,64,0,164,0,0,0,0,0,190,0,107,0,0,0,250,0,39,0,0,0,0,0,179,0,75,0,77,0,50,0,129,0,0,0,69,0,51,0,2,0,0,0,0,0,66,0,79,0,78,0,0,0,178,0,232,0,0,0,0,0,218,0,154,0,185,0,0,0,62,0,133,0,0,0,122,0,33,0,79,0,0,0,0,0,185,0,106,0,130,0,200,0,125,0,79,0,86,0,112,0,42,0,47,0,0,0,0,0,190,0,239,0,86,0,220,0,1,0,0,0,0,0,143,0,155,0,0,0,0,0,207,0,138,0,46,0,68,0,101,0,0,0,5,0,0,0,126,0,155,0,40,0,102,0,3,0,26,0,42,0,92,0,120,0,112,0,94,0,0,0,46,0,126,0,38,0,128,0,75,0,78,0,128,0,77,0,0,0,220,0,3,0,217,0,173,0,138,0,121,0,82,0,120,0,202,0,142,0,208,0,91,0,83,0,159,0,162,0,165,0,227,0,244,0,161,0,71,0,97,0,117,0,243,0,137,0,0,0,59,0,160,0,0,0,38,0,121,0,0,0,0,0,55,0,0,0,208,0,228,0,0,0,0,0,0,0,33,0,0,0,35,0,102,0,6,0,239,0,51,0,74,0,207,0,58,0,74,0,225,0,0,0,74,0,129,0,46,0,18,0,208,0,109,0,8,0,165,0,64,0,110,0,0,0,128,0,227,0,108,0,234,0,0,0,147,0,162,0,36,0,0,0,222,0,60,0,29,0,0,0,40,0,0,0,155,0,83,0,195,0,77,0,0,0,187,0,0,0,167,0,168,0,195,0,173,0,42,0,235,0,233,0,246,0,104,0,0,0,57,0,0,0,58,0,67,0,0,0,86,0,195,0,173,0,121,0,147,0,178,0,238,0,6,0,111,0,136,0,224,0,0,0,216,0,0,0,96,0,0,0,98,0,215,0,89,0,213,0,147,0,1,0,38,0,0,0,156,0,19,0,189,0,19,0,0,0,43,0,10,0,41,0,66,0,11,0,175,0,179,0,162,0,39,0,0,0,0,0,242,0,73,0,0,0,245,0,176,0,140,0,53,0,147,0,236,0,0,0,184,0,108,0,0,0,152,0,31,0,141,0,13,0,86,0,209,0,0,0,0,0,152,0,42,0,94,0,163,0,0,0,97,0,167,0,235,0,207,0,173,0,0,0,93,0,156,0,68,0,49,0,0,0,71,0,145,0,238,0,185,0,19,0,78,0,81,0,91,0,172,0,156,0,0,0,5,0,91,0,129,0,193,0,238,0,0,0,235,0,251,0,25,0,211,0,255,0,92,0,22,0,57,0,118,0,166,0,27,0,38,0,224,0,187,0,217,0,4,0,0,0,153,0,133,0,188,0,74,0,0,0,129,0,20,0,184,0,162,0,4,0,214,0,186,0,0,0,182,0,0,0,187,0,104,0,0,0,69,0,99,0,147,0,33,0,230,0,227,0,160,0,245,0,0,0,150,0,243,0,59,0,0,0,2,0,209,0,217,0,0,0,4,0,179,0,216,0,0,0,83,0,72,0,210,0,103,0,7,0,99,0,205,0,243,0,95,0,0,0,205,0,67,0,43,0,244,0,216,0,102,0,81,0,134,0,23,0,0,0,156,0,163,0,79,0,197,0,76,0,162,0,157,0,151,0,0,0,43,0,255,0,239,0,237,0,248,0,0,0,243,0,175,0,72,0,148,0,0,0,0,0,20,0,133,0,211,0,125,0,133,0,194,0,44,0,121,0,0,0,0,0,186,0,10,0,0,0,240,0,105,0,244,0,0,0,136,0,17,0,203,0,0,0,24,0,120,0,22,0,0,0,138,0,159,0,227,0,17,0,4,0,0,0,178,0,248,0,223,0,227,0,5,0,106,0,0,0,36,0,201,0,175,0,227,0,240,0,99,0,16,0,0,0,53,0,221,0,76,0,151,0,0,0,14,0,59,0,115,0,139,0,108,0,169,0,2,0,70,0,252,0,36,0,42,0,105,0,151,0,158,0,83,0,101,0,0,0,79,0,0,0,0,0,176,0,94,0,187,0,37,0,0,0,181,0,208,0,0,0,255,0,0,0,16,0,137,0,250,0,136,0,147,0,222,0,72,0,43,0,172,0,252,0,65,0,139,0,153,0,0,0,78,0,112,0,0,0,246,0,0,0,188,0,132,0,171,0,12,0,200,0,250,0,215,0,0,0,0,0,50,0,127,0,0,0,0,0,0,0,0,0,122,0,0,0,138,0,217,0,212,0,201,0,0,0,4,0,125,0,79,0,152,0,243,0,129,0,171,0,230,0,0,0,0,0,0,0,0,0,97,0,200,0,189,0,42,0,76,0,110,0,18,0,84,0,22,0,95,0,222,0,0,0,0,0,0,0,90,0,81,0,0,0,62,0,253,0,107,0,100,0,0,0,4,0,10,0,211,0,242,0,72,0,19,0,215,0,205,0,0,0,234,0,153,0,181,0,0,0,154,0,176,0,99,0,76,0,0,0,199,0,47,0,85,0,172,0,78,0,221,0,0,0,72,0,0,0,133,0,179,0,203,0,0,0,128,0,153,0,151,0,151,0,136,0,184,0,35,0,0,0,133,0,0,0,231,0,0,0,0,0,40,0,0,0,116,0,0,0,0,0,143,0,188,0,232,0,0,0,250,0,68,0,28,0,86,0,0,0,148,0,118,0,30,0,142,0,144,0,202,0,190,0,0,0,0,0,125,0,0,0,0,0,97,0,159,0,0,0,6,0,160,0,119,0,0,0,60,0,239,0,169,0,130,0,191,0,0,0,20,0,108,0,190,0,196,0,27,0,51,0,216,0,144,0,216,0,95,0,138,0,42,0,48,0,206,0,18,0,0,0,90,0,111,0,62,0,190,0,0,0,217,0,0,0,46,0,88,0,142,0,78,0,228,0,246,0,43,0,39,0,0,0,206,0,167,0,0,0,213,0,76,0,0,0,134,0,240,0,0,0,189,0,164,0,65,0,161,0,0,0,51,0,0,0,0,0,181,0,23,0,0,0,146,0,130,0,224,0,129,0,36,0,57,0,217,0,43,0,121,0,0,0,225,0,99,0,0,0);
signal scenario_full  : scenario_type := (176,31,85,31,75,31,109,31,42,31,19,31,7,31,7,30,47,31,110,31,252,31,142,31,56,31,200,31,161,31,16,31,16,30,183,31,190,31,103,31,117,31,165,31,173,31,76,31,218,31,58,31,55,31,178,31,20,31,30,31,253,31,39,31,38,31,253,31,155,31,155,30,155,29,124,31,153,31,78,31,205,31,129,31,129,30,129,29,129,28,129,27,69,31,95,31,125,31,175,31,175,30,20,31,74,31,74,30,94,31,94,30,18,31,55,31,238,31,238,30,115,31,188,31,121,31,227,31,143,31,137,31,137,30,9,31,235,31,2,31,188,31,55,31,174,31,106,31,145,31,13,31,232,31,164,31,118,31,226,31,162,31,63,31,44,31,44,30,214,31,214,30,228,31,60,31,60,30,207,31,179,31,179,30,160,31,218,31,139,31,182,31,182,30,184,31,168,31,251,31,131,31,131,30,137,31,83,31,96,31,182,31,249,31,189,31,44,31,44,30,44,29,244,31,53,31,145,31,145,30,149,31,206,31,88,31,88,30,137,31,137,30,137,29,34,31,186,31,107,31,123,31,175,31,110,31,158,31,179,31,181,31,181,30,157,31,157,30,241,31,222,31,50,31,81,31,81,30,241,31,78,31,86,31,86,30,157,31,1,31,1,30,236,31,51,31,200,31,18,31,98,31,230,31,130,31,190,31,63,31,63,30,248,31,33,31,33,30,33,29,33,28,39,31,39,30,116,31,246,31,68,31,88,31,88,30,7,31,92,31,169,31,211,31,50,31,150,31,25,31,25,30,175,31,175,30,91,31,7,31,159,31,189,31,63,31,63,30,63,29,206,31,34,31,8,31,88,31,181,31,148,31,179,31,176,31,97,31,117,31,71,31,71,30,194,31,155,31,25,31,130,31,161,31,161,30,165,31,109,31,109,30,196,31,74,31,74,30,139,31,167,31,162,31,255,31,221,31,102,31,166,31,166,30,112,31,145,31,49,31,187,31,171,31,156,31,176,31,96,31,96,30,235,31,243,31,218,31,136,31,33,31,240,31,205,31,205,30,205,29,92,31,158,31,71,31,71,30,235,31,235,30,235,29,111,31,26,31,203,31,203,30,164,31,151,31,149,31,88,31,130,31,64,31,201,31,201,30,15,31,120,31,134,31,134,30,10,31,140,31,209,31,209,30,227,31,75,31,127,31,127,30,127,29,134,31,134,30,95,31,211,31,138,31,59,31,103,31,243,31,209,31,209,30,32,31,244,31,154,31,154,30,154,29,234,31,222,31,235,31,235,30,15,31,43,31,64,31,164,31,164,30,164,29,190,31,107,31,107,30,250,31,39,31,39,30,39,29,179,31,75,31,77,31,50,31,129,31,129,30,69,31,51,31,2,31,2,30,2,29,66,31,79,31,78,31,78,30,178,31,232,31,232,30,232,29,218,31,154,31,185,31,185,30,62,31,133,31,133,30,122,31,33,31,79,31,79,30,79,29,185,31,106,31,130,31,200,31,125,31,79,31,86,31,112,31,42,31,47,31,47,30,47,29,190,31,239,31,86,31,220,31,1,31,1,30,1,29,143,31,155,31,155,30,155,29,207,31,138,31,46,31,68,31,101,31,101,30,5,31,5,30,126,31,155,31,40,31,102,31,3,31,26,31,42,31,92,31,120,31,112,31,94,31,94,30,46,31,126,31,38,31,128,31,75,31,78,31,128,31,77,31,77,30,220,31,3,31,217,31,173,31,138,31,121,31,82,31,120,31,202,31,142,31,208,31,91,31,83,31,159,31,162,31,165,31,227,31,244,31,161,31,71,31,97,31,117,31,243,31,137,31,137,30,59,31,160,31,160,30,38,31,121,31,121,30,121,29,55,31,55,30,208,31,228,31,228,30,228,29,228,28,33,31,33,30,35,31,102,31,6,31,239,31,51,31,74,31,207,31,58,31,74,31,225,31,225,30,74,31,129,31,46,31,18,31,208,31,109,31,8,31,165,31,64,31,110,31,110,30,128,31,227,31,108,31,234,31,234,30,147,31,162,31,36,31,36,30,222,31,60,31,29,31,29,30,40,31,40,30,155,31,83,31,195,31,77,31,77,30,187,31,187,30,167,31,168,31,195,31,173,31,42,31,235,31,233,31,246,31,104,31,104,30,57,31,57,30,58,31,67,31,67,30,86,31,195,31,173,31,121,31,147,31,178,31,238,31,6,31,111,31,136,31,224,31,224,30,216,31,216,30,96,31,96,30,98,31,215,31,89,31,213,31,147,31,1,31,38,31,38,30,156,31,19,31,189,31,19,31,19,30,43,31,10,31,41,31,66,31,11,31,175,31,179,31,162,31,39,31,39,30,39,29,242,31,73,31,73,30,245,31,176,31,140,31,53,31,147,31,236,31,236,30,184,31,108,31,108,30,152,31,31,31,141,31,13,31,86,31,209,31,209,30,209,29,152,31,42,31,94,31,163,31,163,30,97,31,167,31,235,31,207,31,173,31,173,30,93,31,156,31,68,31,49,31,49,30,71,31,145,31,238,31,185,31,19,31,78,31,81,31,91,31,172,31,156,31,156,30,5,31,91,31,129,31,193,31,238,31,238,30,235,31,251,31,25,31,211,31,255,31,92,31,22,31,57,31,118,31,166,31,27,31,38,31,224,31,187,31,217,31,4,31,4,30,153,31,133,31,188,31,74,31,74,30,129,31,20,31,184,31,162,31,4,31,214,31,186,31,186,30,182,31,182,30,187,31,104,31,104,30,69,31,99,31,147,31,33,31,230,31,227,31,160,31,245,31,245,30,150,31,243,31,59,31,59,30,2,31,209,31,217,31,217,30,4,31,179,31,216,31,216,30,83,31,72,31,210,31,103,31,7,31,99,31,205,31,243,31,95,31,95,30,205,31,67,31,43,31,244,31,216,31,102,31,81,31,134,31,23,31,23,30,156,31,163,31,79,31,197,31,76,31,162,31,157,31,151,31,151,30,43,31,255,31,239,31,237,31,248,31,248,30,243,31,175,31,72,31,148,31,148,30,148,29,20,31,133,31,211,31,125,31,133,31,194,31,44,31,121,31,121,30,121,29,186,31,10,31,10,30,240,31,105,31,244,31,244,30,136,31,17,31,203,31,203,30,24,31,120,31,22,31,22,30,138,31,159,31,227,31,17,31,4,31,4,30,178,31,248,31,223,31,227,31,5,31,106,31,106,30,36,31,201,31,175,31,227,31,240,31,99,31,16,31,16,30,53,31,221,31,76,31,151,31,151,30,14,31,59,31,115,31,139,31,108,31,169,31,2,31,70,31,252,31,36,31,42,31,105,31,151,31,158,31,83,31,101,31,101,30,79,31,79,30,79,29,176,31,94,31,187,31,37,31,37,30,181,31,208,31,208,30,255,31,255,30,16,31,137,31,250,31,136,31,147,31,222,31,72,31,43,31,172,31,252,31,65,31,139,31,153,31,153,30,78,31,112,31,112,30,246,31,246,30,188,31,132,31,171,31,12,31,200,31,250,31,215,31,215,30,215,29,50,31,127,31,127,30,127,29,127,28,127,27,122,31,122,30,138,31,217,31,212,31,201,31,201,30,4,31,125,31,79,31,152,31,243,31,129,31,171,31,230,31,230,30,230,29,230,28,230,27,97,31,200,31,189,31,42,31,76,31,110,31,18,31,84,31,22,31,95,31,222,31,222,30,222,29,222,28,90,31,81,31,81,30,62,31,253,31,107,31,100,31,100,30,4,31,10,31,211,31,242,31,72,31,19,31,215,31,205,31,205,30,234,31,153,31,181,31,181,30,154,31,176,31,99,31,76,31,76,30,199,31,47,31,85,31,172,31,78,31,221,31,221,30,72,31,72,30,133,31,179,31,203,31,203,30,128,31,153,31,151,31,151,31,136,31,184,31,35,31,35,30,133,31,133,30,231,31,231,30,231,29,40,31,40,30,116,31,116,30,116,29,143,31,188,31,232,31,232,30,250,31,68,31,28,31,86,31,86,30,148,31,118,31,30,31,142,31,144,31,202,31,190,31,190,30,190,29,125,31,125,30,125,29,97,31,159,31,159,30,6,31,160,31,119,31,119,30,60,31,239,31,169,31,130,31,191,31,191,30,20,31,108,31,190,31,196,31,27,31,51,31,216,31,144,31,216,31,95,31,138,31,42,31,48,31,206,31,18,31,18,30,90,31,111,31,62,31,190,31,190,30,217,31,217,30,46,31,88,31,142,31,78,31,228,31,246,31,43,31,39,31,39,30,206,31,167,31,167,30,213,31,76,31,76,30,134,31,240,31,240,30,189,31,164,31,65,31,161,31,161,30,51,31,51,30,51,29,181,31,23,31,23,30,146,31,130,31,224,31,129,31,36,31,57,31,217,31,43,31,121,31,121,30,225,31,99,31,99,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
