-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 859;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (31,0,86,0,146,0,188,0,90,0,156,0,40,0,0,0,111,0,145,0,0,0,113,0,223,0,206,0,78,0,249,0,76,0,76,0,118,0,0,0,183,0,54,0,88,0,233,0,87,0,209,0,39,0,149,0,252,0,137,0,217,0,64,0,118,0,89,0,159,0,194,0,238,0,232,0,117,0,34,0,188,0,172,0,116,0,146,0,20,0,178,0,58,0,171,0,0,0,37,0,131,0,219,0,0,0,71,0,251,0,124,0,0,0,225,0,237,0,40,0,179,0,76,0,177,0,61,0,109,0,48,0,35,0,71,0,82,0,0,0,0,0,187,0,176,0,36,0,0,0,146,0,111,0,172,0,123,0,0,0,169,0,190,0,204,0,203,0,0,0,0,0,206,0,255,0,1,0,205,0,222,0,58,0,249,0,187,0,77,0,31,0,148,0,126,0,144,0,12,0,22,0,162,0,0,0,203,0,174,0,43,0,145,0,53,0,83,0,227,0,21,0,115,0,35,0,171,0,116,0,248,0,0,0,149,0,254,0,127,0,200,0,0,0,46,0,105,0,0,0,200,0,148,0,108,0,203,0,121,0,202,0,0,0,8,0,176,0,133,0,35,0,249,0,247,0,219,0,177,0,192,0,134,0,218,0,204,0,0,0,0,0,0,0,147,0,18,0,244,0,202,0,171,0,235,0,69,0,0,0,50,0,160,0,169,0,0,0,25,0,0,0,54,0,153,0,202,0,122,0,100,0,0,0,0,0,202,0,135,0,141,0,156,0,92,0,0,0,0,0,98,0,23,0,216,0,98,0,104,0,0,0,211,0,159,0,92,0,193,0,32,0,197,0,158,0,195,0,47,0,144,0,47,0,0,0,0,0,0,0,0,0,226,0,167,0,56,0,233,0,41,0,236,0,0,0,0,0,3,0,203,0,180,0,91,0,49,0,32,0,48,0,33,0,11,0,71,0,158,0,111,0,14,0,133,0,138,0,88,0,134,0,199,0,116,0,0,0,140,0,127,0,0,0,0,0,72,0,162,0,158,0,188,0,253,0,70,0,97,0,136,0,75,0,35,0,51,0,140,0,144,0,91,0,105,0,188,0,84,0,219,0,38,0,77,0,105,0,0,0,40,0,43,0,144,0,46,0,107,0,184,0,37,0,13,0,92,0,247,0,63,0,0,0,78,0,41,0,79,0,100,0,156,0,0,0,130,0,0,0,160,0,56,0,220,0,248,0,150,0,195,0,0,0,0,0,121,0,92,0,254,0,0,0,227,0,134,0,177,0,167,0,68,0,208,0,0,0,29,0,108,0,106,0,78,0,188,0,30,0,105,0,0,0,205,0,168,0,0,0,0,0,42,0,186,0,33,0,0,0,182,0,189,0,44,0,0,0,0,0,109,0,0,0,0,0,9,0,144,0,89,0,123,0,146,0,0,0,228,0,189,0,22,0,142,0,122,0,198,0,108,0,0,0,131,0,112,0,153,0,251,0,201,0,163,0,102,0,0,0,138,0,144,0,98,0,0,0,5,0,138,0,141,0,130,0,40,0,211,0,0,0,111,0,14,0,249,0,144,0,112,0,0,0,6,0,18,0,121,0,144,0,190,0,9,0,0,0,32,0,27,0,103,0,62,0,127,0,17,0,27,0,255,0,53,0,102,0,100,0,85,0,53,0,0,0,67,0,0,0,207,0,56,0,0,0,30,0,152,0,0,0,0,0,85,0,201,0,54,0,48,0,235,0,46,0,175,0,180,0,180,0,0,0,82,0,0,0,45,0,25,0,0,0,200,0,253,0,138,0,106,0,81,0,182,0,1,0,99,0,222,0,124,0,222,0,24,0,190,0,112,0,5,0,106,0,0,0,238,0,146,0,178,0,0,0,253,0,182,0,220,0,0,0,87,0,227,0,0,0,182,0,130,0,244,0,244,0,0,0,68,0,47,0,34,0,91,0,116,0,0,0,249,0,202,0,159,0,0,0,216,0,63,0,196,0,244,0,192,0,140,0,170,0,123,0,174,0,0,0,0,0,129,0,194,0,165,0,0,0,122,0,4,0,161,0,86,0,230,0,0,0,68,0,71,0,103,0,63,0,0,0,152,0,126,0,55,0,0,0,0,0,177,0,228,0,0,0,217,0,239,0,20,0,200,0,36,0,132,0,206,0,87,0,208,0,170,0,0,0,193,0,101,0,162,0,0,0,191,0,0,0,0,0,163,0,97,0,112,0,69,0,67,0,119,0,222,0,112,0,156,0,124,0,0,0,14,0,134,0,166,0,0,0,204,0,90,0,54,0,165,0,101,0,60,0,106,0,71,0,217,0,0,0,33,0,0,0,43,0,46,0,62,0,197,0,0,0,223,0,107,0,0,0,18,0,0,0,0,0,163,0,246,0,69,0,77,0,201,0,132,0,168,0,133,0,106,0,87,0,52,0,0,0,154,0,143,0,112,0,0,0,5,0,0,0,251,0,76,0,44,0,3,0,122,0,114,0,153,0,0,0,84,0,153,0,0,0,59,0,0,0,210,0,0,0,212,0,19,0,0,0,134,0,107,0,179,0,134,0,146,0,29,0,32,0,53,0,0,0,96,0,0,0,0,0,0,0,154,0,71,0,18,0,89,0,98,0,0,0,216,0,128,0,41,0,189,0,141,0,115,0,202,0,55,0,103,0,52,0,0,0,85,0,239,0,117,0,122,0,167,0,114,0,185,0,89,0,232,0,6,0,0,0,20,0,102,0,102,0,0,0,228,0,40,0,208,0,224,0,58,0,230,0,0,0,209,0,184,0,86,0,171,0,216,0,188,0,79,0,45,0,0,0,101,0,164,0,0,0,3,0,19,0,167,0,254,0,113,0,210,0,166,0,222,0,113,0,43,0,0,0,0,0,0,0,142,0,0,0,0,0,4,0,162,0,0,0,0,0,0,0,0,0,0,0,114,0,58,0,154,0,217,0,132,0,139,0,140,0,185,0,69,0,0,0,0,0,214,0,209,0,77,0,70,0,95,0,58,0,248,0,145,0,149,0,63,0,0,0,20,0,23,0,53,0,212,0,150,0,91,0,23,0,183,0,27,0,0,0,0,0,77,0,0,0,131,0,0,0,79,0,24,0,108,0,123,0,247,0,0,0,8,0,114,0,75,0,118,0,12,0,0,0,209,0,0,0,116,0,206,0,147,0,0,0,226,0,163,0,219,0,11,0,64,0,128,0,202,0,41,0,224,0,12,0,40,0,68,0,180,0,203,0,160,0,91,0,34,0,45,0,0,0,163,0,183,0,34,0,218,0,115,0,220,0,0,0,70,0,0,0,117,0,0,0,0,0,139,0,238,0,3,0,196,0,0,0,64,0,0,0,90,0,0,0,99,0,131,0,128,0,16,0,156,0,0,0,0,0,51,0,51,0,255,0,97,0,70,0,46,0,233,0,88,0,0,0,242,0,126,0,248,0,251,0,2,0,62,0,145,0,242,0,86,0,138,0,10,0,194,0,203,0,15,0,12,0,5,0,23,0,212,0,205,0,0,0,94,0,18,0,62,0,0,0,43,0,117,0,0,0,0,0,0,0,0,0,0,0,25,0,25,0,47,0,0,0,0,0,127,0,0,0,21,0,164,0,226,0,246,0,204,0,178,0,26,0,60,0,0,0,216,0,155,0,116,0,0,0,161,0,0,0,27,0,126,0,218,0,53,0,0,0,0,0,154,0,77,0,192,0,229,0,0,0,221,0,173,0,0,0,0,0,153,0,133,0,166,0,195,0,84,0,0,0,0,0,190,0,126,0,97,0,81,0,14,0,48,0,171,0,155,0,218,0,0,0,1,0,0,0,88,0,242,0,181,0,68,0,61,0,238,0,176,0,230,0);
signal scenario_full  : scenario_type := (31,31,86,31,146,31,188,31,90,31,156,31,40,31,40,30,111,31,145,31,145,30,113,31,223,31,206,31,78,31,249,31,76,31,76,31,118,31,118,30,183,31,54,31,88,31,233,31,87,31,209,31,39,31,149,31,252,31,137,31,217,31,64,31,118,31,89,31,159,31,194,31,238,31,232,31,117,31,34,31,188,31,172,31,116,31,146,31,20,31,178,31,58,31,171,31,171,30,37,31,131,31,219,31,219,30,71,31,251,31,124,31,124,30,225,31,237,31,40,31,179,31,76,31,177,31,61,31,109,31,48,31,35,31,71,31,82,31,82,30,82,29,187,31,176,31,36,31,36,30,146,31,111,31,172,31,123,31,123,30,169,31,190,31,204,31,203,31,203,30,203,29,206,31,255,31,1,31,205,31,222,31,58,31,249,31,187,31,77,31,31,31,148,31,126,31,144,31,12,31,22,31,162,31,162,30,203,31,174,31,43,31,145,31,53,31,83,31,227,31,21,31,115,31,35,31,171,31,116,31,248,31,248,30,149,31,254,31,127,31,200,31,200,30,46,31,105,31,105,30,200,31,148,31,108,31,203,31,121,31,202,31,202,30,8,31,176,31,133,31,35,31,249,31,247,31,219,31,177,31,192,31,134,31,218,31,204,31,204,30,204,29,204,28,147,31,18,31,244,31,202,31,171,31,235,31,69,31,69,30,50,31,160,31,169,31,169,30,25,31,25,30,54,31,153,31,202,31,122,31,100,31,100,30,100,29,202,31,135,31,141,31,156,31,92,31,92,30,92,29,98,31,23,31,216,31,98,31,104,31,104,30,211,31,159,31,92,31,193,31,32,31,197,31,158,31,195,31,47,31,144,31,47,31,47,30,47,29,47,28,47,27,226,31,167,31,56,31,233,31,41,31,236,31,236,30,236,29,3,31,203,31,180,31,91,31,49,31,32,31,48,31,33,31,11,31,71,31,158,31,111,31,14,31,133,31,138,31,88,31,134,31,199,31,116,31,116,30,140,31,127,31,127,30,127,29,72,31,162,31,158,31,188,31,253,31,70,31,97,31,136,31,75,31,35,31,51,31,140,31,144,31,91,31,105,31,188,31,84,31,219,31,38,31,77,31,105,31,105,30,40,31,43,31,144,31,46,31,107,31,184,31,37,31,13,31,92,31,247,31,63,31,63,30,78,31,41,31,79,31,100,31,156,31,156,30,130,31,130,30,160,31,56,31,220,31,248,31,150,31,195,31,195,30,195,29,121,31,92,31,254,31,254,30,227,31,134,31,177,31,167,31,68,31,208,31,208,30,29,31,108,31,106,31,78,31,188,31,30,31,105,31,105,30,205,31,168,31,168,30,168,29,42,31,186,31,33,31,33,30,182,31,189,31,44,31,44,30,44,29,109,31,109,30,109,29,9,31,144,31,89,31,123,31,146,31,146,30,228,31,189,31,22,31,142,31,122,31,198,31,108,31,108,30,131,31,112,31,153,31,251,31,201,31,163,31,102,31,102,30,138,31,144,31,98,31,98,30,5,31,138,31,141,31,130,31,40,31,211,31,211,30,111,31,14,31,249,31,144,31,112,31,112,30,6,31,18,31,121,31,144,31,190,31,9,31,9,30,32,31,27,31,103,31,62,31,127,31,17,31,27,31,255,31,53,31,102,31,100,31,85,31,53,31,53,30,67,31,67,30,207,31,56,31,56,30,30,31,152,31,152,30,152,29,85,31,201,31,54,31,48,31,235,31,46,31,175,31,180,31,180,31,180,30,82,31,82,30,45,31,25,31,25,30,200,31,253,31,138,31,106,31,81,31,182,31,1,31,99,31,222,31,124,31,222,31,24,31,190,31,112,31,5,31,106,31,106,30,238,31,146,31,178,31,178,30,253,31,182,31,220,31,220,30,87,31,227,31,227,30,182,31,130,31,244,31,244,31,244,30,68,31,47,31,34,31,91,31,116,31,116,30,249,31,202,31,159,31,159,30,216,31,63,31,196,31,244,31,192,31,140,31,170,31,123,31,174,31,174,30,174,29,129,31,194,31,165,31,165,30,122,31,4,31,161,31,86,31,230,31,230,30,68,31,71,31,103,31,63,31,63,30,152,31,126,31,55,31,55,30,55,29,177,31,228,31,228,30,217,31,239,31,20,31,200,31,36,31,132,31,206,31,87,31,208,31,170,31,170,30,193,31,101,31,162,31,162,30,191,31,191,30,191,29,163,31,97,31,112,31,69,31,67,31,119,31,222,31,112,31,156,31,124,31,124,30,14,31,134,31,166,31,166,30,204,31,90,31,54,31,165,31,101,31,60,31,106,31,71,31,217,31,217,30,33,31,33,30,43,31,46,31,62,31,197,31,197,30,223,31,107,31,107,30,18,31,18,30,18,29,163,31,246,31,69,31,77,31,201,31,132,31,168,31,133,31,106,31,87,31,52,31,52,30,154,31,143,31,112,31,112,30,5,31,5,30,251,31,76,31,44,31,3,31,122,31,114,31,153,31,153,30,84,31,153,31,153,30,59,31,59,30,210,31,210,30,212,31,19,31,19,30,134,31,107,31,179,31,134,31,146,31,29,31,32,31,53,31,53,30,96,31,96,30,96,29,96,28,154,31,71,31,18,31,89,31,98,31,98,30,216,31,128,31,41,31,189,31,141,31,115,31,202,31,55,31,103,31,52,31,52,30,85,31,239,31,117,31,122,31,167,31,114,31,185,31,89,31,232,31,6,31,6,30,20,31,102,31,102,31,102,30,228,31,40,31,208,31,224,31,58,31,230,31,230,30,209,31,184,31,86,31,171,31,216,31,188,31,79,31,45,31,45,30,101,31,164,31,164,30,3,31,19,31,167,31,254,31,113,31,210,31,166,31,222,31,113,31,43,31,43,30,43,29,43,28,142,31,142,30,142,29,4,31,162,31,162,30,162,29,162,28,162,27,162,26,114,31,58,31,154,31,217,31,132,31,139,31,140,31,185,31,69,31,69,30,69,29,214,31,209,31,77,31,70,31,95,31,58,31,248,31,145,31,149,31,63,31,63,30,20,31,23,31,53,31,212,31,150,31,91,31,23,31,183,31,27,31,27,30,27,29,77,31,77,30,131,31,131,30,79,31,24,31,108,31,123,31,247,31,247,30,8,31,114,31,75,31,118,31,12,31,12,30,209,31,209,30,116,31,206,31,147,31,147,30,226,31,163,31,219,31,11,31,64,31,128,31,202,31,41,31,224,31,12,31,40,31,68,31,180,31,203,31,160,31,91,31,34,31,45,31,45,30,163,31,183,31,34,31,218,31,115,31,220,31,220,30,70,31,70,30,117,31,117,30,117,29,139,31,238,31,3,31,196,31,196,30,64,31,64,30,90,31,90,30,99,31,131,31,128,31,16,31,156,31,156,30,156,29,51,31,51,31,255,31,97,31,70,31,46,31,233,31,88,31,88,30,242,31,126,31,248,31,251,31,2,31,62,31,145,31,242,31,86,31,138,31,10,31,194,31,203,31,15,31,12,31,5,31,23,31,212,31,205,31,205,30,94,31,18,31,62,31,62,30,43,31,117,31,117,30,117,29,117,28,117,27,117,26,25,31,25,31,47,31,47,30,47,29,127,31,127,30,21,31,164,31,226,31,246,31,204,31,178,31,26,31,60,31,60,30,216,31,155,31,116,31,116,30,161,31,161,30,27,31,126,31,218,31,53,31,53,30,53,29,154,31,77,31,192,31,229,31,229,30,221,31,173,31,173,30,173,29,153,31,133,31,166,31,195,31,84,31,84,30,84,29,190,31,126,31,97,31,81,31,14,31,48,31,171,31,155,31,218,31,218,30,1,31,1,30,88,31,242,31,181,31,68,31,61,31,238,31,176,31,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
