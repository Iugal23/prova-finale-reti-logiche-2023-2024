-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 317;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (184,0,241,0,58,0,161,0,162,0,58,0,75,0,73,0,44,0,189,0,0,0,25,0,56,0,181,0,167,0,135,0,0,0,114,0,78,0,122,0,175,0,202,0,229,0,148,0,218,0,0,0,230,0,0,0,167,0,226,0,0,0,4,0,233,0,0,0,0,0,20,0,33,0,0,0,223,0,6,0,0,0,130,0,106,0,239,0,181,0,123,0,109,0,60,0,76,0,0,0,117,0,169,0,221,0,84,0,0,0,90,0,0,0,63,0,135,0,215,0,159,0,217,0,176,0,187,0,0,0,160,0,215,0,47,0,8,0,102,0,0,0,140,0,115,0,23,0,44,0,72,0,101,0,0,0,167,0,56,0,226,0,213,0,132,0,0,0,241,0,0,0,7,0,10,0,14,0,6,0,0,0,202,0,172,0,140,0,38,0,240,0,203,0,165,0,166,0,66,0,116,0,175,0,57,0,88,0,115,0,45,0,128,0,87,0,0,0,188,0,60,0,47,0,39,0,31,0,127,0,131,0,0,0,150,0,190,0,53,0,196,0,6,0,102,0,79,0,234,0,234,0,223,0,163,0,0,0,0,0,188,0,76,0,195,0,175,0,228,0,0,0,0,0,30,0,11,0,0,0,106,0,245,0,166,0,84,0,207,0,179,0,0,0,209,0,199,0,91,0,0,0,140,0,0,0,53,0,202,0,0,0,190,0,132,0,225,0,0,0,54,0,103,0,248,0,76,0,0,0,48,0,0,0,96,0,106,0,163,0,84,0,48,0,0,0,0,0,145,0,110,0,58,0,207,0,26,0,194,0,225,0,153,0,143,0,79,0,142,0,188,0,173,0,60,0,0,0,0,0,203,0,161,0,43,0,139,0,229,0,170,0,161,0,181,0,107,0,159,0,70,0,10,0,188,0,0,0,12,0,158,0,22,0,205,0,0,0,177,0,0,0,0,0,0,0,216,0,178,0,0,0,244,0,235,0,251,0,5,0,132,0,221,0,135,0,242,0,46,0,155,0,174,0,0,0,97,0,187,0,116,0,218,0,205,0,25,0,225,0,31,0,124,0,237,0,188,0,68,0,245,0,56,0,61,0,113,0,173,0,0,0,127,0,187,0,218,0,0,0,125,0,115,0,0,0,156,0,0,0,0,0,199,0,0,0,3,0,240,0,159,0,91,0,50,0,0,0,246,0,218,0,168,0,141,0,0,0,175,0,208,0,243,0,214,0,106,0,238,0,0,0,118,0,143,0,237,0,171,0,139,0,243,0,185,0,57,0,64,0,95,0,0,0,176,0,39,0,0,0,106,0,110,0,0,0,49,0,0,0,21,0,0,0,96,0,71,0,0,0,124,0,42,0,111,0,141,0,144,0,175,0,159,0,48,0,11,0,95,0,90,0,199,0,0,0,23,0,33,0,0,0,230,0);
signal scenario_full  : scenario_type := (184,31,241,31,58,31,161,31,162,31,58,31,75,31,73,31,44,31,189,31,189,30,25,31,56,31,181,31,167,31,135,31,135,30,114,31,78,31,122,31,175,31,202,31,229,31,148,31,218,31,218,30,230,31,230,30,167,31,226,31,226,30,4,31,233,31,233,30,233,29,20,31,33,31,33,30,223,31,6,31,6,30,130,31,106,31,239,31,181,31,123,31,109,31,60,31,76,31,76,30,117,31,169,31,221,31,84,31,84,30,90,31,90,30,63,31,135,31,215,31,159,31,217,31,176,31,187,31,187,30,160,31,215,31,47,31,8,31,102,31,102,30,140,31,115,31,23,31,44,31,72,31,101,31,101,30,167,31,56,31,226,31,213,31,132,31,132,30,241,31,241,30,7,31,10,31,14,31,6,31,6,30,202,31,172,31,140,31,38,31,240,31,203,31,165,31,166,31,66,31,116,31,175,31,57,31,88,31,115,31,45,31,128,31,87,31,87,30,188,31,60,31,47,31,39,31,31,31,127,31,131,31,131,30,150,31,190,31,53,31,196,31,6,31,102,31,79,31,234,31,234,31,223,31,163,31,163,30,163,29,188,31,76,31,195,31,175,31,228,31,228,30,228,29,30,31,11,31,11,30,106,31,245,31,166,31,84,31,207,31,179,31,179,30,209,31,199,31,91,31,91,30,140,31,140,30,53,31,202,31,202,30,190,31,132,31,225,31,225,30,54,31,103,31,248,31,76,31,76,30,48,31,48,30,96,31,106,31,163,31,84,31,48,31,48,30,48,29,145,31,110,31,58,31,207,31,26,31,194,31,225,31,153,31,143,31,79,31,142,31,188,31,173,31,60,31,60,30,60,29,203,31,161,31,43,31,139,31,229,31,170,31,161,31,181,31,107,31,159,31,70,31,10,31,188,31,188,30,12,31,158,31,22,31,205,31,205,30,177,31,177,30,177,29,177,28,216,31,178,31,178,30,244,31,235,31,251,31,5,31,132,31,221,31,135,31,242,31,46,31,155,31,174,31,174,30,97,31,187,31,116,31,218,31,205,31,25,31,225,31,31,31,124,31,237,31,188,31,68,31,245,31,56,31,61,31,113,31,173,31,173,30,127,31,187,31,218,31,218,30,125,31,115,31,115,30,156,31,156,30,156,29,199,31,199,30,3,31,240,31,159,31,91,31,50,31,50,30,246,31,218,31,168,31,141,31,141,30,175,31,208,31,243,31,214,31,106,31,238,31,238,30,118,31,143,31,237,31,171,31,139,31,243,31,185,31,57,31,64,31,95,31,95,30,176,31,39,31,39,30,106,31,110,31,110,30,49,31,49,30,21,31,21,30,96,31,71,31,71,30,124,31,42,31,111,31,141,31,144,31,175,31,159,31,48,31,11,31,95,31,90,31,199,31,199,30,23,31,33,31,33,30,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
