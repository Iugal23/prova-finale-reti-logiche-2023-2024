-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_956 is
end project_tb_956;

architecture project_tb_arch_956 of project_tb_956 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 743;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (108,0,168,0,0,0,228,0,168,0,129,0,0,0,0,0,0,0,0,0,0,0,26,0,142,0,27,0,0,0,116,0,251,0,102,0,13,0,7,0,166,0,241,0,43,0,250,0,0,0,0,0,158,0,186,0,103,0,192,0,0,0,66,0,0,0,128,0,170,0,22,0,44,0,59,0,222,0,123,0,136,0,0,0,34,0,8,0,251,0,0,0,0,0,213,0,148,0,113,0,31,0,153,0,116,0,253,0,27,0,171,0,126,0,164,0,0,0,165,0,0,0,149,0,238,0,77,0,229,0,162,0,66,0,0,0,146,0,148,0,70,0,33,0,154,0,76,0,0,0,60,0,126,0,125,0,106,0,213,0,0,0,72,0,108,0,28,0,58,0,0,0,95,0,71,0,178,0,137,0,178,0,1,0,0,0,0,0,55,0,94,0,120,0,192,0,72,0,67,0,79,0,105,0,0,0,121,0,112,0,0,0,218,0,165,0,0,0,142,0,236,0,18,0,57,0,105,0,214,0,240,0,197,0,0,0,209,0,122,0,127,0,0,0,196,0,31,0,36,0,176,0,116,0,29,0,0,0,0,0,70,0,76,0,0,0,101,0,187,0,73,0,197,0,144,0,126,0,0,0,222,0,251,0,49,0,124,0,47,0,0,0,0,0,0,0,221,0,143,0,0,0,0,0,128,0,120,0,100,0,44,0,99,0,83,0,58,0,117,0,0,0,70,0,113,0,0,0,0,0,105,0,0,0,173,0,33,0,0,0,178,0,183,0,239,0,53,0,125,0,14,0,0,0,206,0,95,0,104,0,115,0,66,0,146,0,110,0,185,0,66,0,180,0,38,0,159,0,105,0,0,0,0,0,245,0,90,0,0,0,120,0,0,0,93,0,223,0,15,0,25,0,61,0,117,0,157,0,106,0,0,0,0,0,156,0,226,0,65,0,0,0,0,0,0,0,226,0,192,0,0,0,221,0,138,0,118,0,98,0,119,0,37,0,0,0,53,0,24,0,3,0,138,0,43,0,190,0,9,0,24,0,250,0,91,0,101,0,92,0,1,0,0,0,159,0,148,0,155,0,92,0,40,0,93,0,231,0,158,0,104,0,64,0,0,0,103,0,250,0,112,0,160,0,227,0,227,0,133,0,45,0,0,0,147,0,146,0,5,0,0,0,0,0,195,0,121,0,75,0,0,0,244,0,182,0,15,0,142,0,140,0,190,0,4,0,201,0,121,0,115,0,246,0,0,0,102,0,104,0,232,0,0,0,99,0,120,0,0,0,0,0,194,0,199,0,0,0,94,0,238,0,190,0,101,0,91,0,0,0,18,0,42,0,251,0,248,0,254,0,218,0,0,0,0,0,179,0,0,0,39,0,112,0,127,0,38,0,242,0,114,0,86,0,108,0,249,0,0,0,178,0,96,0,84,0,0,0,98,0,158,0,0,0,0,0,0,0,192,0,21,0,201,0,92,0,206,0,0,0,0,0,55,0,0,0,137,0,221,0,55,0,70,0,88,0,77,0,0,0,177,0,207,0,155,0,0,0,23,0,238,0,0,0,0,0,71,0,231,0,0,0,140,0,197,0,161,0,35,0,151,0,0,0,161,0,0,0,62,0,132,0,19,0,193,0,0,0,0,0,120,0,164,0,146,0,211,0,0,0,109,0,162,0,0,0,0,0,144,0,48,0,25,0,2,0,206,0,109,0,89,0,0,0,0,0,123,0,79,0,0,0,6,0,212,0,150,0,130,0,48,0,15,0,101,0,0,0,0,0,140,0,248,0,176,0,34,0,147,0,0,0,240,0,164,0,0,0,70,0,91,0,228,0,0,0,101,0,143,0,170,0,81,0,177,0,8,0,5,0,49,0,111,0,151,0,33,0,104,0,0,0,23,0,207,0,153,0,254,0,148,0,77,0,21,0,0,0,66,0,122,0,243,0,72,0,79,0,248,0,0,0,143,0,220,0,252,0,205,0,0,0,118,0,0,0,0,0,123,0,47,0,103,0,114,0,245,0,17,0,223,0,76,0,228,0,193,0,48,0,37,0,144,0,161,0,7,0,57,0,81,0,0,0,209,0,139,0,166,0,0,0,58,0,166,0,6,0,230,0,204,0,237,0,63,0,119,0,97,0,29,0,33,0,166,0,131,0,4,0,255,0,67,0,154,0,230,0,99,0,12,0,62,0,249,0,175,0,55,0,10,0,17,0,53,0,55,0,163,0,0,0,171,0,89,0,112,0,138,0,0,0,165,0,0,0,107,0,18,0,135,0,227,0,229,0,225,0,158,0,212,0,146,0,24,0,0,0,7,0,107,0,0,0,9,0,28,0,234,0,150,0,223,0,50,0,179,0,119,0,237,0,223,0,210,0,211,0,0,0,221,0,0,0,0,0,0,0,47,0,0,0,123,0,121,0,0,0,158,0,0,0,150,0,71,0,6,0,0,0,120,0,187,0,144,0,150,0,94,0,0,0,0,0,166,0,0,0,0,0,26,0,0,0,10,0,92,0,0,0,0,0,0,0,216,0,0,0,248,0,0,0,255,0,162,0,214,0,137,0,0,0,229,0,0,0,176,0,251,0,45,0,0,0,242,0,0,0,0,0,49,0,235,0,196,0,171,0,175,0,204,0,250,0,58,0,0,0,211,0,192,0,62,0,109,0,140,0,38,0,247,0,0,0,0,0,117,0,250,0,56,0,232,0,227,0,169,0,136,0,12,0,58,0,87,0,79,0,119,0,0,0,150,0,0,0,129,0,32,0,159,0,0,0,44,0,183,0,78,0,0,0,236,0,0,0,217,0,226,0,89,0,144,0,118,0,177,0,0,0,63,0,181,0,46,0,24,0,172,0,0,0,186,0,115,0,4,0,56,0,164,0,252,0,235,0,0,0,111,0,0,0,109,0,161,0,63,0,0,0,211,0,50,0,0,0,252,0,219,0,0,0,0,0,0,0,85,0,139,0,148,0,74,0,202,0,198,0,13,0,175,0,165,0,50,0,166,0,236,0,78,0,67,0,167,0,134,0,175,0,114,0,129,0,14,0,188,0,0,0,86,0,0,0,55,0,137,0,169,0,86,0,230,0,64,0,213,0,108,0,0,0,30,0,45,0,195,0,142,0,60,0,125,0,174,0,169,0,113,0,138,0,143,0,228,0,0,0,66,0,44,0,32,0,0,0,7,0,153,0,223,0,48,0,0,0,0,0,126,0,138,0,58,0,0,0,75,0,0,0,0,0,98,0,61,0,191,0,30,0,149,0,34,0,0,0,97,0,229,0,0,0,23,0,0,0,0,0,0,0,216,0,204,0,0,0,220,0,208,0,246,0,96,0,108,0);
signal scenario_full  : scenario_type := (108,31,168,31,168,30,228,31,168,31,129,31,129,30,129,29,129,28,129,27,129,26,26,31,142,31,27,31,27,30,116,31,251,31,102,31,13,31,7,31,166,31,241,31,43,31,250,31,250,30,250,29,158,31,186,31,103,31,192,31,192,30,66,31,66,30,128,31,170,31,22,31,44,31,59,31,222,31,123,31,136,31,136,30,34,31,8,31,251,31,251,30,251,29,213,31,148,31,113,31,31,31,153,31,116,31,253,31,27,31,171,31,126,31,164,31,164,30,165,31,165,30,149,31,238,31,77,31,229,31,162,31,66,31,66,30,146,31,148,31,70,31,33,31,154,31,76,31,76,30,60,31,126,31,125,31,106,31,213,31,213,30,72,31,108,31,28,31,58,31,58,30,95,31,71,31,178,31,137,31,178,31,1,31,1,30,1,29,55,31,94,31,120,31,192,31,72,31,67,31,79,31,105,31,105,30,121,31,112,31,112,30,218,31,165,31,165,30,142,31,236,31,18,31,57,31,105,31,214,31,240,31,197,31,197,30,209,31,122,31,127,31,127,30,196,31,31,31,36,31,176,31,116,31,29,31,29,30,29,29,70,31,76,31,76,30,101,31,187,31,73,31,197,31,144,31,126,31,126,30,222,31,251,31,49,31,124,31,47,31,47,30,47,29,47,28,221,31,143,31,143,30,143,29,128,31,120,31,100,31,44,31,99,31,83,31,58,31,117,31,117,30,70,31,113,31,113,30,113,29,105,31,105,30,173,31,33,31,33,30,178,31,183,31,239,31,53,31,125,31,14,31,14,30,206,31,95,31,104,31,115,31,66,31,146,31,110,31,185,31,66,31,180,31,38,31,159,31,105,31,105,30,105,29,245,31,90,31,90,30,120,31,120,30,93,31,223,31,15,31,25,31,61,31,117,31,157,31,106,31,106,30,106,29,156,31,226,31,65,31,65,30,65,29,65,28,226,31,192,31,192,30,221,31,138,31,118,31,98,31,119,31,37,31,37,30,53,31,24,31,3,31,138,31,43,31,190,31,9,31,24,31,250,31,91,31,101,31,92,31,1,31,1,30,159,31,148,31,155,31,92,31,40,31,93,31,231,31,158,31,104,31,64,31,64,30,103,31,250,31,112,31,160,31,227,31,227,31,133,31,45,31,45,30,147,31,146,31,5,31,5,30,5,29,195,31,121,31,75,31,75,30,244,31,182,31,15,31,142,31,140,31,190,31,4,31,201,31,121,31,115,31,246,31,246,30,102,31,104,31,232,31,232,30,99,31,120,31,120,30,120,29,194,31,199,31,199,30,94,31,238,31,190,31,101,31,91,31,91,30,18,31,42,31,251,31,248,31,254,31,218,31,218,30,218,29,179,31,179,30,39,31,112,31,127,31,38,31,242,31,114,31,86,31,108,31,249,31,249,30,178,31,96,31,84,31,84,30,98,31,158,31,158,30,158,29,158,28,192,31,21,31,201,31,92,31,206,31,206,30,206,29,55,31,55,30,137,31,221,31,55,31,70,31,88,31,77,31,77,30,177,31,207,31,155,31,155,30,23,31,238,31,238,30,238,29,71,31,231,31,231,30,140,31,197,31,161,31,35,31,151,31,151,30,161,31,161,30,62,31,132,31,19,31,193,31,193,30,193,29,120,31,164,31,146,31,211,31,211,30,109,31,162,31,162,30,162,29,144,31,48,31,25,31,2,31,206,31,109,31,89,31,89,30,89,29,123,31,79,31,79,30,6,31,212,31,150,31,130,31,48,31,15,31,101,31,101,30,101,29,140,31,248,31,176,31,34,31,147,31,147,30,240,31,164,31,164,30,70,31,91,31,228,31,228,30,101,31,143,31,170,31,81,31,177,31,8,31,5,31,49,31,111,31,151,31,33,31,104,31,104,30,23,31,207,31,153,31,254,31,148,31,77,31,21,31,21,30,66,31,122,31,243,31,72,31,79,31,248,31,248,30,143,31,220,31,252,31,205,31,205,30,118,31,118,30,118,29,123,31,47,31,103,31,114,31,245,31,17,31,223,31,76,31,228,31,193,31,48,31,37,31,144,31,161,31,7,31,57,31,81,31,81,30,209,31,139,31,166,31,166,30,58,31,166,31,6,31,230,31,204,31,237,31,63,31,119,31,97,31,29,31,33,31,166,31,131,31,4,31,255,31,67,31,154,31,230,31,99,31,12,31,62,31,249,31,175,31,55,31,10,31,17,31,53,31,55,31,163,31,163,30,171,31,89,31,112,31,138,31,138,30,165,31,165,30,107,31,18,31,135,31,227,31,229,31,225,31,158,31,212,31,146,31,24,31,24,30,7,31,107,31,107,30,9,31,28,31,234,31,150,31,223,31,50,31,179,31,119,31,237,31,223,31,210,31,211,31,211,30,221,31,221,30,221,29,221,28,47,31,47,30,123,31,121,31,121,30,158,31,158,30,150,31,71,31,6,31,6,30,120,31,187,31,144,31,150,31,94,31,94,30,94,29,166,31,166,30,166,29,26,31,26,30,10,31,92,31,92,30,92,29,92,28,216,31,216,30,248,31,248,30,255,31,162,31,214,31,137,31,137,30,229,31,229,30,176,31,251,31,45,31,45,30,242,31,242,30,242,29,49,31,235,31,196,31,171,31,175,31,204,31,250,31,58,31,58,30,211,31,192,31,62,31,109,31,140,31,38,31,247,31,247,30,247,29,117,31,250,31,56,31,232,31,227,31,169,31,136,31,12,31,58,31,87,31,79,31,119,31,119,30,150,31,150,30,129,31,32,31,159,31,159,30,44,31,183,31,78,31,78,30,236,31,236,30,217,31,226,31,89,31,144,31,118,31,177,31,177,30,63,31,181,31,46,31,24,31,172,31,172,30,186,31,115,31,4,31,56,31,164,31,252,31,235,31,235,30,111,31,111,30,109,31,161,31,63,31,63,30,211,31,50,31,50,30,252,31,219,31,219,30,219,29,219,28,85,31,139,31,148,31,74,31,202,31,198,31,13,31,175,31,165,31,50,31,166,31,236,31,78,31,67,31,167,31,134,31,175,31,114,31,129,31,14,31,188,31,188,30,86,31,86,30,55,31,137,31,169,31,86,31,230,31,64,31,213,31,108,31,108,30,30,31,45,31,195,31,142,31,60,31,125,31,174,31,169,31,113,31,138,31,143,31,228,31,228,30,66,31,44,31,32,31,32,30,7,31,153,31,223,31,48,31,48,30,48,29,126,31,138,31,58,31,58,30,75,31,75,30,75,29,98,31,61,31,191,31,30,31,149,31,34,31,34,30,97,31,229,31,229,30,23,31,23,30,23,29,23,28,216,31,204,31,204,30,220,31,208,31,246,31,96,31,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
