-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 381;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (211,0,0,0,0,0,173,0,87,0,162,0,252,0,52,0,42,0,184,0,0,0,7,0,59,0,69,0,126,0,92,0,216,0,21,0,123,0,177,0,0,0,204,0,50,0,16,0,241,0,0,0,208,0,124,0,222,0,0,0,248,0,0,0,98,0,0,0,11,0,0,0,98,0,0,0,0,0,0,0,152,0,0,0,135,0,213,0,104,0,81,0,101,0,0,0,0,0,17,0,22,0,0,0,0,0,30,0,208,0,175,0,83,0,63,0,182,0,254,0,78,0,17,0,129,0,241,0,0,0,197,0,0,0,82,0,138,0,98,0,188,0,105,0,50,0,215,0,249,0,0,0,25,0,62,0,127,0,52,0,26,0,202,0,192,0,55,0,243,0,114,0,222,0,172,0,194,0,64,0,102,0,0,0,125,0,66,0,0,0,160,0,235,0,24,0,0,0,126,0,219,0,56,0,19,0,247,0,0,0,209,0,117,0,164,0,0,0,199,0,169,0,46,0,5,0,116,0,192,0,0,0,242,0,224,0,240,0,157,0,113,0,0,0,79,0,184,0,61,0,143,0,79,0,42,0,230,0,8,0,38,0,16,0,0,0,123,0,0,0,191,0,122,0,184,0,0,0,31,0,117,0,147,0,184,0,0,0,231,0,51,0,234,0,243,0,240,0,12,0,60,0,241,0,239,0,0,0,0,0,32,0,233,0,50,0,28,0,112,0,0,0,59,0,0,0,183,0,156,0,0,0,33,0,116,0,253,0,64,0,54,0,164,0,136,0,174,0,36,0,219,0,220,0,117,0,107,0,0,0,85,0,103,0,0,0,121,0,63,0,211,0,46,0,140,0,28,0,240,0,66,0,139,0,53,0,139,0,252,0,189,0,48,0,0,0,113,0,85,0,185,0,73,0,35,0,77,0,212,0,47,0,179,0,167,0,9,0,238,0,102,0,172,0,95,0,9,0,15,0,24,0,224,0,221,0,0,0,158,0,75,0,31,0,187,0,122,0,162,0,111,0,0,0,140,0,68,0,145,0,64,0,8,0,88,0,0,0,16,0,111,0,0,0,218,0,0,0,0,0,0,0,36,0,234,0,190,0,237,0,0,0,0,0,10,0,0,0,32,0,7,0,148,0,168,0,25,0,0,0,0,0,144,0,0,0,13,0,0,0,177,0,0,0,86,0,77,0,224,0,253,0,50,0,233,0,5,0,186,0,204,0,229,0,29,0,22,0,19,0,95,0,203,0,59,0,222,0,159,0,121,0,0,0,38,0,163,0,42,0,34,0,0,0,151,0,230,0,91,0,220,0,6,0,26,0,251,0,0,0,94,0,0,0,0,0,119,0,153,0,0,0,43,0,29,0,212,0,0,0,121,0,97,0,0,0,179,0,234,0,83,0,236,0,119,0,194,0,81,0,148,0,162,0,253,0,0,0,19,0,40,0,150,0,147,0,114,0,49,0,8,0,90,0,16,0,243,0,73,0,210,0,138,0,81,0,252,0,125,0,120,0,160,0,0,0,24,0,36,0,190,0,0,0,16,0,104,0,77,0,61,0,113,0,83,0,137,0,0,0,236,0,219,0,209,0,32,0,25,0,0,0,0,0,0,0,111,0,195,0,48,0,162,0,216,0,85,0,184,0,0,0,26,0,50,0,49,0,236,0,102,0,132,0,215,0,49,0,181,0,0,0,179,0,204,0,0,0,5,0,0,0);
signal scenario_full  : scenario_type := (211,31,211,30,211,29,173,31,87,31,162,31,252,31,52,31,42,31,184,31,184,30,7,31,59,31,69,31,126,31,92,31,216,31,21,31,123,31,177,31,177,30,204,31,50,31,16,31,241,31,241,30,208,31,124,31,222,31,222,30,248,31,248,30,98,31,98,30,11,31,11,30,98,31,98,30,98,29,98,28,152,31,152,30,135,31,213,31,104,31,81,31,101,31,101,30,101,29,17,31,22,31,22,30,22,29,30,31,208,31,175,31,83,31,63,31,182,31,254,31,78,31,17,31,129,31,241,31,241,30,197,31,197,30,82,31,138,31,98,31,188,31,105,31,50,31,215,31,249,31,249,30,25,31,62,31,127,31,52,31,26,31,202,31,192,31,55,31,243,31,114,31,222,31,172,31,194,31,64,31,102,31,102,30,125,31,66,31,66,30,160,31,235,31,24,31,24,30,126,31,219,31,56,31,19,31,247,31,247,30,209,31,117,31,164,31,164,30,199,31,169,31,46,31,5,31,116,31,192,31,192,30,242,31,224,31,240,31,157,31,113,31,113,30,79,31,184,31,61,31,143,31,79,31,42,31,230,31,8,31,38,31,16,31,16,30,123,31,123,30,191,31,122,31,184,31,184,30,31,31,117,31,147,31,184,31,184,30,231,31,51,31,234,31,243,31,240,31,12,31,60,31,241,31,239,31,239,30,239,29,32,31,233,31,50,31,28,31,112,31,112,30,59,31,59,30,183,31,156,31,156,30,33,31,116,31,253,31,64,31,54,31,164,31,136,31,174,31,36,31,219,31,220,31,117,31,107,31,107,30,85,31,103,31,103,30,121,31,63,31,211,31,46,31,140,31,28,31,240,31,66,31,139,31,53,31,139,31,252,31,189,31,48,31,48,30,113,31,85,31,185,31,73,31,35,31,77,31,212,31,47,31,179,31,167,31,9,31,238,31,102,31,172,31,95,31,9,31,15,31,24,31,224,31,221,31,221,30,158,31,75,31,31,31,187,31,122,31,162,31,111,31,111,30,140,31,68,31,145,31,64,31,8,31,88,31,88,30,16,31,111,31,111,30,218,31,218,30,218,29,218,28,36,31,234,31,190,31,237,31,237,30,237,29,10,31,10,30,32,31,7,31,148,31,168,31,25,31,25,30,25,29,144,31,144,30,13,31,13,30,177,31,177,30,86,31,77,31,224,31,253,31,50,31,233,31,5,31,186,31,204,31,229,31,29,31,22,31,19,31,95,31,203,31,59,31,222,31,159,31,121,31,121,30,38,31,163,31,42,31,34,31,34,30,151,31,230,31,91,31,220,31,6,31,26,31,251,31,251,30,94,31,94,30,94,29,119,31,153,31,153,30,43,31,29,31,212,31,212,30,121,31,97,31,97,30,179,31,234,31,83,31,236,31,119,31,194,31,81,31,148,31,162,31,253,31,253,30,19,31,40,31,150,31,147,31,114,31,49,31,8,31,90,31,16,31,243,31,73,31,210,31,138,31,81,31,252,31,125,31,120,31,160,31,160,30,24,31,36,31,190,31,190,30,16,31,104,31,77,31,61,31,113,31,83,31,137,31,137,30,236,31,219,31,209,31,32,31,25,31,25,30,25,29,25,28,111,31,195,31,48,31,162,31,216,31,85,31,184,31,184,30,26,31,50,31,49,31,236,31,102,31,132,31,215,31,49,31,181,31,181,30,179,31,204,31,204,30,5,31,5,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
