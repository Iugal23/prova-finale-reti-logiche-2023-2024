-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 875;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (120,0,0,0,44,0,158,0,92,0,0,0,194,0,215,0,140,0,93,0,0,0,0,0,154,0,168,0,223,0,38,0,78,0,0,0,0,0,125,0,84,0,105,0,0,0,150,0,131,0,0,0,45,0,202,0,96,0,65,0,69,0,0,0,241,0,193,0,169,0,0,0,41,0,134,0,34,0,238,0,115,0,211,0,240,0,184,0,0,0,21,0,90,0,242,0,0,0,58,0,11,0,0,0,0,0,0,0,99,0,126,0,16,0,39,0,243,0,16,0,133,0,16,0,0,0,0,0,154,0,24,0,12,0,196,0,128,0,229,0,96,0,128,0,90,0,162,0,0,0,43,0,71,0,17,0,206,0,12,0,240,0,4,0,19,0,230,0,225,0,81,0,37,0,164,0,232,0,208,0,203,0,145,0,85,0,119,0,0,0,152,0,0,0,62,0,168,0,116,0,47,0,102,0,119,0,60,0,135,0,0,0,198,0,88,0,0,0,109,0,6,0,240,0,54,0,25,0,139,0,0,0,0,0,21,0,51,0,0,0,19,0,0,0,0,0,98,0,219,0,0,0,0,0,0,0,186,0,24,0,112,0,136,0,0,0,0,0,132,0,254,0,216,0,0,0,17,0,215,0,169,0,116,0,106,0,158,0,5,0,54,0,0,0,82,0,122,0,57,0,170,0,27,0,28,0,0,0,211,0,81,0,189,0,227,0,21,0,223,0,192,0,130,0,162,0,45,0,0,0,0,0,23,0,181,0,53,0,23,0,0,0,25,0,0,0,4,0,10,0,36,0,131,0,201,0,235,0,31,0,29,0,200,0,0,0,0,0,44,0,152,0,209,0,237,0,221,0,173,0,193,0,55,0,66,0,0,0,123,0,131,0,175,0,97,0,0,0,169,0,187,0,147,0,0,0,101,0,61,0,0,0,168,0,218,0,0,0,0,0,170,0,252,0,230,0,0,0,123,0,236,0,175,0,113,0,1,0,187,0,149,0,51,0,29,0,84,0,223,0,0,0,8,0,156,0,51,0,19,0,102,0,134,0,116,0,223,0,8,0,115,0,69,0,32,0,240,0,203,0,104,0,145,0,124,0,185,0,236,0,198,0,186,0,15,0,0,0,143,0,179,0,0,0,45,0,188,0,92,0,0,0,202,0,8,0,1,0,186,0,39,0,174,0,199,0,167,0,0,0,89,0,247,0,106,0,229,0,71,0,6,0,111,0,81,0,88,0,124,0,173,0,205,0,193,0,250,0,233,0,193,0,0,0,0,0,200,0,97,0,91,0,0,0,232,0,25,0,0,0,27,0,75,0,196,0,0,0,203,0,174,0,217,0,107,0,181,0,21,0,180,0,70,0,106,0,19,0,152,0,119,0,163,0,149,0,68,0,171,0,0,0,0,0,173,0,41,0,178,0,97,0,60,0,45,0,190,0,0,0,57,0,216,0,236,0,20,0,66,0,76,0,50,0,101,0,0,0,0,0,0,0,189,0,9,0,126,0,169,0,98,0,0,0,0,0,212,0,184,0,50,0,247,0,111,0,173,0,172,0,187,0,186,0,180,0,236,0,215,0,152,0,30,0,0,0,220,0,45,0,246,0,145,0,246,0,144,0,91,0,0,0,134,0,54,0,170,0,0,0,0,0,48,0,0,0,0,0,159,0,32,0,186,0,207,0,32,0,197,0,88,0,0,0,32,0,150,0,180,0,86,0,242,0,194,0,0,0,78,0,5,0,0,0,118,0,101,0,158,0,0,0,39,0,146,0,189,0,209,0,130,0,111,0,204,0,241,0,215,0,168,0,0,0,0,0,0,0,103,0,0,0,16,0,90,0,201,0,192,0,15,0,41,0,78,0,220,0,177,0,106,0,57,0,24,0,147,0,72,0,233,0,215,0,222,0,166,0,144,0,0,0,112,0,4,0,137,0,0,0,195,0,139,0,93,0,93,0,102,0,0,0,44,0,2,0,210,0,0,0,0,0,0,0,25,0,192,0,248,0,37,0,0,0,231,0,220,0,32,0,199,0,227,0,131,0,211,0,20,0,39,0,249,0,196,0,116,0,213,0,80,0,128,0,240,0,0,0,176,0,200,0,0,0,180,0,170,0,199,0,57,0,177,0,8,0,202,0,174,0,170,0,214,0,243,0,148,0,51,0,0,0,189,0,207,0,161,0,103,0,190,0,242,0,216,0,220,0,28,0,65,0,21,0,207,0,123,0,0,0,0,0,197,0,44,0,68,0,163,0,95,0,149,0,250,0,63,0,177,0,215,0,16,0,73,0,68,0,120,0,54,0,101,0,250,0,248,0,12,0,154,0,0,0,7,0,0,0,24,0,60,0,212,0,219,0,214,0,60,0,165,0,210,0,0,0,0,0,23,0,89,0,154,0,0,0,25,0,218,0,134,0,226,0,212,0,185,0,0,0,26,0,96,0,174,0,0,0,0,0,185,0,170,0,185,0,58,0,149,0,217,0,2,0,132,0,44,0,245,0,0,0,210,0,209,0,131,0,245,0,0,0,149,0,144,0,0,0,43,0,156,0,182,0,250,0,82,0,245,0,175,0,0,0,126,0,182,0,98,0,0,0,109,0,56,0,140,0,190,0,35,0,4,0,38,0,209,0,212,0,86,0,175,0,191,0,205,0,109,0,180,0,178,0,210,0,224,0,198,0,37,0,138,0,101,0,211,0,155,0,0,0,36,0,15,0,118,0,0,0,236,0,101,0,188,0,80,0,0,0,75,0,75,0,147,0,46,0,204,0,252,0,187,0,130,0,0,0,42,0,0,0,135,0,38,0,143,0,0,0,4,0,0,0,186,0,0,0,183,0,83,0,78,0,0,0,240,0,230,0,248,0,0,0,58,0,245,0,142,0,190,0,138,0,137,0,235,0,219,0,148,0,56,0,0,0,151,0,17,0,48,0,103,0,123,0,234,0,242,0,74,0,0,0,84,0,0,0,135,0,0,0,254,0,0,0,188,0,0,0,18,0,40,0,253,0,198,0,106,0,167,0,241,0,84,0,177,0,194,0,108,0,0,0,22,0,53,0,204,0,0,0,109,0,0,0,124,0,249,0,103,0,203,0,244,0,161,0,38,0,0,0,171,0,53,0,66,0,188,0,57,0,242,0,125,0,0,0,0,0,208,0,0,0,153,0,108,0,0,0,221,0,91,0,15,0,205,0,53,0,115,0,13,0,42,0,228,0,250,0,154,0,0,0,0,0,243,0,248,0,0,0,119,0,226,0,239,0,117,0,206,0,0,0,158,0,242,0,46,0,0,0,0,0,84,0,0,0,59,0,133,0,195,0,251,0,174,0,0,0,200,0,91,0,186,0,0,0,0,0,0,0,220,0,133,0,74,0,207,0,162,0,70,0,249,0,3,0,124,0,144,0,0,0,46,0,63,0,58,0,145,0,230,0,22,0,43,0,214,0,14,0,154,0,119,0,241,0,254,0,69,0,208,0,132,0,0,0,42,0,0,0,0,0,205,0,219,0,0,0,136,0,89,0,0,0,62,0,249,0,242,0,0,0,115,0,117,0,173,0,177,0,148,0,231,0,123,0,141,0,229,0,30,0,37,0,0,0,100,0,230,0,23,0,0,0,0,0,0,0,98,0,210,0,184,0,41,0,46,0,59,0,79,0,0,0,104,0,77,0,115,0,0,0,91,0,157,0,0,0,167,0,29,0,87,0,140,0,92,0,0,0,0,0,32,0,105,0,100,0,0,0,246,0,111,0,103,0,114,0,0,0,177,0,60,0,139,0,0,0,128,0,89,0,71,0,44,0,0,0,245,0,74,0,106,0,55,0,114,0,52,0,0,0,119,0,0,0,31,0,166,0,139,0,254,0,122,0,95,0,64,0,20,0,232,0,0,0,103,0,99,0,0,0,37,0,69,0,84,0,42,0,9,0,102,0,0,0,236,0);
signal scenario_full  : scenario_type := (120,31,120,30,44,31,158,31,92,31,92,30,194,31,215,31,140,31,93,31,93,30,93,29,154,31,168,31,223,31,38,31,78,31,78,30,78,29,125,31,84,31,105,31,105,30,150,31,131,31,131,30,45,31,202,31,96,31,65,31,69,31,69,30,241,31,193,31,169,31,169,30,41,31,134,31,34,31,238,31,115,31,211,31,240,31,184,31,184,30,21,31,90,31,242,31,242,30,58,31,11,31,11,30,11,29,11,28,99,31,126,31,16,31,39,31,243,31,16,31,133,31,16,31,16,30,16,29,154,31,24,31,12,31,196,31,128,31,229,31,96,31,128,31,90,31,162,31,162,30,43,31,71,31,17,31,206,31,12,31,240,31,4,31,19,31,230,31,225,31,81,31,37,31,164,31,232,31,208,31,203,31,145,31,85,31,119,31,119,30,152,31,152,30,62,31,168,31,116,31,47,31,102,31,119,31,60,31,135,31,135,30,198,31,88,31,88,30,109,31,6,31,240,31,54,31,25,31,139,31,139,30,139,29,21,31,51,31,51,30,19,31,19,30,19,29,98,31,219,31,219,30,219,29,219,28,186,31,24,31,112,31,136,31,136,30,136,29,132,31,254,31,216,31,216,30,17,31,215,31,169,31,116,31,106,31,158,31,5,31,54,31,54,30,82,31,122,31,57,31,170,31,27,31,28,31,28,30,211,31,81,31,189,31,227,31,21,31,223,31,192,31,130,31,162,31,45,31,45,30,45,29,23,31,181,31,53,31,23,31,23,30,25,31,25,30,4,31,10,31,36,31,131,31,201,31,235,31,31,31,29,31,200,31,200,30,200,29,44,31,152,31,209,31,237,31,221,31,173,31,193,31,55,31,66,31,66,30,123,31,131,31,175,31,97,31,97,30,169,31,187,31,147,31,147,30,101,31,61,31,61,30,168,31,218,31,218,30,218,29,170,31,252,31,230,31,230,30,123,31,236,31,175,31,113,31,1,31,187,31,149,31,51,31,29,31,84,31,223,31,223,30,8,31,156,31,51,31,19,31,102,31,134,31,116,31,223,31,8,31,115,31,69,31,32,31,240,31,203,31,104,31,145,31,124,31,185,31,236,31,198,31,186,31,15,31,15,30,143,31,179,31,179,30,45,31,188,31,92,31,92,30,202,31,8,31,1,31,186,31,39,31,174,31,199,31,167,31,167,30,89,31,247,31,106,31,229,31,71,31,6,31,111,31,81,31,88,31,124,31,173,31,205,31,193,31,250,31,233,31,193,31,193,30,193,29,200,31,97,31,91,31,91,30,232,31,25,31,25,30,27,31,75,31,196,31,196,30,203,31,174,31,217,31,107,31,181,31,21,31,180,31,70,31,106,31,19,31,152,31,119,31,163,31,149,31,68,31,171,31,171,30,171,29,173,31,41,31,178,31,97,31,60,31,45,31,190,31,190,30,57,31,216,31,236,31,20,31,66,31,76,31,50,31,101,31,101,30,101,29,101,28,189,31,9,31,126,31,169,31,98,31,98,30,98,29,212,31,184,31,50,31,247,31,111,31,173,31,172,31,187,31,186,31,180,31,236,31,215,31,152,31,30,31,30,30,220,31,45,31,246,31,145,31,246,31,144,31,91,31,91,30,134,31,54,31,170,31,170,30,170,29,48,31,48,30,48,29,159,31,32,31,186,31,207,31,32,31,197,31,88,31,88,30,32,31,150,31,180,31,86,31,242,31,194,31,194,30,78,31,5,31,5,30,118,31,101,31,158,31,158,30,39,31,146,31,189,31,209,31,130,31,111,31,204,31,241,31,215,31,168,31,168,30,168,29,168,28,103,31,103,30,16,31,90,31,201,31,192,31,15,31,41,31,78,31,220,31,177,31,106,31,57,31,24,31,147,31,72,31,233,31,215,31,222,31,166,31,144,31,144,30,112,31,4,31,137,31,137,30,195,31,139,31,93,31,93,31,102,31,102,30,44,31,2,31,210,31,210,30,210,29,210,28,25,31,192,31,248,31,37,31,37,30,231,31,220,31,32,31,199,31,227,31,131,31,211,31,20,31,39,31,249,31,196,31,116,31,213,31,80,31,128,31,240,31,240,30,176,31,200,31,200,30,180,31,170,31,199,31,57,31,177,31,8,31,202,31,174,31,170,31,214,31,243,31,148,31,51,31,51,30,189,31,207,31,161,31,103,31,190,31,242,31,216,31,220,31,28,31,65,31,21,31,207,31,123,31,123,30,123,29,197,31,44,31,68,31,163,31,95,31,149,31,250,31,63,31,177,31,215,31,16,31,73,31,68,31,120,31,54,31,101,31,250,31,248,31,12,31,154,31,154,30,7,31,7,30,24,31,60,31,212,31,219,31,214,31,60,31,165,31,210,31,210,30,210,29,23,31,89,31,154,31,154,30,25,31,218,31,134,31,226,31,212,31,185,31,185,30,26,31,96,31,174,31,174,30,174,29,185,31,170,31,185,31,58,31,149,31,217,31,2,31,132,31,44,31,245,31,245,30,210,31,209,31,131,31,245,31,245,30,149,31,144,31,144,30,43,31,156,31,182,31,250,31,82,31,245,31,175,31,175,30,126,31,182,31,98,31,98,30,109,31,56,31,140,31,190,31,35,31,4,31,38,31,209,31,212,31,86,31,175,31,191,31,205,31,109,31,180,31,178,31,210,31,224,31,198,31,37,31,138,31,101,31,211,31,155,31,155,30,36,31,15,31,118,31,118,30,236,31,101,31,188,31,80,31,80,30,75,31,75,31,147,31,46,31,204,31,252,31,187,31,130,31,130,30,42,31,42,30,135,31,38,31,143,31,143,30,4,31,4,30,186,31,186,30,183,31,83,31,78,31,78,30,240,31,230,31,248,31,248,30,58,31,245,31,142,31,190,31,138,31,137,31,235,31,219,31,148,31,56,31,56,30,151,31,17,31,48,31,103,31,123,31,234,31,242,31,74,31,74,30,84,31,84,30,135,31,135,30,254,31,254,30,188,31,188,30,18,31,40,31,253,31,198,31,106,31,167,31,241,31,84,31,177,31,194,31,108,31,108,30,22,31,53,31,204,31,204,30,109,31,109,30,124,31,249,31,103,31,203,31,244,31,161,31,38,31,38,30,171,31,53,31,66,31,188,31,57,31,242,31,125,31,125,30,125,29,208,31,208,30,153,31,108,31,108,30,221,31,91,31,15,31,205,31,53,31,115,31,13,31,42,31,228,31,250,31,154,31,154,30,154,29,243,31,248,31,248,30,119,31,226,31,239,31,117,31,206,31,206,30,158,31,242,31,46,31,46,30,46,29,84,31,84,30,59,31,133,31,195,31,251,31,174,31,174,30,200,31,91,31,186,31,186,30,186,29,186,28,220,31,133,31,74,31,207,31,162,31,70,31,249,31,3,31,124,31,144,31,144,30,46,31,63,31,58,31,145,31,230,31,22,31,43,31,214,31,14,31,154,31,119,31,241,31,254,31,69,31,208,31,132,31,132,30,42,31,42,30,42,29,205,31,219,31,219,30,136,31,89,31,89,30,62,31,249,31,242,31,242,30,115,31,117,31,173,31,177,31,148,31,231,31,123,31,141,31,229,31,30,31,37,31,37,30,100,31,230,31,23,31,23,30,23,29,23,28,98,31,210,31,184,31,41,31,46,31,59,31,79,31,79,30,104,31,77,31,115,31,115,30,91,31,157,31,157,30,167,31,29,31,87,31,140,31,92,31,92,30,92,29,32,31,105,31,100,31,100,30,246,31,111,31,103,31,114,31,114,30,177,31,60,31,139,31,139,30,128,31,89,31,71,31,44,31,44,30,245,31,74,31,106,31,55,31,114,31,52,31,52,30,119,31,119,30,31,31,166,31,139,31,254,31,122,31,95,31,64,31,20,31,232,31,232,30,103,31,99,31,99,30,37,31,69,31,84,31,42,31,9,31,102,31,102,30,236,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
