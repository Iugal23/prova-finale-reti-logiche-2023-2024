-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 971;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,27,0,41,0,0,0,183,0,221,0,162,0,96,0,119,0,249,0,5,0,123,0,14,0,162,0,0,0,180,0,175,0,64,0,172,0,156,0,0,0,0,0,57,0,82,0,211,0,173,0,155,0,74,0,0,0,216,0,48,0,253,0,112,0,47,0,0,0,206,0,93,0,93,0,196,0,219,0,62,0,207,0,232,0,69,0,97,0,18,0,189,0,40,0,205,0,209,0,8,0,133,0,116,0,8,0,73,0,34,0,220,0,166,0,120,0,0,0,225,0,176,0,0,0,171,0,113,0,61,0,243,0,96,0,0,0,117,0,28,0,42,0,0,0,215,0,0,0,148,0,61,0,212,0,104,0,100,0,240,0,0,0,173,0,236,0,185,0,199,0,119,0,0,0,219,0,194,0,232,0,0,0,234,0,92,0,78,0,157,0,60,0,242,0,172,0,0,0,0,0,0,0,247,0,64,0,40,0,0,0,0,0,113,0,102,0,228,0,95,0,63,0,149,0,132,0,153,0,0,0,0,0,235,0,45,0,91,0,100,0,239,0,0,0,156,0,67,0,25,0,254,0,141,0,242,0,10,0,79,0,84,0,0,0,10,0,94,0,74,0,170,0,104,0,182,0,7,0,148,0,235,0,0,0,23,0,0,0,87,0,106,0,0,0,16,0,185,0,95,0,122,0,0,0,60,0,115,0,178,0,0,0,198,0,224,0,58,0,0,0,0,0,152,0,127,0,160,0,0,0,0,0,236,0,193,0,175,0,203,0,194,0,69,0,182,0,0,0,33,0,33,0,227,0,211,0,89,0,74,0,0,0,0,0,59,0,104,0,140,0,15,0,42,0,250,0,211,0,0,0,121,0,104,0,165,0,114,0,0,0,247,0,48,0,240,0,230,0,131,0,41,0,217,0,77,0,197,0,16,0,181,0,211,0,253,0,178,0,75,0,0,0,0,0,229,0,173,0,185,0,134,0,247,0,165,0,0,0,165,0,0,0,0,0,52,0,13,0,190,0,0,0,51,0,101,0,219,0,171,0,0,0,104,0,202,0,227,0,18,0,141,0,75,0,0,0,210,0,52,0,0,0,157,0,172,0,220,0,139,0,255,0,0,0,0,0,0,0,215,0,170,0,78,0,178,0,29,0,0,0,23,0,0,0,131,0,151,0,0,0,0,0,0,0,147,0,0,0,252,0,71,0,0,0,184,0,0,0,196,0,154,0,12,0,12,0,0,0,8,0,238,0,61,0,107,0,0,0,93,0,194,0,0,0,12,0,173,0,226,0,0,0,0,0,0,0,89,0,172,0,196,0,186,0,64,0,41,0,211,0,176,0,161,0,0,0,59,0,126,0,79,0,43,0,158,0,78,0,119,0,24,0,0,0,0,0,209,0,143,0,171,0,12,0,158,0,234,0,125,0,220,0,0,0,250,0,38,0,215,0,89,0,54,0,134,0,212,0,147,0,0,0,145,0,208,0,200,0,30,0,0,0,0,0,171,0,21,0,168,0,0,0,0,0,193,0,248,0,220,0,0,0,239,0,183,0,0,0,109,0,126,0,226,0,126,0,0,0,226,0,101,0,0,0,207,0,232,0,104,0,120,0,112,0,0,0,171,0,217,0,137,0,133,0,78,0,103,0,97,0,121,0,71,0,177,0,9,0,43,0,208,0,223,0,0,0,187,0,151,0,101,0,107,0,0,0,3,0,61,0,0,0,31,0,180,0,95,0,0,0,130,0,238,0,0,0,0,0,111,0,210,0,223,0,0,0,153,0,5,0,211,0,0,0,156,0,17,0,231,0,198,0,84,0,170,0,141,0,177,0,29,0,161,0,150,0,206,0,160,0,154,0,0,0,154,0,142,0,252,0,157,0,217,0,24,0,62,0,254,0,7,0,167,0,195,0,210,0,63,0,109,0,251,0,212,0,91,0,208,0,223,0,240,0,178,0,180,0,226,0,92,0,0,0,69,0,121,0,0,0,136,0,115,0,129,0,73,0,163,0,0,0,159,0,0,0,39,0,192,0,65,0,125,0,158,0,97,0,0,0,146,0,176,0,45,0,4,0,101,0,244,0,40,0,89,0,133,0,0,0,0,0,235,0,0,0,0,0,107,0,0,0,46,0,0,0,153,0,85,0,6,0,212,0,0,0,238,0,178,0,15,0,82,0,128,0,0,0,0,0,46,0,124,0,227,0,110,0,18,0,162,0,30,0,82,0,186,0,100,0,134,0,12,0,0,0,221,0,204,0,55,0,243,0,168,0,101,0,65,0,222,0,128,0,0,0,225,0,201,0,170,0,200,0,57,0,0,0,0,0,0,0,54,0,0,0,123,0,90,0,0,0,104,0,17,0,208,0,75,0,0,0,79,0,16,0,0,0,14,0,55,0,185,0,0,0,0,0,34,0,234,0,128,0,88,0,200,0,0,0,0,0,4,0,109,0,39,0,41,0,0,0,135,0,54,0,195,0,0,0,0,0,30,0,191,0,5,0,142,0,0,0,0,0,65,0,183,0,20,0,195,0,66,0,9,0,116,0,172,0,89,0,63,0,24,0,0,0,45,0,233,0,0,0,131,0,101,0,104,0,182,0,51,0,197,0,132,0,201,0,0,0,223,0,0,0,229,0,20,0,229,0,112,0,0,0,26,0,209,0,21,0,80,0,37,0,162,0,0,0,243,0,29,0,0,0,188,0,0,0,41,0,169,0,132,0,47,0,99,0,252,0,183,0,127,0,26,0,0,0,0,0,11,0,59,0,76,0,184,0,0,0,198,0,160,0,171,0,195,0,176,0,122,0,0,0,221,0,135,0,186,0,201,0,0,0,237,0,169,0,234,0,78,0,209,0,0,0,198,0,183,0,72,0,187,0,9,0,34,0,48,0,199,0,163,0,138,0,3,0,48,0,191,0,232,0,119,0,161,0,176,0,232,0,96,0,0,0,161,0,148,0,201,0,144,0,93,0,0,0,132,0,99,0,25,0,145,0,149,0,0,0,224,0,0,0,97,0,104,0,190,0,91,0,199,0,138,0,185,0,204,0,49,0,176,0,0,0,40,0,190,0,0,0,0,0,199,0,196,0,53,0,251,0,56,0,111,0,137,0,0,0,133,0,86,0,4,0,247,0,87,0,119,0,0,0,15,0,0,0,107,0,162,0,0,0,254,0,17,0,123,0,8,0,77,0,244,0,0,0,103,0,149,0,198,0,25,0,116,0,115,0,0,0,103,0,158,0,79,0,0,0,166,0,100,0,220,0,38,0,0,0,40,0,0,0,31,0,32,0,169,0,150,0,0,0,83,0,80,0,68,0,0,0,119,0,0,0,64,0,95,0,68,0,2,0,76,0,215,0,0,0,73,0,0,0,0,0,0,0,29,0,0,0,0,0,245,0,101,0,168,0,42,0,38,0,202,0,0,0,0,0,38,0,158,0,64,0,60,0,87,0,251,0,0,0,69,0,0,0,83,0,213,0,146,0,0,0,0,0,137,0,209,0,171,0,196,0,104,0,76,0,64,0,170,0,228,0,37,0,85,0,37,0,180,0,4,0,62,0,241,0,0,0,101,0,0,0,236,0,242,0,0,0,192,0,0,0,0,0,0,0,167,0,151,0,214,0,0,0,249,0,3,0,146,0,204,0,131,0,173,0,60,0,200,0,59,0,125,0,93,0,65,0,64,0,202,0,93,0,85,0,119,0,41,0,0,0,65,0,77,0,0,0,183,0,0,0,16,0,42,0,160,0,0,0,117,0,0,0,245,0,157,0,219,0,228,0,162,0,157,0,128,0,208,0,75,0,229,0,0,0,13,0,124,0,101,0,203,0,0,0,163,0,109,0,187,0,2,0,148,0,0,0,173,0,163,0,0,0,188,0,95,0,61,0,0,0,173,0,0,0,190,0,116,0,35,0,180,0,0,0,0,0,0,0,0,0,0,0,34,0,167,0,220,0,200,0,0,0,112,0,252,0,13,0,0,0,197,0,27,0,194,0,78,0,175,0,90,0,183,0,209,0,0,0,251,0,179,0,209,0,204,0,208,0,41,0,0,0,84,0,4,0,141,0,42,0,62,0,116,0,4,0,120,0,153,0,0,0,0,0,84,0,78,0,203,0,236,0,137,0,133,0,95,0,203,0,0,0,232,0,143,0,0,0,251,0,166,0,0,0,5,0,82,0,26,0,126,0,181,0,235,0,182,0,211,0,218,0,0,0,15,0,149,0,1,0,121,0,132,0,13,0,252,0,0,0,62,0,74,0,0,0,204,0,178,0,189,0,27,0,104,0,131,0,15,0,208,0,129,0,83,0,24,0,75,0,0,0,159,0,0,0,121,0,10,0,140,0,209,0,37,0,250,0,64,0,113,0);
signal scenario_full  : scenario_type := (0,0,27,31,41,31,41,30,183,31,221,31,162,31,96,31,119,31,249,31,5,31,123,31,14,31,162,31,162,30,180,31,175,31,64,31,172,31,156,31,156,30,156,29,57,31,82,31,211,31,173,31,155,31,74,31,74,30,216,31,48,31,253,31,112,31,47,31,47,30,206,31,93,31,93,31,196,31,219,31,62,31,207,31,232,31,69,31,97,31,18,31,189,31,40,31,205,31,209,31,8,31,133,31,116,31,8,31,73,31,34,31,220,31,166,31,120,31,120,30,225,31,176,31,176,30,171,31,113,31,61,31,243,31,96,31,96,30,117,31,28,31,42,31,42,30,215,31,215,30,148,31,61,31,212,31,104,31,100,31,240,31,240,30,173,31,236,31,185,31,199,31,119,31,119,30,219,31,194,31,232,31,232,30,234,31,92,31,78,31,157,31,60,31,242,31,172,31,172,30,172,29,172,28,247,31,64,31,40,31,40,30,40,29,113,31,102,31,228,31,95,31,63,31,149,31,132,31,153,31,153,30,153,29,235,31,45,31,91,31,100,31,239,31,239,30,156,31,67,31,25,31,254,31,141,31,242,31,10,31,79,31,84,31,84,30,10,31,94,31,74,31,170,31,104,31,182,31,7,31,148,31,235,31,235,30,23,31,23,30,87,31,106,31,106,30,16,31,185,31,95,31,122,31,122,30,60,31,115,31,178,31,178,30,198,31,224,31,58,31,58,30,58,29,152,31,127,31,160,31,160,30,160,29,236,31,193,31,175,31,203,31,194,31,69,31,182,31,182,30,33,31,33,31,227,31,211,31,89,31,74,31,74,30,74,29,59,31,104,31,140,31,15,31,42,31,250,31,211,31,211,30,121,31,104,31,165,31,114,31,114,30,247,31,48,31,240,31,230,31,131,31,41,31,217,31,77,31,197,31,16,31,181,31,211,31,253,31,178,31,75,31,75,30,75,29,229,31,173,31,185,31,134,31,247,31,165,31,165,30,165,31,165,30,165,29,52,31,13,31,190,31,190,30,51,31,101,31,219,31,171,31,171,30,104,31,202,31,227,31,18,31,141,31,75,31,75,30,210,31,52,31,52,30,157,31,172,31,220,31,139,31,255,31,255,30,255,29,255,28,215,31,170,31,78,31,178,31,29,31,29,30,23,31,23,30,131,31,151,31,151,30,151,29,151,28,147,31,147,30,252,31,71,31,71,30,184,31,184,30,196,31,154,31,12,31,12,31,12,30,8,31,238,31,61,31,107,31,107,30,93,31,194,31,194,30,12,31,173,31,226,31,226,30,226,29,226,28,89,31,172,31,196,31,186,31,64,31,41,31,211,31,176,31,161,31,161,30,59,31,126,31,79,31,43,31,158,31,78,31,119,31,24,31,24,30,24,29,209,31,143,31,171,31,12,31,158,31,234,31,125,31,220,31,220,30,250,31,38,31,215,31,89,31,54,31,134,31,212,31,147,31,147,30,145,31,208,31,200,31,30,31,30,30,30,29,171,31,21,31,168,31,168,30,168,29,193,31,248,31,220,31,220,30,239,31,183,31,183,30,109,31,126,31,226,31,126,31,126,30,226,31,101,31,101,30,207,31,232,31,104,31,120,31,112,31,112,30,171,31,217,31,137,31,133,31,78,31,103,31,97,31,121,31,71,31,177,31,9,31,43,31,208,31,223,31,223,30,187,31,151,31,101,31,107,31,107,30,3,31,61,31,61,30,31,31,180,31,95,31,95,30,130,31,238,31,238,30,238,29,111,31,210,31,223,31,223,30,153,31,5,31,211,31,211,30,156,31,17,31,231,31,198,31,84,31,170,31,141,31,177,31,29,31,161,31,150,31,206,31,160,31,154,31,154,30,154,31,142,31,252,31,157,31,217,31,24,31,62,31,254,31,7,31,167,31,195,31,210,31,63,31,109,31,251,31,212,31,91,31,208,31,223,31,240,31,178,31,180,31,226,31,92,31,92,30,69,31,121,31,121,30,136,31,115,31,129,31,73,31,163,31,163,30,159,31,159,30,39,31,192,31,65,31,125,31,158,31,97,31,97,30,146,31,176,31,45,31,4,31,101,31,244,31,40,31,89,31,133,31,133,30,133,29,235,31,235,30,235,29,107,31,107,30,46,31,46,30,153,31,85,31,6,31,212,31,212,30,238,31,178,31,15,31,82,31,128,31,128,30,128,29,46,31,124,31,227,31,110,31,18,31,162,31,30,31,82,31,186,31,100,31,134,31,12,31,12,30,221,31,204,31,55,31,243,31,168,31,101,31,65,31,222,31,128,31,128,30,225,31,201,31,170,31,200,31,57,31,57,30,57,29,57,28,54,31,54,30,123,31,90,31,90,30,104,31,17,31,208,31,75,31,75,30,79,31,16,31,16,30,14,31,55,31,185,31,185,30,185,29,34,31,234,31,128,31,88,31,200,31,200,30,200,29,4,31,109,31,39,31,41,31,41,30,135,31,54,31,195,31,195,30,195,29,30,31,191,31,5,31,142,31,142,30,142,29,65,31,183,31,20,31,195,31,66,31,9,31,116,31,172,31,89,31,63,31,24,31,24,30,45,31,233,31,233,30,131,31,101,31,104,31,182,31,51,31,197,31,132,31,201,31,201,30,223,31,223,30,229,31,20,31,229,31,112,31,112,30,26,31,209,31,21,31,80,31,37,31,162,31,162,30,243,31,29,31,29,30,188,31,188,30,41,31,169,31,132,31,47,31,99,31,252,31,183,31,127,31,26,31,26,30,26,29,11,31,59,31,76,31,184,31,184,30,198,31,160,31,171,31,195,31,176,31,122,31,122,30,221,31,135,31,186,31,201,31,201,30,237,31,169,31,234,31,78,31,209,31,209,30,198,31,183,31,72,31,187,31,9,31,34,31,48,31,199,31,163,31,138,31,3,31,48,31,191,31,232,31,119,31,161,31,176,31,232,31,96,31,96,30,161,31,148,31,201,31,144,31,93,31,93,30,132,31,99,31,25,31,145,31,149,31,149,30,224,31,224,30,97,31,104,31,190,31,91,31,199,31,138,31,185,31,204,31,49,31,176,31,176,30,40,31,190,31,190,30,190,29,199,31,196,31,53,31,251,31,56,31,111,31,137,31,137,30,133,31,86,31,4,31,247,31,87,31,119,31,119,30,15,31,15,30,107,31,162,31,162,30,254,31,17,31,123,31,8,31,77,31,244,31,244,30,103,31,149,31,198,31,25,31,116,31,115,31,115,30,103,31,158,31,79,31,79,30,166,31,100,31,220,31,38,31,38,30,40,31,40,30,31,31,32,31,169,31,150,31,150,30,83,31,80,31,68,31,68,30,119,31,119,30,64,31,95,31,68,31,2,31,76,31,215,31,215,30,73,31,73,30,73,29,73,28,29,31,29,30,29,29,245,31,101,31,168,31,42,31,38,31,202,31,202,30,202,29,38,31,158,31,64,31,60,31,87,31,251,31,251,30,69,31,69,30,83,31,213,31,146,31,146,30,146,29,137,31,209,31,171,31,196,31,104,31,76,31,64,31,170,31,228,31,37,31,85,31,37,31,180,31,4,31,62,31,241,31,241,30,101,31,101,30,236,31,242,31,242,30,192,31,192,30,192,29,192,28,167,31,151,31,214,31,214,30,249,31,3,31,146,31,204,31,131,31,173,31,60,31,200,31,59,31,125,31,93,31,65,31,64,31,202,31,93,31,85,31,119,31,41,31,41,30,65,31,77,31,77,30,183,31,183,30,16,31,42,31,160,31,160,30,117,31,117,30,245,31,157,31,219,31,228,31,162,31,157,31,128,31,208,31,75,31,229,31,229,30,13,31,124,31,101,31,203,31,203,30,163,31,109,31,187,31,2,31,148,31,148,30,173,31,163,31,163,30,188,31,95,31,61,31,61,30,173,31,173,30,190,31,116,31,35,31,180,31,180,30,180,29,180,28,180,27,180,26,34,31,167,31,220,31,200,31,200,30,112,31,252,31,13,31,13,30,197,31,27,31,194,31,78,31,175,31,90,31,183,31,209,31,209,30,251,31,179,31,209,31,204,31,208,31,41,31,41,30,84,31,4,31,141,31,42,31,62,31,116,31,4,31,120,31,153,31,153,30,153,29,84,31,78,31,203,31,236,31,137,31,133,31,95,31,203,31,203,30,232,31,143,31,143,30,251,31,166,31,166,30,5,31,82,31,26,31,126,31,181,31,235,31,182,31,211,31,218,31,218,30,15,31,149,31,1,31,121,31,132,31,13,31,252,31,252,30,62,31,74,31,74,30,204,31,178,31,189,31,27,31,104,31,131,31,15,31,208,31,129,31,83,31,24,31,75,31,75,30,159,31,159,30,121,31,10,31,140,31,209,31,37,31,250,31,64,31,113,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
