-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_688 is
end project_tb_688;

architecture project_tb_arch_688 of project_tb_688 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 301;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,126,0,201,0,144,0,0,0,254,0,0,0,123,0,30,0,236,0,0,0,0,0,0,0,58,0,54,0,0,0,0,0,71,0,0,0,13,0,140,0,16,0,216,0,0,0,169,0,3,0,0,0,135,0,17,0,134,0,133,0,206,0,0,0,0,0,57,0,113,0,16,0,143,0,0,0,129,0,108,0,0,0,79,0,245,0,37,0,204,0,0,0,155,0,0,0,0,0,0,0,162,0,12,0,28,0,100,0,57,0,214,0,173,0,0,0,16,0,147,0,205,0,237,0,158,0,0,0,58,0,0,0,238,0,0,0,104,0,236,0,153,0,161,0,158,0,177,0,162,0,168,0,248,0,183,0,0,0,87,0,208,0,110,0,108,0,36,0,94,0,78,0,151,0,0,0,0,0,65,0,235,0,93,0,164,0,192,0,145,0,14,0,1,0,250,0,97,0,91,0,0,0,187,0,62,0,105,0,0,0,133,0,204,0,85,0,70,0,0,0,0,0,79,0,95,0,175,0,129,0,30,0,95,0,149,0,18,0,234,0,95,0,76,0,75,0,131,0,249,0,109,0,44,0,34,0,0,0,175,0,157,0,0,0,74,0,254,0,208,0,65,0,0,0,9,0,217,0,129,0,4,0,14,0,195,0,165,0,0,0,0,0,12,0,23,0,0,0,26,0,33,0,250,0,69,0,123,0,0,0,0,0,0,0,167,0,0,0,1,0,35,0,40,0,93,0,144,0,210,0,84,0,219,0,0,0,219,0,5,0,134,0,178,0,207,0,96,0,217,0,210,0,53,0,1,0,74,0,81,0,58,0,187,0,132,0,68,0,0,0,53,0,236,0,73,0,126,0,0,0,92,0,124,0,136,0,0,0,174,0,107,0,0,0,188,0,223,0,199,0,0,0,174,0,231,0,136,0,196,0,26,0,18,0,224,0,218,0,107,0,234,0,66,0,5,0,182,0,103,0,0,0,16,0,0,0,196,0,57,0,17,0,9,0,20,0,47,0,92,0,143,0,87,0,28,0,0,0,219,0,0,0,79,0,0,0,119,0,80,0,201,0,50,0,78,0,22,0,80,0,3,0,0,0,206,0,188,0,58,0,0,0,119,0,241,0,65,0,107,0,56,0,132,0,0,0,164,0,191,0,23,0,228,0,0,0,152,0,218,0,15,0,0,0,49,0,10,0,115,0,146,0,54,0,67,0,25,0,0,0,88,0,40,0,191,0,49,0,10,0,220,0,83,0,147,0,142,0,153,0,0,0,0,0,98,0,75,0,242,0,45,0,57,0,40,0,9,0,0,0,0,0,13,0,217,0,194,0,9,0,104,0,175,0,214,0,41,0,135,0);
signal scenario_full  : scenario_type := (0,0,126,31,201,31,144,31,144,30,254,31,254,30,123,31,30,31,236,31,236,30,236,29,236,28,58,31,54,31,54,30,54,29,71,31,71,30,13,31,140,31,16,31,216,31,216,30,169,31,3,31,3,30,135,31,17,31,134,31,133,31,206,31,206,30,206,29,57,31,113,31,16,31,143,31,143,30,129,31,108,31,108,30,79,31,245,31,37,31,204,31,204,30,155,31,155,30,155,29,155,28,162,31,12,31,28,31,100,31,57,31,214,31,173,31,173,30,16,31,147,31,205,31,237,31,158,31,158,30,58,31,58,30,238,31,238,30,104,31,236,31,153,31,161,31,158,31,177,31,162,31,168,31,248,31,183,31,183,30,87,31,208,31,110,31,108,31,36,31,94,31,78,31,151,31,151,30,151,29,65,31,235,31,93,31,164,31,192,31,145,31,14,31,1,31,250,31,97,31,91,31,91,30,187,31,62,31,105,31,105,30,133,31,204,31,85,31,70,31,70,30,70,29,79,31,95,31,175,31,129,31,30,31,95,31,149,31,18,31,234,31,95,31,76,31,75,31,131,31,249,31,109,31,44,31,34,31,34,30,175,31,157,31,157,30,74,31,254,31,208,31,65,31,65,30,9,31,217,31,129,31,4,31,14,31,195,31,165,31,165,30,165,29,12,31,23,31,23,30,26,31,33,31,250,31,69,31,123,31,123,30,123,29,123,28,167,31,167,30,1,31,35,31,40,31,93,31,144,31,210,31,84,31,219,31,219,30,219,31,5,31,134,31,178,31,207,31,96,31,217,31,210,31,53,31,1,31,74,31,81,31,58,31,187,31,132,31,68,31,68,30,53,31,236,31,73,31,126,31,126,30,92,31,124,31,136,31,136,30,174,31,107,31,107,30,188,31,223,31,199,31,199,30,174,31,231,31,136,31,196,31,26,31,18,31,224,31,218,31,107,31,234,31,66,31,5,31,182,31,103,31,103,30,16,31,16,30,196,31,57,31,17,31,9,31,20,31,47,31,92,31,143,31,87,31,28,31,28,30,219,31,219,30,79,31,79,30,119,31,80,31,201,31,50,31,78,31,22,31,80,31,3,31,3,30,206,31,188,31,58,31,58,30,119,31,241,31,65,31,107,31,56,31,132,31,132,30,164,31,191,31,23,31,228,31,228,30,152,31,218,31,15,31,15,30,49,31,10,31,115,31,146,31,54,31,67,31,25,31,25,30,88,31,40,31,191,31,49,31,10,31,220,31,83,31,147,31,142,31,153,31,153,30,153,29,98,31,75,31,242,31,45,31,57,31,40,31,9,31,9,30,9,29,13,31,217,31,194,31,9,31,104,31,175,31,214,31,41,31,135,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
