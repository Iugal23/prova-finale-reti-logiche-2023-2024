-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_695 is
end project_tb_695;

architecture project_tb_arch_695 of project_tb_695 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 361;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,20,0,139,0,203,0,194,0,168,0,112,0,2,0,23,0,224,0,84,0,120,0,120,0,161,0,93,0,181,0,1,0,97,0,162,0,26,0,102,0,207,0,72,0,111,0,179,0,192,0,66,0,1,0,0,0,11,0,70,0,188,0,217,0,89,0,206,0,78,0,126,0,26,0,214,0,128,0,0,0,0,0,137,0,0,0,149,0,118,0,0,0,0,0,205,0,137,0,0,0,155,0,0,0,0,0,201,0,118,0,0,0,8,0,51,0,104,0,136,0,38,0,58,0,62,0,149,0,195,0,123,0,160,0,0,0,179,0,36,0,99,0,230,0,150,0,218,0,219,0,134,0,0,0,157,0,18,0,252,0,203,0,183,0,0,0,154,0,35,0,103,0,10,0,9,0,135,0,0,0,210,0,141,0,49,0,0,0,11,0,45,0,0,0,0,0,131,0,110,0,104,0,32,0,251,0,127,0,214,0,53,0,0,0,76,0,60,0,0,0,219,0,28,0,0,0,189,0,164,0,213,0,112,0,63,0,166,0,33,0,14,0,128,0,238,0,132,0,103,0,205,0,62,0,63,0,83,0,20,0,0,0,0,0,14,0,22,0,85,0,218,0,59,0,202,0,215,0,182,0,66,0,160,0,203,0,0,0,0,0,103,0,55,0,183,0,128,0,30,0,171,0,19,0,222,0,133,0,246,0,158,0,245,0,15,0,196,0,89,0,185,0,0,0,53,0,157,0,233,0,0,0,230,0,192,0,81,0,0,0,204,0,0,0,214,0,217,0,109,0,11,0,94,0,112,0,0,0,110,0,0,0,63,0,123,0,106,0,0,0,0,0,18,0,0,0,203,0,91,0,0,0,219,0,91,0,105,0,153,0,0,0,56,0,176,0,228,0,55,0,68,0,33,0,61,0,118,0,6,0,0,0,0,0,3,0,178,0,137,0,11,0,114,0,64,0,141,0,162,0,0,0,43,0,0,0,0,0,252,0,218,0,88,0,213,0,44,0,214,0,194,0,11,0,13,0,176,0,0,0,112,0,0,0,202,0,0,0,62,0,154,0,111,0,0,0,91,0,180,0,42,0,85,0,224,0,52,0,177,0,77,0,129,0,205,0,186,0,0,0,170,0,0,0,141,0,0,0,133,0,111,0,244,0,89,0,189,0,204,0,162,0,41,0,28,0,0,0,103,0,202,0,0,0,204,0,116,0,34,0,231,0,250,0,12,0,171,0,39,0,255,0,186,0,192,0,182,0,154,0,144,0,168,0,0,0,51,0,159,0,0,0,207,0,0,0,81,0,0,0,210,0,222,0,200,0,1,0,0,0,40,0,252,0,96,0,0,0,0,0,0,0,61,0,200,0,0,0,71,0,0,0,164,0,0,0,210,0,182,0,148,0,252,0,89,0,0,0,0,0,118,0,121,0,39,0,194,0,109,0,215,0,52,0,50,0,102,0,5,0,155,0,85,0,144,0,67,0,175,0,0,0,107,0,0,0,48,0,176,0,0,0,154,0,233,0,59,0,28,0,224,0,0,0,206,0,0,0,211,0,219,0,207,0,0,0,147,0,129,0,0,0,152,0,246,0,103,0,55,0,151,0,87,0,63,0,0,0,36,0);
signal scenario_full  : scenario_type := (0,0,20,31,139,31,203,31,194,31,168,31,112,31,2,31,23,31,224,31,84,31,120,31,120,31,161,31,93,31,181,31,1,31,97,31,162,31,26,31,102,31,207,31,72,31,111,31,179,31,192,31,66,31,1,31,1,30,11,31,70,31,188,31,217,31,89,31,206,31,78,31,126,31,26,31,214,31,128,31,128,30,128,29,137,31,137,30,149,31,118,31,118,30,118,29,205,31,137,31,137,30,155,31,155,30,155,29,201,31,118,31,118,30,8,31,51,31,104,31,136,31,38,31,58,31,62,31,149,31,195,31,123,31,160,31,160,30,179,31,36,31,99,31,230,31,150,31,218,31,219,31,134,31,134,30,157,31,18,31,252,31,203,31,183,31,183,30,154,31,35,31,103,31,10,31,9,31,135,31,135,30,210,31,141,31,49,31,49,30,11,31,45,31,45,30,45,29,131,31,110,31,104,31,32,31,251,31,127,31,214,31,53,31,53,30,76,31,60,31,60,30,219,31,28,31,28,30,189,31,164,31,213,31,112,31,63,31,166,31,33,31,14,31,128,31,238,31,132,31,103,31,205,31,62,31,63,31,83,31,20,31,20,30,20,29,14,31,22,31,85,31,218,31,59,31,202,31,215,31,182,31,66,31,160,31,203,31,203,30,203,29,103,31,55,31,183,31,128,31,30,31,171,31,19,31,222,31,133,31,246,31,158,31,245,31,15,31,196,31,89,31,185,31,185,30,53,31,157,31,233,31,233,30,230,31,192,31,81,31,81,30,204,31,204,30,214,31,217,31,109,31,11,31,94,31,112,31,112,30,110,31,110,30,63,31,123,31,106,31,106,30,106,29,18,31,18,30,203,31,91,31,91,30,219,31,91,31,105,31,153,31,153,30,56,31,176,31,228,31,55,31,68,31,33,31,61,31,118,31,6,31,6,30,6,29,3,31,178,31,137,31,11,31,114,31,64,31,141,31,162,31,162,30,43,31,43,30,43,29,252,31,218,31,88,31,213,31,44,31,214,31,194,31,11,31,13,31,176,31,176,30,112,31,112,30,202,31,202,30,62,31,154,31,111,31,111,30,91,31,180,31,42,31,85,31,224,31,52,31,177,31,77,31,129,31,205,31,186,31,186,30,170,31,170,30,141,31,141,30,133,31,111,31,244,31,89,31,189,31,204,31,162,31,41,31,28,31,28,30,103,31,202,31,202,30,204,31,116,31,34,31,231,31,250,31,12,31,171,31,39,31,255,31,186,31,192,31,182,31,154,31,144,31,168,31,168,30,51,31,159,31,159,30,207,31,207,30,81,31,81,30,210,31,222,31,200,31,1,31,1,30,40,31,252,31,96,31,96,30,96,29,96,28,61,31,200,31,200,30,71,31,71,30,164,31,164,30,210,31,182,31,148,31,252,31,89,31,89,30,89,29,118,31,121,31,39,31,194,31,109,31,215,31,52,31,50,31,102,31,5,31,155,31,85,31,144,31,67,31,175,31,175,30,107,31,107,30,48,31,176,31,176,30,154,31,233,31,59,31,28,31,224,31,224,30,206,31,206,30,211,31,219,31,207,31,207,30,147,31,129,31,129,30,152,31,246,31,103,31,55,31,151,31,87,31,63,31,63,30,36,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
