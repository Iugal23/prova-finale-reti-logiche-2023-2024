-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_430 is
end project_tb_430;

architecture project_tb_arch_430 of project_tb_430 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 797;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,253,0,98,0,0,0,0,0,193,0,26,0,220,0,67,0,84,0,107,0,199,0,98,0,240,0,39,0,0,0,34,0,188,0,70,0,164,0,0,0,0,0,204,0,168,0,29,0,0,0,93,0,140,0,170,0,198,0,0,0,192,0,83,0,241,0,103,0,0,0,241,0,0,0,17,0,137,0,0,0,0,0,0,0,64,0,0,0,192,0,44,0,187,0,0,0,1,0,151,0,0,0,107,0,140,0,165,0,134,0,0,0,215,0,0,0,55,0,134,0,102,0,29,0,0,0,70,0,169,0,140,0,0,0,50,0,85,0,92,0,215,0,0,0,206,0,63,0,7,0,104,0,50,0,248,0,142,0,0,0,69,0,221,0,12,0,40,0,241,0,55,0,0,0,78,0,163,0,41,0,31,0,0,0,0,0,120,0,112,0,74,0,55,0,214,0,0,0,36,0,195,0,0,0,131,0,0,0,86,0,219,0,121,0,0,0,97,0,14,0,0,0,190,0,175,0,227,0,11,0,169,0,1,0,0,0,81,0,230,0,154,0,75,0,222,0,0,0,226,0,68,0,0,0,53,0,164,0,176,0,6,0,155,0,134,0,207,0,179,0,101,0,24,0,148,0,143,0,135,0,255,0,128,0,76,0,6,0,143,0,153,0,203,0,19,0,0,0,55,0,14,0,60,0,8,0,90,0,72,0,162,0,137,0,111,0,43,0,39,0,152,0,255,0,11,0,107,0,30,0,0,0,186,0,111,0,154,0,9,0,8,0,225,0,97,0,36,0,12,0,0,0,141,0,112,0,0,0,162,0,0,0,55,0,0,0,117,0,49,0,114,0,211,0,246,0,12,0,228,0,170,0,162,0,0,0,221,0,112,0,231,0,44,0,69,0,185,0,56,0,43,0,0,0,107,0,111,0,35,0,57,0,29,0,198,0,9,0,224,0,0,0,251,0,37,0,50,0,0,0,29,0,0,0,0,0,7,0,156,0,42,0,203,0,0,0,252,0,175,0,171,0,124,0,77,0,0,0,235,0,78,0,0,0,0,0,131,0,0,0,0,0,0,0,0,0,215,0,182,0,0,0,101,0,209,0,118,0,213,0,57,0,19,0,90,0,0,0,22,0,162,0,81,0,97,0,196,0,6,0,214,0,151,0,160,0,196,0,224,0,216,0,32,0,54,0,204,0,0,0,96,0,230,0,72,0,255,0,33,0,214,0,130,0,0,0,0,0,213,0,60,0,202,0,150,0,84,0,117,0,121,0,0,0,59,0,0,0,91,0,5,0,0,0,130,0,228,0,43,0,57,0,138,0,10,0,0,0,0,0,0,0,197,0,85,0,17,0,0,0,219,0,105,0,0,0,33,0,190,0,191,0,237,0,207,0,152,0,208,0,0,0,0,0,62,0,0,0,253,0,3,0,167,0,229,0,165,0,49,0,158,0,218,0,212,0,174,0,0,0,162,0,222,0,247,0,23,0,235,0,254,0,66,0,251,0,181,0,12,0,83,0,21,0,130,0,185,0,213,0,240,0,225,0,151,0,253,0,112,0,237,0,143,0,248,0,0,0,244,0,116,0,212,0,17,0,134,0,0,0,42,0,16,0,8,0,159,0,129,0,155,0,91,0,193,0,200,0,157,0,41,0,0,0,179,0,0,0,0,0,0,0,188,0,0,0,175,0,72,0,54,0,130,0,158,0,19,0,62,0,130,0,135,0,47,0,37,0,192,0,0,0,162,0,85,0,37,0,140,0,0,0,167,0,112,0,0,0,48,0,173,0,49,0,127,0,173,0,202,0,207,0,199,0,63,0,207,0,0,0,27,0,0,0,203,0,238,0,0,0,235,0,232,0,227,0,163,0,90,0,40,0,162,0,172,0,0,0,68,0,196,0,170,0,54,0,80,0,41,0,8,0,193,0,129,0,156,0,113,0,101,0,141,0,71,0,151,0,229,0,0,0,0,0,0,0,0,0,115,0,98,0,45,0,163,0,239,0,91,0,208,0,242,0,0,0,24,0,19,0,29,0,0,0,133,0,149,0,46,0,0,0,104,0,64,0,136,0,202,0,0,0,160,0,0,0,44,0,36,0,78,0,0,0,206,0,0,0,228,0,0,0,184,0,234,0,0,0,20,0,19,0,206,0,69,0,87,0,236,0,190,0,85,0,0,0,74,0,46,0,0,0,0,0,89,0,0,0,187,0,75,0,175,0,0,0,184,0,122,0,93,0,37,0,254,0,0,0,0,0,203,0,0,0,3,0,235,0,186,0,241,0,4,0,132,0,95,0,118,0,24,0,53,0,62,0,119,0,190,0,161,0,181,0,237,0,174,0,0,0,135,0,98,0,45,0,0,0,246,0,198,0,98,0,0,0,176,0,0,0,235,0,0,0,134,0,0,0,25,0,69,0,234,0,0,0,193,0,251,0,146,0,38,0,187,0,180,0,97,0,69,0,212,0,1,0,66,0,162,0,238,0,39,0,0,0,181,0,230,0,215,0,90,0,146,0,0,0,134,0,0,0,183,0,0,0,204,0,244,0,62,0,135,0,2,0,219,0,113,0,81,0,60,0,179,0,122,0,254,0,0,0,0,0,76,0,148,0,235,0,131,0,0,0,0,0,21,0,92,0,91,0,108,0,0,0,0,0,200,0,132,0,116,0,0,0,49,0,79,0,138,0,199,0,208,0,28,0,226,0,252,0,119,0,133,0,10,0,227,0,26,0,0,0,228,0,0,0,182,0,133,0,0,0,0,0,31,0,173,0,0,0,119,0,95,0,210,0,4,0,97,0,183,0,21,0,48,0,138,0,0,0,231,0,78,0,191,0,0,0,55,0,178,0,6,0,25,0,108,0,0,0,136,0,11,0,253,0,62,0,12,0,99,0,191,0,91,0,133,0,148,0,230,0,90,0,0,0,155,0,0,0,5,0,5,0,106,0,170,0,99,0,0,0,0,0,87,0,215,0,5,0,5,0,187,0,0,0,0,0,233,0,222,0,245,0,0,0,173,0,237,0,135,0,16,0,96,0,174,0,143,0,20,0,176,0,216,0,86,0,0,0,152,0,190,0,57,0,167,0,111,0,209,0,101,0,70,0,236,0,0,0,198,0,0,0,107,0,36,0,139,0,22,0,0,0,113,0,0,0,160,0,230,0,238,0,127,0,30,0,0,0,244,0,0,0,68,0,118,0,212,0,20,0,172,0,13,0,210,0,0,0,75,0,87,0,6,0,162,0,63,0,131,0,208,0,98,0,253,0,150,0,24,0,28,0,0,0,199,0,221,0,41,0,0,0,111,0,39,0,0,0,0,0,189,0,37,0,25,0,38,0,113,0,239,0,182,0,114,0,0,0,128,0,203,0,0,0,68,0,49,0,4,0,10,0,229,0,161,0,150,0,0,0,206,0,122,0,254,0,130,0,205,0,115,0,76,0,11,0,133,0,0,0,0,0,93,0,158,0,41,0,157,0,26,0,176,0,85,0,154,0,0,0,0,0,100,0,183,0,26,0,63,0,11,0,0,0,127,0,52,0,253,0,140,0,184,0,228,0,99,0,74,0,117,0,92,0,15,0,236,0);
signal scenario_full  : scenario_type := (195,31,253,31,98,31,98,30,98,29,193,31,26,31,220,31,67,31,84,31,107,31,199,31,98,31,240,31,39,31,39,30,34,31,188,31,70,31,164,31,164,30,164,29,204,31,168,31,29,31,29,30,93,31,140,31,170,31,198,31,198,30,192,31,83,31,241,31,103,31,103,30,241,31,241,30,17,31,137,31,137,30,137,29,137,28,64,31,64,30,192,31,44,31,187,31,187,30,1,31,151,31,151,30,107,31,140,31,165,31,134,31,134,30,215,31,215,30,55,31,134,31,102,31,29,31,29,30,70,31,169,31,140,31,140,30,50,31,85,31,92,31,215,31,215,30,206,31,63,31,7,31,104,31,50,31,248,31,142,31,142,30,69,31,221,31,12,31,40,31,241,31,55,31,55,30,78,31,163,31,41,31,31,31,31,30,31,29,120,31,112,31,74,31,55,31,214,31,214,30,36,31,195,31,195,30,131,31,131,30,86,31,219,31,121,31,121,30,97,31,14,31,14,30,190,31,175,31,227,31,11,31,169,31,1,31,1,30,81,31,230,31,154,31,75,31,222,31,222,30,226,31,68,31,68,30,53,31,164,31,176,31,6,31,155,31,134,31,207,31,179,31,101,31,24,31,148,31,143,31,135,31,255,31,128,31,76,31,6,31,143,31,153,31,203,31,19,31,19,30,55,31,14,31,60,31,8,31,90,31,72,31,162,31,137,31,111,31,43,31,39,31,152,31,255,31,11,31,107,31,30,31,30,30,186,31,111,31,154,31,9,31,8,31,225,31,97,31,36,31,12,31,12,30,141,31,112,31,112,30,162,31,162,30,55,31,55,30,117,31,49,31,114,31,211,31,246,31,12,31,228,31,170,31,162,31,162,30,221,31,112,31,231,31,44,31,69,31,185,31,56,31,43,31,43,30,107,31,111,31,35,31,57,31,29,31,198,31,9,31,224,31,224,30,251,31,37,31,50,31,50,30,29,31,29,30,29,29,7,31,156,31,42,31,203,31,203,30,252,31,175,31,171,31,124,31,77,31,77,30,235,31,78,31,78,30,78,29,131,31,131,30,131,29,131,28,131,27,215,31,182,31,182,30,101,31,209,31,118,31,213,31,57,31,19,31,90,31,90,30,22,31,162,31,81,31,97,31,196,31,6,31,214,31,151,31,160,31,196,31,224,31,216,31,32,31,54,31,204,31,204,30,96,31,230,31,72,31,255,31,33,31,214,31,130,31,130,30,130,29,213,31,60,31,202,31,150,31,84,31,117,31,121,31,121,30,59,31,59,30,91,31,5,31,5,30,130,31,228,31,43,31,57,31,138,31,10,31,10,30,10,29,10,28,197,31,85,31,17,31,17,30,219,31,105,31,105,30,33,31,190,31,191,31,237,31,207,31,152,31,208,31,208,30,208,29,62,31,62,30,253,31,3,31,167,31,229,31,165,31,49,31,158,31,218,31,212,31,174,31,174,30,162,31,222,31,247,31,23,31,235,31,254,31,66,31,251,31,181,31,12,31,83,31,21,31,130,31,185,31,213,31,240,31,225,31,151,31,253,31,112,31,237,31,143,31,248,31,248,30,244,31,116,31,212,31,17,31,134,31,134,30,42,31,16,31,8,31,159,31,129,31,155,31,91,31,193,31,200,31,157,31,41,31,41,30,179,31,179,30,179,29,179,28,188,31,188,30,175,31,72,31,54,31,130,31,158,31,19,31,62,31,130,31,135,31,47,31,37,31,192,31,192,30,162,31,85,31,37,31,140,31,140,30,167,31,112,31,112,30,48,31,173,31,49,31,127,31,173,31,202,31,207,31,199,31,63,31,207,31,207,30,27,31,27,30,203,31,238,31,238,30,235,31,232,31,227,31,163,31,90,31,40,31,162,31,172,31,172,30,68,31,196,31,170,31,54,31,80,31,41,31,8,31,193,31,129,31,156,31,113,31,101,31,141,31,71,31,151,31,229,31,229,30,229,29,229,28,229,27,115,31,98,31,45,31,163,31,239,31,91,31,208,31,242,31,242,30,24,31,19,31,29,31,29,30,133,31,149,31,46,31,46,30,104,31,64,31,136,31,202,31,202,30,160,31,160,30,44,31,36,31,78,31,78,30,206,31,206,30,228,31,228,30,184,31,234,31,234,30,20,31,19,31,206,31,69,31,87,31,236,31,190,31,85,31,85,30,74,31,46,31,46,30,46,29,89,31,89,30,187,31,75,31,175,31,175,30,184,31,122,31,93,31,37,31,254,31,254,30,254,29,203,31,203,30,3,31,235,31,186,31,241,31,4,31,132,31,95,31,118,31,24,31,53,31,62,31,119,31,190,31,161,31,181,31,237,31,174,31,174,30,135,31,98,31,45,31,45,30,246,31,198,31,98,31,98,30,176,31,176,30,235,31,235,30,134,31,134,30,25,31,69,31,234,31,234,30,193,31,251,31,146,31,38,31,187,31,180,31,97,31,69,31,212,31,1,31,66,31,162,31,238,31,39,31,39,30,181,31,230,31,215,31,90,31,146,31,146,30,134,31,134,30,183,31,183,30,204,31,244,31,62,31,135,31,2,31,219,31,113,31,81,31,60,31,179,31,122,31,254,31,254,30,254,29,76,31,148,31,235,31,131,31,131,30,131,29,21,31,92,31,91,31,108,31,108,30,108,29,200,31,132,31,116,31,116,30,49,31,79,31,138,31,199,31,208,31,28,31,226,31,252,31,119,31,133,31,10,31,227,31,26,31,26,30,228,31,228,30,182,31,133,31,133,30,133,29,31,31,173,31,173,30,119,31,95,31,210,31,4,31,97,31,183,31,21,31,48,31,138,31,138,30,231,31,78,31,191,31,191,30,55,31,178,31,6,31,25,31,108,31,108,30,136,31,11,31,253,31,62,31,12,31,99,31,191,31,91,31,133,31,148,31,230,31,90,31,90,30,155,31,155,30,5,31,5,31,106,31,170,31,99,31,99,30,99,29,87,31,215,31,5,31,5,31,187,31,187,30,187,29,233,31,222,31,245,31,245,30,173,31,237,31,135,31,16,31,96,31,174,31,143,31,20,31,176,31,216,31,86,31,86,30,152,31,190,31,57,31,167,31,111,31,209,31,101,31,70,31,236,31,236,30,198,31,198,30,107,31,36,31,139,31,22,31,22,30,113,31,113,30,160,31,230,31,238,31,127,31,30,31,30,30,244,31,244,30,68,31,118,31,212,31,20,31,172,31,13,31,210,31,210,30,75,31,87,31,6,31,162,31,63,31,131,31,208,31,98,31,253,31,150,31,24,31,28,31,28,30,199,31,221,31,41,31,41,30,111,31,39,31,39,30,39,29,189,31,37,31,25,31,38,31,113,31,239,31,182,31,114,31,114,30,128,31,203,31,203,30,68,31,49,31,4,31,10,31,229,31,161,31,150,31,150,30,206,31,122,31,254,31,130,31,205,31,115,31,76,31,11,31,133,31,133,30,133,29,93,31,158,31,41,31,157,31,26,31,176,31,85,31,154,31,154,30,154,29,100,31,183,31,26,31,63,31,11,31,11,30,127,31,52,31,253,31,140,31,184,31,228,31,99,31,74,31,117,31,92,31,15,31,236,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
