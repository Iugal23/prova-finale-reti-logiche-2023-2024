-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 337;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (161,0,0,0,136,0,250,0,122,0,91,0,20,0,12,0,68,0,183,0,0,0,150,0,215,0,124,0,97,0,153,0,0,0,77,0,233,0,0,0,0,0,248,0,152,0,211,0,101,0,104,0,172,0,173,0,0,0,140,0,56,0,0,0,224,0,0,0,215,0,130,0,108,0,134,0,0,0,218,0,0,0,241,0,14,0,220,0,19,0,215,0,0,0,25,0,110,0,201,0,0,0,120,0,215,0,14,0,0,0,207,0,189,0,0,0,109,0,116,0,67,0,0,0,110,0,227,0,96,0,129,0,0,0,2,0,255,0,0,0,86,0,153,0,0,0,0,0,119,0,5,0,44,0,0,0,222,0,49,0,65,0,49,0,199,0,136,0,144,0,247,0,60,0,40,0,0,0,0,0,0,0,230,0,185,0,173,0,0,0,244,0,0,0,61,0,82,0,169,0,44,0,110,0,69,0,208,0,247,0,53,0,0,0,109,0,116,0,201,0,198,0,134,0,65,0,0,0,0,0,0,0,125,0,0,0,102,0,207,0,117,0,29,0,155,0,68,0,84,0,135,0,0,0,238,0,0,0,123,0,236,0,23,0,157,0,43,0,97,0,94,0,50,0,145,0,197,0,251,0,220,0,100,0,0,0,228,0,171,0,187,0,0,0,156,0,0,0,9,0,25,0,0,0,0,0,189,0,183,0,111,0,127,0,176,0,139,0,4,0,0,0,0,0,252,0,9,0,139,0,174,0,244,0,59,0,167,0,60,0,212,0,191,0,0,0,0,0,135,0,181,0,0,0,0,0,209,0,117,0,109,0,0,0,132,0,245,0,26,0,220,0,8,0,85,0,68,0,152,0,137,0,55,0,48,0,199,0,0,0,0,0,53,0,41,0,109,0,117,0,138,0,27,0,129,0,181,0,64,0,0,0,249,0,161,0,0,0,57,0,199,0,144,0,0,0,61,0,230,0,178,0,238,0,214,0,76,0,123,0,150,0,0,0,224,0,0,0,31,0,55,0,0,0,45,0,48,0,186,0,86,0,55,0,252,0,180,0,80,0,0,0,217,0,41,0,44,0,56,0,134,0,240,0,131,0,131,0,118,0,0,0,226,0,211,0,135,0,253,0,181,0,57,0,154,0,0,0,192,0,56,0,0,0,87,0,21,0,0,0,156,0,0,0,67,0,0,0,0,0,103,0,144,0,124,0,0,0,53,0,0,0,151,0,0,0,222,0,43,0,134,0,92,0,31,0,12,0,56,0,185,0,116,0,161,0,0,0,55,0,176,0,0,0,86,0,229,0,133,0,0,0,10,0,122,0,197,0,0,0,149,0,0,0,217,0,1,0,0,0,188,0,0,0,179,0,0,0,6,0,104,0,81,0,44,0,125,0,36,0,83,0,222,0,2,0,216,0,0,0,162,0,11,0,193,0,75,0,193,0,78,0,253,0,135,0,237,0,88,0,219,0,0,0,52,0,0,0,63,0,174,0,0,0,130,0,110,0,69,0,12,0,57,0);
signal scenario_full  : scenario_type := (161,31,161,30,136,31,250,31,122,31,91,31,20,31,12,31,68,31,183,31,183,30,150,31,215,31,124,31,97,31,153,31,153,30,77,31,233,31,233,30,233,29,248,31,152,31,211,31,101,31,104,31,172,31,173,31,173,30,140,31,56,31,56,30,224,31,224,30,215,31,130,31,108,31,134,31,134,30,218,31,218,30,241,31,14,31,220,31,19,31,215,31,215,30,25,31,110,31,201,31,201,30,120,31,215,31,14,31,14,30,207,31,189,31,189,30,109,31,116,31,67,31,67,30,110,31,227,31,96,31,129,31,129,30,2,31,255,31,255,30,86,31,153,31,153,30,153,29,119,31,5,31,44,31,44,30,222,31,49,31,65,31,49,31,199,31,136,31,144,31,247,31,60,31,40,31,40,30,40,29,40,28,230,31,185,31,173,31,173,30,244,31,244,30,61,31,82,31,169,31,44,31,110,31,69,31,208,31,247,31,53,31,53,30,109,31,116,31,201,31,198,31,134,31,65,31,65,30,65,29,65,28,125,31,125,30,102,31,207,31,117,31,29,31,155,31,68,31,84,31,135,31,135,30,238,31,238,30,123,31,236,31,23,31,157,31,43,31,97,31,94,31,50,31,145,31,197,31,251,31,220,31,100,31,100,30,228,31,171,31,187,31,187,30,156,31,156,30,9,31,25,31,25,30,25,29,189,31,183,31,111,31,127,31,176,31,139,31,4,31,4,30,4,29,252,31,9,31,139,31,174,31,244,31,59,31,167,31,60,31,212,31,191,31,191,30,191,29,135,31,181,31,181,30,181,29,209,31,117,31,109,31,109,30,132,31,245,31,26,31,220,31,8,31,85,31,68,31,152,31,137,31,55,31,48,31,199,31,199,30,199,29,53,31,41,31,109,31,117,31,138,31,27,31,129,31,181,31,64,31,64,30,249,31,161,31,161,30,57,31,199,31,144,31,144,30,61,31,230,31,178,31,238,31,214,31,76,31,123,31,150,31,150,30,224,31,224,30,31,31,55,31,55,30,45,31,48,31,186,31,86,31,55,31,252,31,180,31,80,31,80,30,217,31,41,31,44,31,56,31,134,31,240,31,131,31,131,31,118,31,118,30,226,31,211,31,135,31,253,31,181,31,57,31,154,31,154,30,192,31,56,31,56,30,87,31,21,31,21,30,156,31,156,30,67,31,67,30,67,29,103,31,144,31,124,31,124,30,53,31,53,30,151,31,151,30,222,31,43,31,134,31,92,31,31,31,12,31,56,31,185,31,116,31,161,31,161,30,55,31,176,31,176,30,86,31,229,31,133,31,133,30,10,31,122,31,197,31,197,30,149,31,149,30,217,31,1,31,1,30,188,31,188,30,179,31,179,30,6,31,104,31,81,31,44,31,125,31,36,31,83,31,222,31,2,31,216,31,216,30,162,31,11,31,193,31,75,31,193,31,78,31,253,31,135,31,237,31,88,31,219,31,219,30,52,31,52,30,63,31,174,31,174,30,130,31,110,31,69,31,12,31,57,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
