-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_70 is
end project_tb_70;

architecture project_tb_arch_70 of project_tb_70 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 199;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,236,0,82,0,198,0,2,0,119,0,195,0,0,0,0,0,132,0,0,0,249,0,54,0,98,0,165,0,0,0,30,0,0,0,213,0,172,0,97,0,54,0,75,0,0,0,140,0,66,0,147,0,0,0,94,0,146,0,92,0,219,0,0,0,112,0,169,0,112,0,200,0,0,0,228,0,58,0,227,0,126,0,30,0,75,0,115,0,0,0,30,0,112,0,0,0,227,0,194,0,149,0,56,0,0,0,230,0,227,0,3,0,145,0,0,0,0,0,251,0,0,0,173,0,108,0,183,0,0,0,38,0,220,0,141,0,56,0,179,0,20,0,214,0,183,0,249,0,212,0,123,0,117,0,231,0,0,0,244,0,220,0,46,0,236,0,10,0,1,0,83,0,74,0,79,0,249,0,182,0,12,0,38,0,130,0,142,0,107,0,203,0,37,0,44,0,0,0,248,0,117,0,188,0,16,0,49,0,189,0,99,0,125,0,240,0,120,0,144,0,0,0,232,0,152,0,193,0,195,0,166,0,171,0,0,0,127,0,0,0,0,0,132,0,132,0,0,0,178,0,19,0,0,0,179,0,166,0,0,0,9,0,66,0,34,0,110,0,75,0,227,0,94,0,27,0,82,0,178,0,175,0,238,0,57,0,236,0,0,0,253,0,34,0,210,0,153,0,0,0,146,0,61,0,243,0,168,0,13,0,184,0,191,0,51,0,165,0,0,0,93,0,212,0,223,0,0,0,78,0,4,0,0,0,12,0,0,0,0,0,58,0,0,0,144,0,162,0,0,0,110,0,138,0,0,0,119,0,0,0,252,0,0,0,169,0,155,0,71,0,109,0,154,0,0,0,180,0,25,0,0,0,115,0,166,0,222,0,44,0,94,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,236,31,82,31,198,31,2,31,119,31,195,31,195,30,195,29,132,31,132,30,249,31,54,31,98,31,165,31,165,30,30,31,30,30,213,31,172,31,97,31,54,31,75,31,75,30,140,31,66,31,147,31,147,30,94,31,146,31,92,31,219,31,219,30,112,31,169,31,112,31,200,31,200,30,228,31,58,31,227,31,126,31,30,31,75,31,115,31,115,30,30,31,112,31,112,30,227,31,194,31,149,31,56,31,56,30,230,31,227,31,3,31,145,31,145,30,145,29,251,31,251,30,173,31,108,31,183,31,183,30,38,31,220,31,141,31,56,31,179,31,20,31,214,31,183,31,249,31,212,31,123,31,117,31,231,31,231,30,244,31,220,31,46,31,236,31,10,31,1,31,83,31,74,31,79,31,249,31,182,31,12,31,38,31,130,31,142,31,107,31,203,31,37,31,44,31,44,30,248,31,117,31,188,31,16,31,49,31,189,31,99,31,125,31,240,31,120,31,144,31,144,30,232,31,152,31,193,31,195,31,166,31,171,31,171,30,127,31,127,30,127,29,132,31,132,31,132,30,178,31,19,31,19,30,179,31,166,31,166,30,9,31,66,31,34,31,110,31,75,31,227,31,94,31,27,31,82,31,178,31,175,31,238,31,57,31,236,31,236,30,253,31,34,31,210,31,153,31,153,30,146,31,61,31,243,31,168,31,13,31,184,31,191,31,51,31,165,31,165,30,93,31,212,31,223,31,223,30,78,31,4,31,4,30,12,31,12,30,12,29,58,31,58,30,144,31,162,31,162,30,110,31,138,31,138,30,119,31,119,30,252,31,252,30,169,31,155,31,71,31,109,31,154,31,154,30,180,31,25,31,25,30,115,31,166,31,222,31,44,31,94,31,94,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
