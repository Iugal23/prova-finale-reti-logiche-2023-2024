-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 896;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,200,0,0,0,92,0,233,0,229,0,123,0,190,0,228,0,233,0,23,0,150,0,14,0,243,0,74,0,83,0,251,0,240,0,156,0,147,0,60,0,165,0,249,0,0,0,104,0,218,0,79,0,0,0,186,0,200,0,25,0,0,0,100,0,123,0,0,0,17,0,239,0,22,0,233,0,108,0,4,0,0,0,0,0,27,0,0,0,198,0,169,0,113,0,201,0,116,0,126,0,93,0,28,0,246,0,0,0,145,0,166,0,0,0,72,0,59,0,24,0,49,0,209,0,219,0,248,0,230,0,226,0,74,0,214,0,123,0,221,0,0,0,52,0,48,0,0,0,113,0,103,0,230,0,193,0,85,0,128,0,47,0,249,0,247,0,201,0,177,0,0,0,63,0,185,0,0,0,69,0,135,0,0,0,140,0,0,0,164,0,22,0,198,0,108,0,122,0,164,0,0,0,160,0,100,0,139,0,205,0,0,0,0,0,143,0,207,0,83,0,0,0,166,0,158,0,1,0,59,0,0,0,0,0,10,0,166,0,0,0,180,0,0,0,179,0,134,0,107,0,245,0,62,0,172,0,254,0,101,0,0,0,88,0,0,0,35,0,0,0,0,0,3,0,71,0,0,0,191,0,128,0,0,0,247,0,248,0,138,0,0,0,250,0,128,0,117,0,49,0,113,0,168,0,244,0,198,0,84,0,200,0,148,0,0,0,3,0,166,0,0,0,0,0,147,0,219,0,251,0,237,0,238,0,80,0,71,0,0,0,181,0,217,0,0,0,247,0,178,0,0,0,39,0,237,0,99,0,0,0,243,0,90,0,45,0,239,0,100,0,189,0,0,0,0,0,173,0,200,0,43,0,205,0,201,0,171,0,206,0,6,0,152,0,88,0,2,0,115,0,18,0,214,0,173,0,253,0,18,0,118,0,219,0,86,0,35,0,81,0,196,0,164,0,109,0,164,0,185,0,72,0,207,0,0,0,45,0,127,0,79,0,112,0,203,0,178,0,126,0,115,0,104,0,193,0,77,0,213,0,101,0,136,0,0,0,113,0,91,0,20,0,100,0,208,0,197,0,0,0,127,0,231,0,86,0,0,0,15,0,75,0,227,0,142,0,84,0,79,0,51,0,223,0,24,0,127,0,195,0,35,0,79,0,0,0,239,0,198,0,68,0,39,0,0,0,230,0,181,0,224,0,144,0,0,0,160,0,50,0,0,0,0,0,230,0,232,0,157,0,173,0,114,0,0,0,233,0,238,0,36,0,0,0,255,0,222,0,0,0,40,0,9,0,210,0,0,0,24,0,110,0,178,0,133,0,59,0,79,0,16,0,158,0,118,0,204,0,103,0,0,0,253,0,42,0,29,0,80,0,77,0,0,0,81,0,119,0,62,0,0,0,150,0,76,0,13,0,76,0,60,0,255,0,168,0,0,0,255,0,124,0,136,0,252,0,199,0,16,0,142,0,42,0,192,0,139,0,217,0,163,0,65,0,164,0,5,0,108,0,196,0,35,0,148,0,195,0,0,0,178,0,20,0,107,0,51,0,213,0,0,0,222,0,147,0,0,0,104,0,156,0,185,0,115,0,211,0,48,0,255,0,22,0,0,0,201,0,66,0,41,0,91,0,0,0,164,0,140,0,22,0,181,0,58,0,61,0,68,0,84,0,80,0,139,0,79,0,232,0,230,0,0,0,21,0,0,0,82,0,133,0,90,0,77,0,79,0,163,0,9,0,77,0,93,0,56,0,0,0,55,0,142,0,157,0,188,0,82,0,116,0,18,0,102,0,246,0,0,0,28,0,116,0,147,0,41,0,249,0,170,0,12,0,218,0,103,0,80,0,101,0,108,0,44,0,98,0,149,0,83,0,77,0,76,0,0,0,48,0,225,0,253,0,216,0,7,0,202,0,221,0,144,0,108,0,163,0,184,0,0,0,0,0,203,0,120,0,204,0,77,0,126,0,99,0,29,0,248,0,0,0,230,0,0,0,0,0,105,0,90,0,93,0,0,0,0,0,0,0,185,0,255,0,48,0,183,0,70,0,247,0,69,0,104,0,205,0,164,0,0,0,137,0,56,0,0,0,145,0,246,0,233,0,176,0,150,0,0,0,0,0,153,0,76,0,246,0,181,0,57,0,59,0,54,0,0,0,122,0,226,0,22,0,7,0,0,0,0,0,52,0,73,0,0,0,126,0,12,0,127,0,89,0,52,0,148,0,174,0,157,0,168,0,14,0,156,0,175,0,0,0,154,0,54,0,71,0,176,0,135,0,204,0,247,0,166,0,92,0,138,0,108,0,124,0,249,0,24,0,0,0,0,0,150,0,233,0,0,0,165,0,221,0,0,0,0,0,0,0,226,0,158,0,6,0,19,0,226,0,196,0,85,0,5,0,63,0,143,0,49,0,189,0,76,0,163,0,0,0,0,0,37,0,91,0,153,0,151,0,75,0,210,0,0,0,205,0,0,0,130,0,78,0,10,0,0,0,0,0,230,0,110,0,139,0,0,0,27,0,114,0,253,0,138,0,0,0,158,0,0,0,139,0,132,0,236,0,53,0,32,0,124,0,241,0,0,0,0,0,170,0,163,0,186,0,184,0,206,0,0,0,194,0,0,0,0,0,79,0,93,0,187,0,0,0,13,0,0,0,198,0,0,0,240,0,49,0,0,0,157,0,73,0,0,0,130,0,180,0,231,0,202,0,231,0,232,0,100,0,96,0,32,0,113,0,0,0,85,0,148,0,29,0,200,0,179,0,186,0,154,0,71,0,23,0,213,0,108,0,149,0,230,0,219,0,38,0,0,0,142,0,11,0,0,0,0,0,0,0,159,0,9,0,233,0,1,0,243,0,0,0,108,0,0,0,0,0,6,0,97,0,0,0,185,0,0,0,220,0,220,0,65,0,251,0,107,0,89,0,10,0,170,0,35,0,142,0,92,0,100,0,46,0,0,0,123,0,1,0,172,0,100,0,23,0,132,0,22,0,143,0,101,0,177,0,219,0,218,0,5,0,126,0,99,0,252,0,119,0,158,0,249,0,87,0,51,0,0,0,251,0,218,0,246,0,106,0,71,0,204,0,246,0,45,0,190,0,138,0,3,0,208,0,108,0,136,0,179,0,35,0,55,0,47,0,193,0,0,0,176,0,200,0,213,0,123,0,84,0,0,0,2,0,48,0,120,0,50,0,62,0,26,0,239,0,149,0,207,0,158,0,227,0,52,0,124,0,151,0,20,0,144,0,92,0,114,0,170,0,131,0,100,0,0,0,118,0,169,0,76,0,0,0,124,0,160,0,185,0,140,0,17,0,190,0,158,0,35,0,176,0,65,0,234,0,27,0,27,0,172,0,163,0,230,0,97,0,56,0,76,0,136,0,108,0,217,0,141,0,226,0,6,0,49,0,0,0,117,0,36,0,125,0,0,0,34,0,88,0,158,0,42,0,118,0,84,0,150,0,91,0,156,0,143,0,206,0,95,0,0,0,206,0,164,0,0,0,13,0,245,0,29,0,125,0,0,0,0,0,81,0,0,0,158,0,0,0,3,0,0,0,111,0,0,0,95,0,80,0,0,0,35,0,34,0,58,0,145,0,180,0,169,0,20,0,112,0,0,0,167,0,0,0,239,0,152,0,0,0,205,0,0,0,181,0,0,0,70,0,106,0,202,0,0,0,71,0,142,0,23,0,130,0,187,0,249,0,17,0,191,0,46,0,223,0,16,0,255,0,199,0,0,0,0,0,196,0,0,0,30,0,15,0,0,0,38,0,61,0,8,0,62,0,145,0,46,0,160,0,186,0,0,0,0,0,117,0,179,0,0,0,10,0,238,0,133,0,0,0,153,0,47,0,34,0,0,0,120,0,246,0,0,0,0,0,151,0,47,0,237,0,201,0,74,0,195,0,124,0,177,0,121,0,0,0,1,0,6,0,64,0,84,0,188,0,40,0,0,0,62,0,173,0,20,0,23,0,53,0,154,0,83,0,134,0,146,0,81,0,16,0,46,0,0,0,186,0,80,0);
signal scenario_full  : scenario_type := (102,31,200,31,200,30,92,31,233,31,229,31,123,31,190,31,228,31,233,31,23,31,150,31,14,31,243,31,74,31,83,31,251,31,240,31,156,31,147,31,60,31,165,31,249,31,249,30,104,31,218,31,79,31,79,30,186,31,200,31,25,31,25,30,100,31,123,31,123,30,17,31,239,31,22,31,233,31,108,31,4,31,4,30,4,29,27,31,27,30,198,31,169,31,113,31,201,31,116,31,126,31,93,31,28,31,246,31,246,30,145,31,166,31,166,30,72,31,59,31,24,31,49,31,209,31,219,31,248,31,230,31,226,31,74,31,214,31,123,31,221,31,221,30,52,31,48,31,48,30,113,31,103,31,230,31,193,31,85,31,128,31,47,31,249,31,247,31,201,31,177,31,177,30,63,31,185,31,185,30,69,31,135,31,135,30,140,31,140,30,164,31,22,31,198,31,108,31,122,31,164,31,164,30,160,31,100,31,139,31,205,31,205,30,205,29,143,31,207,31,83,31,83,30,166,31,158,31,1,31,59,31,59,30,59,29,10,31,166,31,166,30,180,31,180,30,179,31,134,31,107,31,245,31,62,31,172,31,254,31,101,31,101,30,88,31,88,30,35,31,35,30,35,29,3,31,71,31,71,30,191,31,128,31,128,30,247,31,248,31,138,31,138,30,250,31,128,31,117,31,49,31,113,31,168,31,244,31,198,31,84,31,200,31,148,31,148,30,3,31,166,31,166,30,166,29,147,31,219,31,251,31,237,31,238,31,80,31,71,31,71,30,181,31,217,31,217,30,247,31,178,31,178,30,39,31,237,31,99,31,99,30,243,31,90,31,45,31,239,31,100,31,189,31,189,30,189,29,173,31,200,31,43,31,205,31,201,31,171,31,206,31,6,31,152,31,88,31,2,31,115,31,18,31,214,31,173,31,253,31,18,31,118,31,219,31,86,31,35,31,81,31,196,31,164,31,109,31,164,31,185,31,72,31,207,31,207,30,45,31,127,31,79,31,112,31,203,31,178,31,126,31,115,31,104,31,193,31,77,31,213,31,101,31,136,31,136,30,113,31,91,31,20,31,100,31,208,31,197,31,197,30,127,31,231,31,86,31,86,30,15,31,75,31,227,31,142,31,84,31,79,31,51,31,223,31,24,31,127,31,195,31,35,31,79,31,79,30,239,31,198,31,68,31,39,31,39,30,230,31,181,31,224,31,144,31,144,30,160,31,50,31,50,30,50,29,230,31,232,31,157,31,173,31,114,31,114,30,233,31,238,31,36,31,36,30,255,31,222,31,222,30,40,31,9,31,210,31,210,30,24,31,110,31,178,31,133,31,59,31,79,31,16,31,158,31,118,31,204,31,103,31,103,30,253,31,42,31,29,31,80,31,77,31,77,30,81,31,119,31,62,31,62,30,150,31,76,31,13,31,76,31,60,31,255,31,168,31,168,30,255,31,124,31,136,31,252,31,199,31,16,31,142,31,42,31,192,31,139,31,217,31,163,31,65,31,164,31,5,31,108,31,196,31,35,31,148,31,195,31,195,30,178,31,20,31,107,31,51,31,213,31,213,30,222,31,147,31,147,30,104,31,156,31,185,31,115,31,211,31,48,31,255,31,22,31,22,30,201,31,66,31,41,31,91,31,91,30,164,31,140,31,22,31,181,31,58,31,61,31,68,31,84,31,80,31,139,31,79,31,232,31,230,31,230,30,21,31,21,30,82,31,133,31,90,31,77,31,79,31,163,31,9,31,77,31,93,31,56,31,56,30,55,31,142,31,157,31,188,31,82,31,116,31,18,31,102,31,246,31,246,30,28,31,116,31,147,31,41,31,249,31,170,31,12,31,218,31,103,31,80,31,101,31,108,31,44,31,98,31,149,31,83,31,77,31,76,31,76,30,48,31,225,31,253,31,216,31,7,31,202,31,221,31,144,31,108,31,163,31,184,31,184,30,184,29,203,31,120,31,204,31,77,31,126,31,99,31,29,31,248,31,248,30,230,31,230,30,230,29,105,31,90,31,93,31,93,30,93,29,93,28,185,31,255,31,48,31,183,31,70,31,247,31,69,31,104,31,205,31,164,31,164,30,137,31,56,31,56,30,145,31,246,31,233,31,176,31,150,31,150,30,150,29,153,31,76,31,246,31,181,31,57,31,59,31,54,31,54,30,122,31,226,31,22,31,7,31,7,30,7,29,52,31,73,31,73,30,126,31,12,31,127,31,89,31,52,31,148,31,174,31,157,31,168,31,14,31,156,31,175,31,175,30,154,31,54,31,71,31,176,31,135,31,204,31,247,31,166,31,92,31,138,31,108,31,124,31,249,31,24,31,24,30,24,29,150,31,233,31,233,30,165,31,221,31,221,30,221,29,221,28,226,31,158,31,6,31,19,31,226,31,196,31,85,31,5,31,63,31,143,31,49,31,189,31,76,31,163,31,163,30,163,29,37,31,91,31,153,31,151,31,75,31,210,31,210,30,205,31,205,30,130,31,78,31,10,31,10,30,10,29,230,31,110,31,139,31,139,30,27,31,114,31,253,31,138,31,138,30,158,31,158,30,139,31,132,31,236,31,53,31,32,31,124,31,241,31,241,30,241,29,170,31,163,31,186,31,184,31,206,31,206,30,194,31,194,30,194,29,79,31,93,31,187,31,187,30,13,31,13,30,198,31,198,30,240,31,49,31,49,30,157,31,73,31,73,30,130,31,180,31,231,31,202,31,231,31,232,31,100,31,96,31,32,31,113,31,113,30,85,31,148,31,29,31,200,31,179,31,186,31,154,31,71,31,23,31,213,31,108,31,149,31,230,31,219,31,38,31,38,30,142,31,11,31,11,30,11,29,11,28,159,31,9,31,233,31,1,31,243,31,243,30,108,31,108,30,108,29,6,31,97,31,97,30,185,31,185,30,220,31,220,31,65,31,251,31,107,31,89,31,10,31,170,31,35,31,142,31,92,31,100,31,46,31,46,30,123,31,1,31,172,31,100,31,23,31,132,31,22,31,143,31,101,31,177,31,219,31,218,31,5,31,126,31,99,31,252,31,119,31,158,31,249,31,87,31,51,31,51,30,251,31,218,31,246,31,106,31,71,31,204,31,246,31,45,31,190,31,138,31,3,31,208,31,108,31,136,31,179,31,35,31,55,31,47,31,193,31,193,30,176,31,200,31,213,31,123,31,84,31,84,30,2,31,48,31,120,31,50,31,62,31,26,31,239,31,149,31,207,31,158,31,227,31,52,31,124,31,151,31,20,31,144,31,92,31,114,31,170,31,131,31,100,31,100,30,118,31,169,31,76,31,76,30,124,31,160,31,185,31,140,31,17,31,190,31,158,31,35,31,176,31,65,31,234,31,27,31,27,31,172,31,163,31,230,31,97,31,56,31,76,31,136,31,108,31,217,31,141,31,226,31,6,31,49,31,49,30,117,31,36,31,125,31,125,30,34,31,88,31,158,31,42,31,118,31,84,31,150,31,91,31,156,31,143,31,206,31,95,31,95,30,206,31,164,31,164,30,13,31,245,31,29,31,125,31,125,30,125,29,81,31,81,30,158,31,158,30,3,31,3,30,111,31,111,30,95,31,80,31,80,30,35,31,34,31,58,31,145,31,180,31,169,31,20,31,112,31,112,30,167,31,167,30,239,31,152,31,152,30,205,31,205,30,181,31,181,30,70,31,106,31,202,31,202,30,71,31,142,31,23,31,130,31,187,31,249,31,17,31,191,31,46,31,223,31,16,31,255,31,199,31,199,30,199,29,196,31,196,30,30,31,15,31,15,30,38,31,61,31,8,31,62,31,145,31,46,31,160,31,186,31,186,30,186,29,117,31,179,31,179,30,10,31,238,31,133,31,133,30,153,31,47,31,34,31,34,30,120,31,246,31,246,30,246,29,151,31,47,31,237,31,201,31,74,31,195,31,124,31,177,31,121,31,121,30,1,31,6,31,64,31,84,31,188,31,40,31,40,30,62,31,173,31,20,31,23,31,53,31,154,31,83,31,134,31,146,31,81,31,16,31,46,31,46,30,186,31,80,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
