-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_301 is
end project_tb_301;

architecture project_tb_arch_301 of project_tb_301 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 655;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,251,0,96,0,201,0,0,0,0,0,197,0,0,0,210,0,0,0,100,0,74,0,71,0,184,0,1,0,242,0,187,0,0,0,8,0,80,0,201,0,198,0,77,0,202,0,182,0,251,0,236,0,195,0,172,0,186,0,158,0,8,0,15,0,186,0,8,0,13,0,116,0,151,0,142,0,65,0,0,0,138,0,0,0,151,0,230,0,160,0,173,0,129,0,96,0,216,0,244,0,128,0,236,0,0,0,149,0,72,0,143,0,242,0,101,0,47,0,0,0,254,0,229,0,130,0,0,0,0,0,75,0,99,0,94,0,163,0,173,0,22,0,0,0,225,0,131,0,0,0,254,0,107,0,69,0,93,0,105,0,37,0,77,0,164,0,170,0,195,0,0,0,232,0,0,0,238,0,21,0,53,0,245,0,0,0,146,0,217,0,81,0,134,0,66,0,154,0,0,0,71,0,62,0,0,0,122,0,198,0,253,0,40,0,71,0,156,0,183,0,112,0,0,0,183,0,120,0,54,0,0,0,56,0,23,0,0,0,54,0,123,0,158,0,111,0,203,0,86,0,206,0,207,0,50,0,255,0,73,0,0,0,78,0,167,0,21,0,146,0,110,0,156,0,179,0,158,0,188,0,135,0,0,0,166,0,209,0,247,0,97,0,196,0,106,0,119,0,192,0,74,0,130,0,161,0,119,0,114,0,213,0,179,0,150,0,23,0,0,0,239,0,151,0,0,0,89,0,155,0,167,0,137,0,184,0,154,0,253,0,0,0,0,0,0,0,0,0,244,0,243,0,203,0,37,0,120,0,203,0,227,0,182,0,0,0,135,0,0,0,177,0,230,0,90,0,39,0,0,0,76,0,106,0,57,0,221,0,182,0,21,0,119,0,0,0,0,0,0,0,219,0,194,0,0,0,7,0,166,0,254,0,204,0,0,0,244,0,30,0,51,0,233,0,0,0,247,0,65,0,74,0,171,0,0,0,0,0,170,0,0,0,22,0,249,0,38,0,245,0,214,0,116,0,98,0,184,0,209,0,0,0,134,0,201,0,0,0,0,0,0,0,138,0,119,0,18,0,0,0,215,0,13,0,22,0,110,0,10,0,0,0,0,0,0,0,182,0,0,0,0,0,226,0,115,0,84,0,173,0,126,0,0,0,255,0,242,0,10,0,0,0,3,0,0,0,208,0,200,0,83,0,154,0,79,0,94,0,25,0,94,0,111,0,0,0,23,0,111,0,121,0,0,0,216,0,161,0,243,0,0,0,89,0,80,0,146,0,218,0,198,0,196,0,155,0,248,0,37,0,0,0,165,0,53,0,0,0,113,0,10,0,135,0,178,0,194,0,20,0,0,0,0,0,222,0,0,0,99,0,163,0,124,0,202,0,0,0,96,0,248,0,186,0,241,0,20,0,0,0,193,0,7,0,29,0,38,0,135,0,57,0,145,0,58,0,158,0,0,0,119,0,167,0,100,0,112,0,204,0,115,0,0,0,194,0,52,0,212,0,251,0,37,0,0,0,215,0,0,0,175,0,0,0,69,0,0,0,100,0,11,0,64,0,144,0,18,0,141,0,91,0,77,0,186,0,20,0,176,0,139,0,230,0,0,0,235,0,219,0,0,0,75,0,0,0,157,0,43,0,70,0,195,0,49,0,0,0,59,0,0,0,0,0,227,0,229,0,35,0,255,0,202,0,106,0,178,0,194,0,0,0,0,0,61,0,158,0,0,0,77,0,241,0,160,0,81,0,13,0,0,0,187,0,154,0,92,0,190,0,161,0,168,0,215,0,238,0,0,0,39,0,91,0,49,0,38,0,109,0,117,0,15,0,138,0,57,0,87,0,72,0,217,0,147,0,0,0,249,0,227,0,171,0,32,0,87,0,40,0,243,0,234,0,177,0,212,0,207,0,0,0,64,0,224,0,243,0,167,0,173,0,73,0,105,0,172,0,254,0,216,0,0,0,178,0,228,0,184,0,0,0,106,0,53,0,5,0,155,0,106,0,209,0,1,0,0,0,209,0,77,0,0,0,0,0,192,0,0,0,107,0,27,0,13,0,60,0,63,0,195,0,129,0,47,0,0,0,0,0,216,0,237,0,74,0,175,0,154,0,126,0,0,0,178,0,61,0,175,0,0,0,142,0,116,0,134,0,83,0,0,0,249,0,255,0,0,0,48,0,0,0,0,0,39,0,51,0,17,0,126,0,155,0,236,0,35,0,171,0,168,0,240,0,173,0,44,0,33,0,8,0,0,0,97,0,238,0,192,0,100,0,0,0,109,0,24,0,91,0,152,0,123,0,0,0,109,0,128,0,166,0,0,0,141,0,236,0,23,0,0,0,253,0,44,0,5,0,49,0,44,0,0,0,0,0,206,0,0,0,121,0,125,0,38,0,44,0,37,0,97,0,0,0,248,0,190,0,253,0,219,0,139,0,6,0,173,0,0,0,211,0,0,0,24,0,209,0,150,0,243,0,0,0,105,0,14,0,9,0,190,0,31,0,18,0,2,0,0,0,0,0,21,0,80,0,102,0,210,0,242,0,0,0,201,0,108,0,0,0,33,0,214,0,242,0,17,0,0,0,28,0,254,0,0,0,0,0,122,0,180,0,195,0,157,0,154,0,56,0,86,0,82,0,234,0,203,0,8,0,192,0,123,0,199,0,8,0,0,0,203,0,106,0,227,0,112,0,0,0,0,0,144,0,2,0,131,0,79,0,33,0,67,0,49,0,60,0,56,0,44,0,64,0,127,0,196,0,64,0,66,0,0,0,238,0,154,0,0,0,7,0,0,0,252,0,127,0,179,0,141,0,69,0,214,0,0,0,30,0,0,0,69,0,200,0,94,0,151,0,42,0,161,0,0,0,101,0,172,0,0,0,249,0,0,0,138,0,185,0,67,0,6,0,149,0,179,0,38,0,182,0,51,0,105,0,243,0);
signal scenario_full  : scenario_type := (0,0,251,31,96,31,201,31,201,30,201,29,197,31,197,30,210,31,210,30,100,31,74,31,71,31,184,31,1,31,242,31,187,31,187,30,8,31,80,31,201,31,198,31,77,31,202,31,182,31,251,31,236,31,195,31,172,31,186,31,158,31,8,31,15,31,186,31,8,31,13,31,116,31,151,31,142,31,65,31,65,30,138,31,138,30,151,31,230,31,160,31,173,31,129,31,96,31,216,31,244,31,128,31,236,31,236,30,149,31,72,31,143,31,242,31,101,31,47,31,47,30,254,31,229,31,130,31,130,30,130,29,75,31,99,31,94,31,163,31,173,31,22,31,22,30,225,31,131,31,131,30,254,31,107,31,69,31,93,31,105,31,37,31,77,31,164,31,170,31,195,31,195,30,232,31,232,30,238,31,21,31,53,31,245,31,245,30,146,31,217,31,81,31,134,31,66,31,154,31,154,30,71,31,62,31,62,30,122,31,198,31,253,31,40,31,71,31,156,31,183,31,112,31,112,30,183,31,120,31,54,31,54,30,56,31,23,31,23,30,54,31,123,31,158,31,111,31,203,31,86,31,206,31,207,31,50,31,255,31,73,31,73,30,78,31,167,31,21,31,146,31,110,31,156,31,179,31,158,31,188,31,135,31,135,30,166,31,209,31,247,31,97,31,196,31,106,31,119,31,192,31,74,31,130,31,161,31,119,31,114,31,213,31,179,31,150,31,23,31,23,30,239,31,151,31,151,30,89,31,155,31,167,31,137,31,184,31,154,31,253,31,253,30,253,29,253,28,253,27,244,31,243,31,203,31,37,31,120,31,203,31,227,31,182,31,182,30,135,31,135,30,177,31,230,31,90,31,39,31,39,30,76,31,106,31,57,31,221,31,182,31,21,31,119,31,119,30,119,29,119,28,219,31,194,31,194,30,7,31,166,31,254,31,204,31,204,30,244,31,30,31,51,31,233,31,233,30,247,31,65,31,74,31,171,31,171,30,171,29,170,31,170,30,22,31,249,31,38,31,245,31,214,31,116,31,98,31,184,31,209,31,209,30,134,31,201,31,201,30,201,29,201,28,138,31,119,31,18,31,18,30,215,31,13,31,22,31,110,31,10,31,10,30,10,29,10,28,182,31,182,30,182,29,226,31,115,31,84,31,173,31,126,31,126,30,255,31,242,31,10,31,10,30,3,31,3,30,208,31,200,31,83,31,154,31,79,31,94,31,25,31,94,31,111,31,111,30,23,31,111,31,121,31,121,30,216,31,161,31,243,31,243,30,89,31,80,31,146,31,218,31,198,31,196,31,155,31,248,31,37,31,37,30,165,31,53,31,53,30,113,31,10,31,135,31,178,31,194,31,20,31,20,30,20,29,222,31,222,30,99,31,163,31,124,31,202,31,202,30,96,31,248,31,186,31,241,31,20,31,20,30,193,31,7,31,29,31,38,31,135,31,57,31,145,31,58,31,158,31,158,30,119,31,167,31,100,31,112,31,204,31,115,31,115,30,194,31,52,31,212,31,251,31,37,31,37,30,215,31,215,30,175,31,175,30,69,31,69,30,100,31,11,31,64,31,144,31,18,31,141,31,91,31,77,31,186,31,20,31,176,31,139,31,230,31,230,30,235,31,219,31,219,30,75,31,75,30,157,31,43,31,70,31,195,31,49,31,49,30,59,31,59,30,59,29,227,31,229,31,35,31,255,31,202,31,106,31,178,31,194,31,194,30,194,29,61,31,158,31,158,30,77,31,241,31,160,31,81,31,13,31,13,30,187,31,154,31,92,31,190,31,161,31,168,31,215,31,238,31,238,30,39,31,91,31,49,31,38,31,109,31,117,31,15,31,138,31,57,31,87,31,72,31,217,31,147,31,147,30,249,31,227,31,171,31,32,31,87,31,40,31,243,31,234,31,177,31,212,31,207,31,207,30,64,31,224,31,243,31,167,31,173,31,73,31,105,31,172,31,254,31,216,31,216,30,178,31,228,31,184,31,184,30,106,31,53,31,5,31,155,31,106,31,209,31,1,31,1,30,209,31,77,31,77,30,77,29,192,31,192,30,107,31,27,31,13,31,60,31,63,31,195,31,129,31,47,31,47,30,47,29,216,31,237,31,74,31,175,31,154,31,126,31,126,30,178,31,61,31,175,31,175,30,142,31,116,31,134,31,83,31,83,30,249,31,255,31,255,30,48,31,48,30,48,29,39,31,51,31,17,31,126,31,155,31,236,31,35,31,171,31,168,31,240,31,173,31,44,31,33,31,8,31,8,30,97,31,238,31,192,31,100,31,100,30,109,31,24,31,91,31,152,31,123,31,123,30,109,31,128,31,166,31,166,30,141,31,236,31,23,31,23,30,253,31,44,31,5,31,49,31,44,31,44,30,44,29,206,31,206,30,121,31,125,31,38,31,44,31,37,31,97,31,97,30,248,31,190,31,253,31,219,31,139,31,6,31,173,31,173,30,211,31,211,30,24,31,209,31,150,31,243,31,243,30,105,31,14,31,9,31,190,31,31,31,18,31,2,31,2,30,2,29,21,31,80,31,102,31,210,31,242,31,242,30,201,31,108,31,108,30,33,31,214,31,242,31,17,31,17,30,28,31,254,31,254,30,254,29,122,31,180,31,195,31,157,31,154,31,56,31,86,31,82,31,234,31,203,31,8,31,192,31,123,31,199,31,8,31,8,30,203,31,106,31,227,31,112,31,112,30,112,29,144,31,2,31,131,31,79,31,33,31,67,31,49,31,60,31,56,31,44,31,64,31,127,31,196,31,64,31,66,31,66,30,238,31,154,31,154,30,7,31,7,30,252,31,127,31,179,31,141,31,69,31,214,31,214,30,30,31,30,30,69,31,200,31,94,31,151,31,42,31,161,31,161,30,101,31,172,31,172,30,249,31,249,30,138,31,185,31,67,31,6,31,149,31,179,31,38,31,182,31,51,31,105,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
