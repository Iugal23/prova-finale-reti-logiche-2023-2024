-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 334;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,0,0,56,0,80,0,234,0,0,0,0,0,0,0,132,0,246,0,232,0,151,0,133,0,90,0,0,0,77,0,248,0,213,0,120,0,76,0,74,0,26,0,0,0,206,0,0,0,68,0,34,0,212,0,247,0,220,0,190,0,210,0,41,0,0,0,0,0,51,0,0,0,9,0,122,0,186,0,0,0,103,0,0,0,181,0,0,0,200,0,199,0,2,0,0,0,130,0,43,0,69,0,0,0,239,0,0,0,174,0,62,0,235,0,170,0,39,0,58,0,170,0,68,0,190,0,133,0,178,0,34,0,21,0,44,0,60,0,220,0,183,0,239,0,189,0,0,0,59,0,210,0,89,0,104,0,90,0,13,0,8,0,0,0,0,0,91,0,142,0,240,0,103,0,36,0,0,0,221,0,207,0,0,0,216,0,35,0,146,0,29,0,0,0,2,0,219,0,189,0,186,0,65,0,242,0,117,0,155,0,102,0,184,0,119,0,237,0,10,0,135,0,229,0,231,0,245,0,231,0,0,0,33,0,0,0,66,0,53,0,182,0,218,0,117,0,0,0,134,0,84,0,142,0,196,0,170,0,202,0,93,0,0,0,0,0,10,0,195,0,78,0,210,0,219,0,0,0,7,0,210,0,128,0,0,0,0,0,0,0,111,0,170,0,0,0,35,0,23,0,78,0,243,0,79,0,31,0,251,0,0,0,203,0,182,0,0,0,108,0,251,0,156,0,201,0,0,0,75,0,0,0,29,0,0,0,104,0,145,0,0,0,169,0,255,0,75,0,139,0,66,0,83,0,165,0,115,0,0,0,211,0,228,0,124,0,130,0,21,0,189,0,0,0,187,0,29,0,32,0,67,0,0,0,105,0,229,0,34,0,117,0,151,0,56,0,53,0,250,0,0,0,166,0,82,0,224,0,179,0,143,0,119,0,0,0,147,0,221,0,0,0,228,0,0,0,0,0,181,0,236,0,0,0,43,0,113,0,0,0,53,0,102,0,57,0,51,0,236,0,0,0,54,0,0,0,33,0,44,0,188,0,8,0,0,0,56,0,55,0,0,0,21,0,0,0,193,0,39,0,216,0,17,0,189,0,224,0,102,0,239,0,152,0,189,0,213,0,119,0,183,0,20,0,0,0,212,0,140,0,247,0,94,0,60,0,172,0,0,0,98,0,178,0,45,0,217,0,170,0,30,0,3,0,231,0,197,0,162,0,42,0,51,0,189,0,111,0,16,0,255,0,65,0,27,0,242,0,243,0,197,0,0,0,48,0,27,0,26,0,79,0,116,0,224,0,241,0,100,0,153,0,0,0,177,0,233,0,147,0,74,0,96,0,162,0,243,0,197,0,67,0,105,0,120,0,245,0,0,0,251,0,0,0,0,0,46,0,0,0,93,0,209,0,24,0,0,0,82,0,169,0,169,0,10,0,144,0,180,0,109,0,0,0,233,0,0,0,7,0,197,0,21,0,0,0,229,0,155,0,142,0,200,0,0,0);
signal scenario_full  : scenario_type := (49,31,49,30,56,31,80,31,234,31,234,30,234,29,234,28,132,31,246,31,232,31,151,31,133,31,90,31,90,30,77,31,248,31,213,31,120,31,76,31,74,31,26,31,26,30,206,31,206,30,68,31,34,31,212,31,247,31,220,31,190,31,210,31,41,31,41,30,41,29,51,31,51,30,9,31,122,31,186,31,186,30,103,31,103,30,181,31,181,30,200,31,199,31,2,31,2,30,130,31,43,31,69,31,69,30,239,31,239,30,174,31,62,31,235,31,170,31,39,31,58,31,170,31,68,31,190,31,133,31,178,31,34,31,21,31,44,31,60,31,220,31,183,31,239,31,189,31,189,30,59,31,210,31,89,31,104,31,90,31,13,31,8,31,8,30,8,29,91,31,142,31,240,31,103,31,36,31,36,30,221,31,207,31,207,30,216,31,35,31,146,31,29,31,29,30,2,31,219,31,189,31,186,31,65,31,242,31,117,31,155,31,102,31,184,31,119,31,237,31,10,31,135,31,229,31,231,31,245,31,231,31,231,30,33,31,33,30,66,31,53,31,182,31,218,31,117,31,117,30,134,31,84,31,142,31,196,31,170,31,202,31,93,31,93,30,93,29,10,31,195,31,78,31,210,31,219,31,219,30,7,31,210,31,128,31,128,30,128,29,128,28,111,31,170,31,170,30,35,31,23,31,78,31,243,31,79,31,31,31,251,31,251,30,203,31,182,31,182,30,108,31,251,31,156,31,201,31,201,30,75,31,75,30,29,31,29,30,104,31,145,31,145,30,169,31,255,31,75,31,139,31,66,31,83,31,165,31,115,31,115,30,211,31,228,31,124,31,130,31,21,31,189,31,189,30,187,31,29,31,32,31,67,31,67,30,105,31,229,31,34,31,117,31,151,31,56,31,53,31,250,31,250,30,166,31,82,31,224,31,179,31,143,31,119,31,119,30,147,31,221,31,221,30,228,31,228,30,228,29,181,31,236,31,236,30,43,31,113,31,113,30,53,31,102,31,57,31,51,31,236,31,236,30,54,31,54,30,33,31,44,31,188,31,8,31,8,30,56,31,55,31,55,30,21,31,21,30,193,31,39,31,216,31,17,31,189,31,224,31,102,31,239,31,152,31,189,31,213,31,119,31,183,31,20,31,20,30,212,31,140,31,247,31,94,31,60,31,172,31,172,30,98,31,178,31,45,31,217,31,170,31,30,31,3,31,231,31,197,31,162,31,42,31,51,31,189,31,111,31,16,31,255,31,65,31,27,31,242,31,243,31,197,31,197,30,48,31,27,31,26,31,79,31,116,31,224,31,241,31,100,31,153,31,153,30,177,31,233,31,147,31,74,31,96,31,162,31,243,31,197,31,67,31,105,31,120,31,245,31,245,30,251,31,251,30,251,29,46,31,46,30,93,31,209,31,24,31,24,30,82,31,169,31,169,31,10,31,144,31,180,31,109,31,109,30,233,31,233,30,7,31,197,31,21,31,21,30,229,31,155,31,142,31,200,31,200,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
