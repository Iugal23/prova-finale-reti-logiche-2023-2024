-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 864;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (220,0,137,0,0,0,191,0,0,0,184,0,0,0,173,0,239,0,44,0,27,0,119,0,19,0,213,0,25,0,101,0,225,0,76,0,19,0,47,0,0,0,121,0,230,0,0,0,29,0,151,0,136,0,254,0,217,0,86,0,0,0,0,0,220,0,0,0,131,0,0,0,189,0,218,0,99,0,0,0,126,0,244,0,248,0,0,0,0,0,0,0,0,0,27,0,0,0,0,0,122,0,142,0,183,0,188,0,2,0,0,0,150,0,55,0,158,0,70,0,252,0,107,0,129,0,0,0,48,0,0,0,44,0,228,0,238,0,120,0,31,0,142,0,154,0,136,0,96,0,146,0,0,0,0,0,0,0,107,0,197,0,186,0,91,0,136,0,82,0,204,0,189,0,234,0,133,0,0,0,123,0,0,0,0,0,98,0,0,0,10,0,19,0,40,0,55,0,140,0,23,0,253,0,0,0,169,0,0,0,0,0,129,0,24,0,6,0,157,0,103,0,223,0,170,0,178,0,223,0,91,0,0,0,0,0,70,0,240,0,238,0,92,0,135,0,162,0,183,0,83,0,0,0,226,0,94,0,159,0,105,0,4,0,1,0,102,0,70,0,54,0,170,0,212,0,73,0,160,0,127,0,230,0,222,0,0,0,207,0,185,0,0,0,0,0,219,0,26,0,199,0,42,0,43,0,180,0,249,0,0,0,148,0,244,0,246,0,225,0,136,0,76,0,37,0,106,0,165,0,199,0,236,0,203,0,0,0,38,0,149,0,22,0,42,0,56,0,120,0,221,0,199,0,214,0,239,0,201,0,99,0,0,0,107,0,90,0,0,0,76,0,167,0,126,0,11,0,239,0,129,0,0,0,36,0,95,0,177,0,0,0,119,0,0,0,94,0,113,0,0,0,141,0,171,0,70,0,246,0,7,0,0,0,0,0,0,0,0,0,147,0,0,0,0,0,131,0,54,0,167,0,93,0,218,0,87,0,162,0,69,0,105,0,211,0,220,0,42,0,185,0,129,0,131,0,250,0,31,0,187,0,100,0,133,0,220,0,201,0,186,0,238,0,126,0,0,0,7,0,239,0,217,0,0,0,164,0,204,0,48,0,200,0,242,0,81,0,200,0,39,0,126,0,33,0,131,0,177,0,0,0,74,0,232,0,172,0,0,0,217,0,211,0,69,0,111,0,41,0,82,0,117,0,0,0,10,0,137,0,107,0,249,0,0,0,224,0,0,0,251,0,0,0,0,0,207,0,36,0,131,0,203,0,202,0,197,0,10,0,239,0,125,0,166,0,0,0,232,0,5,0,0,0,213,0,0,0,27,0,38,0,50,0,0,0,92,0,93,0,0,0,148,0,112,0,135,0,0,0,103,0,37,0,212,0,113,0,154,0,106,0,127,0,96,0,203,0,0,0,49,0,0,0,64,0,0,0,157,0,171,0,62,0,218,0,225,0,0,0,79,0,58,0,151,0,216,0,0,0,235,0,251,0,79,0,19,0,166,0,219,0,48,0,0,0,205,0,136,0,113,0,95,0,97,0,54,0,0,0,0,0,96,0,0,0,77,0,26,0,82,0,74,0,0,0,0,0,210,0,236,0,180,0,193,0,106,0,239,0,14,0,118,0,226,0,0,0,0,0,0,0,0,0,33,0,95,0,27,0,0,0,198,0,202,0,101,0,191,0,41,0,183,0,179,0,109,0,55,0,185,0,214,0,185,0,171,0,24,0,106,0,135,0,0,0,97,0,14,0,165,0,69,0,76,0,63,0,0,0,0,0,171,0,194,0,251,0,124,0,61,0,145,0,202,0,47,0,104,0,0,0,0,0,0,0,125,0,242,0,145,0,220,0,209,0,0,0,41,0,102,0,2,0,74,0,155,0,251,0,0,0,0,0,120,0,213,0,130,0,209,0,122,0,85,0,30,0,238,0,0,0,0,0,128,0,241,0,0,0,139,0,228,0,222,0,206,0,0,0,0,0,169,0,111,0,50,0,162,0,255,0,148,0,68,0,122,0,253,0,145,0,29,0,167,0,184,0,216,0,68,0,0,0,158,0,0,0,60,0,8,0,0,0,135,0,114,0,97,0,0,0,61,0,16,0,83,0,130,0,102,0,213,0,127,0,204,0,102,0,78,0,207,0,140,0,77,0,130,0,115,0,113,0,224,0,30,0,192,0,4,0,58,0,144,0,0,0,0,0,253,0,0,0,31,0,65,0,7,0,0,0,9,0,179,0,95,0,147,0,220,0,0,0,129,0,183,0,237,0,0,0,221,0,34,0,78,0,0,0,65,0,58,0,8,0,183,0,243,0,0,0,46,0,126,0,81,0,103,0,23,0,0,0,0,0,247,0,31,0,97,0,160,0,75,0,53,0,60,0,8,0,0,0,65,0,94,0,67,0,115,0,210,0,192,0,13,0,0,0,0,0,247,0,227,0,238,0,0,0,60,0,118,0,254,0,170,0,72,0,250,0,225,0,0,0,0,0,87,0,0,0,10,0,125,0,16,0,145,0,67,0,13,0,152,0,155,0,0,0,0,0,231,0,0,0,152,0,4,0,12,0,117,0,89,0,9,0,0,0,98,0,0,0,50,0,127,0,208,0,54,0,0,0,167,0,137,0,124,0,238,0,151,0,183,0,173,0,0,0,237,0,9,0,72,0,104,0,156,0,196,0,25,0,40,0,100,0,158,0,144,0,102,0,164,0,112,0,204,0,0,0,0,0,94,0,227,0,152,0,171,0,0,0,249,0,58,0,222,0,164,0,19,0,0,0,0,0,46,0,0,0,32,0,83,0,229,0,14,0,215,0,187,0,212,0,230,0,120,0,105,0,0,0,188,0,0,0,139,0,249,0,52,0,106,0,55,0,149,0,22,0,66,0,195,0,126,0,149,0,194,0,190,0,23,0,0,0,62,0,210,0,185,0,197,0,37,0,238,0,122,0,127,0,88,0,54,0,64,0,181,0,24,0,180,0,254,0,167,0,163,0,0,0,0,0,181,0,159,0,128,0,80,0,0,0,161,0,0,0,231,0,0,0,230,0,184,0,0,0,206,0,237,0,0,0,25,0,0,0,117,0,164,0,64,0,0,0,39,0,0,0,172,0,0,0,58,0,225,0,13,0,74,0,142,0,62,0,64,0,95,0,0,0,0,0,233,0,192,0,0,0,154,0,31,0,10,0,230,0,251,0,0,0,0,0,107,0,199,0,93,0,238,0,173,0,243,0,122,0,228,0,61,0,45,0,0,0,33,0,159,0,80,0,0,0,68,0,58,0,202,0,169,0,0,0,91,0,192,0,0,0,128,0,1,0,0,0,0,0,24,0,0,0,127,0,0,0,93,0,0,0,214,0,99,0,88,0,14,0,147,0,245,0,190,0,98,0,0,0,121,0,234,0,25,0,73,0,25,0,215,0,3,0,81,0,0,0,81,0,132,0,127,0,119,0,28,0,89,0,106,0,0,0,231,0,68,0,166,0,39,0,0,0,195,0,0,0,10,0,149,0,0,0,240,0,84,0,0,0,156,0,0,0,0,0,253,0,12,0,31,0,0,0,0,0,53,0,17,0,33,0,103,0,51,0,10,0,254,0,23,0,167,0,150,0,0,0,0,0,25,0,169,0,0,0,10,0,149,0,67,0,40,0,0,0,93,0,194,0,123,0,0,0,231,0,169,0,233,0,210,0,236,0,26,0,90,0,0,0,154,0,238,0,171,0,250,0,193,0,167,0,0,0,0,0,70,0,43,0,81,0,0,0,0,0,37,0,164,0,0,0,7,0,33,0,23,0,169,0,0,0,0,0,174,0,197,0,44,0,187,0,106,0,120,0,207,0,107,0,35,0,77,0,97,0,69,0,0,0,123,0,47,0,0,0,75,0);
signal scenario_full  : scenario_type := (220,31,137,31,137,30,191,31,191,30,184,31,184,30,173,31,239,31,44,31,27,31,119,31,19,31,213,31,25,31,101,31,225,31,76,31,19,31,47,31,47,30,121,31,230,31,230,30,29,31,151,31,136,31,254,31,217,31,86,31,86,30,86,29,220,31,220,30,131,31,131,30,189,31,218,31,99,31,99,30,126,31,244,31,248,31,248,30,248,29,248,28,248,27,27,31,27,30,27,29,122,31,142,31,183,31,188,31,2,31,2,30,150,31,55,31,158,31,70,31,252,31,107,31,129,31,129,30,48,31,48,30,44,31,228,31,238,31,120,31,31,31,142,31,154,31,136,31,96,31,146,31,146,30,146,29,146,28,107,31,197,31,186,31,91,31,136,31,82,31,204,31,189,31,234,31,133,31,133,30,123,31,123,30,123,29,98,31,98,30,10,31,19,31,40,31,55,31,140,31,23,31,253,31,253,30,169,31,169,30,169,29,129,31,24,31,6,31,157,31,103,31,223,31,170,31,178,31,223,31,91,31,91,30,91,29,70,31,240,31,238,31,92,31,135,31,162,31,183,31,83,31,83,30,226,31,94,31,159,31,105,31,4,31,1,31,102,31,70,31,54,31,170,31,212,31,73,31,160,31,127,31,230,31,222,31,222,30,207,31,185,31,185,30,185,29,219,31,26,31,199,31,42,31,43,31,180,31,249,31,249,30,148,31,244,31,246,31,225,31,136,31,76,31,37,31,106,31,165,31,199,31,236,31,203,31,203,30,38,31,149,31,22,31,42,31,56,31,120,31,221,31,199,31,214,31,239,31,201,31,99,31,99,30,107,31,90,31,90,30,76,31,167,31,126,31,11,31,239,31,129,31,129,30,36,31,95,31,177,31,177,30,119,31,119,30,94,31,113,31,113,30,141,31,171,31,70,31,246,31,7,31,7,30,7,29,7,28,7,27,147,31,147,30,147,29,131,31,54,31,167,31,93,31,218,31,87,31,162,31,69,31,105,31,211,31,220,31,42,31,185,31,129,31,131,31,250,31,31,31,187,31,100,31,133,31,220,31,201,31,186,31,238,31,126,31,126,30,7,31,239,31,217,31,217,30,164,31,204,31,48,31,200,31,242,31,81,31,200,31,39,31,126,31,33,31,131,31,177,31,177,30,74,31,232,31,172,31,172,30,217,31,211,31,69,31,111,31,41,31,82,31,117,31,117,30,10,31,137,31,107,31,249,31,249,30,224,31,224,30,251,31,251,30,251,29,207,31,36,31,131,31,203,31,202,31,197,31,10,31,239,31,125,31,166,31,166,30,232,31,5,31,5,30,213,31,213,30,27,31,38,31,50,31,50,30,92,31,93,31,93,30,148,31,112,31,135,31,135,30,103,31,37,31,212,31,113,31,154,31,106,31,127,31,96,31,203,31,203,30,49,31,49,30,64,31,64,30,157,31,171,31,62,31,218,31,225,31,225,30,79,31,58,31,151,31,216,31,216,30,235,31,251,31,79,31,19,31,166,31,219,31,48,31,48,30,205,31,136,31,113,31,95,31,97,31,54,31,54,30,54,29,96,31,96,30,77,31,26,31,82,31,74,31,74,30,74,29,210,31,236,31,180,31,193,31,106,31,239,31,14,31,118,31,226,31,226,30,226,29,226,28,226,27,33,31,95,31,27,31,27,30,198,31,202,31,101,31,191,31,41,31,183,31,179,31,109,31,55,31,185,31,214,31,185,31,171,31,24,31,106,31,135,31,135,30,97,31,14,31,165,31,69,31,76,31,63,31,63,30,63,29,171,31,194,31,251,31,124,31,61,31,145,31,202,31,47,31,104,31,104,30,104,29,104,28,125,31,242,31,145,31,220,31,209,31,209,30,41,31,102,31,2,31,74,31,155,31,251,31,251,30,251,29,120,31,213,31,130,31,209,31,122,31,85,31,30,31,238,31,238,30,238,29,128,31,241,31,241,30,139,31,228,31,222,31,206,31,206,30,206,29,169,31,111,31,50,31,162,31,255,31,148,31,68,31,122,31,253,31,145,31,29,31,167,31,184,31,216,31,68,31,68,30,158,31,158,30,60,31,8,31,8,30,135,31,114,31,97,31,97,30,61,31,16,31,83,31,130,31,102,31,213,31,127,31,204,31,102,31,78,31,207,31,140,31,77,31,130,31,115,31,113,31,224,31,30,31,192,31,4,31,58,31,144,31,144,30,144,29,253,31,253,30,31,31,65,31,7,31,7,30,9,31,179,31,95,31,147,31,220,31,220,30,129,31,183,31,237,31,237,30,221,31,34,31,78,31,78,30,65,31,58,31,8,31,183,31,243,31,243,30,46,31,126,31,81,31,103,31,23,31,23,30,23,29,247,31,31,31,97,31,160,31,75,31,53,31,60,31,8,31,8,30,65,31,94,31,67,31,115,31,210,31,192,31,13,31,13,30,13,29,247,31,227,31,238,31,238,30,60,31,118,31,254,31,170,31,72,31,250,31,225,31,225,30,225,29,87,31,87,30,10,31,125,31,16,31,145,31,67,31,13,31,152,31,155,31,155,30,155,29,231,31,231,30,152,31,4,31,12,31,117,31,89,31,9,31,9,30,98,31,98,30,50,31,127,31,208,31,54,31,54,30,167,31,137,31,124,31,238,31,151,31,183,31,173,31,173,30,237,31,9,31,72,31,104,31,156,31,196,31,25,31,40,31,100,31,158,31,144,31,102,31,164,31,112,31,204,31,204,30,204,29,94,31,227,31,152,31,171,31,171,30,249,31,58,31,222,31,164,31,19,31,19,30,19,29,46,31,46,30,32,31,83,31,229,31,14,31,215,31,187,31,212,31,230,31,120,31,105,31,105,30,188,31,188,30,139,31,249,31,52,31,106,31,55,31,149,31,22,31,66,31,195,31,126,31,149,31,194,31,190,31,23,31,23,30,62,31,210,31,185,31,197,31,37,31,238,31,122,31,127,31,88,31,54,31,64,31,181,31,24,31,180,31,254,31,167,31,163,31,163,30,163,29,181,31,159,31,128,31,80,31,80,30,161,31,161,30,231,31,231,30,230,31,184,31,184,30,206,31,237,31,237,30,25,31,25,30,117,31,164,31,64,31,64,30,39,31,39,30,172,31,172,30,58,31,225,31,13,31,74,31,142,31,62,31,64,31,95,31,95,30,95,29,233,31,192,31,192,30,154,31,31,31,10,31,230,31,251,31,251,30,251,29,107,31,199,31,93,31,238,31,173,31,243,31,122,31,228,31,61,31,45,31,45,30,33,31,159,31,80,31,80,30,68,31,58,31,202,31,169,31,169,30,91,31,192,31,192,30,128,31,1,31,1,30,1,29,24,31,24,30,127,31,127,30,93,31,93,30,214,31,99,31,88,31,14,31,147,31,245,31,190,31,98,31,98,30,121,31,234,31,25,31,73,31,25,31,215,31,3,31,81,31,81,30,81,31,132,31,127,31,119,31,28,31,89,31,106,31,106,30,231,31,68,31,166,31,39,31,39,30,195,31,195,30,10,31,149,31,149,30,240,31,84,31,84,30,156,31,156,30,156,29,253,31,12,31,31,31,31,30,31,29,53,31,17,31,33,31,103,31,51,31,10,31,254,31,23,31,167,31,150,31,150,30,150,29,25,31,169,31,169,30,10,31,149,31,67,31,40,31,40,30,93,31,194,31,123,31,123,30,231,31,169,31,233,31,210,31,236,31,26,31,90,31,90,30,154,31,238,31,171,31,250,31,193,31,167,31,167,30,167,29,70,31,43,31,81,31,81,30,81,29,37,31,164,31,164,30,7,31,33,31,23,31,169,31,169,30,169,29,174,31,197,31,44,31,187,31,106,31,120,31,207,31,107,31,35,31,77,31,97,31,69,31,69,30,123,31,47,31,47,30,75,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
