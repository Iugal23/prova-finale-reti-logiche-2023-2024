-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_133 is
end project_tb_133;

architecture project_tb_arch_133 of project_tb_133 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 263;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,0,0,86,0,74,0,186,0,0,0,201,0,86,0,155,0,205,0,255,0,158,0,219,0,0,0,22,0,235,0,65,0,213,0,85,0,27,0,0,0,127,0,244,0,94,0,166,0,181,0,0,0,140,0,202,0,174,0,181,0,0,0,208,0,47,0,196,0,54,0,19,0,216,0,33,0,45,0,55,0,63,0,69,0,109,0,217,0,0,0,208,0,0,0,242,0,169,0,25,0,194,0,37,0,146,0,120,0,0,0,215,0,12,0,214,0,0,0,173,0,249,0,168,0,33,0,76,0,170,0,141,0,186,0,220,0,0,0,0,0,11,0,211,0,251,0,118,0,157,0,51,0,229,0,165,0,176,0,45,0,97,0,248,0,32,0,0,0,33,0,6,0,116,0,0,0,0,0,84,0,153,0,74,0,228,0,19,0,136,0,0,0,86,0,221,0,185,0,18,0,95,0,186,0,61,0,140,0,120,0,0,0,29,0,13,0,17,0,59,0,183,0,0,0,47,0,133,0,129,0,251,0,146,0,168,0,0,0,0,0,72,0,0,0,0,0,202,0,0,0,49,0,66,0,0,0,0,0,0,0,249,0,33,0,209,0,72,0,0,0,242,0,143,0,199,0,0,0,0,0,143,0,161,0,0,0,0,0,94,0,15,0,233,0,104,0,123,0,249,0,222,0,34,0,170,0,211,0,23,0,0,0,0,0,95,0,250,0,252,0,0,0,69,0,189,0,0,0,237,0,0,0,81,0,85,0,130,0,69,0,4,0,215,0,76,0,126,0,201,0,82,0,24,0,210,0,0,0,0,0,0,0,53,0,0,0,52,0,192,0,89,0,150,0,189,0,253,0,78,0,9,0,66,0,0,0,0,0,134,0,0,0,235,0,0,0,129,0,141,0,196,0,81,0,16,0,207,0,207,0,107,0,207,0,101,0,0,0,82,0,46,0,37,0,64,0,215,0,69,0,0,0,0,0,25,0,61,0,0,0,143,0,96,0,211,0,176,0,208,0,75,0,225,0,155,0,220,0,68,0,151,0,157,0,221,0,237,0,123,0,35,0,0,0,190,0,92,0,200,0,188,0,0,0,0,0,0,0,0,0,0,0,88,0,180,0,42,0,0,0,97,0,179,0,37,0,122,0,212,0,49,0,151,0,0,0,112,0,183,0,120,0,0,0);
signal scenario_full  : scenario_type := (214,31,214,30,86,31,74,31,186,31,186,30,201,31,86,31,155,31,205,31,255,31,158,31,219,31,219,30,22,31,235,31,65,31,213,31,85,31,27,31,27,30,127,31,244,31,94,31,166,31,181,31,181,30,140,31,202,31,174,31,181,31,181,30,208,31,47,31,196,31,54,31,19,31,216,31,33,31,45,31,55,31,63,31,69,31,109,31,217,31,217,30,208,31,208,30,242,31,169,31,25,31,194,31,37,31,146,31,120,31,120,30,215,31,12,31,214,31,214,30,173,31,249,31,168,31,33,31,76,31,170,31,141,31,186,31,220,31,220,30,220,29,11,31,211,31,251,31,118,31,157,31,51,31,229,31,165,31,176,31,45,31,97,31,248,31,32,31,32,30,33,31,6,31,116,31,116,30,116,29,84,31,153,31,74,31,228,31,19,31,136,31,136,30,86,31,221,31,185,31,18,31,95,31,186,31,61,31,140,31,120,31,120,30,29,31,13,31,17,31,59,31,183,31,183,30,47,31,133,31,129,31,251,31,146,31,168,31,168,30,168,29,72,31,72,30,72,29,202,31,202,30,49,31,66,31,66,30,66,29,66,28,249,31,33,31,209,31,72,31,72,30,242,31,143,31,199,31,199,30,199,29,143,31,161,31,161,30,161,29,94,31,15,31,233,31,104,31,123,31,249,31,222,31,34,31,170,31,211,31,23,31,23,30,23,29,95,31,250,31,252,31,252,30,69,31,189,31,189,30,237,31,237,30,81,31,85,31,130,31,69,31,4,31,215,31,76,31,126,31,201,31,82,31,24,31,210,31,210,30,210,29,210,28,53,31,53,30,52,31,192,31,89,31,150,31,189,31,253,31,78,31,9,31,66,31,66,30,66,29,134,31,134,30,235,31,235,30,129,31,141,31,196,31,81,31,16,31,207,31,207,31,107,31,207,31,101,31,101,30,82,31,46,31,37,31,64,31,215,31,69,31,69,30,69,29,25,31,61,31,61,30,143,31,96,31,211,31,176,31,208,31,75,31,225,31,155,31,220,31,68,31,151,31,157,31,221,31,237,31,123,31,35,31,35,30,190,31,92,31,200,31,188,31,188,30,188,29,188,28,188,27,188,26,88,31,180,31,42,31,42,30,97,31,179,31,37,31,122,31,212,31,49,31,151,31,151,30,112,31,183,31,120,31,120,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
