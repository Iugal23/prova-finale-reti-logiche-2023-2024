-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_302 is
end project_tb_302;

architecture project_tb_arch_302 of project_tb_302 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 259;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,64,0,247,0,151,0,62,0,20,0,3,0,0,0,0,0,73,0,22,0,238,0,233,0,200,0,105,0,253,0,38,0,135,0,28,0,71,0,177,0,163,0,247,0,143,0,0,0,133,0,244,0,0,0,186,0,152,0,0,0,154,0,220,0,0,0,79,0,218,0,225,0,226,0,155,0,0,0,184,0,199,0,237,0,151,0,32,0,0,0,60,0,207,0,223,0,32,0,0,0,235,0,0,0,34,0,1,0,0,0,0,0,150,0,196,0,182,0,170,0,0,0,199,0,78,0,90,0,0,0,49,0,147,0,116,0,186,0,23,0,70,0,154,0,0,0,0,0,0,0,213,0,51,0,140,0,83,0,12,0,23,0,172,0,191,0,51,0,225,0,122,0,144,0,157,0,108,0,32,0,16,0,25,0,0,0,5,0,232,0,15,0,189,0,26,0,17,0,0,0,17,0,154,0,151,0,37,0,134,0,0,0,0,0,0,0,0,0,45,0,1,0,150,0,244,0,154,0,47,0,0,0,0,0,76,0,50,0,144,0,0,0,201,0,230,0,231,0,86,0,0,0,0,0,0,0,50,0,184,0,151,0,0,0,0,0,240,0,115,0,190,0,254,0,0,0,0,0,0,0,99,0,212,0,132,0,178,0,0,0,167,0,123,0,247,0,100,0,254,0,97,0,108,0,9,0,0,0,2,0,0,0,50,0,89,0,132,0,4,0,189,0,222,0,10,0,2,0,148,0,27,0,24,0,47,0,83,0,192,0,184,0,65,0,151,0,173,0,0,0,161,0,212,0,220,0,30,0,40,0,155,0,168,0,227,0,129,0,217,0,233,0,0,0,242,0,0,0,90,0,67,0,121,0,0,0,20,0,197,0,210,0,198,0,236,0,204,0,125,0,239,0,36,0,113,0,0,0,170,0,175,0,65,0,242,0,181,0,177,0,37,0,222,0,18,0,59,0,0,0,157,0,18,0,6,0,22,0,167,0,114,0,213,0,138,0,156,0,237,0,0,0,46,0,38,0,112,0,116,0,0,0,218,0,226,0,242,0,209,0,179,0,143,0,232,0,10,0,75,0,80,0,0,0,254,0,19,0,137,0,198,0,151,0,132,0,20,0,0,0,27,0,134,0,0,0,29,0,208,0,119,0,236,0,0,0);
signal scenario_full  : scenario_type := (36,31,64,31,247,31,151,31,62,31,20,31,3,31,3,30,3,29,73,31,22,31,238,31,233,31,200,31,105,31,253,31,38,31,135,31,28,31,71,31,177,31,163,31,247,31,143,31,143,30,133,31,244,31,244,30,186,31,152,31,152,30,154,31,220,31,220,30,79,31,218,31,225,31,226,31,155,31,155,30,184,31,199,31,237,31,151,31,32,31,32,30,60,31,207,31,223,31,32,31,32,30,235,31,235,30,34,31,1,31,1,30,1,29,150,31,196,31,182,31,170,31,170,30,199,31,78,31,90,31,90,30,49,31,147,31,116,31,186,31,23,31,70,31,154,31,154,30,154,29,154,28,213,31,51,31,140,31,83,31,12,31,23,31,172,31,191,31,51,31,225,31,122,31,144,31,157,31,108,31,32,31,16,31,25,31,25,30,5,31,232,31,15,31,189,31,26,31,17,31,17,30,17,31,154,31,151,31,37,31,134,31,134,30,134,29,134,28,134,27,45,31,1,31,150,31,244,31,154,31,47,31,47,30,47,29,76,31,50,31,144,31,144,30,201,31,230,31,231,31,86,31,86,30,86,29,86,28,50,31,184,31,151,31,151,30,151,29,240,31,115,31,190,31,254,31,254,30,254,29,254,28,99,31,212,31,132,31,178,31,178,30,167,31,123,31,247,31,100,31,254,31,97,31,108,31,9,31,9,30,2,31,2,30,50,31,89,31,132,31,4,31,189,31,222,31,10,31,2,31,148,31,27,31,24,31,47,31,83,31,192,31,184,31,65,31,151,31,173,31,173,30,161,31,212,31,220,31,30,31,40,31,155,31,168,31,227,31,129,31,217,31,233,31,233,30,242,31,242,30,90,31,67,31,121,31,121,30,20,31,197,31,210,31,198,31,236,31,204,31,125,31,239,31,36,31,113,31,113,30,170,31,175,31,65,31,242,31,181,31,177,31,37,31,222,31,18,31,59,31,59,30,157,31,18,31,6,31,22,31,167,31,114,31,213,31,138,31,156,31,237,31,237,30,46,31,38,31,112,31,116,31,116,30,218,31,226,31,242,31,209,31,179,31,143,31,232,31,10,31,75,31,80,31,80,30,254,31,19,31,137,31,198,31,151,31,132,31,20,31,20,30,27,31,134,31,134,30,29,31,208,31,119,31,236,31,236,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
