-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 205;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (171,0,29,0,88,0,104,0,153,0,122,0,69,0,0,0,174,0,146,0,63,0,0,0,244,0,248,0,207,0,172,0,0,0,94,0,131,0,7,0,178,0,103,0,0,0,87,0,75,0,191,0,96,0,145,0,0,0,0,0,0,0,0,0,0,0,46,0,216,0,184,0,6,0,0,0,78,0,0,0,0,0,22,0,18,0,246,0,0,0,101,0,2,0,35,0,0,0,197,0,100,0,200,0,135,0,170,0,199,0,14,0,117,0,125,0,0,0,0,0,0,0,74,0,46,0,126,0,0,0,220,0,110,0,116,0,124,0,0,0,176,0,252,0,93,0,104,0,116,0,65,0,0,0,101,0,176,0,0,0,204,0,120,0,28,0,113,0,62,0,46,0,0,0,0,0,0,0,33,0,206,0,182,0,228,0,225,0,128,0,215,0,151,0,78,0,0,0,0,0,48,0,191,0,81,0,81,0,232,0,239,0,201,0,178,0,0,0,211,0,74,0,30,0,0,0,183,0,0,0,201,0,88,0,48,0,111,0,98,0,197,0,161,0,155,0,8,0,160,0,41,0,245,0,0,0,43,0,182,0,178,0,91,0,141,0,226,0,210,0,187,0,125,0,235,0,0,0,46,0,165,0,201,0,2,0,0,0,121,0,124,0,110,0,49,0,22,0,82,0,170,0,141,0,165,0,133,0,0,0,156,0,9,0,135,0,247,0,181,0,0,0,0,0,230,0,0,0,252,0,17,0,45,0,76,0,99,0,0,0,5,0,0,0,193,0,0,0,70,0,175,0,236,0,0,0,29,0,248,0,176,0,0,0,102,0,178,0,62,0,241,0,218,0,185,0,0,0,162,0,0,0,125,0,134,0,225,0,0,0,0,0,120,0,215,0,230,0,169,0,121,0,15,0,0,0,66,0,107,0);
signal scenario_full  : scenario_type := (171,31,29,31,88,31,104,31,153,31,122,31,69,31,69,30,174,31,146,31,63,31,63,30,244,31,248,31,207,31,172,31,172,30,94,31,131,31,7,31,178,31,103,31,103,30,87,31,75,31,191,31,96,31,145,31,145,30,145,29,145,28,145,27,145,26,46,31,216,31,184,31,6,31,6,30,78,31,78,30,78,29,22,31,18,31,246,31,246,30,101,31,2,31,35,31,35,30,197,31,100,31,200,31,135,31,170,31,199,31,14,31,117,31,125,31,125,30,125,29,125,28,74,31,46,31,126,31,126,30,220,31,110,31,116,31,124,31,124,30,176,31,252,31,93,31,104,31,116,31,65,31,65,30,101,31,176,31,176,30,204,31,120,31,28,31,113,31,62,31,46,31,46,30,46,29,46,28,33,31,206,31,182,31,228,31,225,31,128,31,215,31,151,31,78,31,78,30,78,29,48,31,191,31,81,31,81,31,232,31,239,31,201,31,178,31,178,30,211,31,74,31,30,31,30,30,183,31,183,30,201,31,88,31,48,31,111,31,98,31,197,31,161,31,155,31,8,31,160,31,41,31,245,31,245,30,43,31,182,31,178,31,91,31,141,31,226,31,210,31,187,31,125,31,235,31,235,30,46,31,165,31,201,31,2,31,2,30,121,31,124,31,110,31,49,31,22,31,82,31,170,31,141,31,165,31,133,31,133,30,156,31,9,31,135,31,247,31,181,31,181,30,181,29,230,31,230,30,252,31,17,31,45,31,76,31,99,31,99,30,5,31,5,30,193,31,193,30,70,31,175,31,236,31,236,30,29,31,248,31,176,31,176,30,102,31,178,31,62,31,241,31,218,31,185,31,185,30,162,31,162,30,125,31,134,31,225,31,225,30,225,29,120,31,215,31,230,31,169,31,121,31,15,31,15,30,66,31,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
