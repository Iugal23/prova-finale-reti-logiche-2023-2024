-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 618;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (145,0,78,0,164,0,80,0,44,0,129,0,25,0,217,0,0,0,128,0,25,0,0,0,65,0,193,0,157,0,15,0,87,0,59,0,8,0,56,0,147,0,120,0,176,0,0,0,90,0,16,0,216,0,216,0,7,0,87,0,71,0,74,0,9,0,62,0,0,0,22,0,131,0,37,0,96,0,117,0,159,0,67,0,72,0,138,0,35,0,137,0,0,0,0,0,0,0,146,0,228,0,163,0,0,0,143,0,0,0,148,0,87,0,111,0,80,0,0,0,194,0,0,0,0,0,226,0,49,0,75,0,0,0,0,0,48,0,204,0,90,0,188,0,58,0,0,0,245,0,245,0,118,0,172,0,25,0,23,0,109,0,103,0,3,0,89,0,0,0,136,0,37,0,66,0,0,0,232,0,66,0,88,0,0,0,157,0,2,0,88,0,173,0,191,0,126,0,242,0,74,0,233,0,23,0,220,0,84,0,132,0,250,0,151,0,174,0,114,0,0,0,0,0,34,0,92,0,108,0,195,0,171,0,245,0,0,0,2,0,66,0,0,0,197,0,108,0,154,0,68,0,0,0,173,0,0,0,172,0,189,0,201,0,52,0,27,0,201,0,235,0,8,0,155,0,108,0,110,0,0,0,22,0,0,0,184,0,164,0,145,0,32,0,240,0,253,0,0,0,0,0,170,0,157,0,54,0,0,0,185,0,0,0,187,0,95,0,72,0,224,0,119,0,193,0,170,0,91,0,0,0,98,0,36,0,204,0,13,0,253,0,142,0,72,0,132,0,139,0,144,0,141,0,141,0,173,0,38,0,169,0,208,0,142,0,209,0,1,0,228,0,42,0,67,0,28,0,220,0,0,0,209,0,211,0,67,0,113,0,47,0,71,0,83,0,56,0,17,0,227,0,84,0,0,0,170,0,24,0,0,0,0,0,173,0,16,0,5,0,26,0,0,0,104,0,87,0,232,0,141,0,235,0,210,0,125,0,14,0,179,0,0,0,240,0,152,0,254,0,115,0,4,0,14,0,255,0,175,0,108,0,2,0,153,0,235,0,220,0,104,0,248,0,194,0,148,0,159,0,0,0,233,0,46,0,16,0,125,0,60,0,233,0,242,0,3,0,43,0,118,0,92,0,170,0,0,0,0,0,198,0,201,0,19,0,136,0,206,0,104,0,0,0,0,0,214,0,58,0,135,0,26,0,86,0,0,0,41,0,165,0,151,0,144,0,86,0,0,0,0,0,202,0,0,0,156,0,141,0,55,0,16,0,0,0,223,0,67,0,0,0,18,0,105,0,207,0,51,0,0,0,0,0,244,0,0,0,135,0,216,0,0,0,65,0,0,0,248,0,165,0,17,0,0,0,63,0,0,0,120,0,93,0,161,0,132,0,120,0,83,0,222,0,195,0,38,0,0,0,66,0,26,0,100,0,5,0,20,0,221,0,177,0,0,0,30,0,185,0,128,0,135,0,214,0,0,0,174,0,28,0,178,0,47,0,0,0,207,0,101,0,126,0,176,0,0,0,131,0,113,0,35,0,0,0,241,0,80,0,0,0,116,0,30,0,0,0,127,0,87,0,151,0,0,0,187,0,224,0,0,0,233,0,0,0,40,0,111,0,62,0,249,0,0,0,20,0,180,0,0,0,137,0,0,0,240,0,234,0,69,0,4,0,70,0,238,0,24,0,135,0,69,0,131,0,125,0,1,0,93,0,52,0,34,0,0,0,89,0,74,0,0,0,77,0,192,0,19,0,162,0,200,0,140,0,247,0,86,0,15,0,225,0,24,0,17,0,48,0,206,0,37,0,95,0,102,0,93,0,204,0,25,0,0,0,231,0,210,0,212,0,10,0,194,0,0,0,0,0,0,0,184,0,107,0,20,0,0,0,104,0,30,0,0,0,150,0,149,0,72,0,128,0,0,0,70,0,128,0,0,0,81,0,0,0,225,0,15,0,150,0,175,0,96,0,52,0,32,0,156,0,12,0,224,0,173,0,111,0,41,0,0,0,247,0,27,0,31,0,216,0,123,0,46,0,171,0,109,0,34,0,0,0,0,0,74,0,36,0,71,0,97,0,0,0,255,0,237,0,183,0,65,0,146,0,92,0,137,0,0,0,56,0,53,0,211,0,203,0,0,0,153,0,206,0,6,0,89,0,110,0,67,0,162,0,85,0,0,0,0,0,0,0,70,0,41,0,103,0,121,0,129,0,175,0,197,0,238,0,84,0,247,0,70,0,0,0,15,0,182,0,0,0,241,0,225,0,0,0,0,0,0,0,137,0,45,0,0,0,105,0,53,0,142,0,222,0,22,0,0,0,173,0,29,0,0,0,124,0,0,0,106,0,105,0,218,0,124,0,218,0,237,0,0,0,70,0,201,0,186,0,23,0,186,0,0,0,52,0,0,0,0,0,0,0,95,0,94,0,152,0,224,0,137,0,240,0,146,0,46,0,14,0,64,0,176,0,145,0,187,0,136,0,213,0,0,0,105,0,158,0,218,0,0,0,46,0,149,0,0,0,4,0,8,0,16,0,0,0,252,0,102,0,87,0,56,0,0,0,44,0,21,0,243,0,47,0,0,0,0,0,171,0,55,0,15,0,214,0,220,0,14,0,137,0,121,0,129,0,58,0,248,0,42,0,240,0,0,0,0,0,0,0,198,0,51,0,185,0,124,0,0,0,67,0,250,0,192,0,62,0,73,0,0,0,233,0,9,0,37,0,0,0,87,0,133,0,60,0,178,0,127,0,232,0,48,0,254,0,41,0,0,0,84,0);
signal scenario_full  : scenario_type := (145,31,78,31,164,31,80,31,44,31,129,31,25,31,217,31,217,30,128,31,25,31,25,30,65,31,193,31,157,31,15,31,87,31,59,31,8,31,56,31,147,31,120,31,176,31,176,30,90,31,16,31,216,31,216,31,7,31,87,31,71,31,74,31,9,31,62,31,62,30,22,31,131,31,37,31,96,31,117,31,159,31,67,31,72,31,138,31,35,31,137,31,137,30,137,29,137,28,146,31,228,31,163,31,163,30,143,31,143,30,148,31,87,31,111,31,80,31,80,30,194,31,194,30,194,29,226,31,49,31,75,31,75,30,75,29,48,31,204,31,90,31,188,31,58,31,58,30,245,31,245,31,118,31,172,31,25,31,23,31,109,31,103,31,3,31,89,31,89,30,136,31,37,31,66,31,66,30,232,31,66,31,88,31,88,30,157,31,2,31,88,31,173,31,191,31,126,31,242,31,74,31,233,31,23,31,220,31,84,31,132,31,250,31,151,31,174,31,114,31,114,30,114,29,34,31,92,31,108,31,195,31,171,31,245,31,245,30,2,31,66,31,66,30,197,31,108,31,154,31,68,31,68,30,173,31,173,30,172,31,189,31,201,31,52,31,27,31,201,31,235,31,8,31,155,31,108,31,110,31,110,30,22,31,22,30,184,31,164,31,145,31,32,31,240,31,253,31,253,30,253,29,170,31,157,31,54,31,54,30,185,31,185,30,187,31,95,31,72,31,224,31,119,31,193,31,170,31,91,31,91,30,98,31,36,31,204,31,13,31,253,31,142,31,72,31,132,31,139,31,144,31,141,31,141,31,173,31,38,31,169,31,208,31,142,31,209,31,1,31,228,31,42,31,67,31,28,31,220,31,220,30,209,31,211,31,67,31,113,31,47,31,71,31,83,31,56,31,17,31,227,31,84,31,84,30,170,31,24,31,24,30,24,29,173,31,16,31,5,31,26,31,26,30,104,31,87,31,232,31,141,31,235,31,210,31,125,31,14,31,179,31,179,30,240,31,152,31,254,31,115,31,4,31,14,31,255,31,175,31,108,31,2,31,153,31,235,31,220,31,104,31,248,31,194,31,148,31,159,31,159,30,233,31,46,31,16,31,125,31,60,31,233,31,242,31,3,31,43,31,118,31,92,31,170,31,170,30,170,29,198,31,201,31,19,31,136,31,206,31,104,31,104,30,104,29,214,31,58,31,135,31,26,31,86,31,86,30,41,31,165,31,151,31,144,31,86,31,86,30,86,29,202,31,202,30,156,31,141,31,55,31,16,31,16,30,223,31,67,31,67,30,18,31,105,31,207,31,51,31,51,30,51,29,244,31,244,30,135,31,216,31,216,30,65,31,65,30,248,31,165,31,17,31,17,30,63,31,63,30,120,31,93,31,161,31,132,31,120,31,83,31,222,31,195,31,38,31,38,30,66,31,26,31,100,31,5,31,20,31,221,31,177,31,177,30,30,31,185,31,128,31,135,31,214,31,214,30,174,31,28,31,178,31,47,31,47,30,207,31,101,31,126,31,176,31,176,30,131,31,113,31,35,31,35,30,241,31,80,31,80,30,116,31,30,31,30,30,127,31,87,31,151,31,151,30,187,31,224,31,224,30,233,31,233,30,40,31,111,31,62,31,249,31,249,30,20,31,180,31,180,30,137,31,137,30,240,31,234,31,69,31,4,31,70,31,238,31,24,31,135,31,69,31,131,31,125,31,1,31,93,31,52,31,34,31,34,30,89,31,74,31,74,30,77,31,192,31,19,31,162,31,200,31,140,31,247,31,86,31,15,31,225,31,24,31,17,31,48,31,206,31,37,31,95,31,102,31,93,31,204,31,25,31,25,30,231,31,210,31,212,31,10,31,194,31,194,30,194,29,194,28,184,31,107,31,20,31,20,30,104,31,30,31,30,30,150,31,149,31,72,31,128,31,128,30,70,31,128,31,128,30,81,31,81,30,225,31,15,31,150,31,175,31,96,31,52,31,32,31,156,31,12,31,224,31,173,31,111,31,41,31,41,30,247,31,27,31,31,31,216,31,123,31,46,31,171,31,109,31,34,31,34,30,34,29,74,31,36,31,71,31,97,31,97,30,255,31,237,31,183,31,65,31,146,31,92,31,137,31,137,30,56,31,53,31,211,31,203,31,203,30,153,31,206,31,6,31,89,31,110,31,67,31,162,31,85,31,85,30,85,29,85,28,70,31,41,31,103,31,121,31,129,31,175,31,197,31,238,31,84,31,247,31,70,31,70,30,15,31,182,31,182,30,241,31,225,31,225,30,225,29,225,28,137,31,45,31,45,30,105,31,53,31,142,31,222,31,22,31,22,30,173,31,29,31,29,30,124,31,124,30,106,31,105,31,218,31,124,31,218,31,237,31,237,30,70,31,201,31,186,31,23,31,186,31,186,30,52,31,52,30,52,29,52,28,95,31,94,31,152,31,224,31,137,31,240,31,146,31,46,31,14,31,64,31,176,31,145,31,187,31,136,31,213,31,213,30,105,31,158,31,218,31,218,30,46,31,149,31,149,30,4,31,8,31,16,31,16,30,252,31,102,31,87,31,56,31,56,30,44,31,21,31,243,31,47,31,47,30,47,29,171,31,55,31,15,31,214,31,220,31,14,31,137,31,121,31,129,31,58,31,248,31,42,31,240,31,240,30,240,29,240,28,198,31,51,31,185,31,124,31,124,30,67,31,250,31,192,31,62,31,73,31,73,30,233,31,9,31,37,31,37,30,87,31,133,31,60,31,178,31,127,31,232,31,48,31,254,31,41,31,41,30,84,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
