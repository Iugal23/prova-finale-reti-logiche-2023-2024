-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_25 is
end project_tb_25;

architecture project_tb_arch_25 of project_tb_25 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 910;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,90,0,231,0,68,0,11,0,226,0,73,0,35,0,97,0,167,0,0,0,0,0,13,0,41,0,33,0,152,0,244,0,93,0,178,0,223,0,198,0,164,0,242,0,109,0,7,0,0,0,0,0,0,0,182,0,67,0,190,0,23,0,30,0,236,0,107,0,39,0,52,0,194,0,155,0,0,0,34,0,0,0,237,0,200,0,0,0,99,0,0,0,23,0,41,0,209,0,22,0,35,0,0,0,47,0,152,0,1,0,68,0,173,0,0,0,0,0,56,0,226,0,34,0,45,0,179,0,215,0,211,0,221,0,0,0,236,0,109,0,218,0,238,0,36,0,78,0,8,0,70,0,159,0,233,0,78,0,24,0,196,0,107,0,182,0,65,0,183,0,35,0,0,0,0,0,0,0,255,0,221,0,222,0,197,0,136,0,0,0,16,0,42,0,0,0,0,0,10,0,142,0,251,0,114,0,0,0,203,0,218,0,245,0,0,0,0,0,145,0,239,0,100,0,181,0,190,0,108,0,86,0,37,0,89,0,56,0,0,0,0,0,72,0,229,0,244,0,83,0,121,0,0,0,170,0,174,0,108,0,0,0,0,0,134,0,165,0,54,0,0,0,243,0,119,0,195,0,166,0,8,0,101,0,226,0,77,0,41,0,130,0,58,0,104,0,90,0,12,0,61,0,179,0,88,0,211,0,0,0,0,0,25,0,140,0,26,0,28,0,28,0,31,0,171,0,174,0,222,0,43,0,15,0,247,0,212,0,211,0,179,0,0,0,30,0,12,0,138,0,0,0,0,0,106,0,226,0,172,0,215,0,84,0,4,0,0,0,14,0,0,0,249,0,181,0,0,0,235,0,182,0,0,0,170,0,143,0,74,0,241,0,113,0,0,0,0,0,0,0,140,0,11,0,197,0,72,0,143,0,248,0,216,0,244,0,46,0,133,0,33,0,216,0,48,0,18,0,129,0,229,0,0,0,19,0,0,0,0,0,61,0,61,0,46,0,202,0,212,0,62,0,183,0,9,0,70,0,38,0,46,0,144,0,0,0,68,0,73,0,54,0,224,0,32,0,223,0,33,0,58,0,59,0,0,0,0,0,252,0,0,0,105,0,103,0,0,0,202,0,195,0,0,0,28,0,117,0,35,0,168,0,57,0,143,0,174,0,0,0,33,0,180,0,78,0,0,0,15,0,0,0,0,0,0,0,134,0,79,0,187,0,55,0,152,0,0,0,132,0,167,0,121,0,0,0,84,0,14,0,92,0,82,0,109,0,220,0,0,0,47,0,145,0,0,0,0,0,19,0,0,0,246,0,0,0,233,0,198,0,196,0,179,0,148,0,41,0,0,0,30,0,172,0,170,0,66,0,179,0,56,0,21,0,34,0,136,0,200,0,0,0,62,0,158,0,43,0,250,0,12,0,255,0,88,0,96,0,0,0,179,0,179,0,79,0,0,0,115,0,252,0,91,0,106,0,60,0,95,0,21,0,132,0,243,0,176,0,182,0,229,0,179,0,185,0,66,0,22,0,228,0,71,0,107,0,78,0,89,0,102,0,0,0,138,0,58,0,154,0,248,0,79,0,234,0,0,0,60,0,0,0,147,0,82,0,119,0,94,0,0,0,190,0,149,0,2,0,0,0,122,0,147,0,235,0,91,0,91,0,186,0,102,0,183,0,0,0,0,0,97,0,206,0,18,0,0,0,44,0,204,0,235,0,84,0,234,0,211,0,0,0,220,0,173,0,111,0,198,0,78,0,170,0,158,0,230,0,0,0,146,0,145,0,0,0,58,0,21,0,174,0,236,0,150,0,172,0,31,0,190,0,242,0,228,0,21,0,64,0,0,0,156,0,33,0,109,0,190,0,2,0,248,0,83,0,0,0,27,0,0,0,189,0,33,0,68,0,113,0,119,0,97,0,253,0,0,0,68,0,152,0,189,0,0,0,0,0,116,0,0,0,0,0,36,0,95,0,0,0,176,0,48,0,86,0,137,0,5,0,178,0,6,0,1,0,167,0,147,0,134,0,73,0,240,0,168,0,121,0,135,0,223,0,246,0,75,0,0,0,165,0,0,0,114,0,48,0,178,0,234,0,0,0,0,0,10,0,37,0,123,0,51,0,17,0,174,0,129,0,74,0,200,0,56,0,37,0,90,0,51,0,0,0,70,0,124,0,0,0,155,0,243,0,163,0,252,0,0,0,148,0,39,0,237,0,178,0,0,0,0,0,12,0,56,0,0,0,203,0,32,0,89,0,247,0,0,0,44,0,137,0,153,0,0,0,116,0,0,0,189,0,211,0,17,0,0,0,202,0,56,0,0,0,0,0,145,0,212,0,0,0,228,0,12,0,130,0,128,0,0,0,148,0,112,0,125,0,13,0,254,0,12,0,209,0,51,0,169,0,11,0,190,0,83,0,69,0,177,0,7,0,134,0,182,0,8,0,62,0,44,0,38,0,9,0,120,0,127,0,154,0,51,0,30,0,60,0,245,0,97,0,0,0,0,0,159,0,193,0,0,0,181,0,96,0,193,0,152,0,96,0,83,0,73,0,183,0,51,0,0,0,185,0,215,0,169,0,0,0,165,0,0,0,217,0,103,0,145,0,78,0,11,0,54,0,75,0,61,0,227,0,190,0,156,0,101,0,255,0,90,0,171,0,102,0,17,0,232,0,136,0,26,0,31,0,125,0,103,0,226,0,146,0,173,0,220,0,225,0,146,0,115,0,77,0,65,0,0,0,115,0,69,0,108,0,0,0,0,0,36,0,0,0,11,0,0,0,8,0,34,0,249,0,60,0,208,0,0,0,94,0,180,0,30,0,142,0,92,0,135,0,183,0,33,0,206,0,132,0,0,0,0,0,178,0,0,0,107,0,140,0,133,0,0,0,66,0,0,0,86,0,51,0,249,0,34,0,33,0,0,0,240,0,220,0,15,0,155,0,241,0,0,0,102,0,159,0,222,0,209,0,155,0,41,0,185,0,163,0,51,0,0,0,241,0,42,0,0,0,70,0,0,0,59,0,0,0,158,0,70,0,138,0,179,0,173,0,22,0,39,0,8,0,0,0,128,0,96,0,251,0,253,0,140,0,0,0,174,0,125,0,75,0,28,0,33,0,86,0,159,0,115,0,169,0,49,0,106,0,0,0,167,0,38,0,84,0,242,0,0,0,0,0,98,0,9,0,87,0,69,0,0,0,174,0,218,0,177,0,80,0,0,0,0,0,0,0,0,0,224,0,108,0,0,0,0,0,233,0,232,0,254,0,0,0,6,0,181,0,146,0,185,0,3,0,26,0,23,0,149,0,0,0,77,0,7,0,55,0,86,0,232,0,122,0,0,0,163,0,113,0,200,0,255,0,73,0,76,0,197,0,220,0,130,0,0,0,27,0,45,0,110,0,97,0,142,0,115,0,57,0,64,0,221,0,0,0,47,0,171,0,182,0,0,0,248,0,102,0,180,0,52,0,122,0,152,0,194,0,90,0,106,0,221,0,238,0,0,0,111,0,156,0,113,0,0,0,166,0,81,0,57,0,81,0,189,0,106,0,0,0,174,0,70,0,202,0,132,0,62,0,105,0,13,0,206,0,0,0,90,0,242,0,0,0,170,0,77,0,236,0,0,0,0,0,0,0,107,0,61,0,214,0,242,0,82,0,183,0,0,0,99,0,214,0,253,0,184,0,142,0,81,0,31,0,132,0,216,0,0,0,133,0,137,0,134,0,92,0,91,0,115,0,109,0,242,0,13,0,248,0,0,0,100,0,67,0,74,0,195,0,0,0,69,0,86,0,64,0,0,0,0,0,108,0,131,0,133,0,160,0,0,0,3,0,61,0,107,0,0,0,241,0,5,0,250,0,53,0,5,0,152,0,175,0,72,0,15,0,1,0,24,0,158,0,0,0,0,0,222,0,109,0,69,0,226,0,17,0,0,0,184,0,4,0,14,0,96,0,43,0,172,0,0,0,224,0,119,0,175,0,238,0,42,0,166,0,159,0,72,0,147,0,245,0,249,0,0,0,48,0,0,0,4,0,130,0,177,0,0,0,128,0,170,0,0,0,221,0,87,0,126,0,0,0,16,0);
signal scenario_full  : scenario_type := (0,0,90,31,231,31,68,31,11,31,226,31,73,31,35,31,97,31,167,31,167,30,167,29,13,31,41,31,33,31,152,31,244,31,93,31,178,31,223,31,198,31,164,31,242,31,109,31,7,31,7,30,7,29,7,28,182,31,67,31,190,31,23,31,30,31,236,31,107,31,39,31,52,31,194,31,155,31,155,30,34,31,34,30,237,31,200,31,200,30,99,31,99,30,23,31,41,31,209,31,22,31,35,31,35,30,47,31,152,31,1,31,68,31,173,31,173,30,173,29,56,31,226,31,34,31,45,31,179,31,215,31,211,31,221,31,221,30,236,31,109,31,218,31,238,31,36,31,78,31,8,31,70,31,159,31,233,31,78,31,24,31,196,31,107,31,182,31,65,31,183,31,35,31,35,30,35,29,35,28,255,31,221,31,222,31,197,31,136,31,136,30,16,31,42,31,42,30,42,29,10,31,142,31,251,31,114,31,114,30,203,31,218,31,245,31,245,30,245,29,145,31,239,31,100,31,181,31,190,31,108,31,86,31,37,31,89,31,56,31,56,30,56,29,72,31,229,31,244,31,83,31,121,31,121,30,170,31,174,31,108,31,108,30,108,29,134,31,165,31,54,31,54,30,243,31,119,31,195,31,166,31,8,31,101,31,226,31,77,31,41,31,130,31,58,31,104,31,90,31,12,31,61,31,179,31,88,31,211,31,211,30,211,29,25,31,140,31,26,31,28,31,28,31,31,31,171,31,174,31,222,31,43,31,15,31,247,31,212,31,211,31,179,31,179,30,30,31,12,31,138,31,138,30,138,29,106,31,226,31,172,31,215,31,84,31,4,31,4,30,14,31,14,30,249,31,181,31,181,30,235,31,182,31,182,30,170,31,143,31,74,31,241,31,113,31,113,30,113,29,113,28,140,31,11,31,197,31,72,31,143,31,248,31,216,31,244,31,46,31,133,31,33,31,216,31,48,31,18,31,129,31,229,31,229,30,19,31,19,30,19,29,61,31,61,31,46,31,202,31,212,31,62,31,183,31,9,31,70,31,38,31,46,31,144,31,144,30,68,31,73,31,54,31,224,31,32,31,223,31,33,31,58,31,59,31,59,30,59,29,252,31,252,30,105,31,103,31,103,30,202,31,195,31,195,30,28,31,117,31,35,31,168,31,57,31,143,31,174,31,174,30,33,31,180,31,78,31,78,30,15,31,15,30,15,29,15,28,134,31,79,31,187,31,55,31,152,31,152,30,132,31,167,31,121,31,121,30,84,31,14,31,92,31,82,31,109,31,220,31,220,30,47,31,145,31,145,30,145,29,19,31,19,30,246,31,246,30,233,31,198,31,196,31,179,31,148,31,41,31,41,30,30,31,172,31,170,31,66,31,179,31,56,31,21,31,34,31,136,31,200,31,200,30,62,31,158,31,43,31,250,31,12,31,255,31,88,31,96,31,96,30,179,31,179,31,79,31,79,30,115,31,252,31,91,31,106,31,60,31,95,31,21,31,132,31,243,31,176,31,182,31,229,31,179,31,185,31,66,31,22,31,228,31,71,31,107,31,78,31,89,31,102,31,102,30,138,31,58,31,154,31,248,31,79,31,234,31,234,30,60,31,60,30,147,31,82,31,119,31,94,31,94,30,190,31,149,31,2,31,2,30,122,31,147,31,235,31,91,31,91,31,186,31,102,31,183,31,183,30,183,29,97,31,206,31,18,31,18,30,44,31,204,31,235,31,84,31,234,31,211,31,211,30,220,31,173,31,111,31,198,31,78,31,170,31,158,31,230,31,230,30,146,31,145,31,145,30,58,31,21,31,174,31,236,31,150,31,172,31,31,31,190,31,242,31,228,31,21,31,64,31,64,30,156,31,33,31,109,31,190,31,2,31,248,31,83,31,83,30,27,31,27,30,189,31,33,31,68,31,113,31,119,31,97,31,253,31,253,30,68,31,152,31,189,31,189,30,189,29,116,31,116,30,116,29,36,31,95,31,95,30,176,31,48,31,86,31,137,31,5,31,178,31,6,31,1,31,167,31,147,31,134,31,73,31,240,31,168,31,121,31,135,31,223,31,246,31,75,31,75,30,165,31,165,30,114,31,48,31,178,31,234,31,234,30,234,29,10,31,37,31,123,31,51,31,17,31,174,31,129,31,74,31,200,31,56,31,37,31,90,31,51,31,51,30,70,31,124,31,124,30,155,31,243,31,163,31,252,31,252,30,148,31,39,31,237,31,178,31,178,30,178,29,12,31,56,31,56,30,203,31,32,31,89,31,247,31,247,30,44,31,137,31,153,31,153,30,116,31,116,30,189,31,211,31,17,31,17,30,202,31,56,31,56,30,56,29,145,31,212,31,212,30,228,31,12,31,130,31,128,31,128,30,148,31,112,31,125,31,13,31,254,31,12,31,209,31,51,31,169,31,11,31,190,31,83,31,69,31,177,31,7,31,134,31,182,31,8,31,62,31,44,31,38,31,9,31,120,31,127,31,154,31,51,31,30,31,60,31,245,31,97,31,97,30,97,29,159,31,193,31,193,30,181,31,96,31,193,31,152,31,96,31,83,31,73,31,183,31,51,31,51,30,185,31,215,31,169,31,169,30,165,31,165,30,217,31,103,31,145,31,78,31,11,31,54,31,75,31,61,31,227,31,190,31,156,31,101,31,255,31,90,31,171,31,102,31,17,31,232,31,136,31,26,31,31,31,125,31,103,31,226,31,146,31,173,31,220,31,225,31,146,31,115,31,77,31,65,31,65,30,115,31,69,31,108,31,108,30,108,29,36,31,36,30,11,31,11,30,8,31,34,31,249,31,60,31,208,31,208,30,94,31,180,31,30,31,142,31,92,31,135,31,183,31,33,31,206,31,132,31,132,30,132,29,178,31,178,30,107,31,140,31,133,31,133,30,66,31,66,30,86,31,51,31,249,31,34,31,33,31,33,30,240,31,220,31,15,31,155,31,241,31,241,30,102,31,159,31,222,31,209,31,155,31,41,31,185,31,163,31,51,31,51,30,241,31,42,31,42,30,70,31,70,30,59,31,59,30,158,31,70,31,138,31,179,31,173,31,22,31,39,31,8,31,8,30,128,31,96,31,251,31,253,31,140,31,140,30,174,31,125,31,75,31,28,31,33,31,86,31,159,31,115,31,169,31,49,31,106,31,106,30,167,31,38,31,84,31,242,31,242,30,242,29,98,31,9,31,87,31,69,31,69,30,174,31,218,31,177,31,80,31,80,30,80,29,80,28,80,27,224,31,108,31,108,30,108,29,233,31,232,31,254,31,254,30,6,31,181,31,146,31,185,31,3,31,26,31,23,31,149,31,149,30,77,31,7,31,55,31,86,31,232,31,122,31,122,30,163,31,113,31,200,31,255,31,73,31,76,31,197,31,220,31,130,31,130,30,27,31,45,31,110,31,97,31,142,31,115,31,57,31,64,31,221,31,221,30,47,31,171,31,182,31,182,30,248,31,102,31,180,31,52,31,122,31,152,31,194,31,90,31,106,31,221,31,238,31,238,30,111,31,156,31,113,31,113,30,166,31,81,31,57,31,81,31,189,31,106,31,106,30,174,31,70,31,202,31,132,31,62,31,105,31,13,31,206,31,206,30,90,31,242,31,242,30,170,31,77,31,236,31,236,30,236,29,236,28,107,31,61,31,214,31,242,31,82,31,183,31,183,30,99,31,214,31,253,31,184,31,142,31,81,31,31,31,132,31,216,31,216,30,133,31,137,31,134,31,92,31,91,31,115,31,109,31,242,31,13,31,248,31,248,30,100,31,67,31,74,31,195,31,195,30,69,31,86,31,64,31,64,30,64,29,108,31,131,31,133,31,160,31,160,30,3,31,61,31,107,31,107,30,241,31,5,31,250,31,53,31,5,31,152,31,175,31,72,31,15,31,1,31,24,31,158,31,158,30,158,29,222,31,109,31,69,31,226,31,17,31,17,30,184,31,4,31,14,31,96,31,43,31,172,31,172,30,224,31,119,31,175,31,238,31,42,31,166,31,159,31,72,31,147,31,245,31,249,31,249,30,48,31,48,30,4,31,130,31,177,31,177,30,128,31,170,31,170,30,221,31,87,31,126,31,126,30,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
