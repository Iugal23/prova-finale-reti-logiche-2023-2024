-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 382;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (123,0,208,0,118,0,49,0,42,0,243,0,27,0,102,0,238,0,62,0,149,0,104,0,240,0,136,0,83,0,192,0,81,0,185,0,170,0,112,0,0,0,142,0,0,0,8,0,92,0,0,0,83,0,0,0,221,0,24,0,161,0,203,0,20,0,13,0,68,0,179,0,124,0,177,0,118,0,68,0,222,0,129,0,204,0,242,0,205,0,185,0,0,0,143,0,152,0,60,0,171,0,121,0,42,0,115,0,151,0,15,0,139,0,89,0,64,0,100,0,40,0,0,0,138,0,251,0,54,0,172,0,81,0,171,0,41,0,236,0,241,0,162,0,97,0,58,0,0,0,175,0,194,0,0,0,49,0,50,0,153,0,0,0,227,0,62,0,145,0,240,0,204,0,205,0,176,0,242,0,0,0,147,0,57,0,155,0,116,0,112,0,98,0,130,0,255,0,0,0,101,0,68,0,91,0,85,0,106,0,227,0,0,0,6,0,192,0,0,0,168,0,147,0,141,0,255,0,176,0,194,0,111,0,179,0,53,0,227,0,239,0,62,0,84,0,181,0,222,0,245,0,130,0,165,0,87,0,0,0,43,0,0,0,101,0,0,0,236,0,112,0,0,0,165,0,114,0,0,0,224,0,29,0,171,0,0,0,142,0,0,0,7,0,0,0,0,0,121,0,0,0,72,0,244,0,0,0,23,0,212,0,0,0,63,0,67,0,193,0,0,0,3,0,161,0,196,0,163,0,87,0,33,0,35,0,203,0,33,0,65,0,76,0,143,0,0,0,142,0,0,0,39,0,0,0,76,0,114,0,113,0,248,0,251,0,217,0,57,0,0,0,44,0,39,0,91,0,0,0,0,0,206,0,60,0,13,0,216,0,190,0,142,0,37,0,171,0,215,0,225,0,72,0,0,0,174,0,89,0,160,0,72,0,0,0,187,0,145,0,50,0,0,0,194,0,227,0,237,0,107,0,115,0,0,0,248,0,65,0,244,0,97,0,0,0,158,0,99,0,134,0,207,0,215,0,229,0,74,0,101,0,0,0,19,0,31,0,61,0,73,0,0,0,100,0,0,0,157,0,28,0,135,0,155,0,0,0,218,0,184,0,0,0,96,0,5,0,227,0,89,0,0,0,31,0,54,0,0,0,204,0,166,0,181,0,0,0,0,0,179,0,0,0,227,0,55,0,26,0,254,0,7,0,208,0,99,0,0,0,122,0,247,0,0,0,99,0,0,0,127,0,252,0,0,0,216,0,209,0,248,0,60,0,13,0,46,0,90,0,0,0,85,0,32,0,167,0,0,0,0,0,0,0,151,0,11,0,207,0,238,0,218,0,70,0,0,0,200,0,116,0,205,0,46,0,0,0,224,0,194,0,243,0,38,0,0,0,0,0,0,0,0,0,201,0,191,0,100,0,86,0,0,0,0,0,129,0,219,0,228,0,31,0,75,0,0,0,0,0,216,0,0,0,146,0,16,0,178,0,255,0,142,0,105,0,120,0,245,0,32,0,15,0,73,0,181,0,242,0,132,0,112,0,41,0,0,0,254,0,110,0,178,0,0,0,75,0,165,0,0,0,178,0,24,0,31,0,0,0,156,0,19,0,156,0,43,0,45,0,237,0,235,0,0,0,242,0,0,0,0,0,255,0,224,0,122,0,0,0,16,0,0,0,62,0,0,0,246,0,177,0,219,0,125,0,0,0,128,0,139,0,124,0);
signal scenario_full  : scenario_type := (123,31,208,31,118,31,49,31,42,31,243,31,27,31,102,31,238,31,62,31,149,31,104,31,240,31,136,31,83,31,192,31,81,31,185,31,170,31,112,31,112,30,142,31,142,30,8,31,92,31,92,30,83,31,83,30,221,31,24,31,161,31,203,31,20,31,13,31,68,31,179,31,124,31,177,31,118,31,68,31,222,31,129,31,204,31,242,31,205,31,185,31,185,30,143,31,152,31,60,31,171,31,121,31,42,31,115,31,151,31,15,31,139,31,89,31,64,31,100,31,40,31,40,30,138,31,251,31,54,31,172,31,81,31,171,31,41,31,236,31,241,31,162,31,97,31,58,31,58,30,175,31,194,31,194,30,49,31,50,31,153,31,153,30,227,31,62,31,145,31,240,31,204,31,205,31,176,31,242,31,242,30,147,31,57,31,155,31,116,31,112,31,98,31,130,31,255,31,255,30,101,31,68,31,91,31,85,31,106,31,227,31,227,30,6,31,192,31,192,30,168,31,147,31,141,31,255,31,176,31,194,31,111,31,179,31,53,31,227,31,239,31,62,31,84,31,181,31,222,31,245,31,130,31,165,31,87,31,87,30,43,31,43,30,101,31,101,30,236,31,112,31,112,30,165,31,114,31,114,30,224,31,29,31,171,31,171,30,142,31,142,30,7,31,7,30,7,29,121,31,121,30,72,31,244,31,244,30,23,31,212,31,212,30,63,31,67,31,193,31,193,30,3,31,161,31,196,31,163,31,87,31,33,31,35,31,203,31,33,31,65,31,76,31,143,31,143,30,142,31,142,30,39,31,39,30,76,31,114,31,113,31,248,31,251,31,217,31,57,31,57,30,44,31,39,31,91,31,91,30,91,29,206,31,60,31,13,31,216,31,190,31,142,31,37,31,171,31,215,31,225,31,72,31,72,30,174,31,89,31,160,31,72,31,72,30,187,31,145,31,50,31,50,30,194,31,227,31,237,31,107,31,115,31,115,30,248,31,65,31,244,31,97,31,97,30,158,31,99,31,134,31,207,31,215,31,229,31,74,31,101,31,101,30,19,31,31,31,61,31,73,31,73,30,100,31,100,30,157,31,28,31,135,31,155,31,155,30,218,31,184,31,184,30,96,31,5,31,227,31,89,31,89,30,31,31,54,31,54,30,204,31,166,31,181,31,181,30,181,29,179,31,179,30,227,31,55,31,26,31,254,31,7,31,208,31,99,31,99,30,122,31,247,31,247,30,99,31,99,30,127,31,252,31,252,30,216,31,209,31,248,31,60,31,13,31,46,31,90,31,90,30,85,31,32,31,167,31,167,30,167,29,167,28,151,31,11,31,207,31,238,31,218,31,70,31,70,30,200,31,116,31,205,31,46,31,46,30,224,31,194,31,243,31,38,31,38,30,38,29,38,28,38,27,201,31,191,31,100,31,86,31,86,30,86,29,129,31,219,31,228,31,31,31,75,31,75,30,75,29,216,31,216,30,146,31,16,31,178,31,255,31,142,31,105,31,120,31,245,31,32,31,15,31,73,31,181,31,242,31,132,31,112,31,41,31,41,30,254,31,110,31,178,31,178,30,75,31,165,31,165,30,178,31,24,31,31,31,31,30,156,31,19,31,156,31,43,31,45,31,237,31,235,31,235,30,242,31,242,30,242,29,255,31,224,31,122,31,122,30,16,31,16,30,62,31,62,30,246,31,177,31,219,31,125,31,125,30,128,31,139,31,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
