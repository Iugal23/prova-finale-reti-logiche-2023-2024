-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 945;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (119,0,210,0,36,0,0,0,75,0,50,0,76,0,75,0,212,0,252,0,169,0,210,0,0,0,217,0,38,0,144,0,0,0,23,0,168,0,247,0,0,0,168,0,0,0,0,0,236,0,189,0,10,0,43,0,154,0,219,0,179,0,86,0,112,0,15,0,0,0,10,0,39,0,102,0,209,0,118,0,133,0,76,0,0,0,0,0,209,0,8,0,86,0,250,0,172,0,63,0,122,0,254,0,18,0,0,0,101,0,39,0,107,0,24,0,48,0,42,0,216,0,61,0,40,0,254,0,140,0,102,0,166,0,135,0,31,0,114,0,43,0,124,0,62,0,102,0,128,0,218,0,42,0,124,0,172,0,211,0,0,0,214,0,0,0,147,0,7,0,123,0,199,0,0,0,115,0,110,0,0,0,5,0,232,0,179,0,242,0,0,0,188,0,0,0,67,0,212,0,63,0,39,0,70,0,66,0,71,0,104,0,0,0,126,0,16,0,109,0,206,0,159,0,75,0,0,0,251,0,15,0,116,0,63,0,0,0,210,0,226,0,0,0,187,0,201,0,60,0,12,0,27,0,104,0,117,0,89,0,26,0,61,0,21,0,31,0,0,0,69,0,183,0,97,0,37,0,206,0,118,0,71,0,13,0,0,0,86,0,0,0,0,0,8,0,246,0,133,0,30,0,89,0,197,0,99,0,51,0,183,0,0,0,137,0,161,0,66,0,28,0,28,0,0,0,0,0,184,0,0,0,47,0,219,0,0,0,112,0,138,0,152,0,148,0,242,0,0,0,94,0,96,0,72,0,85,0,56,0,0,0,0,0,98,0,0,0,40,0,90,0,12,0,148,0,0,0,147,0,0,0,35,0,114,0,114,0,74,0,88,0,235,0,129,0,76,0,62,0,212,0,13,0,213,0,0,0,250,0,0,0,226,0,131,0,71,0,189,0,129,0,138,0,74,0,84,0,166,0,115,0,11,0,0,0,8,0,87,0,182,0,0,0,21,0,255,0,2,0,165,0,197,0,98,0,65,0,23,0,116,0,0,0,14,0,76,0,136,0,246,0,232,0,35,0,144,0,57,0,0,0,88,0,56,0,66,0,30,0,0,0,206,0,161,0,40,0,95,0,0,0,43,0,51,0,225,0,0,0,6,0,213,0,117,0,159,0,247,0,92,0,197,0,23,0,0,0,139,0,0,0,252,0,0,0,0,0,213,0,0,0,56,0,49,0,0,0,250,0,146,0,15,0,196,0,0,0,209,0,96,0,178,0,181,0,0,0,226,0,224,0,87,0,191,0,48,0,12,0,77,0,235,0,0,0,249,0,77,0,65,0,89,0,255,0,60,0,25,0,204,0,64,0,110,0,148,0,150,0,159,0,103,0,58,0,73,0,0,0,0,0,0,0,51,0,0,0,39,0,79,0,0,0,0,0,239,0,147,0,30,0,0,0,97,0,13,0,75,0,106,0,81,0,223,0,0,0,107,0,74,0,108,0,0,0,112,0,241,0,196,0,195,0,210,0,221,0,188,0,213,0,113,0,200,0,113,0,201,0,1,0,0,0,117,0,0,0,4,0,75,0,129,0,231,0,0,0,172,0,3,0,0,0,0,0,0,0,83,0,0,0,198,0,0,0,176,0,193,0,211,0,32,0,51,0,252,0,0,0,37,0,0,0,136,0,157,0,193,0,242,0,0,0,0,0,160,0,178,0,150,0,64,0,165,0,223,0,209,0,43,0,146,0,0,0,107,0,42,0,218,0,0,0,105,0,134,0,113,0,47,0,0,0,63,0,69,0,143,0,16,0,46,0,62,0,71,0,64,0,0,0,0,0,195,0,62,0,212,0,209,0,44,0,156,0,128,0,18,0,215,0,86,0,167,0,189,0,109,0,108,0,22,0,202,0,76,0,0,0,150,0,103,0,31,0,179,0,92,0,232,0,0,0,142,0,25,0,179,0,78,0,53,0,71,0,192,0,4,0,117,0,73,0,12,0,42,0,42,0,124,0,109,0,56,0,0,0,0,0,219,0,0,0,0,0,13,0,0,0,25,0,53,0,174,0,0,0,22,0,183,0,113,0,149,0,128,0,7,0,51,0,227,0,247,0,119,0,155,0,51,0,223,0,144,0,245,0,135,0,185,0,0,0,68,0,100,0,246,0,0,0,205,0,140,0,86,0,195,0,0,0,165,0,29,0,146,0,251,0,0,0,68,0,234,0,5,0,2,0,121,0,0,0,96,0,95,0,223,0,0,0,63,0,38,0,0,0,0,0,240,0,191,0,235,0,72,0,123,0,64,0,111,0,205,0,187,0,167,0,235,0,160,0,38,0,130,0,222,0,0,0,98,0,0,0,4,0,21,0,11,0,48,0,204,0,132,0,166,0,207,0,0,0,0,0,0,0,0,0,193,0,197,0,3,0,33,0,106,0,0,0,28,0,225,0,117,0,224,0,56,0,120,0,142,0,0,0,175,0,68,0,72,0,94,0,82,0,75,0,0,0,0,0,72,0,106,0,121,0,226,0,55,0,144,0,175,0,141,0,117,0,0,0,94,0,105,0,163,0,215,0,243,0,136,0,208,0,27,0,0,0,0,0,223,0,0,0,214,0,117,0,16,0,1,0,208,0,215,0,0,0,148,0,0,0,26,0,116,0,0,0,166,0,29,0,116,0,0,0,203,0,252,0,91,0,0,0,235,0,168,0,94,0,24,0,116,0,135,0,47,0,224,0,28,0,65,0,255,0,15,0,180,0,0,0,1,0,0,0,145,0,184,0,205,0,118,0,219,0,29,0,50,0,0,0,89,0,98,0,179,0,42,0,23,0,69,0,74,0,17,0,117,0,104,0,207,0,73,0,0,0,34,0,21,0,201,0,0,0,0,0,0,0,34,0,242,0,143,0,95,0,21,0,0,0,93,0,94,0,110,0,0,0,172,0,114,0,150,0,185,0,0,0,39,0,192,0,27,0,145,0,236,0,221,0,67,0,0,0,106,0,102,0,228,0,247,0,5,0,63,0,70,0,84,0,155,0,154,0,121,0,0,0,109,0,180,0,0,0,46,0,0,0,91,0,182,0,114,0,0,0,233,0,85,0,149,0,95,0,0,0,80,0,208,0,0,0,95,0,132,0,102,0,170,0,29,0,70,0,0,0,55,0,203,0,232,0,0,0,61,0,54,0,119,0,232,0,61,0,0,0,249,0,101,0,0,0,197,0,115,0,37,0,128,0,197,0,105,0,161,0,123,0,246,0,133,0,174,0,0,0,220,0,91,0,218,0,66,0,253,0,0,0,0,0,165,0,39,0,0,0,162,0,93,0,0,0,62,0,103,0,49,0,150,0,4,0,250,0,175,0,0,0,221,0,94,0,0,0,162,0,44,0,59,0,46,0,102,0,161,0,0,0,108,0,135,0,0,0,235,0,199,0,133,0,192,0,0,0,223,0,168,0,85,0,0,0,107,0,190,0,178,0,219,0,112,0,47,0,159,0,191,0,0,0,6,0,239,0,61,0,141,0,163,0,50,0,208,0,0,0,232,0,213,0,12,0,164,0,134,0,0,0,189,0,219,0,101,0,13,0,131,0,200,0,23,0,44,0,179,0,0,0,106,0,122,0,25,0,243,0,84,0,127,0,153,0,130,0,167,0,255,0,40,0,163,0,216,0,129,0,155,0,0,0,53,0,150,0,44,0,0,0,55,0,0,0,163,0,0,0,197,0,15,0,0,0,213,0,193,0,83,0,220,0,181,0,102,0,12,0,105,0,70,0,0,0,177,0,209,0,0,0,68,0,194,0,0,0,155,0,44,0,0,0,38,0,197,0,12,0,156,0,0,0,95,0,3,0,188,0,58,0,178,0,0,0,229,0,245,0,21,0,2,0,24,0,62,0,230,0,174,0,180,0,79,0,77,0,0,0,196,0,77,0,0,0,103,0,22,0,0,0,146,0,0,0,33,0,220,0,225,0,0,0,38,0,6,0,239,0,0,0,1,0,40,0,181,0,53,0,38,0,16,0,182,0,0,0,206,0,55,0,231,0,0,0,0,0,0,0,107,0,235,0,194,0,184,0,147,0,0,0,182,0,173,0,152,0,192,0,0,0,49,0,0,0,132,0,180,0,238,0,43,0,40,0,206,0,0,0,36,0,44,0,0,0,0,0,81,0,163,0,89,0,190,0,0,0,89,0,195,0,103,0,0,0,30,0,6,0,0,0,0,0,191,0,209,0,33,0,123,0,0,0,149,0,124,0);
signal scenario_full  : scenario_type := (119,31,210,31,36,31,36,30,75,31,50,31,76,31,75,31,212,31,252,31,169,31,210,31,210,30,217,31,38,31,144,31,144,30,23,31,168,31,247,31,247,30,168,31,168,30,168,29,236,31,189,31,10,31,43,31,154,31,219,31,179,31,86,31,112,31,15,31,15,30,10,31,39,31,102,31,209,31,118,31,133,31,76,31,76,30,76,29,209,31,8,31,86,31,250,31,172,31,63,31,122,31,254,31,18,31,18,30,101,31,39,31,107,31,24,31,48,31,42,31,216,31,61,31,40,31,254,31,140,31,102,31,166,31,135,31,31,31,114,31,43,31,124,31,62,31,102,31,128,31,218,31,42,31,124,31,172,31,211,31,211,30,214,31,214,30,147,31,7,31,123,31,199,31,199,30,115,31,110,31,110,30,5,31,232,31,179,31,242,31,242,30,188,31,188,30,67,31,212,31,63,31,39,31,70,31,66,31,71,31,104,31,104,30,126,31,16,31,109,31,206,31,159,31,75,31,75,30,251,31,15,31,116,31,63,31,63,30,210,31,226,31,226,30,187,31,201,31,60,31,12,31,27,31,104,31,117,31,89,31,26,31,61,31,21,31,31,31,31,30,69,31,183,31,97,31,37,31,206,31,118,31,71,31,13,31,13,30,86,31,86,30,86,29,8,31,246,31,133,31,30,31,89,31,197,31,99,31,51,31,183,31,183,30,137,31,161,31,66,31,28,31,28,31,28,30,28,29,184,31,184,30,47,31,219,31,219,30,112,31,138,31,152,31,148,31,242,31,242,30,94,31,96,31,72,31,85,31,56,31,56,30,56,29,98,31,98,30,40,31,90,31,12,31,148,31,148,30,147,31,147,30,35,31,114,31,114,31,74,31,88,31,235,31,129,31,76,31,62,31,212,31,13,31,213,31,213,30,250,31,250,30,226,31,131,31,71,31,189,31,129,31,138,31,74,31,84,31,166,31,115,31,11,31,11,30,8,31,87,31,182,31,182,30,21,31,255,31,2,31,165,31,197,31,98,31,65,31,23,31,116,31,116,30,14,31,76,31,136,31,246,31,232,31,35,31,144,31,57,31,57,30,88,31,56,31,66,31,30,31,30,30,206,31,161,31,40,31,95,31,95,30,43,31,51,31,225,31,225,30,6,31,213,31,117,31,159,31,247,31,92,31,197,31,23,31,23,30,139,31,139,30,252,31,252,30,252,29,213,31,213,30,56,31,49,31,49,30,250,31,146,31,15,31,196,31,196,30,209,31,96,31,178,31,181,31,181,30,226,31,224,31,87,31,191,31,48,31,12,31,77,31,235,31,235,30,249,31,77,31,65,31,89,31,255,31,60,31,25,31,204,31,64,31,110,31,148,31,150,31,159,31,103,31,58,31,73,31,73,30,73,29,73,28,51,31,51,30,39,31,79,31,79,30,79,29,239,31,147,31,30,31,30,30,97,31,13,31,75,31,106,31,81,31,223,31,223,30,107,31,74,31,108,31,108,30,112,31,241,31,196,31,195,31,210,31,221,31,188,31,213,31,113,31,200,31,113,31,201,31,1,31,1,30,117,31,117,30,4,31,75,31,129,31,231,31,231,30,172,31,3,31,3,30,3,29,3,28,83,31,83,30,198,31,198,30,176,31,193,31,211,31,32,31,51,31,252,31,252,30,37,31,37,30,136,31,157,31,193,31,242,31,242,30,242,29,160,31,178,31,150,31,64,31,165,31,223,31,209,31,43,31,146,31,146,30,107,31,42,31,218,31,218,30,105,31,134,31,113,31,47,31,47,30,63,31,69,31,143,31,16,31,46,31,62,31,71,31,64,31,64,30,64,29,195,31,62,31,212,31,209,31,44,31,156,31,128,31,18,31,215,31,86,31,167,31,189,31,109,31,108,31,22,31,202,31,76,31,76,30,150,31,103,31,31,31,179,31,92,31,232,31,232,30,142,31,25,31,179,31,78,31,53,31,71,31,192,31,4,31,117,31,73,31,12,31,42,31,42,31,124,31,109,31,56,31,56,30,56,29,219,31,219,30,219,29,13,31,13,30,25,31,53,31,174,31,174,30,22,31,183,31,113,31,149,31,128,31,7,31,51,31,227,31,247,31,119,31,155,31,51,31,223,31,144,31,245,31,135,31,185,31,185,30,68,31,100,31,246,31,246,30,205,31,140,31,86,31,195,31,195,30,165,31,29,31,146,31,251,31,251,30,68,31,234,31,5,31,2,31,121,31,121,30,96,31,95,31,223,31,223,30,63,31,38,31,38,30,38,29,240,31,191,31,235,31,72,31,123,31,64,31,111,31,205,31,187,31,167,31,235,31,160,31,38,31,130,31,222,31,222,30,98,31,98,30,4,31,21,31,11,31,48,31,204,31,132,31,166,31,207,31,207,30,207,29,207,28,207,27,193,31,197,31,3,31,33,31,106,31,106,30,28,31,225,31,117,31,224,31,56,31,120,31,142,31,142,30,175,31,68,31,72,31,94,31,82,31,75,31,75,30,75,29,72,31,106,31,121,31,226,31,55,31,144,31,175,31,141,31,117,31,117,30,94,31,105,31,163,31,215,31,243,31,136,31,208,31,27,31,27,30,27,29,223,31,223,30,214,31,117,31,16,31,1,31,208,31,215,31,215,30,148,31,148,30,26,31,116,31,116,30,166,31,29,31,116,31,116,30,203,31,252,31,91,31,91,30,235,31,168,31,94,31,24,31,116,31,135,31,47,31,224,31,28,31,65,31,255,31,15,31,180,31,180,30,1,31,1,30,145,31,184,31,205,31,118,31,219,31,29,31,50,31,50,30,89,31,98,31,179,31,42,31,23,31,69,31,74,31,17,31,117,31,104,31,207,31,73,31,73,30,34,31,21,31,201,31,201,30,201,29,201,28,34,31,242,31,143,31,95,31,21,31,21,30,93,31,94,31,110,31,110,30,172,31,114,31,150,31,185,31,185,30,39,31,192,31,27,31,145,31,236,31,221,31,67,31,67,30,106,31,102,31,228,31,247,31,5,31,63,31,70,31,84,31,155,31,154,31,121,31,121,30,109,31,180,31,180,30,46,31,46,30,91,31,182,31,114,31,114,30,233,31,85,31,149,31,95,31,95,30,80,31,208,31,208,30,95,31,132,31,102,31,170,31,29,31,70,31,70,30,55,31,203,31,232,31,232,30,61,31,54,31,119,31,232,31,61,31,61,30,249,31,101,31,101,30,197,31,115,31,37,31,128,31,197,31,105,31,161,31,123,31,246,31,133,31,174,31,174,30,220,31,91,31,218,31,66,31,253,31,253,30,253,29,165,31,39,31,39,30,162,31,93,31,93,30,62,31,103,31,49,31,150,31,4,31,250,31,175,31,175,30,221,31,94,31,94,30,162,31,44,31,59,31,46,31,102,31,161,31,161,30,108,31,135,31,135,30,235,31,199,31,133,31,192,31,192,30,223,31,168,31,85,31,85,30,107,31,190,31,178,31,219,31,112,31,47,31,159,31,191,31,191,30,6,31,239,31,61,31,141,31,163,31,50,31,208,31,208,30,232,31,213,31,12,31,164,31,134,31,134,30,189,31,219,31,101,31,13,31,131,31,200,31,23,31,44,31,179,31,179,30,106,31,122,31,25,31,243,31,84,31,127,31,153,31,130,31,167,31,255,31,40,31,163,31,216,31,129,31,155,31,155,30,53,31,150,31,44,31,44,30,55,31,55,30,163,31,163,30,197,31,15,31,15,30,213,31,193,31,83,31,220,31,181,31,102,31,12,31,105,31,70,31,70,30,177,31,209,31,209,30,68,31,194,31,194,30,155,31,44,31,44,30,38,31,197,31,12,31,156,31,156,30,95,31,3,31,188,31,58,31,178,31,178,30,229,31,245,31,21,31,2,31,24,31,62,31,230,31,174,31,180,31,79,31,77,31,77,30,196,31,77,31,77,30,103,31,22,31,22,30,146,31,146,30,33,31,220,31,225,31,225,30,38,31,6,31,239,31,239,30,1,31,40,31,181,31,53,31,38,31,16,31,182,31,182,30,206,31,55,31,231,31,231,30,231,29,231,28,107,31,235,31,194,31,184,31,147,31,147,30,182,31,173,31,152,31,192,31,192,30,49,31,49,30,132,31,180,31,238,31,43,31,40,31,206,31,206,30,36,31,44,31,44,30,44,29,81,31,163,31,89,31,190,31,190,30,89,31,195,31,103,31,103,30,30,31,6,31,6,30,6,29,191,31,209,31,33,31,123,31,123,30,149,31,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
