-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 429;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (208,0,96,0,81,0,0,0,194,0,44,0,157,0,177,0,194,0,27,0,7,0,188,0,155,0,161,0,0,0,38,0,0,0,161,0,0,0,44,0,0,0,124,0,0,0,175,0,136,0,212,0,155,0,174,0,73,0,191,0,13,0,0,0,163,0,125,0,67,0,66,0,38,0,19,0,131,0,226,0,0,0,130,0,20,0,120,0,98,0,253,0,49,0,93,0,159,0,0,0,234,0,165,0,0,0,179,0,0,0,28,0,57,0,0,0,0,0,111,0,105,0,0,0,0,0,184,0,204,0,176,0,206,0,174,0,193,0,0,0,34,0,190,0,81,0,102,0,90,0,143,0,62,0,34,0,254,0,177,0,126,0,0,0,205,0,0,0,152,0,71,0,0,0,0,0,218,0,136,0,0,0,168,0,54,0,152,0,79,0,211,0,209,0,69,0,226,0,210,0,0,0,208,0,149,0,211,0,135,0,94,0,150,0,0,0,186,0,174,0,59,0,0,0,161,0,183,0,0,0,130,0,0,0,55,0,0,0,199,0,241,0,146,0,24,0,92,0,209,0,61,0,126,0,224,0,144,0,214,0,47,0,54,0,85,0,62,0,108,0,60,0,231,0,12,0,108,0,34,0,160,0,126,0,208,0,82,0,70,0,161,0,1,0,153,0,127,0,145,0,103,0,0,0,0,0,229,0,96,0,152,0,66,0,141,0,0,0,0,0,83,0,204,0,34,0,0,0,82,0,0,0,195,0,65,0,99,0,0,0,83,0,90,0,215,0,0,0,107,0,176,0,0,0,134,0,55,0,0,0,0,0,104,0,99,0,158,0,72,0,132,0,236,0,119,0,0,0,108,0,22,0,0,0,87,0,27,0,238,0,77,0,0,0,28,0,0,0,51,0,165,0,230,0,205,0,253,0,0,0,227,0,188,0,2,0,45,0,0,0,37,0,0,0,0,0,253,0,188,0,149,0,200,0,51,0,213,0,0,0,11,0,177,0,132,0,168,0,227,0,0,0,0,0,0,0,171,0,25,0,32,0,203,0,177,0,0,0,63,0,109,0,210,0,107,0,171,0,154,0,250,0,118,0,129,0,142,0,0,0,178,0,240,0,154,0,4,0,171,0,239,0,0,0,0,0,221,0,199,0,154,0,0,0,27,0,13,0,248,0,37,0,194,0,232,0,162,0,40,0,208,0,116,0,32,0,0,0,121,0,63,0,95,0,11,0,1,0,0,0,0,0,116,0,178,0,15,0,4,0,238,0,85,0,255,0,112,0,181,0,166,0,0,0,51,0,70,0,237,0,0,0,174,0,0,0,201,0,143,0,101,0,89,0,132,0,37,0,52,0,0,0,35,0,4,0,253,0,102,0,128,0,0,0,88,0,225,0,151,0,0,0,237,0,87,0,248,0,58,0,45,0,63,0,125,0,150,0,57,0,142,0,101,0,42,0,0,0,146,0,102,0,240,0,209,0,56,0,37,0,120,0,166,0,198,0,28,0,254,0,114,0,229,0,122,0,0,0,113,0,61,0,143,0,218,0,39,0,212,0,87,0,54,0,51,0,49,0,109,0,1,0,32,0,0,0,208,0,179,0,215,0,0,0,0,0,0,0,81,0,224,0,49,0,102,0,72,0,0,0,187,0,226,0,0,0,254,0,207,0,254,0,4,0,87,0,0,0,26,0,13,0,140,0,151,0,8,0,157,0,71,0,127,0,93,0,0,0,247,0,223,0,14,0,93,0,116,0,171,0,0,0,47,0,157,0,42,0,103,0,249,0,182,0,74,0,176,0,0,0,0,0,15,0,229,0,69,0,48,0,209,0,34,0,127,0,153,0,219,0,0,0,197,0,186,0,129,0,120,0,149,0,87,0,9,0,67,0,0,0,113,0,0,0,0,0,169,0,138,0,0,0,157,0,116,0,61,0);
signal scenario_full  : scenario_type := (208,31,96,31,81,31,81,30,194,31,44,31,157,31,177,31,194,31,27,31,7,31,188,31,155,31,161,31,161,30,38,31,38,30,161,31,161,30,44,31,44,30,124,31,124,30,175,31,136,31,212,31,155,31,174,31,73,31,191,31,13,31,13,30,163,31,125,31,67,31,66,31,38,31,19,31,131,31,226,31,226,30,130,31,20,31,120,31,98,31,253,31,49,31,93,31,159,31,159,30,234,31,165,31,165,30,179,31,179,30,28,31,57,31,57,30,57,29,111,31,105,31,105,30,105,29,184,31,204,31,176,31,206,31,174,31,193,31,193,30,34,31,190,31,81,31,102,31,90,31,143,31,62,31,34,31,254,31,177,31,126,31,126,30,205,31,205,30,152,31,71,31,71,30,71,29,218,31,136,31,136,30,168,31,54,31,152,31,79,31,211,31,209,31,69,31,226,31,210,31,210,30,208,31,149,31,211,31,135,31,94,31,150,31,150,30,186,31,174,31,59,31,59,30,161,31,183,31,183,30,130,31,130,30,55,31,55,30,199,31,241,31,146,31,24,31,92,31,209,31,61,31,126,31,224,31,144,31,214,31,47,31,54,31,85,31,62,31,108,31,60,31,231,31,12,31,108,31,34,31,160,31,126,31,208,31,82,31,70,31,161,31,1,31,153,31,127,31,145,31,103,31,103,30,103,29,229,31,96,31,152,31,66,31,141,31,141,30,141,29,83,31,204,31,34,31,34,30,82,31,82,30,195,31,65,31,99,31,99,30,83,31,90,31,215,31,215,30,107,31,176,31,176,30,134,31,55,31,55,30,55,29,104,31,99,31,158,31,72,31,132,31,236,31,119,31,119,30,108,31,22,31,22,30,87,31,27,31,238,31,77,31,77,30,28,31,28,30,51,31,165,31,230,31,205,31,253,31,253,30,227,31,188,31,2,31,45,31,45,30,37,31,37,30,37,29,253,31,188,31,149,31,200,31,51,31,213,31,213,30,11,31,177,31,132,31,168,31,227,31,227,30,227,29,227,28,171,31,25,31,32,31,203,31,177,31,177,30,63,31,109,31,210,31,107,31,171,31,154,31,250,31,118,31,129,31,142,31,142,30,178,31,240,31,154,31,4,31,171,31,239,31,239,30,239,29,221,31,199,31,154,31,154,30,27,31,13,31,248,31,37,31,194,31,232,31,162,31,40,31,208,31,116,31,32,31,32,30,121,31,63,31,95,31,11,31,1,31,1,30,1,29,116,31,178,31,15,31,4,31,238,31,85,31,255,31,112,31,181,31,166,31,166,30,51,31,70,31,237,31,237,30,174,31,174,30,201,31,143,31,101,31,89,31,132,31,37,31,52,31,52,30,35,31,4,31,253,31,102,31,128,31,128,30,88,31,225,31,151,31,151,30,237,31,87,31,248,31,58,31,45,31,63,31,125,31,150,31,57,31,142,31,101,31,42,31,42,30,146,31,102,31,240,31,209,31,56,31,37,31,120,31,166,31,198,31,28,31,254,31,114,31,229,31,122,31,122,30,113,31,61,31,143,31,218,31,39,31,212,31,87,31,54,31,51,31,49,31,109,31,1,31,32,31,32,30,208,31,179,31,215,31,215,30,215,29,215,28,81,31,224,31,49,31,102,31,72,31,72,30,187,31,226,31,226,30,254,31,207,31,254,31,4,31,87,31,87,30,26,31,13,31,140,31,151,31,8,31,157,31,71,31,127,31,93,31,93,30,247,31,223,31,14,31,93,31,116,31,171,31,171,30,47,31,157,31,42,31,103,31,249,31,182,31,74,31,176,31,176,30,176,29,15,31,229,31,69,31,48,31,209,31,34,31,127,31,153,31,219,31,219,30,197,31,186,31,129,31,120,31,149,31,87,31,9,31,67,31,67,30,113,31,113,30,113,29,169,31,138,31,138,30,157,31,116,31,61,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
