-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 944;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (67,0,145,0,187,0,0,0,90,0,242,0,195,0,228,0,177,0,0,0,159,0,33,0,136,0,121,0,236,0,91,0,117,0,254,0,209,0,174,0,255,0,0,0,0,0,147,0,255,0,3,0,128,0,105,0,184,0,0,0,35,0,235,0,0,0,8,0,56,0,0,0,0,0,118,0,0,0,53,0,59,0,77,0,0,0,89,0,212,0,254,0,7,0,236,0,8,0,102,0,29,0,42,0,235,0,123,0,0,0,248,0,35,0,156,0,242,0,172,0,0,0,164,0,205,0,0,0,137,0,91,0,254,0,232,0,52,0,139,0,0,0,38,0,105,0,0,0,0,0,0,0,0,0,183,0,178,0,0,0,45,0,79,0,61,0,129,0,222,0,13,0,0,0,0,0,147,0,0,0,0,0,18,0,89,0,82,0,255,0,38,0,62,0,0,0,98,0,160,0,0,0,58,0,254,0,118,0,123,0,174,0,69,0,229,0,68,0,236,0,78,0,14,0,71,0,24,0,178,0,43,0,146,0,29,0,5,0,250,0,0,0,60,0,57,0,190,0,175,0,56,0,0,0,145,0,28,0,210,0,215,0,115,0,230,0,47,0,81,0,54,0,210,0,136,0,23,0,238,0,75,0,111,0,221,0,90,0,97,0,160,0,13,0,218,0,0,0,200,0,0,0,0,0,144,0,84,0,29,0,61,0,141,0,170,0,184,0,177,0,44,0,15,0,107,0,73,0,222,0,231,0,132,0,163,0,218,0,21,0,160,0,230,0,56,0,226,0,0,0,131,0,226,0,25,0,0,0,247,0,0,0,36,0,174,0,123,0,29,0,50,0,124,0,159,0,6,0,179,0,3,0,86,0,180,0,0,0,0,0,66,0,167,0,193,0,68,0,92,0,221,0,125,0,74,0,123,0,40,0,0,0,0,0,0,0,178,0,26,0,0,0,0,0,59,0,0,0,0,0,0,0,132,0,75,0,0,0,54,0,114,0,227,0,33,0,0,0,114,0,21,0,106,0,115,0,51,0,191,0,125,0,48,0,108,0,142,0,191,0,0,0,0,0,0,0,39,0,151,0,135,0,81,0,156,0,199,0,0,0,234,0,37,0,220,0,206,0,167,0,68,0,10,0,0,0,0,0,32,0,251,0,181,0,166,0,111,0,0,0,57,0,13,0,194,0,177,0,59,0,0,0,89,0,25,0,0,0,0,0,238,0,46,0,98,0,200,0,191,0,0,0,159,0,129,0,240,0,164,0,59,0,115,0,0,0,9,0,32,0,0,0,0,0,131,0,146,0,16,0,138,0,0,0,0,0,33,0,166,0,0,0,0,0,169,0,71,0,154,0,251,0,0,0,59,0,140,0,81,0,175,0,103,0,0,0,102,0,0,0,0,0,30,0,234,0,158,0,0,0,255,0,0,0,0,0,174,0,244,0,44,0,0,0,96,0,253,0,77,0,102,0,92,0,105,0,106,0,233,0,10,0,102,0,54,0,99,0,0,0,0,0,247,0,255,0,68,0,64,0,0,0,0,0,245,0,165,0,0,0,0,0,167,0,250,0,62,0,238,0,21,0,234,0,71,0,135,0,0,0,0,0,206,0,0,0,41,0,88,0,240,0,113,0,0,0,90,0,93,0,0,0,118,0,0,0,63,0,72,0,84,0,84,0,77,0,145,0,134,0,229,0,0,0,0,0,0,0,253,0,28,0,100,0,41,0,140,0,75,0,3,0,90,0,22,0,83,0,90,0,209,0,180,0,50,0,159,0,44,0,12,0,0,0,115,0,241,0,60,0,190,0,39,0,46,0,161,0,138,0,165,0,34,0,5,0,32,0,116,0,126,0,213,0,102,0,246,0,18,0,46,0,0,0,0,0,121,0,232,0,155,0,0,0,243,0,173,0,227,0,65,0,31,0,250,0,227,0,176,0,0,0,0,0,89,0,184,0,163,0,0,0,251,0,0,0,81,0,146,0,140,0,0,0,0,0,178,0,0,0,99,0,0,0,20,0,229,0,190,0,76,0,170,0,114,0,0,0,196,0,174,0,164,0,216,0,134,0,246,0,135,0,0,0,29,0,122,0,242,0,248,0,47,0,69,0,222,0,209,0,17,0,199,0,47,0,149,0,0,0,236,0,21,0,17,0,215,0,51,0,199,0,182,0,246,0,90,0,203,0,87,0,138,0,0,0,62,0,0,0,74,0,42,0,0,0,11,0,91,0,211,0,193,0,98,0,255,0,80,0,0,0,26,0,215,0,0,0,247,0,140,0,3,0,190,0,25,0,177,0,11,0,62,0,125,0,0,0,192,0,51,0,23,0,20,0,161,0,124,0,7,0,193,0,146,0,162,0,164,0,123,0,0,0,102,0,175,0,195,0,68,0,246,0,165,0,2,0,240,0,0,0,188,0,0,0,137,0,177,0,0,0,136,0,15,0,211,0,0,0,146,0,209,0,251,0,195,0,0,0,224,0,124,0,26,0,224,0,0,0,225,0,0,0,124,0,115,0,173,0,191,0,139,0,65,0,144,0,171,0,0,0,0,0,0,0,143,0,1,0,123,0,0,0,203,0,60,0,206,0,128,0,80,0,151,0,20,0,28,0,212,0,160,0,0,0,0,0,224,0,0,0,188,0,54,0,0,0,0,0,206,0,165,0,88,0,0,0,215,0,0,0,201,0,0,0,81,0,92,0,138,0,221,0,57,0,2,0,119,0,0,0,82,0,18,0,114,0,210,0,0,0,169,0,0,0,121,0,196,0,103,0,96,0,138,0,35,0,57,0,52,0,112,0,4,0,128,0,176,0,135,0,151,0,0,0,255,0,50,0,125,0,0,0,3,0,183,0,110,0,199,0,210,0,0,0,0,0,0,0,0,0,20,0,0,0,173,0,0,0,0,0,216,0,0,0,250,0,31,0,149,0,0,0,151,0,139,0,175,0,12,0,86,0,219,0,0,0,0,0,79,0,0,0,0,0,194,0,219,0,231,0,88,0,186,0,125,0,22,0,0,0,136,0,86,0,0,0,95,0,0,0,0,0,0,0,203,0,255,0,248,0,71,0,49,0,0,0,70,0,82,0,0,0,115,0,115,0,191,0,58,0,0,0,81,0,88,0,0,0,34,0,0,0,133,0,231,0,178,0,0,0,0,0,0,0,91,0,161,0,220,0,0,0,106,0,70,0,55,0,189,0,155,0,213,0,136,0,43,0,0,0,247,0,168,0,206,0,66,0,81,0,183,0,92,0,231,0,203,0,222,0,126,0,254,0,39,0,164,0,32,0,145,0,159,0,129,0,133,0,0,0,191,0,91,0,58,0,89,0,254,0,204,0,20,0,0,0,0,0,0,0,145,0,0,0,0,0,254,0,134,0,2,0,138,0,204,0,86,0,246,0,9,0,103,0,83,0,0,0,210,0,20,0,231,0,167,0,76,0,78,0,64,0,0,0,33,0,150,0,59,0,126,0,125,0,98,0,193,0,21,0,221,0,63,0,213,0,93,0,18,0,0,0,180,0,92,0,33,0,34,0,0,0,202,0,161,0,249,0,0,0,70,0,54,0,28,0,62,0,87,0,0,0,196,0,125,0,134,0,239,0,14,0,247,0,57,0,51,0,165,0,99,0,76,0,0,0,49,0,0,0,117,0,223,0,77,0,250,0,0,0,150,0,173,0,254,0,0,0,89,0,161,0,202,0,236,0,0,0,190,0,99,0,103,0,89,0,117,0,65,0,206,0,79,0,172,0,226,0,200,0,0,0,39,0,0,0,117,0,126,0,152,0,58,0,34,0,186,0,115,0,184,0,22,0,114,0,161,0,0,0,101,0,17,0,0,0,165,0,171,0,193,0,0,0,254,0,0,0,187,0,25,0,222,0,88,0,1,0,127,0,195,0,93,0,0,0,231,0,206,0,184,0,106,0,98,0,55,0,0,0,232,0,0,0,102,0,0,0,237,0,35,0,0,0,0,0,83,0,116,0,129,0,90,0,179,0,8,0,0,0,0,0,124,0,149,0,157,0,35,0,238,0,74,0,234,0,38,0,144,0,14,0,192,0,0,0,0,0,50,0,49,0,14,0,0,0,147,0,0,0,7,0,76,0,235,0,235,0,215,0,0,0,170,0,217,0,177,0,0,0,252,0,61,0,29,0,80,0,86,0,0,0,62,0,0,0,37,0,171,0,168,0,243,0,40,0,119,0,82,0,80,0,48,0,236,0,129,0,0,0,86,0,176,0,128,0);
signal scenario_full  : scenario_type := (67,31,145,31,187,31,187,30,90,31,242,31,195,31,228,31,177,31,177,30,159,31,33,31,136,31,121,31,236,31,91,31,117,31,254,31,209,31,174,31,255,31,255,30,255,29,147,31,255,31,3,31,128,31,105,31,184,31,184,30,35,31,235,31,235,30,8,31,56,31,56,30,56,29,118,31,118,30,53,31,59,31,77,31,77,30,89,31,212,31,254,31,7,31,236,31,8,31,102,31,29,31,42,31,235,31,123,31,123,30,248,31,35,31,156,31,242,31,172,31,172,30,164,31,205,31,205,30,137,31,91,31,254,31,232,31,52,31,139,31,139,30,38,31,105,31,105,30,105,29,105,28,105,27,183,31,178,31,178,30,45,31,79,31,61,31,129,31,222,31,13,31,13,30,13,29,147,31,147,30,147,29,18,31,89,31,82,31,255,31,38,31,62,31,62,30,98,31,160,31,160,30,58,31,254,31,118,31,123,31,174,31,69,31,229,31,68,31,236,31,78,31,14,31,71,31,24,31,178,31,43,31,146,31,29,31,5,31,250,31,250,30,60,31,57,31,190,31,175,31,56,31,56,30,145,31,28,31,210,31,215,31,115,31,230,31,47,31,81,31,54,31,210,31,136,31,23,31,238,31,75,31,111,31,221,31,90,31,97,31,160,31,13,31,218,31,218,30,200,31,200,30,200,29,144,31,84,31,29,31,61,31,141,31,170,31,184,31,177,31,44,31,15,31,107,31,73,31,222,31,231,31,132,31,163,31,218,31,21,31,160,31,230,31,56,31,226,31,226,30,131,31,226,31,25,31,25,30,247,31,247,30,36,31,174,31,123,31,29,31,50,31,124,31,159,31,6,31,179,31,3,31,86,31,180,31,180,30,180,29,66,31,167,31,193,31,68,31,92,31,221,31,125,31,74,31,123,31,40,31,40,30,40,29,40,28,178,31,26,31,26,30,26,29,59,31,59,30,59,29,59,28,132,31,75,31,75,30,54,31,114,31,227,31,33,31,33,30,114,31,21,31,106,31,115,31,51,31,191,31,125,31,48,31,108,31,142,31,191,31,191,30,191,29,191,28,39,31,151,31,135,31,81,31,156,31,199,31,199,30,234,31,37,31,220,31,206,31,167,31,68,31,10,31,10,30,10,29,32,31,251,31,181,31,166,31,111,31,111,30,57,31,13,31,194,31,177,31,59,31,59,30,89,31,25,31,25,30,25,29,238,31,46,31,98,31,200,31,191,31,191,30,159,31,129,31,240,31,164,31,59,31,115,31,115,30,9,31,32,31,32,30,32,29,131,31,146,31,16,31,138,31,138,30,138,29,33,31,166,31,166,30,166,29,169,31,71,31,154,31,251,31,251,30,59,31,140,31,81,31,175,31,103,31,103,30,102,31,102,30,102,29,30,31,234,31,158,31,158,30,255,31,255,30,255,29,174,31,244,31,44,31,44,30,96,31,253,31,77,31,102,31,92,31,105,31,106,31,233,31,10,31,102,31,54,31,99,31,99,30,99,29,247,31,255,31,68,31,64,31,64,30,64,29,245,31,165,31,165,30,165,29,167,31,250,31,62,31,238,31,21,31,234,31,71,31,135,31,135,30,135,29,206,31,206,30,41,31,88,31,240,31,113,31,113,30,90,31,93,31,93,30,118,31,118,30,63,31,72,31,84,31,84,31,77,31,145,31,134,31,229,31,229,30,229,29,229,28,253,31,28,31,100,31,41,31,140,31,75,31,3,31,90,31,22,31,83,31,90,31,209,31,180,31,50,31,159,31,44,31,12,31,12,30,115,31,241,31,60,31,190,31,39,31,46,31,161,31,138,31,165,31,34,31,5,31,32,31,116,31,126,31,213,31,102,31,246,31,18,31,46,31,46,30,46,29,121,31,232,31,155,31,155,30,243,31,173,31,227,31,65,31,31,31,250,31,227,31,176,31,176,30,176,29,89,31,184,31,163,31,163,30,251,31,251,30,81,31,146,31,140,31,140,30,140,29,178,31,178,30,99,31,99,30,20,31,229,31,190,31,76,31,170,31,114,31,114,30,196,31,174,31,164,31,216,31,134,31,246,31,135,31,135,30,29,31,122,31,242,31,248,31,47,31,69,31,222,31,209,31,17,31,199,31,47,31,149,31,149,30,236,31,21,31,17,31,215,31,51,31,199,31,182,31,246,31,90,31,203,31,87,31,138,31,138,30,62,31,62,30,74,31,42,31,42,30,11,31,91,31,211,31,193,31,98,31,255,31,80,31,80,30,26,31,215,31,215,30,247,31,140,31,3,31,190,31,25,31,177,31,11,31,62,31,125,31,125,30,192,31,51,31,23,31,20,31,161,31,124,31,7,31,193,31,146,31,162,31,164,31,123,31,123,30,102,31,175,31,195,31,68,31,246,31,165,31,2,31,240,31,240,30,188,31,188,30,137,31,177,31,177,30,136,31,15,31,211,31,211,30,146,31,209,31,251,31,195,31,195,30,224,31,124,31,26,31,224,31,224,30,225,31,225,30,124,31,115,31,173,31,191,31,139,31,65,31,144,31,171,31,171,30,171,29,171,28,143,31,1,31,123,31,123,30,203,31,60,31,206,31,128,31,80,31,151,31,20,31,28,31,212,31,160,31,160,30,160,29,224,31,224,30,188,31,54,31,54,30,54,29,206,31,165,31,88,31,88,30,215,31,215,30,201,31,201,30,81,31,92,31,138,31,221,31,57,31,2,31,119,31,119,30,82,31,18,31,114,31,210,31,210,30,169,31,169,30,121,31,196,31,103,31,96,31,138,31,35,31,57,31,52,31,112,31,4,31,128,31,176,31,135,31,151,31,151,30,255,31,50,31,125,31,125,30,3,31,183,31,110,31,199,31,210,31,210,30,210,29,210,28,210,27,20,31,20,30,173,31,173,30,173,29,216,31,216,30,250,31,31,31,149,31,149,30,151,31,139,31,175,31,12,31,86,31,219,31,219,30,219,29,79,31,79,30,79,29,194,31,219,31,231,31,88,31,186,31,125,31,22,31,22,30,136,31,86,31,86,30,95,31,95,30,95,29,95,28,203,31,255,31,248,31,71,31,49,31,49,30,70,31,82,31,82,30,115,31,115,31,191,31,58,31,58,30,81,31,88,31,88,30,34,31,34,30,133,31,231,31,178,31,178,30,178,29,178,28,91,31,161,31,220,31,220,30,106,31,70,31,55,31,189,31,155,31,213,31,136,31,43,31,43,30,247,31,168,31,206,31,66,31,81,31,183,31,92,31,231,31,203,31,222,31,126,31,254,31,39,31,164,31,32,31,145,31,159,31,129,31,133,31,133,30,191,31,91,31,58,31,89,31,254,31,204,31,20,31,20,30,20,29,20,28,145,31,145,30,145,29,254,31,134,31,2,31,138,31,204,31,86,31,246,31,9,31,103,31,83,31,83,30,210,31,20,31,231,31,167,31,76,31,78,31,64,31,64,30,33,31,150,31,59,31,126,31,125,31,98,31,193,31,21,31,221,31,63,31,213,31,93,31,18,31,18,30,180,31,92,31,33,31,34,31,34,30,202,31,161,31,249,31,249,30,70,31,54,31,28,31,62,31,87,31,87,30,196,31,125,31,134,31,239,31,14,31,247,31,57,31,51,31,165,31,99,31,76,31,76,30,49,31,49,30,117,31,223,31,77,31,250,31,250,30,150,31,173,31,254,31,254,30,89,31,161,31,202,31,236,31,236,30,190,31,99,31,103,31,89,31,117,31,65,31,206,31,79,31,172,31,226,31,200,31,200,30,39,31,39,30,117,31,126,31,152,31,58,31,34,31,186,31,115,31,184,31,22,31,114,31,161,31,161,30,101,31,17,31,17,30,165,31,171,31,193,31,193,30,254,31,254,30,187,31,25,31,222,31,88,31,1,31,127,31,195,31,93,31,93,30,231,31,206,31,184,31,106,31,98,31,55,31,55,30,232,31,232,30,102,31,102,30,237,31,35,31,35,30,35,29,83,31,116,31,129,31,90,31,179,31,8,31,8,30,8,29,124,31,149,31,157,31,35,31,238,31,74,31,234,31,38,31,144,31,14,31,192,31,192,30,192,29,50,31,49,31,14,31,14,30,147,31,147,30,7,31,76,31,235,31,235,31,215,31,215,30,170,31,217,31,177,31,177,30,252,31,61,31,29,31,80,31,86,31,86,30,62,31,62,30,37,31,171,31,168,31,243,31,40,31,119,31,82,31,80,31,48,31,236,31,129,31,129,30,86,31,176,31,128,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
