-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_53 is
end project_tb_53;

architecture project_tb_arch_53 of project_tb_53 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 991;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,147,0,178,0,0,0,144,0,157,0,237,0,38,0,241,0,117,0,48,0,232,0,138,0,19,0,0,0,97,0,64,0,0,0,14,0,131,0,164,0,17,0,90,0,195,0,198,0,221,0,0,0,14,0,72,0,216,0,96,0,0,0,140,0,0,0,182,0,25,0,0,0,5,0,145,0,223,0,175,0,135,0,250,0,219,0,173,0,134,0,233,0,80,0,229,0,0,0,86,0,26,0,201,0,215,0,240,0,74,0,0,0,0,0,0,0,230,0,19,0,0,0,129,0,61,0,128,0,101,0,0,0,12,0,107,0,54,0,245,0,100,0,117,0,225,0,127,0,128,0,0,0,21,0,0,0,143,0,0,0,139,0,171,0,0,0,146,0,162,0,0,0,0,0,212,0,83,0,0,0,0,0,164,0,165,0,154,0,36,0,106,0,120,0,0,0,245,0,18,0,62,0,213,0,122,0,102,0,0,0,0,0,121,0,0,0,184,0,233,0,98,0,77,0,0,0,66,0,117,0,82,0,203,0,125,0,104,0,41,0,0,0,240,0,23,0,13,0,47,0,192,0,0,0,83,0,49,0,0,0,123,0,0,0,9,0,111,0,63,0,28,0,0,0,0,0,96,0,0,0,110,0,0,0,110,0,0,0,218,0,58,0,148,0,27,0,198,0,0,0,127,0,173,0,166,0,233,0,9,0,206,0,227,0,107,0,164,0,73,0,196,0,0,0,0,0,64,0,226,0,169,0,108,0,7,0,32,0,63,0,174,0,108,0,183,0,14,0,114,0,0,0,0,0,48,0,163,0,128,0,174,0,27,0,221,0,59,0,104,0,152,0,47,0,236,0,15,0,36,0,175,0,141,0,140,0,37,0,0,0,109,0,49,0,0,0,0,0,145,0,200,0,252,0,252,0,78,0,137,0,253,0,179,0,162,0,252,0,135,0,43,0,126,0,149,0,0,0,63,0,77,0,0,0,231,0,38,0,197,0,68,0,207,0,0,0,153,0,88,0,123,0,162,0,0,0,0,0,126,0,0,0,0,0,82,0,170,0,0,0,0,0,1,0,45,0,100,0,245,0,113,0,83,0,199,0,16,0,67,0,124,0,164,0,20,0,124,0,79,0,118,0,23,0,82,0,192,0,0,0,161,0,11,0,14,0,97,0,203,0,110,0,44,0,30,0,0,0,74,0,133,0,28,0,0,0,254,0,0,0,142,0,0,0,133,0,14,0,200,0,208,0,0,0,207,0,0,0,162,0,143,0,0,0,126,0,0,0,59,0,235,0,83,0,0,0,55,0,31,0,67,0,242,0,149,0,166,0,252,0,149,0,218,0,144,0,0,0,232,0,195,0,14,0,135,0,13,0,0,0,31,0,0,0,204,0,17,0,241,0,0,0,141,0,31,0,3,0,227,0,0,0,111,0,32,0,247,0,103,0,100,0,158,0,0,0,0,0,77,0,21,0,61,0,68,0,58,0,0,0,249,0,216,0,45,0,112,0,55,0,0,0,18,0,134,0,0,0,44,0,18,0,41,0,172,0,141,0,137,0,173,0,241,0,161,0,187,0,0,0,103,0,0,0,252,0,186,0,218,0,185,0,199,0,241,0,33,0,97,0,31,0,122,0,122,0,140,0,40,0,22,0,226,0,250,0,100,0,50,0,115,0,91,0,94,0,145,0,137,0,60,0,234,0,255,0,0,0,221,0,46,0,39,0,203,0,225,0,0,0,86,0,223,0,41,0,228,0,13,0,0,0,190,0,45,0,53,0,179,0,197,0,161,0,0,0,162,0,124,0,174,0,139,0,168,0,0,0,241,0,143,0,200,0,0,0,54,0,243,0,195,0,243,0,128,0,203,0,25,0,53,0,203,0,0,0,29,0,74,0,150,0,200,0,57,0,52,0,0,0,0,0,210,0,98,0,232,0,132,0,159,0,112,0,117,0,161,0,83,0,30,0,33,0,249,0,0,0,181,0,214,0,73,0,0,0,67,0,41,0,253,0,0,0,150,0,23,0,190,0,129,0,0,0,43,0,18,0,51,0,11,0,1,0,209,0,55,0,0,0,153,0,125,0,17,0,24,0,149,0,254,0,240,0,253,0,144,0,175,0,0,0,176,0,0,0,0,0,245,0,7,0,0,0,243,0,30,0,53,0,127,0,91,0,23,0,24,0,173,0,8,0,131,0,134,0,0,0,72,0,238,0,0,0,221,0,36,0,187,0,156,0,20,0,46,0,242,0,25,0,31,0,216,0,149,0,56,0,161,0,38,0,201,0,64,0,0,0,14,0,0,0,156,0,133,0,171,0,85,0,101,0,6,0,57,0,118,0,23,0,0,0,46,0,0,0,206,0,0,0,172,0,129,0,50,0,200,0,0,0,0,0,0,0,62,0,121,0,48,0,0,0,188,0,0,0,141,0,189,0,114,0,237,0,101,0,29,0,0,0,99,0,85,0,244,0,26,0,0,0,172,0,107,0,0,0,112,0,173,0,0,0,169,0,0,0,92,0,252,0,0,0,12,0,68,0,187,0,0,0,17,0,0,0,54,0,43,0,86,0,0,0,4,0,116,0,141,0,0,0,92,0,5,0,230,0,201,0,224,0,227,0,0,0,0,0,95,0,246,0,144,0,61,0,117,0,175,0,85,0,226,0,176,0,220,0,175,0,255,0,214,0,120,0,167,0,205,0,123,0,128,0,0,0,39,0,188,0,124,0,105,0,205,0,0,0,12,0,95,0,187,0,119,0,45,0,11,0,80,0,246,0,5,0,32,0,0,0,150,0,3,0,0,0,22,0,221,0,0,0,196,0,166,0,247,0,243,0,165,0,143,0,111,0,204,0,46,0,27,0,186,0,59,0,84,0,197,0,0,0,215,0,0,0,47,0,130,0,116,0,174,0,0,0,160,0,219,0,96,0,147,0,92,0,37,0,0,0,64,0,70,0,121,0,114,0,201,0,0,0,126,0,100,0,211,0,127,0,253,0,118,0,0,0,92,0,83,0,56,0,127,0,0,0,98,0,213,0,179,0,142,0,0,0,136,0,33,0,0,0,78,0,170,0,192,0,146,0,113,0,211,0,22,0,5,0,241,0,217,0,159,0,89,0,228,0,2,0,198,0,81,0,207,0,104,0,119,0,9,0,68,0,8,0,246,0,249,0,134,0,224,0,73,0,11,0,109,0,0,0,0,0,194,0,30,0,31,0,0,0,62,0,25,0,0,0,0,0,127,0,108,0,50,0,237,0,182,0,226,0,15,0,227,0,254,0,30,0,216,0,3,0,0,0,44,0,254,0,0,0,160,0,103,0,105,0,97,0,0,0,187,0,10,0,231,0,0,0,62,0,0,0,198,0,0,0,228,0,124,0,167,0,181,0,184,0,145,0,241,0,76,0,126,0,0,0,201,0,254,0,62,0,181,0,107,0,0,0,162,0,0,0,249,0,225,0,178,0,53,0,0,0,197,0,70,0,239,0,220,0,47,0,0,0,69,0,94,0,119,0,237,0,131,0,182,0,59,0,42,0,246,0,17,0,154,0,34,0,0,0,186,0,85,0,97,0,49,0,190,0,20,0,183,0,125,0,239,0,246,0,61,0,23,0,29,0,197,0,225,0,0,0,0,0,165,0,80,0,210,0,0,0,120,0,239,0,56,0,0,0,195,0,5,0,37,0,202,0,174,0,0,0,188,0,52,0,105,0,0,0,62,0,39,0,221,0,0,0,74,0,252,0,0,0,133,0,33,0,251,0,145,0,212,0,121,0,0,0,127,0,33,0,168,0,21,0,156,0,208,0,216,0,0,0,222,0,19,0,156,0,0,0,186,0,6,0,90,0,69,0,201,0,199,0,34,0,0,0,124,0,98,0,0,0,240,0,51,0,158,0,0,0,0,0,15,0,174,0,242,0,151,0,208,0,148,0,115,0,0,0,42,0,249,0,25,0,114,0,0,0,26,0,118,0,35,0,0,0,222,0,209,0,130,0,70,0,96,0,0,0,28,0,65,0,130,0,0,0,252,0,229,0,170,0,83,0,55,0,96,0,199,0,115,0,61,0,100,0,161,0,164,0,110,0,51,0,74,0,42,0,0,0,174,0,0,0,78,0,0,0,0,0,0,0,245,0,11,0,59,0,0,0,206,0,0,0,0,0,224,0,156,0,185,0,178,0,143,0,81,0,231,0,190,0,229,0,102,0,225,0,199,0,135,0,96,0,6,0,36,0,148,0,4,0,40,0,134,0,34,0,0,0,4,0,254,0,102,0,117,0,92,0,11,0,13,0,29,0,122,0,91,0,14,0,139,0,158,0,0,0,60,0,163,0,0,0,154,0,90,0,0,0,94,0,0,0,0,0,221,0,124,0,135,0,0,0,44,0,0,0,184,0,132,0,66,0,243,0,25,0,170,0,18,0,120,0,0,0,131,0,254,0,26,0,98,0,98,0,179,0);
signal scenario_full  : scenario_type := (16,31,147,31,178,31,178,30,144,31,157,31,237,31,38,31,241,31,117,31,48,31,232,31,138,31,19,31,19,30,97,31,64,31,64,30,14,31,131,31,164,31,17,31,90,31,195,31,198,31,221,31,221,30,14,31,72,31,216,31,96,31,96,30,140,31,140,30,182,31,25,31,25,30,5,31,145,31,223,31,175,31,135,31,250,31,219,31,173,31,134,31,233,31,80,31,229,31,229,30,86,31,26,31,201,31,215,31,240,31,74,31,74,30,74,29,74,28,230,31,19,31,19,30,129,31,61,31,128,31,101,31,101,30,12,31,107,31,54,31,245,31,100,31,117,31,225,31,127,31,128,31,128,30,21,31,21,30,143,31,143,30,139,31,171,31,171,30,146,31,162,31,162,30,162,29,212,31,83,31,83,30,83,29,164,31,165,31,154,31,36,31,106,31,120,31,120,30,245,31,18,31,62,31,213,31,122,31,102,31,102,30,102,29,121,31,121,30,184,31,233,31,98,31,77,31,77,30,66,31,117,31,82,31,203,31,125,31,104,31,41,31,41,30,240,31,23,31,13,31,47,31,192,31,192,30,83,31,49,31,49,30,123,31,123,30,9,31,111,31,63,31,28,31,28,30,28,29,96,31,96,30,110,31,110,30,110,31,110,30,218,31,58,31,148,31,27,31,198,31,198,30,127,31,173,31,166,31,233,31,9,31,206,31,227,31,107,31,164,31,73,31,196,31,196,30,196,29,64,31,226,31,169,31,108,31,7,31,32,31,63,31,174,31,108,31,183,31,14,31,114,31,114,30,114,29,48,31,163,31,128,31,174,31,27,31,221,31,59,31,104,31,152,31,47,31,236,31,15,31,36,31,175,31,141,31,140,31,37,31,37,30,109,31,49,31,49,30,49,29,145,31,200,31,252,31,252,31,78,31,137,31,253,31,179,31,162,31,252,31,135,31,43,31,126,31,149,31,149,30,63,31,77,31,77,30,231,31,38,31,197,31,68,31,207,31,207,30,153,31,88,31,123,31,162,31,162,30,162,29,126,31,126,30,126,29,82,31,170,31,170,30,170,29,1,31,45,31,100,31,245,31,113,31,83,31,199,31,16,31,67,31,124,31,164,31,20,31,124,31,79,31,118,31,23,31,82,31,192,31,192,30,161,31,11,31,14,31,97,31,203,31,110,31,44,31,30,31,30,30,74,31,133,31,28,31,28,30,254,31,254,30,142,31,142,30,133,31,14,31,200,31,208,31,208,30,207,31,207,30,162,31,143,31,143,30,126,31,126,30,59,31,235,31,83,31,83,30,55,31,31,31,67,31,242,31,149,31,166,31,252,31,149,31,218,31,144,31,144,30,232,31,195,31,14,31,135,31,13,31,13,30,31,31,31,30,204,31,17,31,241,31,241,30,141,31,31,31,3,31,227,31,227,30,111,31,32,31,247,31,103,31,100,31,158,31,158,30,158,29,77,31,21,31,61,31,68,31,58,31,58,30,249,31,216,31,45,31,112,31,55,31,55,30,18,31,134,31,134,30,44,31,18,31,41,31,172,31,141,31,137,31,173,31,241,31,161,31,187,31,187,30,103,31,103,30,252,31,186,31,218,31,185,31,199,31,241,31,33,31,97,31,31,31,122,31,122,31,140,31,40,31,22,31,226,31,250,31,100,31,50,31,115,31,91,31,94,31,145,31,137,31,60,31,234,31,255,31,255,30,221,31,46,31,39,31,203,31,225,31,225,30,86,31,223,31,41,31,228,31,13,31,13,30,190,31,45,31,53,31,179,31,197,31,161,31,161,30,162,31,124,31,174,31,139,31,168,31,168,30,241,31,143,31,200,31,200,30,54,31,243,31,195,31,243,31,128,31,203,31,25,31,53,31,203,31,203,30,29,31,74,31,150,31,200,31,57,31,52,31,52,30,52,29,210,31,98,31,232,31,132,31,159,31,112,31,117,31,161,31,83,31,30,31,33,31,249,31,249,30,181,31,214,31,73,31,73,30,67,31,41,31,253,31,253,30,150,31,23,31,190,31,129,31,129,30,43,31,18,31,51,31,11,31,1,31,209,31,55,31,55,30,153,31,125,31,17,31,24,31,149,31,254,31,240,31,253,31,144,31,175,31,175,30,176,31,176,30,176,29,245,31,7,31,7,30,243,31,30,31,53,31,127,31,91,31,23,31,24,31,173,31,8,31,131,31,134,31,134,30,72,31,238,31,238,30,221,31,36,31,187,31,156,31,20,31,46,31,242,31,25,31,31,31,216,31,149,31,56,31,161,31,38,31,201,31,64,31,64,30,14,31,14,30,156,31,133,31,171,31,85,31,101,31,6,31,57,31,118,31,23,31,23,30,46,31,46,30,206,31,206,30,172,31,129,31,50,31,200,31,200,30,200,29,200,28,62,31,121,31,48,31,48,30,188,31,188,30,141,31,189,31,114,31,237,31,101,31,29,31,29,30,99,31,85,31,244,31,26,31,26,30,172,31,107,31,107,30,112,31,173,31,173,30,169,31,169,30,92,31,252,31,252,30,12,31,68,31,187,31,187,30,17,31,17,30,54,31,43,31,86,31,86,30,4,31,116,31,141,31,141,30,92,31,5,31,230,31,201,31,224,31,227,31,227,30,227,29,95,31,246,31,144,31,61,31,117,31,175,31,85,31,226,31,176,31,220,31,175,31,255,31,214,31,120,31,167,31,205,31,123,31,128,31,128,30,39,31,188,31,124,31,105,31,205,31,205,30,12,31,95,31,187,31,119,31,45,31,11,31,80,31,246,31,5,31,32,31,32,30,150,31,3,31,3,30,22,31,221,31,221,30,196,31,166,31,247,31,243,31,165,31,143,31,111,31,204,31,46,31,27,31,186,31,59,31,84,31,197,31,197,30,215,31,215,30,47,31,130,31,116,31,174,31,174,30,160,31,219,31,96,31,147,31,92,31,37,31,37,30,64,31,70,31,121,31,114,31,201,31,201,30,126,31,100,31,211,31,127,31,253,31,118,31,118,30,92,31,83,31,56,31,127,31,127,30,98,31,213,31,179,31,142,31,142,30,136,31,33,31,33,30,78,31,170,31,192,31,146,31,113,31,211,31,22,31,5,31,241,31,217,31,159,31,89,31,228,31,2,31,198,31,81,31,207,31,104,31,119,31,9,31,68,31,8,31,246,31,249,31,134,31,224,31,73,31,11,31,109,31,109,30,109,29,194,31,30,31,31,31,31,30,62,31,25,31,25,30,25,29,127,31,108,31,50,31,237,31,182,31,226,31,15,31,227,31,254,31,30,31,216,31,3,31,3,30,44,31,254,31,254,30,160,31,103,31,105,31,97,31,97,30,187,31,10,31,231,31,231,30,62,31,62,30,198,31,198,30,228,31,124,31,167,31,181,31,184,31,145,31,241,31,76,31,126,31,126,30,201,31,254,31,62,31,181,31,107,31,107,30,162,31,162,30,249,31,225,31,178,31,53,31,53,30,197,31,70,31,239,31,220,31,47,31,47,30,69,31,94,31,119,31,237,31,131,31,182,31,59,31,42,31,246,31,17,31,154,31,34,31,34,30,186,31,85,31,97,31,49,31,190,31,20,31,183,31,125,31,239,31,246,31,61,31,23,31,29,31,197,31,225,31,225,30,225,29,165,31,80,31,210,31,210,30,120,31,239,31,56,31,56,30,195,31,5,31,37,31,202,31,174,31,174,30,188,31,52,31,105,31,105,30,62,31,39,31,221,31,221,30,74,31,252,31,252,30,133,31,33,31,251,31,145,31,212,31,121,31,121,30,127,31,33,31,168,31,21,31,156,31,208,31,216,31,216,30,222,31,19,31,156,31,156,30,186,31,6,31,90,31,69,31,201,31,199,31,34,31,34,30,124,31,98,31,98,30,240,31,51,31,158,31,158,30,158,29,15,31,174,31,242,31,151,31,208,31,148,31,115,31,115,30,42,31,249,31,25,31,114,31,114,30,26,31,118,31,35,31,35,30,222,31,209,31,130,31,70,31,96,31,96,30,28,31,65,31,130,31,130,30,252,31,229,31,170,31,83,31,55,31,96,31,199,31,115,31,61,31,100,31,161,31,164,31,110,31,51,31,74,31,42,31,42,30,174,31,174,30,78,31,78,30,78,29,78,28,245,31,11,31,59,31,59,30,206,31,206,30,206,29,224,31,156,31,185,31,178,31,143,31,81,31,231,31,190,31,229,31,102,31,225,31,199,31,135,31,96,31,6,31,36,31,148,31,4,31,40,31,134,31,34,31,34,30,4,31,254,31,102,31,117,31,92,31,11,31,13,31,29,31,122,31,91,31,14,31,139,31,158,31,158,30,60,31,163,31,163,30,154,31,90,31,90,30,94,31,94,30,94,29,221,31,124,31,135,31,135,30,44,31,44,30,184,31,132,31,66,31,243,31,25,31,170,31,18,31,120,31,120,30,131,31,254,31,26,31,98,31,98,31,179,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
