-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 547;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,168,0,144,0,64,0,204,0,0,0,161,0,151,0,226,0,16,0,0,0,238,0,0,0,66,0,51,0,172,0,81,0,81,0,0,0,0,0,198,0,0,0,180,0,91,0,190,0,0,0,82,0,0,0,0,0,0,0,14,0,1,0,235,0,22,0,0,0,30,0,247,0,142,0,210,0,77,0,92,0,205,0,193,0,117,0,55,0,163,0,49,0,65,0,124,0,189,0,84,0,180,0,0,0,26,0,144,0,129,0,15,0,0,0,208,0,159,0,60,0,14,0,160,0,0,0,252,0,147,0,0,0,43,0,0,0,218,0,87,0,0,0,70,0,246,0,130,0,17,0,116,0,78,0,225,0,0,0,230,0,5,0,119,0,177,0,86,0,54,0,0,0,214,0,238,0,224,0,150,0,138,0,196,0,31,0,35,0,242,0,0,0,212,0,114,0,204,0,0,0,150,0,133,0,236,0,0,0,47,0,78,0,122,0,64,0,233,0,180,0,0,0,0,0,0,0,12,0,108,0,0,0,0,0,0,0,88,0,213,0,0,0,98,0,126,0,0,0,199,0,0,0,120,0,0,0,174,0,0,0,25,0,98,0,11,0,1,0,87,0,74,0,242,0,226,0,152,0,254,0,0,0,103,0,0,0,0,0,100,0,101,0,0,0,252,0,70,0,208,0,87,0,233,0,0,0,57,0,0,0,7,0,0,0,63,0,26,0,100,0,96,0,32,0,0,0,0,0,171,0,0,0,61,0,169,0,0,0,131,0,210,0,244,0,99,0,140,0,23,0,0,0,0,0,115,0,57,0,176,0,0,0,12,0,100,0,0,0,123,0,9,0,190,0,247,0,186,0,215,0,229,0,111,0,58,0,97,0,0,0,157,0,101,0,246,0,14,0,1,0,11,0,85,0,47,0,0,0,0,0,0,0,207,0,0,0,251,0,50,0,237,0,41,0,182,0,0,0,0,0,218,0,210,0,42,0,0,0,246,0,0,0,0,0,166,0,252,0,222,0,204,0,0,0,13,0,42,0,183,0,253,0,231,0,232,0,58,0,68,0,252,0,0,0,90,0,209,0,229,0,0,0,219,0,154,0,193,0,73,0,92,0,0,0,0,0,230,0,0,0,24,0,115,0,105,0,58,0,93,0,230,0,240,0,143,0,203,0,245,0,36,0,107,0,130,0,198,0,124,0,101,0,150,0,66,0,84,0,134,0,0,0,255,0,13,0,245,0,38,0,176,0,162,0,190,0,18,0,171,0,60,0,0,0,184,0,185,0,231,0,139,0,120,0,226,0,121,0,221,0,156,0,0,0,195,0,11,0,50,0,20,0,84,0,243,0,126,0,0,0,7,0,29,0,162,0,5,0,84,0,0,0,113,0,38,0,26,0,16,0,178,0,0,0,198,0,223,0,0,0,174,0,31,0,50,0,254,0,231,0,129,0,0,0,236,0,0,0,175,0,82,0,0,0,0,0,10,0,0,0,235,0,123,0,0,0,135,0,160,0,110,0,233,0,0,0,104,0,101,0,112,0,0,0,0,0,78,0,0,0,0,0,187,0,162,0,154,0,172,0,96,0,0,0,51,0,173,0,0,0,0,0,0,0,223,0,133,0,28,0,141,0,0,0,143,0,15,0,26,0,163,0,83,0,59,0,52,0,170,0,89,0,214,0,92,0,78,0,0,0,181,0,245,0,0,0,0,0,108,0,225,0,39,0,54,0,44,0,167,0,214,0,23,0,152,0,135,0,92,0,0,0,179,0,82,0,57,0,187,0,168,0,166,0,41,0,0,0,32,0,201,0,188,0,210,0,138,0,240,0,233,0,105,0,0,0,0,0,14,0,0,0,195,0,65,0,204,0,0,0,202,0,123,0,0,0,0,0,163,0,138,0,0,0,50,0,90,0,56,0,88,0,138,0,84,0,230,0,170,0,97,0,227,0,100,0,106,0,163,0,17,0,0,0,0,0,123,0,0,0,144,0,25,0,0,0,0,0,85,0,0,0,0,0,130,0,177,0,206,0,93,0,43,0,46,0,0,0,33,0,0,0,0,0,232,0,0,0,72,0,23,0,152,0,83,0,97,0,0,0,147,0,16,0,180,0,195,0,14,0,160,0,240,0,99,0,25,0,79,0,0,0,17,0,0,0,115,0,0,0,164,0,83,0,190,0,227,0,0,0,228,0,212,0,149,0,185,0,187,0,29,0,155,0,255,0,243,0,199,0,180,0,211,0,240,0,139,0,0,0,0,0,47,0,42,0,0,0,138,0,46,0,63,0,59,0,6,0,160,0,181,0,168,0,163,0,111,0,15,0,17,0,183,0,68,0,0,0,193,0,0,0,246,0,150,0,14,0,22,0,206,0,0,0,154,0,95,0,201,0,0,0,112,0,45,0,174,0,48,0,240,0,188,0,0,0,131,0,0,0,96,0,54,0,210,0,165,0,0,0,0,0);
signal scenario_full  : scenario_type := (214,31,168,31,144,31,64,31,204,31,204,30,161,31,151,31,226,31,16,31,16,30,238,31,238,30,66,31,51,31,172,31,81,31,81,31,81,30,81,29,198,31,198,30,180,31,91,31,190,31,190,30,82,31,82,30,82,29,82,28,14,31,1,31,235,31,22,31,22,30,30,31,247,31,142,31,210,31,77,31,92,31,205,31,193,31,117,31,55,31,163,31,49,31,65,31,124,31,189,31,84,31,180,31,180,30,26,31,144,31,129,31,15,31,15,30,208,31,159,31,60,31,14,31,160,31,160,30,252,31,147,31,147,30,43,31,43,30,218,31,87,31,87,30,70,31,246,31,130,31,17,31,116,31,78,31,225,31,225,30,230,31,5,31,119,31,177,31,86,31,54,31,54,30,214,31,238,31,224,31,150,31,138,31,196,31,31,31,35,31,242,31,242,30,212,31,114,31,204,31,204,30,150,31,133,31,236,31,236,30,47,31,78,31,122,31,64,31,233,31,180,31,180,30,180,29,180,28,12,31,108,31,108,30,108,29,108,28,88,31,213,31,213,30,98,31,126,31,126,30,199,31,199,30,120,31,120,30,174,31,174,30,25,31,98,31,11,31,1,31,87,31,74,31,242,31,226,31,152,31,254,31,254,30,103,31,103,30,103,29,100,31,101,31,101,30,252,31,70,31,208,31,87,31,233,31,233,30,57,31,57,30,7,31,7,30,63,31,26,31,100,31,96,31,32,31,32,30,32,29,171,31,171,30,61,31,169,31,169,30,131,31,210,31,244,31,99,31,140,31,23,31,23,30,23,29,115,31,57,31,176,31,176,30,12,31,100,31,100,30,123,31,9,31,190,31,247,31,186,31,215,31,229,31,111,31,58,31,97,31,97,30,157,31,101,31,246,31,14,31,1,31,11,31,85,31,47,31,47,30,47,29,47,28,207,31,207,30,251,31,50,31,237,31,41,31,182,31,182,30,182,29,218,31,210,31,42,31,42,30,246,31,246,30,246,29,166,31,252,31,222,31,204,31,204,30,13,31,42,31,183,31,253,31,231,31,232,31,58,31,68,31,252,31,252,30,90,31,209,31,229,31,229,30,219,31,154,31,193,31,73,31,92,31,92,30,92,29,230,31,230,30,24,31,115,31,105,31,58,31,93,31,230,31,240,31,143,31,203,31,245,31,36,31,107,31,130,31,198,31,124,31,101,31,150,31,66,31,84,31,134,31,134,30,255,31,13,31,245,31,38,31,176,31,162,31,190,31,18,31,171,31,60,31,60,30,184,31,185,31,231,31,139,31,120,31,226,31,121,31,221,31,156,31,156,30,195,31,11,31,50,31,20,31,84,31,243,31,126,31,126,30,7,31,29,31,162,31,5,31,84,31,84,30,113,31,38,31,26,31,16,31,178,31,178,30,198,31,223,31,223,30,174,31,31,31,50,31,254,31,231,31,129,31,129,30,236,31,236,30,175,31,82,31,82,30,82,29,10,31,10,30,235,31,123,31,123,30,135,31,160,31,110,31,233,31,233,30,104,31,101,31,112,31,112,30,112,29,78,31,78,30,78,29,187,31,162,31,154,31,172,31,96,31,96,30,51,31,173,31,173,30,173,29,173,28,223,31,133,31,28,31,141,31,141,30,143,31,15,31,26,31,163,31,83,31,59,31,52,31,170,31,89,31,214,31,92,31,78,31,78,30,181,31,245,31,245,30,245,29,108,31,225,31,39,31,54,31,44,31,167,31,214,31,23,31,152,31,135,31,92,31,92,30,179,31,82,31,57,31,187,31,168,31,166,31,41,31,41,30,32,31,201,31,188,31,210,31,138,31,240,31,233,31,105,31,105,30,105,29,14,31,14,30,195,31,65,31,204,31,204,30,202,31,123,31,123,30,123,29,163,31,138,31,138,30,50,31,90,31,56,31,88,31,138,31,84,31,230,31,170,31,97,31,227,31,100,31,106,31,163,31,17,31,17,30,17,29,123,31,123,30,144,31,25,31,25,30,25,29,85,31,85,30,85,29,130,31,177,31,206,31,93,31,43,31,46,31,46,30,33,31,33,30,33,29,232,31,232,30,72,31,23,31,152,31,83,31,97,31,97,30,147,31,16,31,180,31,195,31,14,31,160,31,240,31,99,31,25,31,79,31,79,30,17,31,17,30,115,31,115,30,164,31,83,31,190,31,227,31,227,30,228,31,212,31,149,31,185,31,187,31,29,31,155,31,255,31,243,31,199,31,180,31,211,31,240,31,139,31,139,30,139,29,47,31,42,31,42,30,138,31,46,31,63,31,59,31,6,31,160,31,181,31,168,31,163,31,111,31,15,31,17,31,183,31,68,31,68,30,193,31,193,30,246,31,150,31,14,31,22,31,206,31,206,30,154,31,95,31,201,31,201,30,112,31,45,31,174,31,48,31,240,31,188,31,188,30,131,31,131,30,96,31,54,31,210,31,165,31,165,30,165,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
