-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 680;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (47,0,47,0,193,0,201,0,195,0,220,0,27,0,141,0,96,0,0,0,230,0,218,0,14,0,243,0,244,0,153,0,21,0,0,0,79,0,0,0,110,0,194,0,34,0,0,0,165,0,244,0,161,0,234,0,44,0,165,0,82,0,43,0,0,0,229,0,49,0,51,0,116,0,240,0,148,0,90,0,99,0,112,0,64,0,0,0,157,0,67,0,223,0,183,0,255,0,26,0,116,0,107,0,222,0,0,0,132,0,125,0,8,0,127,0,23,0,0,0,138,0,210,0,0,0,50,0,112,0,123,0,0,0,86,0,174,0,247,0,194,0,175,0,253,0,154,0,29,0,189,0,118,0,0,0,209,0,0,0,244,0,0,0,11,0,19,0,73,0,53,0,164,0,57,0,86,0,3,0,20,0,171,0,0,0,135,0,88,0,0,0,69,0,245,0,64,0,154,0,222,0,70,0,34,0,252,0,137,0,247,0,56,0,0,0,74,0,77,0,0,0,198,0,0,0,0,0,35,0,236,0,223,0,182,0,162,0,64,0,241,0,142,0,192,0,225,0,79,0,218,0,99,0,0,0,12,0,193,0,77,0,0,0,0,0,159,0,226,0,22,0,63,0,40,0,133,0,0,0,69,0,0,0,69,0,195,0,233,0,74,0,0,0,196,0,91,0,16,0,73,0,124,0,249,0,108,0,78,0,157,0,0,0,26,0,144,0,184,0,0,0,199,0,0,0,194,0,180,0,0,0,40,0,2,0,43,0,0,0,70,0,180,0,0,0,48,0,232,0,16,0,211,0,0,0,91,0,57,0,102,0,0,0,142,0,0,0,115,0,70,0,200,0,148,0,246,0,88,0,28,0,31,0,66,0,163,0,0,0,2,0,72,0,57,0,236,0,181,0,0,0,185,0,19,0,226,0,224,0,242,0,236,0,107,0,180,0,122,0,240,0,128,0,66,0,112,0,238,0,35,0,126,0,152,0,9,0,51,0,81,0,174,0,98,0,237,0,247,0,0,0,42,0,77,0,121,0,101,0,12,0,103,0,121,0,39,0,147,0,106,0,146,0,0,0,128,0,0,0,15,0,0,0,208,0,245,0,87,0,13,0,241,0,9,0,179,0,171,0,13,0,136,0,0,0,255,0,93,0,165,0,198,0,106,0,134,0,51,0,88,0,0,0,162,0,0,0,181,0,74,0,215,0,28,0,195,0,113,0,39,0,194,0,144,0,162,0,0,0,130,0,0,0,113,0,228,0,192,0,171,0,0,0,191,0,0,0,153,0,97,0,125,0,73,0,245,0,0,0,171,0,0,0,193,0,139,0,194,0,115,0,0,0,0,0,183,0,214,0,82,0,179,0,81,0,105,0,0,0,0,0,0,0,0,0,247,0,255,0,60,0,45,0,206,0,207,0,81,0,59,0,250,0,0,0,0,0,185,0,0,0,249,0,0,0,101,0,0,0,197,0,161,0,0,0,38,0,157,0,201,0,0,0,158,0,98,0,128,0,53,0,27,0,131,0,241,0,0,0,134,0,74,0,193,0,83,0,217,0,0,0,14,0,196,0,197,0,168,0,0,0,64,0,135,0,141,0,56,0,43,0,93,0,19,0,8,0,178,0,122,0,210,0,134,0,15,0,201,0,0,0,42,0,49,0,0,0,122,0,184,0,89,0,46,0,170,0,130,0,0,0,251,0,181,0,59,0,233,0,84,0,255,0,201,0,72,0,43,0,248,0,229,0,100,0,156,0,242,0,150,0,255,0,80,0,0,0,254,0,144,0,6,0,179,0,228,0,154,0,223,0,0,0,224,0,175,0,101,0,0,0,197,0,87,0,209,0,16,0,83,0,183,0,73,0,218,0,0,0,164,0,214,0,0,0,128,0,0,0,228,0,5,0,65,0,129,0,60,0,85,0,0,0,199,0,213,0,212,0,117,0,0,0,157,0,242,0,0,0,115,0,83,0,16,0,145,0,147,0,0,0,150,0,169,0,143,0,204,0,128,0,209,0,9,0,48,0,4,0,0,0,1,0,109,0,116,0,0,0,6,0,0,0,0,0,204,0,47,0,0,0,192,0,0,0,39,0,60,0,0,0,161,0,223,0,43,0,159,0,0,0,240,0,246,0,238,0,176,0,0,0,167,0,255,0,63,0,14,0,215,0,0,0,91,0,178,0,16,0,0,0,118,0,21,0,144,0,0,0,0,0,66,0,0,0,0,0,221,0,107,0,5,0,187,0,61,0,83,0,0,0,76,0,0,0,183,0,139,0,232,0,10,0,90,0,0,0,72,0,0,0,195,0,31,0,108,0,55,0,198,0,84,0,54,0,39,0,0,0,33,0,172,0,125,0,136,0,173,0,110,0,19,0,0,0,38,0,0,0,122,0,41,0,0,0,106,0,202,0,207,0,79,0,241,0,0,0,0,0,0,0,119,0,245,0,170,0,188,0,131,0,0,0,67,0,1,0,6,0,75,0,127,0,211,0,155,0,0,0,134,0,7,0,66,0,212,0,45,0,212,0,41,0,26,0,89,0,41,0,0,0,149,0,6,0,0,0,112,0,184,0,127,0,29,0,0,0,137,0,70,0,176,0,107,0,170,0,73,0,56,0,119,0,0,0,245,0,0,0,0,0,252,0,43,0,209,0,22,0,69,0,61,0,191,0,158,0,0,0,88,0,90,0,17,0,252,0,252,0,170,0,108,0,42,0,56,0,0,0,8,0,0,0,96,0,247,0,40,0,0,0,0,0,6,0,139,0,35,0,241,0,121,0,0,0,163,0,228,0,6,0,0,0,148,0,160,0,125,0,0,0,66,0,42,0,171,0,119,0,79,0,0,0,235,0,32,0,0,0,228,0,139,0,219,0,121,0,174,0,126,0,50,0,163,0,228,0,0,0,198,0,131,0,0,0,173,0,0,0,234,0,247,0,0,0,49,0,52,0,174,0,182,0,0,0,25,0,190,0,193,0,0,0,37,0,133,0,0,0,132,0,142,0,110,0,19,0,248,0,184,0,43,0,201,0,245,0,171,0,36,0,16,0,0,0,71,0,44,0);
signal scenario_full  : scenario_type := (47,31,47,31,193,31,201,31,195,31,220,31,27,31,141,31,96,31,96,30,230,31,218,31,14,31,243,31,244,31,153,31,21,31,21,30,79,31,79,30,110,31,194,31,34,31,34,30,165,31,244,31,161,31,234,31,44,31,165,31,82,31,43,31,43,30,229,31,49,31,51,31,116,31,240,31,148,31,90,31,99,31,112,31,64,31,64,30,157,31,67,31,223,31,183,31,255,31,26,31,116,31,107,31,222,31,222,30,132,31,125,31,8,31,127,31,23,31,23,30,138,31,210,31,210,30,50,31,112,31,123,31,123,30,86,31,174,31,247,31,194,31,175,31,253,31,154,31,29,31,189,31,118,31,118,30,209,31,209,30,244,31,244,30,11,31,19,31,73,31,53,31,164,31,57,31,86,31,3,31,20,31,171,31,171,30,135,31,88,31,88,30,69,31,245,31,64,31,154,31,222,31,70,31,34,31,252,31,137,31,247,31,56,31,56,30,74,31,77,31,77,30,198,31,198,30,198,29,35,31,236,31,223,31,182,31,162,31,64,31,241,31,142,31,192,31,225,31,79,31,218,31,99,31,99,30,12,31,193,31,77,31,77,30,77,29,159,31,226,31,22,31,63,31,40,31,133,31,133,30,69,31,69,30,69,31,195,31,233,31,74,31,74,30,196,31,91,31,16,31,73,31,124,31,249,31,108,31,78,31,157,31,157,30,26,31,144,31,184,31,184,30,199,31,199,30,194,31,180,31,180,30,40,31,2,31,43,31,43,30,70,31,180,31,180,30,48,31,232,31,16,31,211,31,211,30,91,31,57,31,102,31,102,30,142,31,142,30,115,31,70,31,200,31,148,31,246,31,88,31,28,31,31,31,66,31,163,31,163,30,2,31,72,31,57,31,236,31,181,31,181,30,185,31,19,31,226,31,224,31,242,31,236,31,107,31,180,31,122,31,240,31,128,31,66,31,112,31,238,31,35,31,126,31,152,31,9,31,51,31,81,31,174,31,98,31,237,31,247,31,247,30,42,31,77,31,121,31,101,31,12,31,103,31,121,31,39,31,147,31,106,31,146,31,146,30,128,31,128,30,15,31,15,30,208,31,245,31,87,31,13,31,241,31,9,31,179,31,171,31,13,31,136,31,136,30,255,31,93,31,165,31,198,31,106,31,134,31,51,31,88,31,88,30,162,31,162,30,181,31,74,31,215,31,28,31,195,31,113,31,39,31,194,31,144,31,162,31,162,30,130,31,130,30,113,31,228,31,192,31,171,31,171,30,191,31,191,30,153,31,97,31,125,31,73,31,245,31,245,30,171,31,171,30,193,31,139,31,194,31,115,31,115,30,115,29,183,31,214,31,82,31,179,31,81,31,105,31,105,30,105,29,105,28,105,27,247,31,255,31,60,31,45,31,206,31,207,31,81,31,59,31,250,31,250,30,250,29,185,31,185,30,249,31,249,30,101,31,101,30,197,31,161,31,161,30,38,31,157,31,201,31,201,30,158,31,98,31,128,31,53,31,27,31,131,31,241,31,241,30,134,31,74,31,193,31,83,31,217,31,217,30,14,31,196,31,197,31,168,31,168,30,64,31,135,31,141,31,56,31,43,31,93,31,19,31,8,31,178,31,122,31,210,31,134,31,15,31,201,31,201,30,42,31,49,31,49,30,122,31,184,31,89,31,46,31,170,31,130,31,130,30,251,31,181,31,59,31,233,31,84,31,255,31,201,31,72,31,43,31,248,31,229,31,100,31,156,31,242,31,150,31,255,31,80,31,80,30,254,31,144,31,6,31,179,31,228,31,154,31,223,31,223,30,224,31,175,31,101,31,101,30,197,31,87,31,209,31,16,31,83,31,183,31,73,31,218,31,218,30,164,31,214,31,214,30,128,31,128,30,228,31,5,31,65,31,129,31,60,31,85,31,85,30,199,31,213,31,212,31,117,31,117,30,157,31,242,31,242,30,115,31,83,31,16,31,145,31,147,31,147,30,150,31,169,31,143,31,204,31,128,31,209,31,9,31,48,31,4,31,4,30,1,31,109,31,116,31,116,30,6,31,6,30,6,29,204,31,47,31,47,30,192,31,192,30,39,31,60,31,60,30,161,31,223,31,43,31,159,31,159,30,240,31,246,31,238,31,176,31,176,30,167,31,255,31,63,31,14,31,215,31,215,30,91,31,178,31,16,31,16,30,118,31,21,31,144,31,144,30,144,29,66,31,66,30,66,29,221,31,107,31,5,31,187,31,61,31,83,31,83,30,76,31,76,30,183,31,139,31,232,31,10,31,90,31,90,30,72,31,72,30,195,31,31,31,108,31,55,31,198,31,84,31,54,31,39,31,39,30,33,31,172,31,125,31,136,31,173,31,110,31,19,31,19,30,38,31,38,30,122,31,41,31,41,30,106,31,202,31,207,31,79,31,241,31,241,30,241,29,241,28,119,31,245,31,170,31,188,31,131,31,131,30,67,31,1,31,6,31,75,31,127,31,211,31,155,31,155,30,134,31,7,31,66,31,212,31,45,31,212,31,41,31,26,31,89,31,41,31,41,30,149,31,6,31,6,30,112,31,184,31,127,31,29,31,29,30,137,31,70,31,176,31,107,31,170,31,73,31,56,31,119,31,119,30,245,31,245,30,245,29,252,31,43,31,209,31,22,31,69,31,61,31,191,31,158,31,158,30,88,31,90,31,17,31,252,31,252,31,170,31,108,31,42,31,56,31,56,30,8,31,8,30,96,31,247,31,40,31,40,30,40,29,6,31,139,31,35,31,241,31,121,31,121,30,163,31,228,31,6,31,6,30,148,31,160,31,125,31,125,30,66,31,42,31,171,31,119,31,79,31,79,30,235,31,32,31,32,30,228,31,139,31,219,31,121,31,174,31,126,31,50,31,163,31,228,31,228,30,198,31,131,31,131,30,173,31,173,30,234,31,247,31,247,30,49,31,52,31,174,31,182,31,182,30,25,31,190,31,193,31,193,30,37,31,133,31,133,30,132,31,142,31,110,31,19,31,248,31,184,31,43,31,201,31,245,31,171,31,36,31,16,31,16,30,71,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
