-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_509 is
end project_tb_509;

architecture project_tb_arch_509 of project_tb_509 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 675;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (77,0,45,0,0,0,68,0,0,0,122,0,22,0,59,0,14,0,233,0,197,0,117,0,0,0,14,0,0,0,0,0,138,0,217,0,0,0,25,0,0,0,74,0,156,0,145,0,147,0,39,0,107,0,246,0,179,0,224,0,0,0,0,0,0,0,217,0,52,0,191,0,21,0,2,0,165,0,84,0,217,0,0,0,121,0,159,0,104,0,131,0,53,0,184,0,0,0,0,0,18,0,196,0,202,0,53,0,0,0,172,0,0,0,163,0,240,0,141,0,251,0,0,0,214,0,234,0,229,0,72,0,159,0,125,0,185,0,127,0,147,0,231,0,171,0,31,0,1,0,128,0,69,0,106,0,0,0,77,0,167,0,96,0,69,0,0,0,189,0,0,0,187,0,0,0,253,0,216,0,144,0,215,0,26,0,0,0,209,0,21,0,152,0,0,0,69,0,182,0,0,0,152,0,198,0,255,0,182,0,205,0,207,0,168,0,0,0,96,0,135,0,234,0,189,0,87,0,226,0,106,0,137,0,120,0,168,0,184,0,64,0,0,0,182,0,124,0,13,0,111,0,123,0,179,0,37,0,40,0,92,0,59,0,35,0,34,0,0,0,103,0,210,0,250,0,217,0,0,0,0,0,168,0,147,0,203,0,33,0,88,0,245,0,0,0,191,0,147,0,103,0,105,0,7,0,0,0,46,0,141,0,40,0,43,0,157,0,138,0,253,0,113,0,189,0,43,0,178,0,19,0,216,0,243,0,18,0,0,0,95,0,58,0,101,0,180,0,0,0,122,0,150,0,204,0,0,0,14,0,0,0,0,0,241,0,98,0,0,0,150,0,68,0,214,0,234,0,0,0,106,0,0,0,27,0,0,0,203,0,169,0,92,0,222,0,79,0,79,0,255,0,0,0,200,0,22,0,125,0,0,0,139,0,153,0,194,0,228,0,0,0,33,0,128,0,58,0,236,0,64,0,159,0,158,0,0,0,229,0,0,0,255,0,91,0,112,0,0,0,107,0,155,0,0,0,0,0,121,0,15,0,22,0,248,0,158,0,0,0,73,0,0,0,23,0,59,0,178,0,178,0,143,0,0,0,0,0,155,0,179,0,45,0,251,0,208,0,150,0,105,0,196,0,253,0,0,0,59,0,184,0,0,0,147,0,0,0,129,0,24,0,4,0,144,0,106,0,17,0,60,0,170,0,0,0,0,0,64,0,185,0,0,0,0,0,230,0,129,0,151,0,62,0,0,0,69,0,74,0,4,0,65,0,110,0,207,0,134,0,4,0,141,0,0,0,176,0,116,0,88,0,43,0,207,0,0,0,239,0,0,0,134,0,166,0,126,0,44,0,66,0,0,0,10,0,215,0,232,0,53,0,147,0,245,0,126,0,180,0,70,0,21,0,195,0,245,0,101,0,152,0,110,0,13,0,75,0,0,0,117,0,195,0,95,0,98,0,123,0,232,0,157,0,98,0,131,0,74,0,79,0,128,0,14,0,157,0,83,0,0,0,150,0,179,0,0,0,6,0,87,0,133,0,220,0,85,0,76,0,152,0,183,0,205,0,50,0,19,0,106,0,203,0,97,0,0,0,74,0,247,0,49,0,219,0,0,0,189,0,153,0,216,0,63,0,164,0,0,0,40,0,147,0,121,0,0,0,0,0,0,0,249,0,41,0,189,0,29,0,64,0,123,0,52,0,135,0,211,0,106,0,84,0,86,0,206,0,253,0,38,0,179,0,0,0,231,0,133,0,26,0,90,0,253,0,0,0,5,0,115,0,0,0,31,0,174,0,0,0,0,0,38,0,42,0,144,0,49,0,185,0,117,0,0,0,122,0,141,0,95,0,191,0,172,0,119,0,151,0,205,0,14,0,181,0,38,0,215,0,4,0,234,0,96,0,83,0,181,0,208,0,189,0,0,0,90,0,162,0,0,0,181,0,0,0,14,0,132,0,196,0,22,0,200,0,170,0,0,0,163,0,0,0,0,0,16,0,122,0,35,0,29,0,0,0,51,0,186,0,36,0,117,0,0,0,23,0,59,0,0,0,85,0,113,0,73,0,74,0,144,0,235,0,144,0,20,0,158,0,0,0,0,0,71,0,195,0,0,0,0,0,168,0,0,0,128,0,0,0,0,0,232,0,231,0,118,0,0,0,223,0,227,0,0,0,0,0,9,0,63,0,218,0,0,0,0,0,0,0,203,0,106,0,236,0,3,0,159,0,253,0,0,0,130,0,222,0,22,0,0,0,200,0,46,0,120,0,157,0,11,0,89,0,144,0,120,0,113,0,185,0,215,0,148,0,199,0,49,0,0,0,92,0,40,0,0,0,38,0,151,0,0,0,146,0,233,0,121,0,101,0,153,0,97,0,2,0,32,0,111,0,0,0,8,0,174,0,245,0,0,0,0,0,4,0,97,0,204,0,162,0,86,0,49,0,0,0,165,0,235,0,173,0,0,0,150,0,162,0,67,0,56,0,0,0,82,0,0,0,187,0,191,0,30,0,244,0,218,0,0,0,141,0,0,0,201,0,105,0,29,0,201,0,153,0,149,0,31,0,0,0,160,0,28,0,112,0,116,0,125,0,172,0,0,0,200,0,44,0,155,0,0,0,213,0,57,0,14,0,0,0,172,0,86,0,195,0,0,0,193,0,0,0,214,0,241,0,163,0,244,0,160,0,52,0,53,0,154,0,142,0,225,0,0,0,98,0,121,0,19,0,0,0,0,0,38,0,216,0,0,0,9,0,136,0,157,0,174,0,188,0,13,0,0,0,149,0,221,0,60,0,165,0,101,0,101,0,32,0,157,0,20,0,214,0,17,0,159,0,49,0,0,0,86,0,225,0,48,0,139,0,206,0,0,0,0,0,7,0,0,0,74,0,47,0,105,0,123,0,72,0,174,0,181,0,233,0,186,0,226,0,45,0,131,0,219,0,212,0,2,0,30,0,227,0,28,0,1,0,236,0,198,0,202,0,0,0,114,0,152,0,132,0,11,0,148,0,0,0,159,0,116,0,128,0,224,0,200,0);
signal scenario_full  : scenario_type := (77,31,45,31,45,30,68,31,68,30,122,31,22,31,59,31,14,31,233,31,197,31,117,31,117,30,14,31,14,30,14,29,138,31,217,31,217,30,25,31,25,30,74,31,156,31,145,31,147,31,39,31,107,31,246,31,179,31,224,31,224,30,224,29,224,28,217,31,52,31,191,31,21,31,2,31,165,31,84,31,217,31,217,30,121,31,159,31,104,31,131,31,53,31,184,31,184,30,184,29,18,31,196,31,202,31,53,31,53,30,172,31,172,30,163,31,240,31,141,31,251,31,251,30,214,31,234,31,229,31,72,31,159,31,125,31,185,31,127,31,147,31,231,31,171,31,31,31,1,31,128,31,69,31,106,31,106,30,77,31,167,31,96,31,69,31,69,30,189,31,189,30,187,31,187,30,253,31,216,31,144,31,215,31,26,31,26,30,209,31,21,31,152,31,152,30,69,31,182,31,182,30,152,31,198,31,255,31,182,31,205,31,207,31,168,31,168,30,96,31,135,31,234,31,189,31,87,31,226,31,106,31,137,31,120,31,168,31,184,31,64,31,64,30,182,31,124,31,13,31,111,31,123,31,179,31,37,31,40,31,92,31,59,31,35,31,34,31,34,30,103,31,210,31,250,31,217,31,217,30,217,29,168,31,147,31,203,31,33,31,88,31,245,31,245,30,191,31,147,31,103,31,105,31,7,31,7,30,46,31,141,31,40,31,43,31,157,31,138,31,253,31,113,31,189,31,43,31,178,31,19,31,216,31,243,31,18,31,18,30,95,31,58,31,101,31,180,31,180,30,122,31,150,31,204,31,204,30,14,31,14,30,14,29,241,31,98,31,98,30,150,31,68,31,214,31,234,31,234,30,106,31,106,30,27,31,27,30,203,31,169,31,92,31,222,31,79,31,79,31,255,31,255,30,200,31,22,31,125,31,125,30,139,31,153,31,194,31,228,31,228,30,33,31,128,31,58,31,236,31,64,31,159,31,158,31,158,30,229,31,229,30,255,31,91,31,112,31,112,30,107,31,155,31,155,30,155,29,121,31,15,31,22,31,248,31,158,31,158,30,73,31,73,30,23,31,59,31,178,31,178,31,143,31,143,30,143,29,155,31,179,31,45,31,251,31,208,31,150,31,105,31,196,31,253,31,253,30,59,31,184,31,184,30,147,31,147,30,129,31,24,31,4,31,144,31,106,31,17,31,60,31,170,31,170,30,170,29,64,31,185,31,185,30,185,29,230,31,129,31,151,31,62,31,62,30,69,31,74,31,4,31,65,31,110,31,207,31,134,31,4,31,141,31,141,30,176,31,116,31,88,31,43,31,207,31,207,30,239,31,239,30,134,31,166,31,126,31,44,31,66,31,66,30,10,31,215,31,232,31,53,31,147,31,245,31,126,31,180,31,70,31,21,31,195,31,245,31,101,31,152,31,110,31,13,31,75,31,75,30,117,31,195,31,95,31,98,31,123,31,232,31,157,31,98,31,131,31,74,31,79,31,128,31,14,31,157,31,83,31,83,30,150,31,179,31,179,30,6,31,87,31,133,31,220,31,85,31,76,31,152,31,183,31,205,31,50,31,19,31,106,31,203,31,97,31,97,30,74,31,247,31,49,31,219,31,219,30,189,31,153,31,216,31,63,31,164,31,164,30,40,31,147,31,121,31,121,30,121,29,121,28,249,31,41,31,189,31,29,31,64,31,123,31,52,31,135,31,211,31,106,31,84,31,86,31,206,31,253,31,38,31,179,31,179,30,231,31,133,31,26,31,90,31,253,31,253,30,5,31,115,31,115,30,31,31,174,31,174,30,174,29,38,31,42,31,144,31,49,31,185,31,117,31,117,30,122,31,141,31,95,31,191,31,172,31,119,31,151,31,205,31,14,31,181,31,38,31,215,31,4,31,234,31,96,31,83,31,181,31,208,31,189,31,189,30,90,31,162,31,162,30,181,31,181,30,14,31,132,31,196,31,22,31,200,31,170,31,170,30,163,31,163,30,163,29,16,31,122,31,35,31,29,31,29,30,51,31,186,31,36,31,117,31,117,30,23,31,59,31,59,30,85,31,113,31,73,31,74,31,144,31,235,31,144,31,20,31,158,31,158,30,158,29,71,31,195,31,195,30,195,29,168,31,168,30,128,31,128,30,128,29,232,31,231,31,118,31,118,30,223,31,227,31,227,30,227,29,9,31,63,31,218,31,218,30,218,29,218,28,203,31,106,31,236,31,3,31,159,31,253,31,253,30,130,31,222,31,22,31,22,30,200,31,46,31,120,31,157,31,11,31,89,31,144,31,120,31,113,31,185,31,215,31,148,31,199,31,49,31,49,30,92,31,40,31,40,30,38,31,151,31,151,30,146,31,233,31,121,31,101,31,153,31,97,31,2,31,32,31,111,31,111,30,8,31,174,31,245,31,245,30,245,29,4,31,97,31,204,31,162,31,86,31,49,31,49,30,165,31,235,31,173,31,173,30,150,31,162,31,67,31,56,31,56,30,82,31,82,30,187,31,191,31,30,31,244,31,218,31,218,30,141,31,141,30,201,31,105,31,29,31,201,31,153,31,149,31,31,31,31,30,160,31,28,31,112,31,116,31,125,31,172,31,172,30,200,31,44,31,155,31,155,30,213,31,57,31,14,31,14,30,172,31,86,31,195,31,195,30,193,31,193,30,214,31,241,31,163,31,244,31,160,31,52,31,53,31,154,31,142,31,225,31,225,30,98,31,121,31,19,31,19,30,19,29,38,31,216,31,216,30,9,31,136,31,157,31,174,31,188,31,13,31,13,30,149,31,221,31,60,31,165,31,101,31,101,31,32,31,157,31,20,31,214,31,17,31,159,31,49,31,49,30,86,31,225,31,48,31,139,31,206,31,206,30,206,29,7,31,7,30,74,31,47,31,105,31,123,31,72,31,174,31,181,31,233,31,186,31,226,31,45,31,131,31,219,31,212,31,2,31,30,31,227,31,28,31,1,31,236,31,198,31,202,31,202,30,114,31,152,31,132,31,11,31,148,31,148,30,159,31,116,31,128,31,224,31,200,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
