-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_664 is
end project_tb_664;

architecture project_tb_arch_664 of project_tb_664 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 861;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,234,0,197,0,201,0,191,0,71,0,124,0,161,0,17,0,43,0,102,0,65,0,97,0,126,0,0,0,73,0,199,0,60,0,128,0,59,0,220,0,0,0,189,0,0,0,0,0,0,0,42,0,114,0,253,0,0,0,61,0,0,0,42,0,117,0,221,0,181,0,172,0,31,0,18,0,127,0,164,0,18,0,82,0,218,0,117,0,248,0,21,0,199,0,231,0,159,0,91,0,163,0,31,0,207,0,27,0,109,0,6,0,196,0,121,0,223,0,245,0,200,0,242,0,168,0,128,0,113,0,64,0,0,0,76,0,115,0,128,0,0,0,13,0,158,0,0,0,208,0,116,0,0,0,0,0,32,0,136,0,226,0,46,0,0,0,95,0,43,0,109,0,240,0,144,0,73,0,84,0,35,0,239,0,26,0,89,0,139,0,196,0,34,0,171,0,23,0,136,0,144,0,0,0,39,0,165,0,46,0,0,0,207,0,255,0,110,0,195,0,66,0,154,0,0,0,0,0,48,0,131,0,54,0,213,0,0,0,103,0,0,0,51,0,0,0,219,0,104,0,35,0,106,0,177,0,111,0,183,0,182,0,101,0,0,0,63,0,0,0,198,0,106,0,62,0,0,0,67,0,107,0,41,0,189,0,199,0,0,0,130,0,173,0,179,0,218,0,8,0,200,0,64,0,218,0,153,0,106,0,186,0,223,0,17,0,51,0,159,0,247,0,0,0,139,0,202,0,239,0,182,0,0,0,34,0,152,0,34,0,134,0,0,0,84,0,107,0,215,0,50,0,235,0,38,0,172,0,0,0,186,0,197,0,0,0,0,0,90,0,155,0,178,0,0,0,89,0,79,0,0,0,191,0,0,0,60,0,0,0,20,0,224,0,106,0,139,0,68,0,98,0,0,0,135,0,228,0,206,0,131,0,85,0,130,0,172,0,0,0,12,0,57,0,0,0,127,0,75,0,90,0,89,0,16,0,72,0,46,0,255,0,239,0,70,0,224,0,39,0,65,0,184,0,106,0,73,0,168,0,0,0,7,0,128,0,202,0,3,0,64,0,221,0,239,0,169,0,37,0,104,0,144,0,0,0,195,0,0,0,193,0,203,0,193,0,67,0,226,0,186,0,50,0,0,0,0,0,125,0,119,0,54,0,84,0,0,0,38,0,0,0,134,0,0,0,38,0,173,0,223,0,141,0,161,0,139,0,0,0,193,0,72,0,0,0,106,0,105,0,112,0,65,0,163,0,148,0,74,0,0,0,228,0,210,0,3,0,124,0,90,0,0,0,15,0,83,0,212,0,137,0,142,0,191,0,26,0,9,0,181,0,143,0,0,0,215,0,85,0,0,0,66,0,0,0,20,0,0,0,53,0,0,0,173,0,135,0,60,0,111,0,106,0,0,0,169,0,242,0,102,0,0,0,0,0,231,0,204,0,0,0,96,0,54,0,51,0,226,0,209,0,160,0,147,0,86,0,30,0,224,0,0,0,193,0,5,0,139,0,0,0,164,0,4,0,135,0,222,0,226,0,162,0,179,0,61,0,153,0,0,0,188,0,26,0,9,0,141,0,63,0,0,0,174,0,45,0,97,0,17,0,79,0,35,0,0,0,240,0,173,0,0,0,0,0,188,0,7,0,234,0,90,0,8,0,201,0,12,0,229,0,93,0,253,0,219,0,99,0,18,0,18,0,137,0,0,0,162,0,76,0,0,0,240,0,68,0,169,0,0,0,26,0,92,0,250,0,0,0,126,0,252,0,228,0,155,0,213,0,186,0,202,0,154,0,0,0,86,0,0,0,38,0,92,0,101,0,81,0,20,0,69,0,107,0,105,0,241,0,83,0,65,0,93,0,14,0,182,0,166,0,0,0,135,0,253,0,0,0,0,0,216,0,164,0,75,0,114,0,33,0,219,0,145,0,61,0,20,0,133,0,175,0,248,0,244,0,81,0,206,0,253,0,32,0,0,0,205,0,91,0,190,0,108,0,42,0,55,0,100,0,193,0,233,0,63,0,173,0,253,0,211,0,116,0,0,0,89,0,105,0,29,0,0,0,108,0,114,0,172,0,0,0,188,0,180,0,244,0,40,0,30,0,0,0,116,0,197,0,222,0,71,0,4,0,198,0,27,0,0,0,0,0,43,0,135,0,0,0,32,0,0,0,159,0,110,0,31,0,242,0,174,0,77,0,206,0,236,0,191,0,242,0,183,0,245,0,65,0,200,0,164,0,108,0,99,0,0,0,117,0,53,0,78,0,131,0,151,0,197,0,127,0,0,0,193,0,133,0,180,0,136,0,221,0,244,0,189,0,8,0,0,0,157,0,0,0,212,0,30,0,0,0,203,0,56,0,47,0,231,0,244,0,0,0,227,0,0,0,87,0,190,0,0,0,98,0,30,0,205,0,212,0,0,0,75,0,0,0,163,0,207,0,62,0,114,0,84,0,213,0,0,0,0,0,0,0,183,0,111,0,214,0,59,0,220,0,11,0,57,0,240,0,39,0,124,0,127,0,0,0,122,0,15,0,7,0,0,0,0,0,85,0,50,0,201,0,147,0,86,0,99,0,75,0,190,0,20,0,176,0,0,0,10,0,228,0,181,0,34,0,84,0,46,0,230,0,229,0,0,0,113,0,0,0,129,0,225,0,150,0,98,0,187,0,185,0,0,0,116,0,0,0,0,0,232,0,62,0,0,0,11,0,193,0,192,0,126,0,69,0,229,0,148,0,239,0,185,0,165,0,0,0,188,0,0,0,111,0,189,0,55,0,182,0,160,0,0,0,165,0,65,0,223,0,169,0,26,0,146,0,246,0,0,0,0,0,0,0,0,0,58,0,123,0,0,0,116,0,0,0,94,0,150,0,103,0,240,0,127,0,0,0,0,0,31,0,113,0,13,0,0,0,44,0,104,0,0,0,66,0,0,0,94,0,243,0,187,0,32,0,230,0,0,0,66,0,0,0,0,0,0,0,0,0,198,0,55,0,83,0,0,0,214,0,0,0,164,0,0,0,34,0,79,0,130,0,0,0,35,0,122,0,243,0,186,0,60,0,44,0,39,0,67,0,124,0,0,0,101,0,0,0,182,0,9,0,165,0,241,0,117,0,90,0,34,0,147,0,142,0,161,0,222,0,0,0,40,0,0,0,177,0,4,0,0,0,138,0,0,0,0,0,147,0,199,0,0,0,183,0,0,0,116,0,227,0,216,0,206,0,0,0,42,0,106,0,117,0,242,0,136,0,147,0,19,0,167,0,78,0,0,0,198,0,96,0,226,0,0,0,9,0,52,0,225,0,0,0,61,0,225,0,71,0,34,0,69,0,49,0,248,0,196,0,96,0,135,0,75,0,65,0,232,0,94,0,146,0,140,0,118,0,247,0,0,0,203,0,85,0,131,0,89,0,0,0,153,0,108,0,123,0,41,0,178,0,108,0,215,0,116,0,87,0,114,0,199,0,95,0,225,0,0,0,159,0,0,0,24,0,245,0,143,0,13,0,244,0,132,0,136,0,179,0,181,0,0,0,219,0,78,0,147,0,101,0,239,0,8,0,0,0,76,0,0,0,0,0,87,0,55,0,49,0,29,0,252,0,212,0,236,0,186,0,67,0,138,0,222,0,239,0,120,0,188,0,173,0,0,0,0,0,92,0,240,0,0,0,161,0,252,0,143,0,0,0,7,0,99,0,0,0,3,0,26,0,0,0,46,0,107,0,106,0,0,0,219,0,0,0,2,0,154,0,0,0,0,0,176,0,147,0,147,0,26,0,206,0,50,0,217,0,225,0,203,0,47,0,79,0,101,0,6,0,73,0,249,0,14,0,47,0,221,0,251,0,230,0,226,0,189,0,214,0,0,0,0,0);
signal scenario_full  : scenario_type := (195,31,234,31,197,31,201,31,191,31,71,31,124,31,161,31,17,31,43,31,102,31,65,31,97,31,126,31,126,30,73,31,199,31,60,31,128,31,59,31,220,31,220,30,189,31,189,30,189,29,189,28,42,31,114,31,253,31,253,30,61,31,61,30,42,31,117,31,221,31,181,31,172,31,31,31,18,31,127,31,164,31,18,31,82,31,218,31,117,31,248,31,21,31,199,31,231,31,159,31,91,31,163,31,31,31,207,31,27,31,109,31,6,31,196,31,121,31,223,31,245,31,200,31,242,31,168,31,128,31,113,31,64,31,64,30,76,31,115,31,128,31,128,30,13,31,158,31,158,30,208,31,116,31,116,30,116,29,32,31,136,31,226,31,46,31,46,30,95,31,43,31,109,31,240,31,144,31,73,31,84,31,35,31,239,31,26,31,89,31,139,31,196,31,34,31,171,31,23,31,136,31,144,31,144,30,39,31,165,31,46,31,46,30,207,31,255,31,110,31,195,31,66,31,154,31,154,30,154,29,48,31,131,31,54,31,213,31,213,30,103,31,103,30,51,31,51,30,219,31,104,31,35,31,106,31,177,31,111,31,183,31,182,31,101,31,101,30,63,31,63,30,198,31,106,31,62,31,62,30,67,31,107,31,41,31,189,31,199,31,199,30,130,31,173,31,179,31,218,31,8,31,200,31,64,31,218,31,153,31,106,31,186,31,223,31,17,31,51,31,159,31,247,31,247,30,139,31,202,31,239,31,182,31,182,30,34,31,152,31,34,31,134,31,134,30,84,31,107,31,215,31,50,31,235,31,38,31,172,31,172,30,186,31,197,31,197,30,197,29,90,31,155,31,178,31,178,30,89,31,79,31,79,30,191,31,191,30,60,31,60,30,20,31,224,31,106,31,139,31,68,31,98,31,98,30,135,31,228,31,206,31,131,31,85,31,130,31,172,31,172,30,12,31,57,31,57,30,127,31,75,31,90,31,89,31,16,31,72,31,46,31,255,31,239,31,70,31,224,31,39,31,65,31,184,31,106,31,73,31,168,31,168,30,7,31,128,31,202,31,3,31,64,31,221,31,239,31,169,31,37,31,104,31,144,31,144,30,195,31,195,30,193,31,203,31,193,31,67,31,226,31,186,31,50,31,50,30,50,29,125,31,119,31,54,31,84,31,84,30,38,31,38,30,134,31,134,30,38,31,173,31,223,31,141,31,161,31,139,31,139,30,193,31,72,31,72,30,106,31,105,31,112,31,65,31,163,31,148,31,74,31,74,30,228,31,210,31,3,31,124,31,90,31,90,30,15,31,83,31,212,31,137,31,142,31,191,31,26,31,9,31,181,31,143,31,143,30,215,31,85,31,85,30,66,31,66,30,20,31,20,30,53,31,53,30,173,31,135,31,60,31,111,31,106,31,106,30,169,31,242,31,102,31,102,30,102,29,231,31,204,31,204,30,96,31,54,31,51,31,226,31,209,31,160,31,147,31,86,31,30,31,224,31,224,30,193,31,5,31,139,31,139,30,164,31,4,31,135,31,222,31,226,31,162,31,179,31,61,31,153,31,153,30,188,31,26,31,9,31,141,31,63,31,63,30,174,31,45,31,97,31,17,31,79,31,35,31,35,30,240,31,173,31,173,30,173,29,188,31,7,31,234,31,90,31,8,31,201,31,12,31,229,31,93,31,253,31,219,31,99,31,18,31,18,31,137,31,137,30,162,31,76,31,76,30,240,31,68,31,169,31,169,30,26,31,92,31,250,31,250,30,126,31,252,31,228,31,155,31,213,31,186,31,202,31,154,31,154,30,86,31,86,30,38,31,92,31,101,31,81,31,20,31,69,31,107,31,105,31,241,31,83,31,65,31,93,31,14,31,182,31,166,31,166,30,135,31,253,31,253,30,253,29,216,31,164,31,75,31,114,31,33,31,219,31,145,31,61,31,20,31,133,31,175,31,248,31,244,31,81,31,206,31,253,31,32,31,32,30,205,31,91,31,190,31,108,31,42,31,55,31,100,31,193,31,233,31,63,31,173,31,253,31,211,31,116,31,116,30,89,31,105,31,29,31,29,30,108,31,114,31,172,31,172,30,188,31,180,31,244,31,40,31,30,31,30,30,116,31,197,31,222,31,71,31,4,31,198,31,27,31,27,30,27,29,43,31,135,31,135,30,32,31,32,30,159,31,110,31,31,31,242,31,174,31,77,31,206,31,236,31,191,31,242,31,183,31,245,31,65,31,200,31,164,31,108,31,99,31,99,30,117,31,53,31,78,31,131,31,151,31,197,31,127,31,127,30,193,31,133,31,180,31,136,31,221,31,244,31,189,31,8,31,8,30,157,31,157,30,212,31,30,31,30,30,203,31,56,31,47,31,231,31,244,31,244,30,227,31,227,30,87,31,190,31,190,30,98,31,30,31,205,31,212,31,212,30,75,31,75,30,163,31,207,31,62,31,114,31,84,31,213,31,213,30,213,29,213,28,183,31,111,31,214,31,59,31,220,31,11,31,57,31,240,31,39,31,124,31,127,31,127,30,122,31,15,31,7,31,7,30,7,29,85,31,50,31,201,31,147,31,86,31,99,31,75,31,190,31,20,31,176,31,176,30,10,31,228,31,181,31,34,31,84,31,46,31,230,31,229,31,229,30,113,31,113,30,129,31,225,31,150,31,98,31,187,31,185,31,185,30,116,31,116,30,116,29,232,31,62,31,62,30,11,31,193,31,192,31,126,31,69,31,229,31,148,31,239,31,185,31,165,31,165,30,188,31,188,30,111,31,189,31,55,31,182,31,160,31,160,30,165,31,65,31,223,31,169,31,26,31,146,31,246,31,246,30,246,29,246,28,246,27,58,31,123,31,123,30,116,31,116,30,94,31,150,31,103,31,240,31,127,31,127,30,127,29,31,31,113,31,13,31,13,30,44,31,104,31,104,30,66,31,66,30,94,31,243,31,187,31,32,31,230,31,230,30,66,31,66,30,66,29,66,28,66,27,198,31,55,31,83,31,83,30,214,31,214,30,164,31,164,30,34,31,79,31,130,31,130,30,35,31,122,31,243,31,186,31,60,31,44,31,39,31,67,31,124,31,124,30,101,31,101,30,182,31,9,31,165,31,241,31,117,31,90,31,34,31,147,31,142,31,161,31,222,31,222,30,40,31,40,30,177,31,4,31,4,30,138,31,138,30,138,29,147,31,199,31,199,30,183,31,183,30,116,31,227,31,216,31,206,31,206,30,42,31,106,31,117,31,242,31,136,31,147,31,19,31,167,31,78,31,78,30,198,31,96,31,226,31,226,30,9,31,52,31,225,31,225,30,61,31,225,31,71,31,34,31,69,31,49,31,248,31,196,31,96,31,135,31,75,31,65,31,232,31,94,31,146,31,140,31,118,31,247,31,247,30,203,31,85,31,131,31,89,31,89,30,153,31,108,31,123,31,41,31,178,31,108,31,215,31,116,31,87,31,114,31,199,31,95,31,225,31,225,30,159,31,159,30,24,31,245,31,143,31,13,31,244,31,132,31,136,31,179,31,181,31,181,30,219,31,78,31,147,31,101,31,239,31,8,31,8,30,76,31,76,30,76,29,87,31,55,31,49,31,29,31,252,31,212,31,236,31,186,31,67,31,138,31,222,31,239,31,120,31,188,31,173,31,173,30,173,29,92,31,240,31,240,30,161,31,252,31,143,31,143,30,7,31,99,31,99,30,3,31,26,31,26,30,46,31,107,31,106,31,106,30,219,31,219,30,2,31,154,31,154,30,154,29,176,31,147,31,147,31,26,31,206,31,50,31,217,31,225,31,203,31,47,31,79,31,101,31,6,31,73,31,249,31,14,31,47,31,221,31,251,31,230,31,226,31,189,31,214,31,214,30,214,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
