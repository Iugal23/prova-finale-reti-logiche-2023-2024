-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 180;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,107,0,0,0,147,0,44,0,250,0,0,0,93,0,59,0,200,0,0,0,249,0,165,0,0,0,220,0,205,0,45,0,82,0,187,0,92,0,0,0,71,0,0,0,0,0,75,0,0,0,115,0,213,0,245,0,179,0,175,0,209,0,28,0,146,0,26,0,128,0,225,0,68,0,66,0,195,0,0,0,22,0,33,0,4,0,0,0,24,0,0,0,191,0,174,0,239,0,0,0,135,0,250,0,155,0,175,0,146,0,234,0,81,0,58,0,134,0,187,0,0,0,238,0,10,0,0,0,79,0,203,0,249,0,19,0,246,0,254,0,217,0,32,0,125,0,154,0,113,0,52,0,238,0,189,0,0,0,0,0,227,0,27,0,41,0,22,0,222,0,21,0,0,0,105,0,0,0,24,0,176,0,215,0,0,0,0,0,126,0,81,0,151,0,226,0,131,0,0,0,234,0,0,0,81,0,170,0,1,0,174,0,29,0,18,0,134,0,167,0,235,0,142,0,253,0,208,0,30,0,0,0,126,0,5,0,253,0,169,0,249,0,165,0,224,0,75,0,253,0,172,0,133,0,58,0,20,0,22,0,17,0,54,0,130,0,0,0,0,0,0,0,117,0,172,0,0,0,182,0,36,0,140,0,87,0,107,0,170,0,0,0,127,0,0,0,255,0,206,0,45,0,16,0,112,0,114,0,104,0,201,0,160,0,167,0,16,0,246,0,236,0,146,0,237,0,36,0,0,0,0,0,54,0,0,0,55,0,0,0,213,0,14,0,181,0,213,0,250,0,124,0,178,0,0,0,216,0);
signal scenario_full  : scenario_type := (250,31,107,31,107,30,147,31,44,31,250,31,250,30,93,31,59,31,200,31,200,30,249,31,165,31,165,30,220,31,205,31,45,31,82,31,187,31,92,31,92,30,71,31,71,30,71,29,75,31,75,30,115,31,213,31,245,31,179,31,175,31,209,31,28,31,146,31,26,31,128,31,225,31,68,31,66,31,195,31,195,30,22,31,33,31,4,31,4,30,24,31,24,30,191,31,174,31,239,31,239,30,135,31,250,31,155,31,175,31,146,31,234,31,81,31,58,31,134,31,187,31,187,30,238,31,10,31,10,30,79,31,203,31,249,31,19,31,246,31,254,31,217,31,32,31,125,31,154,31,113,31,52,31,238,31,189,31,189,30,189,29,227,31,27,31,41,31,22,31,222,31,21,31,21,30,105,31,105,30,24,31,176,31,215,31,215,30,215,29,126,31,81,31,151,31,226,31,131,31,131,30,234,31,234,30,81,31,170,31,1,31,174,31,29,31,18,31,134,31,167,31,235,31,142,31,253,31,208,31,30,31,30,30,126,31,5,31,253,31,169,31,249,31,165,31,224,31,75,31,253,31,172,31,133,31,58,31,20,31,22,31,17,31,54,31,130,31,130,30,130,29,130,28,117,31,172,31,172,30,182,31,36,31,140,31,87,31,107,31,170,31,170,30,127,31,127,30,255,31,206,31,45,31,16,31,112,31,114,31,104,31,201,31,160,31,167,31,16,31,246,31,236,31,146,31,237,31,36,31,36,30,36,29,54,31,54,30,55,31,55,30,213,31,14,31,181,31,213,31,250,31,124,31,178,31,178,30,216,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
