-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 643;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,218,0,0,0,50,0,0,0,234,0,41,0,131,0,235,0,0,0,15,0,0,0,0,0,217,0,0,0,151,0,112,0,0,0,40,0,124,0,210,0,111,0,0,0,0,0,11,0,98,0,227,0,223,0,219,0,80,0,182,0,30,0,190,0,5,0,5,0,92,0,64,0,189,0,168,0,101,0,0,0,0,0,245,0,20,0,24,0,196,0,0,0,121,0,0,0,40,0,105,0,190,0,0,0,145,0,183,0,33,0,0,0,0,0,255,0,107,0,71,0,217,0,77,0,221,0,56,0,0,0,6,0,0,0,142,0,255,0,238,0,7,0,0,0,28,0,45,0,28,0,0,0,0,0,120,0,0,0,108,0,246,0,161,0,0,0,53,0,0,0,0,0,100,0,0,0,100,0,243,0,0,0,113,0,203,0,149,0,59,0,166,0,120,0,55,0,16,0,0,0,53,0,62,0,226,0,192,0,18,0,144,0,230,0,0,0,130,0,182,0,69,0,0,0,18,0,248,0,212,0,124,0,59,0,60,0,255,0,0,0,250,0,102,0,147,0,49,0,6,0,0,0,0,0,217,0,0,0,35,0,0,0,0,0,194,0,0,0,16,0,131,0,0,0,177,0,220,0,19,0,230,0,121,0,0,0,0,0,90,0,89,0,182,0,104,0,107,0,93,0,0,0,0,0,40,0,0,0,0,0,72,0,35,0,181,0,0,0,0,0,11,0,0,0,0,0,64,0,0,0,10,0,0,0,28,0,0,0,164,0,133,0,144,0,252,0,35,0,53,0,118,0,11,0,0,0,58,0,161,0,0,0,0,0,56,0,229,0,139,0,204,0,144,0,11,0,92,0,23,0,2,0,0,0,183,0,67,0,173,0,104,0,242,0,141,0,0,0,0,0,52,0,74,0,21,0,219,0,66,0,189,0,250,0,0,0,207,0,111,0,122,0,61,0,0,0,125,0,14,0,67,0,210,0,160,0,150,0,0,0,52,0,0,0,24,0,136,0,15,0,246,0,236,0,41,0,0,0,88,0,44,0,203,0,220,0,243,0,144,0,86,0,99,0,0,0,116,0,166,0,83,0,0,0,0,0,219,0,81,0,220,0,229,0,238,0,246,0,147,0,12,0,0,0,206,0,0,0,0,0,187,0,136,0,149,0,2,0,19,0,175,0,95,0,118,0,227,0,231,0,0,0,157,0,136,0,80,0,187,0,0,0,63,0,214,0,71,0,0,0,141,0,0,0,0,0,0,0,239,0,50,0,230,0,73,0,0,0,0,0,0,0,0,0,228,0,212,0,44,0,218,0,113,0,57,0,7,0,10,0,213,0,246,0,152,0,0,0,105,0,144,0,165,0,99,0,68,0,85,0,0,0,163,0,171,0,69,0,158,0,0,0,50,0,72,0,29,0,193,0,52,0,42,0,50,0,60,0,215,0,153,0,25,0,187,0,121,0,131,0,0,0,212,0,69,0,147,0,138,0,175,0,20,0,116,0,0,0,236,0,0,0,147,0,0,0,0,0,161,0,99,0,14,0,240,0,72,0,250,0,0,0,211,0,153,0,0,0,135,0,0,0,185,0,0,0,69,0,20,0,108,0,0,0,109,0,174,0,187,0,219,0,17,0,21,0,123,0,116,0,125,0,209,0,0,0,0,0,64,0,199,0,0,0,245,0,35,0,0,0,0,0,183,0,191,0,183,0,49,0,45,0,189,0,135,0,152,0,0,0,0,0,254,0,152,0,200,0,205,0,2,0,0,0,222,0,13,0,159,0,223,0,155,0,102,0,252,0,150,0,25,0,0,0,190,0,0,0,0,0,154,0,56,0,105,0,82,0,0,0,141,0,0,0,0,0,94,0,139,0,232,0,219,0,0,0,169,0,98,0,95,0,0,0,132,0,6,0,0,0,253,0,157,0,105,0,23,0,103,0,0,0,123,0,135,0,240,0,202,0,185,0,0,0,0,0,204,0,136,0,135,0,164,0,0,0,148,0,81,0,223,0,95,0,8,0,222,0,147,0,189,0,59,0,86,0,253,0,224,0,232,0,14,0,34,0,156,0,14,0,97,0,14,0,117,0,2,0,58,0,136,0,74,0,144,0,152,0,0,0,0,0,47,0,158,0,51,0,242,0,0,0,218,0,12,0,235,0,84,0,193,0,0,0,135,0,157,0,165,0,0,0,188,0,0,0,244,0,21,0,96,0,94,0,248,0,0,0,104,0,113,0,8,0,127,0,223,0,206,0,79,0,247,0,0,0,254,0,196,0,187,0,131,0,0,0,195,0,3,0,99,0,213,0,16,0,44,0,0,0,52,0,0,0,0,0,234,0,70,0,0,0,80,0,58,0,25,0,153,0,149,0,0,0,9,0,118,0,31,0,215,0,139,0,37,0,15,0,163,0,13,0,2,0,213,0,0,0,209,0,0,0,14,0,152,0,0,0,217,0,108,0,0,0,139,0,92,0,105,0,101,0,100,0,0,0,0,0,180,0,205,0,238,0,157,0,0,0,154,0,188,0,0,0,181,0,130,0,0,0,249,0,223,0,223,0,223,0,130,0,231,0,199,0,142,0,160,0,0,0,88,0,98,0,0,0,112,0,167,0,187,0,95,0,139,0,204,0,0,0,112,0,122,0,143,0,229,0,31,0,162,0,18,0,5,0,95,0,146,0,11,0,250,0,107,0,0,0,211,0,42,0,0,0,121,0,240,0,0,0,0,0,0,0,39,0,85,0,157,0,21,0,190,0,9,0,194,0,118,0,0,0,0,0,12,0,0,0,0,0,78,0,69,0,151,0,234,0,226,0,29,0,98,0,91,0,0,0,0,0,0,0,0,0,226,0,133,0,129,0,0,0,0,0,101,0,0,0,35,0,251,0);
signal scenario_full  : scenario_type := (0,0,0,0,218,31,218,30,50,31,50,30,234,31,41,31,131,31,235,31,235,30,15,31,15,30,15,29,217,31,217,30,151,31,112,31,112,30,40,31,124,31,210,31,111,31,111,30,111,29,11,31,98,31,227,31,223,31,219,31,80,31,182,31,30,31,190,31,5,31,5,31,92,31,64,31,189,31,168,31,101,31,101,30,101,29,245,31,20,31,24,31,196,31,196,30,121,31,121,30,40,31,105,31,190,31,190,30,145,31,183,31,33,31,33,30,33,29,255,31,107,31,71,31,217,31,77,31,221,31,56,31,56,30,6,31,6,30,142,31,255,31,238,31,7,31,7,30,28,31,45,31,28,31,28,30,28,29,120,31,120,30,108,31,246,31,161,31,161,30,53,31,53,30,53,29,100,31,100,30,100,31,243,31,243,30,113,31,203,31,149,31,59,31,166,31,120,31,55,31,16,31,16,30,53,31,62,31,226,31,192,31,18,31,144,31,230,31,230,30,130,31,182,31,69,31,69,30,18,31,248,31,212,31,124,31,59,31,60,31,255,31,255,30,250,31,102,31,147,31,49,31,6,31,6,30,6,29,217,31,217,30,35,31,35,30,35,29,194,31,194,30,16,31,131,31,131,30,177,31,220,31,19,31,230,31,121,31,121,30,121,29,90,31,89,31,182,31,104,31,107,31,93,31,93,30,93,29,40,31,40,30,40,29,72,31,35,31,181,31,181,30,181,29,11,31,11,30,11,29,64,31,64,30,10,31,10,30,28,31,28,30,164,31,133,31,144,31,252,31,35,31,53,31,118,31,11,31,11,30,58,31,161,31,161,30,161,29,56,31,229,31,139,31,204,31,144,31,11,31,92,31,23,31,2,31,2,30,183,31,67,31,173,31,104,31,242,31,141,31,141,30,141,29,52,31,74,31,21,31,219,31,66,31,189,31,250,31,250,30,207,31,111,31,122,31,61,31,61,30,125,31,14,31,67,31,210,31,160,31,150,31,150,30,52,31,52,30,24,31,136,31,15,31,246,31,236,31,41,31,41,30,88,31,44,31,203,31,220,31,243,31,144,31,86,31,99,31,99,30,116,31,166,31,83,31,83,30,83,29,219,31,81,31,220,31,229,31,238,31,246,31,147,31,12,31,12,30,206,31,206,30,206,29,187,31,136,31,149,31,2,31,19,31,175,31,95,31,118,31,227,31,231,31,231,30,157,31,136,31,80,31,187,31,187,30,63,31,214,31,71,31,71,30,141,31,141,30,141,29,141,28,239,31,50,31,230,31,73,31,73,30,73,29,73,28,73,27,228,31,212,31,44,31,218,31,113,31,57,31,7,31,10,31,213,31,246,31,152,31,152,30,105,31,144,31,165,31,99,31,68,31,85,31,85,30,163,31,171,31,69,31,158,31,158,30,50,31,72,31,29,31,193,31,52,31,42,31,50,31,60,31,215,31,153,31,25,31,187,31,121,31,131,31,131,30,212,31,69,31,147,31,138,31,175,31,20,31,116,31,116,30,236,31,236,30,147,31,147,30,147,29,161,31,99,31,14,31,240,31,72,31,250,31,250,30,211,31,153,31,153,30,135,31,135,30,185,31,185,30,69,31,20,31,108,31,108,30,109,31,174,31,187,31,219,31,17,31,21,31,123,31,116,31,125,31,209,31,209,30,209,29,64,31,199,31,199,30,245,31,35,31,35,30,35,29,183,31,191,31,183,31,49,31,45,31,189,31,135,31,152,31,152,30,152,29,254,31,152,31,200,31,205,31,2,31,2,30,222,31,13,31,159,31,223,31,155,31,102,31,252,31,150,31,25,31,25,30,190,31,190,30,190,29,154,31,56,31,105,31,82,31,82,30,141,31,141,30,141,29,94,31,139,31,232,31,219,31,219,30,169,31,98,31,95,31,95,30,132,31,6,31,6,30,253,31,157,31,105,31,23,31,103,31,103,30,123,31,135,31,240,31,202,31,185,31,185,30,185,29,204,31,136,31,135,31,164,31,164,30,148,31,81,31,223,31,95,31,8,31,222,31,147,31,189,31,59,31,86,31,253,31,224,31,232,31,14,31,34,31,156,31,14,31,97,31,14,31,117,31,2,31,58,31,136,31,74,31,144,31,152,31,152,30,152,29,47,31,158,31,51,31,242,31,242,30,218,31,12,31,235,31,84,31,193,31,193,30,135,31,157,31,165,31,165,30,188,31,188,30,244,31,21,31,96,31,94,31,248,31,248,30,104,31,113,31,8,31,127,31,223,31,206,31,79,31,247,31,247,30,254,31,196,31,187,31,131,31,131,30,195,31,3,31,99,31,213,31,16,31,44,31,44,30,52,31,52,30,52,29,234,31,70,31,70,30,80,31,58,31,25,31,153,31,149,31,149,30,9,31,118,31,31,31,215,31,139,31,37,31,15,31,163,31,13,31,2,31,213,31,213,30,209,31,209,30,14,31,152,31,152,30,217,31,108,31,108,30,139,31,92,31,105,31,101,31,100,31,100,30,100,29,180,31,205,31,238,31,157,31,157,30,154,31,188,31,188,30,181,31,130,31,130,30,249,31,223,31,223,31,223,31,130,31,231,31,199,31,142,31,160,31,160,30,88,31,98,31,98,30,112,31,167,31,187,31,95,31,139,31,204,31,204,30,112,31,122,31,143,31,229,31,31,31,162,31,18,31,5,31,95,31,146,31,11,31,250,31,107,31,107,30,211,31,42,31,42,30,121,31,240,31,240,30,240,29,240,28,39,31,85,31,157,31,21,31,190,31,9,31,194,31,118,31,118,30,118,29,12,31,12,30,12,29,78,31,69,31,151,31,234,31,226,31,29,31,98,31,91,31,91,30,91,29,91,28,91,27,226,31,133,31,129,31,129,30,129,29,101,31,101,30,35,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
