-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 660;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (158,0,0,0,139,0,84,0,0,0,209,0,0,0,0,0,188,0,178,0,0,0,0,0,11,0,103,0,48,0,150,0,159,0,0,0,94,0,0,0,153,0,0,0,145,0,217,0,158,0,138,0,0,0,230,0,241,0,79,0,182,0,85,0,149,0,0,0,250,0,120,0,209,0,244,0,253,0,8,0,27,0,81,0,237,0,0,0,186,0,0,0,117,0,146,0,7,0,219,0,51,0,0,0,151,0,190,0,143,0,25,0,0,0,35,0,110,0,86,0,196,0,218,0,203,0,0,0,229,0,0,0,0,0,42,0,196,0,32,0,189,0,54,0,158,0,142,0,66,0,142,0,189,0,0,0,152,0,150,0,148,0,196,0,152,0,17,0,211,0,0,0,0,0,35,0,145,0,217,0,25,0,59,0,200,0,205,0,23,0,63,0,104,0,197,0,53,0,40,0,93,0,170,0,157,0,54,0,132,0,126,0,134,0,48,0,12,0,135,0,0,0,245,0,228,0,147,0,241,0,8,0,95,0,57,0,219,0,14,0,0,0,0,0,117,0,147,0,0,0,200,0,2,0,17,0,0,0,168,0,169,0,133,0,85,0,124,0,175,0,0,0,214,0,201,0,222,0,126,0,152,0,0,0,62,0,214,0,234,0,61,0,49,0,58,0,220,0,134,0,17,0,50,0,230,0,48,0,55,0,0,0,24,0,216,0,37,0,118,0,201,0,27,0,11,0,160,0,175,0,15,0,126,0,198,0,89,0,0,0,243,0,0,0,82,0,68,0,0,0,101,0,204,0,88,0,170,0,10,0,0,0,56,0,243,0,0,0,208,0,71,0,154,0,201,0,97,0,46,0,163,0,119,0,214,0,0,0,87,0,0,0,0,0,58,0,68,0,132,0,120,0,0,0,209,0,0,0,0,0,0,0,195,0,0,0,0,0,0,0,221,0,0,0,0,0,183,0,5,0,0,0,0,0,12,0,244,0,67,0,69,0,11,0,0,0,0,0,0,0,47,0,71,0,14,0,227,0,251,0,0,0,39,0,131,0,0,0,41,0,124,0,203,0,39,0,253,0,51,0,142,0,210,0,130,0,163,0,223,0,127,0,27,0,0,0,228,0,221,0,69,0,102,0,3,0,218,0,90,0,0,0,226,0,246,0,106,0,11,0,185,0,121,0,220,0,178,0,215,0,182,0,0,0,188,0,18,0,0,0,218,0,39,0,177,0,238,0,203,0,24,0,127,0,65,0,0,0,218,0,30,0,0,0,206,0,202,0,0,0,20,0,0,0,156,0,238,0,90,0,209,0,168,0,65,0,0,0,0,0,233,0,236,0,0,0,9,0,212,0,204,0,32,0,228,0,51,0,250,0,0,0,130,0,126,0,137,0,3,0,92,0,39,0,132,0,111,0,2,0,245,0,252,0,146,0,72,0,12,0,17,0,98,0,0,0,12,0,0,0,70,0,241,0,75,0,105,0,18,0,0,0,247,0,50,0,158,0,238,0,27,0,7,0,0,0,190,0,0,0,0,0,0,0,107,0,73,0,0,0,17,0,62,0,154,0,129,0,88,0,155,0,42,0,20,0,254,0,0,0,131,0,68,0,0,0,66,0,59,0,129,0,235,0,92,0,197,0,77,0,147,0,0,0,242,0,90,0,78,0,242,0,64,0,212,0,131,0,253,0,147,0,212,0,4,0,112,0,93,0,145,0,0,0,0,0,123,0,19,0,168,0,80,0,227,0,213,0,131,0,83,0,86,0,87,0,194,0,33,0,0,0,0,0,0,0,75,0,217,0,91,0,0,0,150,0,96,0,229,0,193,0,208,0,69,0,165,0,198,0,0,0,118,0,57,0,172,0,0,0,242,0,195,0,213,0,87,0,128,0,48,0,138,0,0,0,0,0,145,0,90,0,152,0,138,0,94,0,66,0,28,0,90,0,99,0,0,0,0,0,155,0,0,0,3,0,0,0,0,0,247,0,232,0,102,0,252,0,12,0,0,0,193,0,118,0,161,0,76,0,236,0,162,0,0,0,138,0,0,0,1,0,175,0,23,0,97,0,216,0,220,0,0,0,44,0,18,0,176,0,68,0,201,0,250,0,163,0,69,0,164,0,56,0,26,0,62,0,102,0,0,0,6,0,0,0,127,0,0,0,0,0,0,0,133,0,0,0,73,0,24,0,213,0,134,0,9,0,0,0,63,0,0,0,156,0,234,0,214,0,223,0,109,0,2,0,208,0,232,0,0,0,0,0,6,0,135,0,119,0,136,0,252,0,20,0,242,0,35,0,252,0,0,0,160,0,252,0,80,0,0,0,255,0,248,0,252,0,78,0,206,0,147,0,0,0,35,0,157,0,218,0,0,0,74,0,8,0,0,0,58,0,132,0,179,0,114,0,206,0,67,0,169,0,246,0,0,0,36,0,0,0,210,0,144,0,98,0,42,0,172,0,249,0,246,0,217,0,228,0,50,0,210,0,177,0,240,0,0,0,87,0,0,0,174,0,28,0,145,0,116,0,201,0,113,0,55,0,22,0,96,0,40,0,211,0,40,0,18,0,140,0,227,0,141,0,85,0,78,0,0,0,9,0,122,0,120,0,0,0,197,0,35,0,213,0,0,0,0,0,0,0,145,0,161,0,184,0,140,0,145,0,191,0,0,0,234,0,67,0,165,0,119,0,45,0,99,0,80,0,103,0,115,0,223,0,159,0,196,0,168,0,189,0,63,0,201,0,41,0,36,0,0,0,0,0,56,0,187,0,0,0,228,0,228,0,176,0,0,0,123,0,0,0,79,0,88,0,73,0,203,0,75,0,41,0,46,0,133,0,61,0,222,0,223,0,181,0,9,0,0,0,0,0,144,0,178,0,138,0,151,0,189,0,164,0,198,0,37,0,195,0,251,0,225,0,165,0,110,0,177,0,253,0,193,0,82,0,210,0,182,0,57,0,161,0,68,0,0,0);
signal scenario_full  : scenario_type := (158,31,158,30,139,31,84,31,84,30,209,31,209,30,209,29,188,31,178,31,178,30,178,29,11,31,103,31,48,31,150,31,159,31,159,30,94,31,94,30,153,31,153,30,145,31,217,31,158,31,138,31,138,30,230,31,241,31,79,31,182,31,85,31,149,31,149,30,250,31,120,31,209,31,244,31,253,31,8,31,27,31,81,31,237,31,237,30,186,31,186,30,117,31,146,31,7,31,219,31,51,31,51,30,151,31,190,31,143,31,25,31,25,30,35,31,110,31,86,31,196,31,218,31,203,31,203,30,229,31,229,30,229,29,42,31,196,31,32,31,189,31,54,31,158,31,142,31,66,31,142,31,189,31,189,30,152,31,150,31,148,31,196,31,152,31,17,31,211,31,211,30,211,29,35,31,145,31,217,31,25,31,59,31,200,31,205,31,23,31,63,31,104,31,197,31,53,31,40,31,93,31,170,31,157,31,54,31,132,31,126,31,134,31,48,31,12,31,135,31,135,30,245,31,228,31,147,31,241,31,8,31,95,31,57,31,219,31,14,31,14,30,14,29,117,31,147,31,147,30,200,31,2,31,17,31,17,30,168,31,169,31,133,31,85,31,124,31,175,31,175,30,214,31,201,31,222,31,126,31,152,31,152,30,62,31,214,31,234,31,61,31,49,31,58,31,220,31,134,31,17,31,50,31,230,31,48,31,55,31,55,30,24,31,216,31,37,31,118,31,201,31,27,31,11,31,160,31,175,31,15,31,126,31,198,31,89,31,89,30,243,31,243,30,82,31,68,31,68,30,101,31,204,31,88,31,170,31,10,31,10,30,56,31,243,31,243,30,208,31,71,31,154,31,201,31,97,31,46,31,163,31,119,31,214,31,214,30,87,31,87,30,87,29,58,31,68,31,132,31,120,31,120,30,209,31,209,30,209,29,209,28,195,31,195,30,195,29,195,28,221,31,221,30,221,29,183,31,5,31,5,30,5,29,12,31,244,31,67,31,69,31,11,31,11,30,11,29,11,28,47,31,71,31,14,31,227,31,251,31,251,30,39,31,131,31,131,30,41,31,124,31,203,31,39,31,253,31,51,31,142,31,210,31,130,31,163,31,223,31,127,31,27,31,27,30,228,31,221,31,69,31,102,31,3,31,218,31,90,31,90,30,226,31,246,31,106,31,11,31,185,31,121,31,220,31,178,31,215,31,182,31,182,30,188,31,18,31,18,30,218,31,39,31,177,31,238,31,203,31,24,31,127,31,65,31,65,30,218,31,30,31,30,30,206,31,202,31,202,30,20,31,20,30,156,31,238,31,90,31,209,31,168,31,65,31,65,30,65,29,233,31,236,31,236,30,9,31,212,31,204,31,32,31,228,31,51,31,250,31,250,30,130,31,126,31,137,31,3,31,92,31,39,31,132,31,111,31,2,31,245,31,252,31,146,31,72,31,12,31,17,31,98,31,98,30,12,31,12,30,70,31,241,31,75,31,105,31,18,31,18,30,247,31,50,31,158,31,238,31,27,31,7,31,7,30,190,31,190,30,190,29,190,28,107,31,73,31,73,30,17,31,62,31,154,31,129,31,88,31,155,31,42,31,20,31,254,31,254,30,131,31,68,31,68,30,66,31,59,31,129,31,235,31,92,31,197,31,77,31,147,31,147,30,242,31,90,31,78,31,242,31,64,31,212,31,131,31,253,31,147,31,212,31,4,31,112,31,93,31,145,31,145,30,145,29,123,31,19,31,168,31,80,31,227,31,213,31,131,31,83,31,86,31,87,31,194,31,33,31,33,30,33,29,33,28,75,31,217,31,91,31,91,30,150,31,96,31,229,31,193,31,208,31,69,31,165,31,198,31,198,30,118,31,57,31,172,31,172,30,242,31,195,31,213,31,87,31,128,31,48,31,138,31,138,30,138,29,145,31,90,31,152,31,138,31,94,31,66,31,28,31,90,31,99,31,99,30,99,29,155,31,155,30,3,31,3,30,3,29,247,31,232,31,102,31,252,31,12,31,12,30,193,31,118,31,161,31,76,31,236,31,162,31,162,30,138,31,138,30,1,31,175,31,23,31,97,31,216,31,220,31,220,30,44,31,18,31,176,31,68,31,201,31,250,31,163,31,69,31,164,31,56,31,26,31,62,31,102,31,102,30,6,31,6,30,127,31,127,30,127,29,127,28,133,31,133,30,73,31,24,31,213,31,134,31,9,31,9,30,63,31,63,30,156,31,234,31,214,31,223,31,109,31,2,31,208,31,232,31,232,30,232,29,6,31,135,31,119,31,136,31,252,31,20,31,242,31,35,31,252,31,252,30,160,31,252,31,80,31,80,30,255,31,248,31,252,31,78,31,206,31,147,31,147,30,35,31,157,31,218,31,218,30,74,31,8,31,8,30,58,31,132,31,179,31,114,31,206,31,67,31,169,31,246,31,246,30,36,31,36,30,210,31,144,31,98,31,42,31,172,31,249,31,246,31,217,31,228,31,50,31,210,31,177,31,240,31,240,30,87,31,87,30,174,31,28,31,145,31,116,31,201,31,113,31,55,31,22,31,96,31,40,31,211,31,40,31,18,31,140,31,227,31,141,31,85,31,78,31,78,30,9,31,122,31,120,31,120,30,197,31,35,31,213,31,213,30,213,29,213,28,145,31,161,31,184,31,140,31,145,31,191,31,191,30,234,31,67,31,165,31,119,31,45,31,99,31,80,31,103,31,115,31,223,31,159,31,196,31,168,31,189,31,63,31,201,31,41,31,36,31,36,30,36,29,56,31,187,31,187,30,228,31,228,31,176,31,176,30,123,31,123,30,79,31,88,31,73,31,203,31,75,31,41,31,46,31,133,31,61,31,222,31,223,31,181,31,9,31,9,30,9,29,144,31,178,31,138,31,151,31,189,31,164,31,198,31,37,31,195,31,251,31,225,31,165,31,110,31,177,31,253,31,193,31,82,31,210,31,182,31,57,31,161,31,68,31,68,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
