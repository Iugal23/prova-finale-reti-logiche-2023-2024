-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 504;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (25,0,234,0,133,0,239,0,188,0,0,0,169,0,159,0,178,0,174,0,211,0,69,0,20,0,0,0,0,0,0,0,0,0,44,0,164,0,5,0,0,0,177,0,0,0,181,0,0,0,0,0,117,0,78,0,60,0,106,0,251,0,120,0,203,0,156,0,0,0,0,0,160,0,32,0,38,0,0,0,99,0,162,0,242,0,249,0,125,0,164,0,98,0,196,0,216,0,42,0,217,0,185,0,120,0,24,0,85,0,0,0,238,0,235,0,77,0,61,0,0,0,153,0,108,0,30,0,170,0,0,0,131,0,70,0,160,0,23,0,0,0,0,0,82,0,116,0,0,0,188,0,60,0,49,0,0,0,0,0,124,0,146,0,160,0,105,0,244,0,0,0,234,0,0,0,180,0,84,0,231,0,75,0,0,0,0,0,175,0,122,0,252,0,163,0,138,0,229,0,252,0,26,0,144,0,97,0,169,0,72,0,159,0,0,0,54,0,0,0,93,0,46,0,25,0,0,0,242,0,68,0,112,0,134,0,48,0,221,0,0,0,27,0,127,0,243,0,0,0,237,0,114,0,164,0,0,0,228,0,16,0,169,0,0,0,0,0,0,0,168,0,224,0,212,0,217,0,248,0,84,0,108,0,0,0,48,0,30,0,255,0,112,0,8,0,63,0,222,0,79,0,0,0,52,0,0,0,229,0,148,0,169,0,211,0,190,0,29,0,170,0,8,0,69,0,212,0,0,0,68,0,0,0,171,0,151,0,0,0,163,0,0,0,254,0,185,0,129,0,75,0,0,0,81,0,15,0,123,0,142,0,0,0,161,0,0,0,168,0,0,0,214,0,177,0,235,0,0,0,232,0,211,0,0,0,11,0,243,0,54,0,65,0,167,0,160,0,148,0,164,0,176,0,100,0,0,0,186,0,147,0,0,0,210,0,95,0,131,0,27,0,162,0,0,0,70,0,233,0,76,0,50,0,105,0,186,0,208,0,0,0,38,0,0,0,251,0,0,0,73,0,56,0,213,0,33,0,37,0,0,0,168,0,157,0,6,0,198,0,0,0,59,0,0,0,0,0,35,0,117,0,0,0,110,0,252,0,62,0,105,0,125,0,0,0,199,0,197,0,0,0,14,0,173,0,35,0,201,0,161,0,241,0,178,0,0,0,72,0,193,0,247,0,222,0,107,0,53,0,97,0,206,0,146,0,46,0,34,0,0,0,122,0,172,0,146,0,0,0,90,0,1,0,231,0,89,0,33,0,80,0,0,0,239,0,143,0,38,0,0,0,223,0,50,0,62,0,12,0,13,0,79,0,64,0,92,0,66,0,249,0,55,0,0,0,31,0,58,0,231,0,42,0,184,0,199,0,234,0,3,0,0,0,11,0,36,0,0,0,225,0,75,0,151,0,83,0,109,0,77,0,247,0,23,0,217,0,177,0,243,0,100,0,19,0,110,0,57,0,186,0,0,0,35,0,123,0,0,0,0,0,0,0,154,0,163,0,4,0,0,0,238,0,0,0,0,0,240,0,36,0,204,0,0,0,0,0,106,0,165,0,44,0,0,0,252,0,9,0,207,0,0,0,75,0,0,0,0,0,0,0,154,0,41,0,10,0,69,0,209,0,243,0,0,0,200,0,176,0,141,0,38,0,64,0,106,0,169,0,0,0,161,0,51,0,171,0,0,0,0,0,0,0,0,0,133,0,153,0,161,0,0,0,170,0,0,0,0,0,238,0,125,0,251,0,0,0,209,0,149,0,103,0,132,0,177,0,0,0,140,0,0,0,14,0,50,0,51,0,141,0,0,0,173,0,14,0,0,0,225,0,162,0,0,0,166,0,156,0,90,0,205,0,0,0,0,0,242,0,0,0,72,0,207,0,231,0,141,0,80,0,207,0,165,0,18,0,204,0,101,0,0,0,0,0,0,0,123,0,0,0,0,0,24,0,0,0,227,0,120,0,225,0,0,0,0,0,233,0,0,0,0,0,0,0,0,0,232,0,19,0,202,0,130,0,73,0,107,0,0,0,141,0,2,0,0,0,215,0,0,0,130,0,118,0,88,0,0,0,63,0,183,0,41,0,237,0,21,0,190,0,124,0,119,0,39,0,73,0,132,0,161,0,243,0,124,0,58,0,144,0,138,0,31,0,0,0,235,0,79,0,181,0,59,0,197,0,0,0,173,0,66,0,60,0,148,0,0,0,139,0,72,0,250,0,119,0,0,0,167,0,192,0,24,0,171,0,0,0,11,0,72,0,120,0,37,0);
signal scenario_full  : scenario_type := (25,31,234,31,133,31,239,31,188,31,188,30,169,31,159,31,178,31,174,31,211,31,69,31,20,31,20,30,20,29,20,28,20,27,44,31,164,31,5,31,5,30,177,31,177,30,181,31,181,30,181,29,117,31,78,31,60,31,106,31,251,31,120,31,203,31,156,31,156,30,156,29,160,31,32,31,38,31,38,30,99,31,162,31,242,31,249,31,125,31,164,31,98,31,196,31,216,31,42,31,217,31,185,31,120,31,24,31,85,31,85,30,238,31,235,31,77,31,61,31,61,30,153,31,108,31,30,31,170,31,170,30,131,31,70,31,160,31,23,31,23,30,23,29,82,31,116,31,116,30,188,31,60,31,49,31,49,30,49,29,124,31,146,31,160,31,105,31,244,31,244,30,234,31,234,30,180,31,84,31,231,31,75,31,75,30,75,29,175,31,122,31,252,31,163,31,138,31,229,31,252,31,26,31,144,31,97,31,169,31,72,31,159,31,159,30,54,31,54,30,93,31,46,31,25,31,25,30,242,31,68,31,112,31,134,31,48,31,221,31,221,30,27,31,127,31,243,31,243,30,237,31,114,31,164,31,164,30,228,31,16,31,169,31,169,30,169,29,169,28,168,31,224,31,212,31,217,31,248,31,84,31,108,31,108,30,48,31,30,31,255,31,112,31,8,31,63,31,222,31,79,31,79,30,52,31,52,30,229,31,148,31,169,31,211,31,190,31,29,31,170,31,8,31,69,31,212,31,212,30,68,31,68,30,171,31,151,31,151,30,163,31,163,30,254,31,185,31,129,31,75,31,75,30,81,31,15,31,123,31,142,31,142,30,161,31,161,30,168,31,168,30,214,31,177,31,235,31,235,30,232,31,211,31,211,30,11,31,243,31,54,31,65,31,167,31,160,31,148,31,164,31,176,31,100,31,100,30,186,31,147,31,147,30,210,31,95,31,131,31,27,31,162,31,162,30,70,31,233,31,76,31,50,31,105,31,186,31,208,31,208,30,38,31,38,30,251,31,251,30,73,31,56,31,213,31,33,31,37,31,37,30,168,31,157,31,6,31,198,31,198,30,59,31,59,30,59,29,35,31,117,31,117,30,110,31,252,31,62,31,105,31,125,31,125,30,199,31,197,31,197,30,14,31,173,31,35,31,201,31,161,31,241,31,178,31,178,30,72,31,193,31,247,31,222,31,107,31,53,31,97,31,206,31,146,31,46,31,34,31,34,30,122,31,172,31,146,31,146,30,90,31,1,31,231,31,89,31,33,31,80,31,80,30,239,31,143,31,38,31,38,30,223,31,50,31,62,31,12,31,13,31,79,31,64,31,92,31,66,31,249,31,55,31,55,30,31,31,58,31,231,31,42,31,184,31,199,31,234,31,3,31,3,30,11,31,36,31,36,30,225,31,75,31,151,31,83,31,109,31,77,31,247,31,23,31,217,31,177,31,243,31,100,31,19,31,110,31,57,31,186,31,186,30,35,31,123,31,123,30,123,29,123,28,154,31,163,31,4,31,4,30,238,31,238,30,238,29,240,31,36,31,204,31,204,30,204,29,106,31,165,31,44,31,44,30,252,31,9,31,207,31,207,30,75,31,75,30,75,29,75,28,154,31,41,31,10,31,69,31,209,31,243,31,243,30,200,31,176,31,141,31,38,31,64,31,106,31,169,31,169,30,161,31,51,31,171,31,171,30,171,29,171,28,171,27,133,31,153,31,161,31,161,30,170,31,170,30,170,29,238,31,125,31,251,31,251,30,209,31,149,31,103,31,132,31,177,31,177,30,140,31,140,30,14,31,50,31,51,31,141,31,141,30,173,31,14,31,14,30,225,31,162,31,162,30,166,31,156,31,90,31,205,31,205,30,205,29,242,31,242,30,72,31,207,31,231,31,141,31,80,31,207,31,165,31,18,31,204,31,101,31,101,30,101,29,101,28,123,31,123,30,123,29,24,31,24,30,227,31,120,31,225,31,225,30,225,29,233,31,233,30,233,29,233,28,233,27,232,31,19,31,202,31,130,31,73,31,107,31,107,30,141,31,2,31,2,30,215,31,215,30,130,31,118,31,88,31,88,30,63,31,183,31,41,31,237,31,21,31,190,31,124,31,119,31,39,31,73,31,132,31,161,31,243,31,124,31,58,31,144,31,138,31,31,31,31,30,235,31,79,31,181,31,59,31,197,31,197,30,173,31,66,31,60,31,148,31,148,30,139,31,72,31,250,31,119,31,119,30,167,31,192,31,24,31,171,31,171,30,11,31,72,31,120,31,37,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
