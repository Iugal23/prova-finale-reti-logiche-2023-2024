-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 166;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,30,0,247,0,186,0,96,0,204,0,67,0,0,0,76,0,230,0,149,0,163,0,126,0,0,0,213,0,240,0,198,0,182,0,202,0,180,0,0,0,0,0,66,0,22,0,0,0,180,0,39,0,154,0,194,0,21,0,163,0,15,0,111,0,150,0,10,0,183,0,251,0,103,0,243,0,96,0,0,0,80,0,161,0,114,0,155,0,225,0,233,0,232,0,8,0,225,0,139,0,126,0,159,0,171,0,131,0,105,0,118,0,88,0,102,0,57,0,67,0,129,0,16,0,245,0,0,0,44,0,0,0,0,0,108,0,233,0,142,0,57,0,132,0,240,0,0,0,212,0,126,0,170,0,0,0,198,0,115,0,172,0,129,0,233,0,129,0,109,0,147,0,126,0,238,0,165,0,11,0,173,0,136,0,181,0,196,0,9,0,0,0,230,0,135,0,163,0,198,0,0,0,42,0,255,0,0,0,0,0,29,0,127,0,166,0,181,0,169,0,97,0,106,0,0,0,24,0,0,0,106,0,171,0,21,0,169,0,0,0,57,0,216,0,9,0,79,0,194,0,129,0,172,0,0,0,179,0,225,0,100,0,82,0,145,0,202,0,0,0,163,0,0,0,12,0,58,0,0,0,0,0,188,0,163,0,170,0,0,0,15,0,0,0,224,0,0,0,210,0,199,0,160,0,41,0,188,0,0,0,93,0,250,0,218,0,231,0,174,0,0,0,56,0,77,0,210,0,0,0);
signal scenario_full  : scenario_type := (0,0,30,31,247,31,186,31,96,31,204,31,67,31,67,30,76,31,230,31,149,31,163,31,126,31,126,30,213,31,240,31,198,31,182,31,202,31,180,31,180,30,180,29,66,31,22,31,22,30,180,31,39,31,154,31,194,31,21,31,163,31,15,31,111,31,150,31,10,31,183,31,251,31,103,31,243,31,96,31,96,30,80,31,161,31,114,31,155,31,225,31,233,31,232,31,8,31,225,31,139,31,126,31,159,31,171,31,131,31,105,31,118,31,88,31,102,31,57,31,67,31,129,31,16,31,245,31,245,30,44,31,44,30,44,29,108,31,233,31,142,31,57,31,132,31,240,31,240,30,212,31,126,31,170,31,170,30,198,31,115,31,172,31,129,31,233,31,129,31,109,31,147,31,126,31,238,31,165,31,11,31,173,31,136,31,181,31,196,31,9,31,9,30,230,31,135,31,163,31,198,31,198,30,42,31,255,31,255,30,255,29,29,31,127,31,166,31,181,31,169,31,97,31,106,31,106,30,24,31,24,30,106,31,171,31,21,31,169,31,169,30,57,31,216,31,9,31,79,31,194,31,129,31,172,31,172,30,179,31,225,31,100,31,82,31,145,31,202,31,202,30,163,31,163,30,12,31,58,31,58,30,58,29,188,31,163,31,170,31,170,30,15,31,15,30,224,31,224,30,210,31,199,31,160,31,41,31,188,31,188,30,93,31,250,31,218,31,231,31,174,31,174,30,56,31,77,31,210,31,210,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
