-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 196;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,168,0,149,0,0,0,0,0,12,0,210,0,0,0,50,0,224,0,51,0,220,0,98,0,0,0,43,0,245,0,209,0,24,0,0,0,76,0,107,0,0,0,143,0,187,0,166,0,113,0,84,0,0,0,0,0,19,0,116,0,0,0,40,0,0,0,176,0,122,0,155,0,133,0,88,0,241,0,245,0,170,0,0,0,0,0,118,0,113,0,5,0,189,0,0,0,0,0,42,0,67,0,0,0,160,0,0,0,19,0,74,0,248,0,33,0,198,0,79,0,0,0,0,0,105,0,240,0,38,0,90,0,101,0,247,0,0,0,251,0,38,0,107,0,192,0,76,0,0,0,214,0,229,0,55,0,0,0,0,0,131,0,106,0,220,0,0,0,0,0,0,0,0,0,93,0,92,0,186,0,141,0,0,0,251,0,182,0,85,0,247,0,0,0,169,0,238,0,61,0,238,0,7,0,212,0,10,0,50,0,151,0,0,0,0,0,246,0,131,0,252,0,207,0,27,0,53,0,0,0,235,0,118,0,0,0,141,0,73,0,0,0,223,0,18,0,31,0,26,0,93,0,46,0,110,0,43,0,0,0,0,0,135,0,0,0,35,0,0,0,2,0,0,0,166,0,0,0,49,0,253,0,86,0,76,0,166,0,203,0,14,0,197,0,4,0,94,0,0,0,0,0,203,0,236,0,0,0,231,0,103,0,149,0,91,0,206,0,152,0,64,0,131,0,74,0,0,0,63,0,150,0,0,0,0,0,182,0,0,0,102,0,0,0,159,0,200,0,166,0,38,0,46,0,92,0,140,0,117,0,0,0,22,0,89,0,50,0,0,0,201,0,167,0,0,0,72,0,0,0,83,0,130,0,200,0,118,0,0,0);
signal scenario_full  : scenario_type := (250,31,168,31,149,31,149,30,149,29,12,31,210,31,210,30,50,31,224,31,51,31,220,31,98,31,98,30,43,31,245,31,209,31,24,31,24,30,76,31,107,31,107,30,143,31,187,31,166,31,113,31,84,31,84,30,84,29,19,31,116,31,116,30,40,31,40,30,176,31,122,31,155,31,133,31,88,31,241,31,245,31,170,31,170,30,170,29,118,31,113,31,5,31,189,31,189,30,189,29,42,31,67,31,67,30,160,31,160,30,19,31,74,31,248,31,33,31,198,31,79,31,79,30,79,29,105,31,240,31,38,31,90,31,101,31,247,31,247,30,251,31,38,31,107,31,192,31,76,31,76,30,214,31,229,31,55,31,55,30,55,29,131,31,106,31,220,31,220,30,220,29,220,28,220,27,93,31,92,31,186,31,141,31,141,30,251,31,182,31,85,31,247,31,247,30,169,31,238,31,61,31,238,31,7,31,212,31,10,31,50,31,151,31,151,30,151,29,246,31,131,31,252,31,207,31,27,31,53,31,53,30,235,31,118,31,118,30,141,31,73,31,73,30,223,31,18,31,31,31,26,31,93,31,46,31,110,31,43,31,43,30,43,29,135,31,135,30,35,31,35,30,2,31,2,30,166,31,166,30,49,31,253,31,86,31,76,31,166,31,203,31,14,31,197,31,4,31,94,31,94,30,94,29,203,31,236,31,236,30,231,31,103,31,149,31,91,31,206,31,152,31,64,31,131,31,74,31,74,30,63,31,150,31,150,30,150,29,182,31,182,30,102,31,102,30,159,31,200,31,166,31,38,31,46,31,92,31,140,31,117,31,117,30,22,31,89,31,50,31,50,30,201,31,167,31,167,30,72,31,72,30,83,31,130,31,200,31,118,31,118,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
