-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 775;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,0,0,0,0,255,0,128,0,99,0,0,0,146,0,88,0,225,0,47,0,210,0,0,0,0,0,84,0,192,0,244,0,232,0,23,0,153,0,232,0,65,0,208,0,0,0,0,0,238,0,0,0,240,0,0,0,0,0,0,0,22,0,253,0,0,0,0,0,234,0,171,0,11,0,31,0,0,0,141,0,245,0,65,0,0,0,129,0,0,0,71,0,20,0,165,0,96,0,0,0,246,0,90,0,8,0,137,0,0,0,0,0,0,0,70,0,68,0,13,0,50,0,209,0,66,0,176,0,9,0,217,0,0,0,0,0,135,0,228,0,229,0,145,0,0,0,128,0,18,0,63,0,0,0,238,0,39,0,172,0,79,0,116,0,112,0,0,0,43,0,197,0,0,0,143,0,0,0,167,0,0,0,0,0,51,0,222,0,177,0,0,0,75,0,98,0,189,0,0,0,98,0,7,0,236,0,27,0,77,0,225,0,83,0,179,0,0,0,241,0,217,0,159,0,252,0,27,0,0,0,0,0,11,0,91,0,95,0,225,0,237,0,0,0,211,0,73,0,96,0,168,0,0,0,74,0,248,0,249,0,101,0,106,0,119,0,113,0,0,0,0,0,169,0,0,0,225,0,225,0,11,0,201,0,85,0,0,0,17,0,85,0,12,0,166,0,253,0,0,0,0,0,138,0,34,0,0,0,246,0,182,0,120,0,243,0,190,0,148,0,52,0,73,0,26,0,11,0,213,0,0,0,0,0,12,0,22,0,45,0,85,0,129,0,72,0,220,0,134,0,221,0,210,0,247,0,110,0,245,0,130,0,33,0,68,0,191,0,249,0,156,0,146,0,252,0,49,0,83,0,252,0,159,0,93,0,28,0,154,0,12,0,164,0,44,0,234,0,14,0,211,0,199,0,28,0,239,0,0,0,0,0,83,0,155,0,209,0,98,0,0,0,37,0,206,0,0,0,0,0,0,0,25,0,168,0,102,0,0,0,30,0,28,0,121,0,236,0,160,0,184,0,110,0,25,0,27,0,162,0,0,0,186,0,103,0,59,0,105,0,0,0,3,0,149,0,29,0,112,0,70,0,238,0,0,0,201,0,181,0,236,0,14,0,64,0,33,0,55,0,112,0,118,0,0,0,226,0,0,0,228,0,0,0,7,0,32,0,176,0,0,0,239,0,193,0,54,0,210,0,116,0,0,0,162,0,225,0,241,0,13,0,0,0,83,0,222,0,132,0,44,0,234,0,45,0,143,0,0,0,172,0,251,0,0,0,49,0,232,0,183,0,215,0,0,0,139,0,0,0,234,0,22,0,91,0,206,0,79,0,112,0,0,0,58,0,192,0,139,0,206,0,134,0,64,0,141,0,104,0,157,0,194,0,106,0,0,0,0,0,146,0,110,0,157,0,179,0,109,0,0,0,202,0,204,0,13,0,50,0,239,0,212,0,192,0,32,0,36,0,21,0,116,0,89,0,207,0,234,0,137,0,0,0,12,0,177,0,0,0,114,0,0,0,245,0,0,0,42,0,186,0,86,0,37,0,244,0,196,0,0,0,73,0,0,0,64,0,194,0,148,0,180,0,11,0,0,0,119,0,90,0,118,0,58,0,0,0,93,0,181,0,163,0,111,0,83,0,60,0,46,0,0,0,176,0,34,0,209,0,167,0,165,0,75,0,23,0,0,0,189,0,143,0,0,0,0,0,246,0,0,0,0,0,0,0,0,0,128,0,207,0,0,0,148,0,0,0,98,0,129,0,32,0,147,0,164,0,13,0,95,0,127,0,196,0,86,0,190,0,223,0,126,0,0,0,69,0,37,0,0,0,173,0,6,0,0,0,0,0,0,0,40,0,156,0,252,0,207,0,135,0,74,0,124,0,177,0,161,0,76,0,150,0,95,0,180,0,225,0,136,0,122,0,0,0,168,0,107,0,220,0,0,0,157,0,9,0,1,0,135,0,186,0,68,0,54,0,200,0,214,0,12,0,139,0,12,0,160,0,0,0,99,0,167,0,0,0,60,0,240,0,104,0,225,0,0,0,145,0,184,0,4,0,223,0,17,0,6,0,155,0,0,0,40,0,26,0,86,0,54,0,175,0,0,0,0,0,0,0,77,0,116,0,208,0,0,0,14,0,91,0,84,0,48,0,103,0,154,0,83,0,9,0,170,0,212,0,0,0,171,0,189,0,81,0,184,0,72,0,160,0,43,0,119,0,0,0,112,0,168,0,223,0,87,0,231,0,111,0,130,0,251,0,73,0,87,0,184,0,135,0,111,0,0,0,126,0,0,0,0,0,179,0,30,0,216,0,0,0,54,0,0,0,98,0,203,0,229,0,0,0,0,0,157,0,141,0,0,0,201,0,0,0,0,0,160,0,0,0,0,0,0,0,37,0,24,0,175,0,73,0,179,0,144,0,0,0,241,0,0,0,95,0,33,0,183,0,193,0,140,0,154,0,0,0,224,0,0,0,219,0,0,0,0,0,21,0,169,0,187,0,0,0,133,0,0,0,206,0,24,0,237,0,189,0,116,0,127,0,135,0,8,0,0,0,73,0,24,0,115,0,247,0,224,0,83,0,105,0,87,0,247,0,0,0,149,0,176,0,157,0,0,0,32,0,0,0,203,0,215,0,119,0,176,0,90,0,37,0,207,0,109,0,121,0,140,0,0,0,108,0,35,0,0,0,0,0,184,0,142,0,205,0,0,0,221,0,0,0,177,0,243,0,243,0,134,0,0,0,61,0,0,0,0,0,232,0,196,0,192,0,0,0,0,0,101,0,153,0,82,0,0,0,231,0,131,0,80,0,79,0,0,0,86,0,246,0,0,0,163,0,125,0,87,0,42,0,149,0,117,0,0,0,119,0,106,0,108,0,0,0,204,0,120,0,113,0,181,0,0,0,221,0,101,0,151,0,218,0,165,0,6,0,212,0,197,0,70,0,107,0,30,0,123,0,215,0,64,0,0,0,21,0,106,0,90,0,65,0,63,0,10,0,149,0,142,0,50,0,0,0,94,0,186,0,9,0,148,0,13,0,40,0,108,0,184,0,94,0,83,0,249,0,142,0,139,0,55,0,172,0,168,0,100,0,0,0,182,0,0,0,119,0,59,0,0,0,247,0,0,0,130,0,65,0,0,0,18,0,0,0,220,0,207,0,0,0,0,0,1,0,100,0,132,0,47,0,191,0,171,0,189,0,0,0,192,0,105,0,163,0,0,0,0,0,193,0,54,0,252,0,70,0,0,0,130,0,252,0,143,0,194,0,203,0,226,0,71,0,0,0,191,0,37,0,211,0,38,0,231,0,104,0,100,0,36,0,36,0,97,0,230,0,0,0,242,0,219,0,53,0,148,0,239,0,108,0,109,0,0,0,0,0,123,0,240,0,95,0,176,0,80,0,114,0,27,0,0,0,0,0,93,0,78,0,230,0,196,0,0,0,0,0,38,0,0,0,172,0,238,0,119,0,68,0,255,0);
signal scenario_full  : scenario_type := (95,31,95,30,95,29,255,31,128,31,99,31,99,30,146,31,88,31,225,31,47,31,210,31,210,30,210,29,84,31,192,31,244,31,232,31,23,31,153,31,232,31,65,31,208,31,208,30,208,29,238,31,238,30,240,31,240,30,240,29,240,28,22,31,253,31,253,30,253,29,234,31,171,31,11,31,31,31,31,30,141,31,245,31,65,31,65,30,129,31,129,30,71,31,20,31,165,31,96,31,96,30,246,31,90,31,8,31,137,31,137,30,137,29,137,28,70,31,68,31,13,31,50,31,209,31,66,31,176,31,9,31,217,31,217,30,217,29,135,31,228,31,229,31,145,31,145,30,128,31,18,31,63,31,63,30,238,31,39,31,172,31,79,31,116,31,112,31,112,30,43,31,197,31,197,30,143,31,143,30,167,31,167,30,167,29,51,31,222,31,177,31,177,30,75,31,98,31,189,31,189,30,98,31,7,31,236,31,27,31,77,31,225,31,83,31,179,31,179,30,241,31,217,31,159,31,252,31,27,31,27,30,27,29,11,31,91,31,95,31,225,31,237,31,237,30,211,31,73,31,96,31,168,31,168,30,74,31,248,31,249,31,101,31,106,31,119,31,113,31,113,30,113,29,169,31,169,30,225,31,225,31,11,31,201,31,85,31,85,30,17,31,85,31,12,31,166,31,253,31,253,30,253,29,138,31,34,31,34,30,246,31,182,31,120,31,243,31,190,31,148,31,52,31,73,31,26,31,11,31,213,31,213,30,213,29,12,31,22,31,45,31,85,31,129,31,72,31,220,31,134,31,221,31,210,31,247,31,110,31,245,31,130,31,33,31,68,31,191,31,249,31,156,31,146,31,252,31,49,31,83,31,252,31,159,31,93,31,28,31,154,31,12,31,164,31,44,31,234,31,14,31,211,31,199,31,28,31,239,31,239,30,239,29,83,31,155,31,209,31,98,31,98,30,37,31,206,31,206,30,206,29,206,28,25,31,168,31,102,31,102,30,30,31,28,31,121,31,236,31,160,31,184,31,110,31,25,31,27,31,162,31,162,30,186,31,103,31,59,31,105,31,105,30,3,31,149,31,29,31,112,31,70,31,238,31,238,30,201,31,181,31,236,31,14,31,64,31,33,31,55,31,112,31,118,31,118,30,226,31,226,30,228,31,228,30,7,31,32,31,176,31,176,30,239,31,193,31,54,31,210,31,116,31,116,30,162,31,225,31,241,31,13,31,13,30,83,31,222,31,132,31,44,31,234,31,45,31,143,31,143,30,172,31,251,31,251,30,49,31,232,31,183,31,215,31,215,30,139,31,139,30,234,31,22,31,91,31,206,31,79,31,112,31,112,30,58,31,192,31,139,31,206,31,134,31,64,31,141,31,104,31,157,31,194,31,106,31,106,30,106,29,146,31,110,31,157,31,179,31,109,31,109,30,202,31,204,31,13,31,50,31,239,31,212,31,192,31,32,31,36,31,21,31,116,31,89,31,207,31,234,31,137,31,137,30,12,31,177,31,177,30,114,31,114,30,245,31,245,30,42,31,186,31,86,31,37,31,244,31,196,31,196,30,73,31,73,30,64,31,194,31,148,31,180,31,11,31,11,30,119,31,90,31,118,31,58,31,58,30,93,31,181,31,163,31,111,31,83,31,60,31,46,31,46,30,176,31,34,31,209,31,167,31,165,31,75,31,23,31,23,30,189,31,143,31,143,30,143,29,246,31,246,30,246,29,246,28,246,27,128,31,207,31,207,30,148,31,148,30,98,31,129,31,32,31,147,31,164,31,13,31,95,31,127,31,196,31,86,31,190,31,223,31,126,31,126,30,69,31,37,31,37,30,173,31,6,31,6,30,6,29,6,28,40,31,156,31,252,31,207,31,135,31,74,31,124,31,177,31,161,31,76,31,150,31,95,31,180,31,225,31,136,31,122,31,122,30,168,31,107,31,220,31,220,30,157,31,9,31,1,31,135,31,186,31,68,31,54,31,200,31,214,31,12,31,139,31,12,31,160,31,160,30,99,31,167,31,167,30,60,31,240,31,104,31,225,31,225,30,145,31,184,31,4,31,223,31,17,31,6,31,155,31,155,30,40,31,26,31,86,31,54,31,175,31,175,30,175,29,175,28,77,31,116,31,208,31,208,30,14,31,91,31,84,31,48,31,103,31,154,31,83,31,9,31,170,31,212,31,212,30,171,31,189,31,81,31,184,31,72,31,160,31,43,31,119,31,119,30,112,31,168,31,223,31,87,31,231,31,111,31,130,31,251,31,73,31,87,31,184,31,135,31,111,31,111,30,126,31,126,30,126,29,179,31,30,31,216,31,216,30,54,31,54,30,98,31,203,31,229,31,229,30,229,29,157,31,141,31,141,30,201,31,201,30,201,29,160,31,160,30,160,29,160,28,37,31,24,31,175,31,73,31,179,31,144,31,144,30,241,31,241,30,95,31,33,31,183,31,193,31,140,31,154,31,154,30,224,31,224,30,219,31,219,30,219,29,21,31,169,31,187,31,187,30,133,31,133,30,206,31,24,31,237,31,189,31,116,31,127,31,135,31,8,31,8,30,73,31,24,31,115,31,247,31,224,31,83,31,105,31,87,31,247,31,247,30,149,31,176,31,157,31,157,30,32,31,32,30,203,31,215,31,119,31,176,31,90,31,37,31,207,31,109,31,121,31,140,31,140,30,108,31,35,31,35,30,35,29,184,31,142,31,205,31,205,30,221,31,221,30,177,31,243,31,243,31,134,31,134,30,61,31,61,30,61,29,232,31,196,31,192,31,192,30,192,29,101,31,153,31,82,31,82,30,231,31,131,31,80,31,79,31,79,30,86,31,246,31,246,30,163,31,125,31,87,31,42,31,149,31,117,31,117,30,119,31,106,31,108,31,108,30,204,31,120,31,113,31,181,31,181,30,221,31,101,31,151,31,218,31,165,31,6,31,212,31,197,31,70,31,107,31,30,31,123,31,215,31,64,31,64,30,21,31,106,31,90,31,65,31,63,31,10,31,149,31,142,31,50,31,50,30,94,31,186,31,9,31,148,31,13,31,40,31,108,31,184,31,94,31,83,31,249,31,142,31,139,31,55,31,172,31,168,31,100,31,100,30,182,31,182,30,119,31,59,31,59,30,247,31,247,30,130,31,65,31,65,30,18,31,18,30,220,31,207,31,207,30,207,29,1,31,100,31,132,31,47,31,191,31,171,31,189,31,189,30,192,31,105,31,163,31,163,30,163,29,193,31,54,31,252,31,70,31,70,30,130,31,252,31,143,31,194,31,203,31,226,31,71,31,71,30,191,31,37,31,211,31,38,31,231,31,104,31,100,31,36,31,36,31,97,31,230,31,230,30,242,31,219,31,53,31,148,31,239,31,108,31,109,31,109,30,109,29,123,31,240,31,95,31,176,31,80,31,114,31,27,31,27,30,27,29,93,31,78,31,230,31,196,31,196,30,196,29,38,31,38,30,172,31,238,31,119,31,68,31,255,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
