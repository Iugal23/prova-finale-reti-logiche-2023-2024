-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (108,0,164,0,245,0,8,0,0,0,0,0,37,0,45,0,0,0,156,0,166,0,107,0,83,0,208,0,0,0,250,0,42,0,25,0,0,0,11,0,171,0,85,0,158,0,118,0,146,0,186,0,162,0,106,0,0,0,0,0,184,0,61,0,223,0,132,0,157,0,180,0,41,0,230,0,172,0,71,0,74,0,221,0,27,0,189,0,58,0,162,0,0,0,27,0,39,0,244,0,0,0,0,0,157,0,82,0,0,0,38,0,173,0,131,0,223,0,241,0,0,0,0,0,167,0,162,0,133,0,123,0,176,0,0,0,163,0,231,0,69,0,139,0,28,0,137,0,87,0,217,0,167,0,0,0,219,0,195,0,95,0,242,0,220,0,23,0,36,0,130,0,29,0,149,0,171,0,128,0,229,0,32,0,250,0,133,0,0,0,211,0,119,0,99,0,233,0,252,0,33,0,59,0,0,0,233,0,198,0,95,0,111,0,41,0,0,0,106,0,0,0,68,0,53,0,144,0,193,0,110,0,99,0,58,0,145,0,175,0,94,0,46,0,194,0,130,0,0,0,159,0,220,0,102,0,241,0,0,0,0,0,77,0,98,0,155,0,0,0,224,0,14,0,56,0,200,0,185,0,181,0,107,0,202,0,0,0,0,0,71,0,36,0,0,0,241,0,0,0,0,0,116,0,159,0,189,0,0,0,194,0,194,0,14,0,148,0,130,0,225,0,200,0,158,0,0,0,216,0,150,0,20,0,203,0,0,0,105,0,41,0,18,0,107,0,53,0,189,0,13,0,10,0,182,0,76,0,134,0,190,0,79,0,0,0,197,0,138,0,40,0,97,0,182,0,0,0,207,0,169,0,20,0,50,0,242,0,44,0,214,0,14,0,60,0,96,0,129,0,32,0,75,0,144,0,173,0,0,0,0,0,160,0,93,0,11,0,6,0,73,0,81,0,199,0,227,0,114,0,0,0,0,0,138,0,35,0,138,0,185,0,116,0,150,0,49,0,253,0,254,0,0,0,75,0,6,0,66,0,109,0,18,0,197,0,227,0,209,0,122,0,168,0,0,0,48,0,0,0,0,0,152,0,89,0,0,0,0,0,212,0,221,0,191,0,42,0,45,0,3,0,126,0,67,0,130,0,0,0,205,0,133,0,168,0,0,0,20,0,134,0,125,0,231,0,244,0,193,0,31,0,229,0,0,0,115,0,180,0,0,0,0,0,0,0,39,0,111,0,238,0,176,0,45,0,233,0,123,0,153,0,0,0,0,0,51,0,56,0,169,0,237,0,117,0,229,0,0,0,150,0,132,0,96,0,182,0,0,0,162,0,241,0,192,0,216,0,54,0,166,0,129,0,182,0,21,0,156,0,119,0,0,0,33,0,0,0,211,0,137,0,207,0,18,0,129,0,156,0,36,0,111,0,170,0,134,0,0,0,0,0,181,0,225,0,64,0,0,0,0,0,0,0,48,0,247,0,27,0,37,0,63,0,24,0,167,0,235,0,141,0,171,0,148,0,0,0,159,0,82,0,125,0,0,0,0,0,217,0,212,0,95,0,0,0,228,0,213,0,122,0,102,0,125,0,224,0,178,0,8,0,41,0,144,0,35,0,198,0,25,0,244,0,3,0,37,0,231,0,68,0,0,0,205,0,117,0,24,0,117,0,0,0,182,0,245,0,0,0,145,0,0,0,217,0,100,0,181,0,148,0,97,0,254,0,252,0,126,0,74,0,242,0,200,0,43,0,25,0,229,0,126,0,153,0,198,0,209,0,192,0,236,0,218,0,11,0,125,0,115,0,221,0,210,0,0,0,108,0,0,0,45,0,197,0,0,0,241,0,0,0,28,0,202,0,0,0,170,0,114,0,165,0,0,0,147,0,23,0,107,0,0,0,106,0,0,0,121,0,0,0,246,0,108,0,0,0,230,0,100,0,194,0,0,0,232,0,0,0,114,0,77,0,55,0,221,0,0,0,108,0,52,0,112,0,119,0,211,0,0,0,183,0,27,0,0,0,32,0,13,0,0,0,192,0,0,0,22,0,0,0,64,0,137,0,39,0,141,0,222,0,3,0,0,0,180,0,0,0,77,0,0,0,7,0,250,0,244,0,170,0,13,0,65,0,255,0,222,0,0,0,65,0,0,0,0,0,68,0,67,0,227,0,0,0,59,0,82,0,99,0,0,0,76,0,156,0,200,0,91,0,0,0,181,0,196,0,81,0,0,0,25,0,0,0,38,0,198,0,101,0,228,0,107,0,17,0,160,0,242,0,126,0,176,0,41,0,23,0,0,0,27,0,33,0,56,0,0,0,97,0,0,0,0,0,5,0,168,0,150,0,77,0,0,0,221,0,0,0,245,0,219,0,0,0,162,0,232,0,189,0,0,0,219,0,30,0,6,0,222,0,25,0,211,0,188,0,0,0,0,0,161,0,124,0,238,0,76,0,215,0,238,0,234,0,213,0,232,0,63,0,0,0,142,0,153,0,190,0,129,0,71,0,0,0,61,0,197,0,86,0,180,0,158,0,96,0,234,0,229,0,0,0,208,0,138,0,19,0,0,0,70,0,62,0,217,0,23,0,254,0,123,0,144,0,0,0,133,0,0,0,0,0,214,0,148,0,70,0,204,0,206,0,208,0,248,0,71,0,85,0,249,0,212,0,10,0,180,0,188,0,245,0,135,0,77,0,231,0,4,0,0,0,95,0,22,0,200,0,42,0,236,0,190,0,128,0,180,0,175,0,209,0,84,0,28,0,134,0,122,0,168,0,207,0,253,0,0,0,192,0,129,0,113,0,200,0,45,0,65,0,212,0,128,0,1,0,216,0,57,0,0,0,20,0,175,0,89,0,52,0,174,0,24,0,192,0,84,0,103,0,37,0,0,0,37,0,163,0,253,0,45,0,180,0,27,0,0,0,247,0,35,0,109,0,25,0,252,0,4,0,128,0,0,0,0,0,178,0,154,0,100,0,138,0,204,0,15,0,240,0,0,0,221,0,215,0,201,0,39,0,212,0,0,0,77,0,219,0,23,0,0,0,66,0,174,0,145,0,0,0,0,0,0,0,123,0,0,0,55,0,224,0,119,0,222,0,111,0,129,0,225,0,240,0,41,0,123,0,251,0,94,0,142,0,244,0,213,0,122,0,218,0,102,0,142,0,14,0,115,0,0,0,223,0,165,0,9,0,62,0,0,0,58,0,0,0,76,0,0,0,200,0,159,0,20,0,0,0,72,0,0,0,248,0,234,0,134,0,15,0,164,0,0,0,193,0,169,0,115,0,213,0,91,0,239,0,9,0,104,0,36,0,180,0,218,0,0,0,236,0,0,0,213,0,163,0,0,0,236,0,192,0,107,0,28,0,245,0,0,0,215,0,33,0,47,0,65,0,18,0,26,0,75,0,142,0,58,0,0,0,0,0,78,0,253,0,0,0,196,0,0,0,128,0,0,0,52,0,15,0,43,0,142,0,72,0,0,0,88,0,103,0,0,0,0,0,66,0,69,0,25,0,0,0,0,0,134,0,66,0,138,0,42,0,94,0,0,0,0,0,39,0,137,0,86,0,124,0,70,0,33,0,0,0,175,0,109,0,123,0,32,0,144,0,0,0,250,0,0,0,0,0,90,0,40,0,0,0,211,0,22,0,0,0,0,0,140,0,63,0,2,0,199,0,205,0,0,0,0,0,39,0,12,0,2,0,106,0,0,0,69,0,10,0,197,0,7,0,0,0,185,0,0,0,218,0,0,0,0,0,132,0,115,0,255,0,24,0,0,0,0,0,25,0,54,0,221,0,0,0,0,0,99,0,6,0,73,0,57,0,176,0,150,0,137,0,135,0,27,0,226,0);
signal scenario_full  : scenario_type := (108,31,164,31,245,31,8,31,8,30,8,29,37,31,45,31,45,30,156,31,166,31,107,31,83,31,208,31,208,30,250,31,42,31,25,31,25,30,11,31,171,31,85,31,158,31,118,31,146,31,186,31,162,31,106,31,106,30,106,29,184,31,61,31,223,31,132,31,157,31,180,31,41,31,230,31,172,31,71,31,74,31,221,31,27,31,189,31,58,31,162,31,162,30,27,31,39,31,244,31,244,30,244,29,157,31,82,31,82,30,38,31,173,31,131,31,223,31,241,31,241,30,241,29,167,31,162,31,133,31,123,31,176,31,176,30,163,31,231,31,69,31,139,31,28,31,137,31,87,31,217,31,167,31,167,30,219,31,195,31,95,31,242,31,220,31,23,31,36,31,130,31,29,31,149,31,171,31,128,31,229,31,32,31,250,31,133,31,133,30,211,31,119,31,99,31,233,31,252,31,33,31,59,31,59,30,233,31,198,31,95,31,111,31,41,31,41,30,106,31,106,30,68,31,53,31,144,31,193,31,110,31,99,31,58,31,145,31,175,31,94,31,46,31,194,31,130,31,130,30,159,31,220,31,102,31,241,31,241,30,241,29,77,31,98,31,155,31,155,30,224,31,14,31,56,31,200,31,185,31,181,31,107,31,202,31,202,30,202,29,71,31,36,31,36,30,241,31,241,30,241,29,116,31,159,31,189,31,189,30,194,31,194,31,14,31,148,31,130,31,225,31,200,31,158,31,158,30,216,31,150,31,20,31,203,31,203,30,105,31,41,31,18,31,107,31,53,31,189,31,13,31,10,31,182,31,76,31,134,31,190,31,79,31,79,30,197,31,138,31,40,31,97,31,182,31,182,30,207,31,169,31,20,31,50,31,242,31,44,31,214,31,14,31,60,31,96,31,129,31,32,31,75,31,144,31,173,31,173,30,173,29,160,31,93,31,11,31,6,31,73,31,81,31,199,31,227,31,114,31,114,30,114,29,138,31,35,31,138,31,185,31,116,31,150,31,49,31,253,31,254,31,254,30,75,31,6,31,66,31,109,31,18,31,197,31,227,31,209,31,122,31,168,31,168,30,48,31,48,30,48,29,152,31,89,31,89,30,89,29,212,31,221,31,191,31,42,31,45,31,3,31,126,31,67,31,130,31,130,30,205,31,133,31,168,31,168,30,20,31,134,31,125,31,231,31,244,31,193,31,31,31,229,31,229,30,115,31,180,31,180,30,180,29,180,28,39,31,111,31,238,31,176,31,45,31,233,31,123,31,153,31,153,30,153,29,51,31,56,31,169,31,237,31,117,31,229,31,229,30,150,31,132,31,96,31,182,31,182,30,162,31,241,31,192,31,216,31,54,31,166,31,129,31,182,31,21,31,156,31,119,31,119,30,33,31,33,30,211,31,137,31,207,31,18,31,129,31,156,31,36,31,111,31,170,31,134,31,134,30,134,29,181,31,225,31,64,31,64,30,64,29,64,28,48,31,247,31,27,31,37,31,63,31,24,31,167,31,235,31,141,31,171,31,148,31,148,30,159,31,82,31,125,31,125,30,125,29,217,31,212,31,95,31,95,30,228,31,213,31,122,31,102,31,125,31,224,31,178,31,8,31,41,31,144,31,35,31,198,31,25,31,244,31,3,31,37,31,231,31,68,31,68,30,205,31,117,31,24,31,117,31,117,30,182,31,245,31,245,30,145,31,145,30,217,31,100,31,181,31,148,31,97,31,254,31,252,31,126,31,74,31,242,31,200,31,43,31,25,31,229,31,126,31,153,31,198,31,209,31,192,31,236,31,218,31,11,31,125,31,115,31,221,31,210,31,210,30,108,31,108,30,45,31,197,31,197,30,241,31,241,30,28,31,202,31,202,30,170,31,114,31,165,31,165,30,147,31,23,31,107,31,107,30,106,31,106,30,121,31,121,30,246,31,108,31,108,30,230,31,100,31,194,31,194,30,232,31,232,30,114,31,77,31,55,31,221,31,221,30,108,31,52,31,112,31,119,31,211,31,211,30,183,31,27,31,27,30,32,31,13,31,13,30,192,31,192,30,22,31,22,30,64,31,137,31,39,31,141,31,222,31,3,31,3,30,180,31,180,30,77,31,77,30,7,31,250,31,244,31,170,31,13,31,65,31,255,31,222,31,222,30,65,31,65,30,65,29,68,31,67,31,227,31,227,30,59,31,82,31,99,31,99,30,76,31,156,31,200,31,91,31,91,30,181,31,196,31,81,31,81,30,25,31,25,30,38,31,198,31,101,31,228,31,107,31,17,31,160,31,242,31,126,31,176,31,41,31,23,31,23,30,27,31,33,31,56,31,56,30,97,31,97,30,97,29,5,31,168,31,150,31,77,31,77,30,221,31,221,30,245,31,219,31,219,30,162,31,232,31,189,31,189,30,219,31,30,31,6,31,222,31,25,31,211,31,188,31,188,30,188,29,161,31,124,31,238,31,76,31,215,31,238,31,234,31,213,31,232,31,63,31,63,30,142,31,153,31,190,31,129,31,71,31,71,30,61,31,197,31,86,31,180,31,158,31,96,31,234,31,229,31,229,30,208,31,138,31,19,31,19,30,70,31,62,31,217,31,23,31,254,31,123,31,144,31,144,30,133,31,133,30,133,29,214,31,148,31,70,31,204,31,206,31,208,31,248,31,71,31,85,31,249,31,212,31,10,31,180,31,188,31,245,31,135,31,77,31,231,31,4,31,4,30,95,31,22,31,200,31,42,31,236,31,190,31,128,31,180,31,175,31,209,31,84,31,28,31,134,31,122,31,168,31,207,31,253,31,253,30,192,31,129,31,113,31,200,31,45,31,65,31,212,31,128,31,1,31,216,31,57,31,57,30,20,31,175,31,89,31,52,31,174,31,24,31,192,31,84,31,103,31,37,31,37,30,37,31,163,31,253,31,45,31,180,31,27,31,27,30,247,31,35,31,109,31,25,31,252,31,4,31,128,31,128,30,128,29,178,31,154,31,100,31,138,31,204,31,15,31,240,31,240,30,221,31,215,31,201,31,39,31,212,31,212,30,77,31,219,31,23,31,23,30,66,31,174,31,145,31,145,30,145,29,145,28,123,31,123,30,55,31,224,31,119,31,222,31,111,31,129,31,225,31,240,31,41,31,123,31,251,31,94,31,142,31,244,31,213,31,122,31,218,31,102,31,142,31,14,31,115,31,115,30,223,31,165,31,9,31,62,31,62,30,58,31,58,30,76,31,76,30,200,31,159,31,20,31,20,30,72,31,72,30,248,31,234,31,134,31,15,31,164,31,164,30,193,31,169,31,115,31,213,31,91,31,239,31,9,31,104,31,36,31,180,31,218,31,218,30,236,31,236,30,213,31,163,31,163,30,236,31,192,31,107,31,28,31,245,31,245,30,215,31,33,31,47,31,65,31,18,31,26,31,75,31,142,31,58,31,58,30,58,29,78,31,253,31,253,30,196,31,196,30,128,31,128,30,52,31,15,31,43,31,142,31,72,31,72,30,88,31,103,31,103,30,103,29,66,31,69,31,25,31,25,30,25,29,134,31,66,31,138,31,42,31,94,31,94,30,94,29,39,31,137,31,86,31,124,31,70,31,33,31,33,30,175,31,109,31,123,31,32,31,144,31,144,30,250,31,250,30,250,29,90,31,40,31,40,30,211,31,22,31,22,30,22,29,140,31,63,31,2,31,199,31,205,31,205,30,205,29,39,31,12,31,2,31,106,31,106,30,69,31,10,31,197,31,7,31,7,30,185,31,185,30,218,31,218,30,218,29,132,31,115,31,255,31,24,31,24,30,24,29,25,31,54,31,221,31,221,30,221,29,99,31,6,31,73,31,57,31,176,31,150,31,137,31,135,31,27,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
