-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 837;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (104,0,114,0,0,0,0,0,236,0,177,0,109,0,7,0,255,0,127,0,10,0,156,0,161,0,232,0,31,0,37,0,128,0,234,0,18,0,0,0,102,0,54,0,0,0,34,0,19,0,186,0,0,0,129,0,130,0,103,0,131,0,177,0,144,0,51,0,217,0,19,0,0,0,242,0,122,0,196,0,165,0,157,0,140,0,78,0,89,0,0,0,7,0,179,0,248,0,33,0,206,0,0,0,180,0,250,0,66,0,0,0,0,0,167,0,0,0,0,0,207,0,0,0,34,0,110,0,218,0,218,0,14,0,0,0,0,0,219,0,0,0,100,0,188,0,0,0,210,0,110,0,182,0,75,0,146,0,0,0,0,0,0,0,159,0,135,0,83,0,0,0,240,0,250,0,113,0,92,0,56,0,107,0,0,0,107,0,246,0,100,0,0,0,0,0,156,0,5,0,153,0,248,0,181,0,0,0,179,0,69,0,127,0,160,0,244,0,0,0,203,0,37,0,198,0,49,0,89,0,143,0,74,0,183,0,56,0,0,0,173,0,244,0,0,0,230,0,229,0,214,0,233,0,78,0,167,0,203,0,64,0,0,0,142,0,139,0,220,0,0,0,167,0,23,0,39,0,0,0,38,0,179,0,0,0,227,0,90,0,182,0,64,0,122,0,104,0,178,0,0,0,103,0,0,0,83,0,122,0,165,0,80,0,239,0,216,0,100,0,206,0,97,0,240,0,172,0,231,0,6,0,0,0,34,0,0,0,0,0,218,0,163,0,0,0,131,0,0,0,249,0,56,0,0,0,10,0,64,0,142,0,11,0,129,0,77,0,63,0,111,0,110,0,0,0,249,0,100,0,139,0,204,0,209,0,0,0,251,0,79,0,103,0,82,0,0,0,171,0,203,0,99,0,84,0,217,0,13,0,66,0,89,0,201,0,162,0,184,0,230,0,45,0,116,0,1,0,166,0,61,0,103,0,239,0,0,0,173,0,198,0,158,0,0,0,173,0,178,0,152,0,219,0,78,0,178,0,249,0,151,0,0,0,53,0,6,0,16,0,99,0,214,0,0,0,85,0,0,0,130,0,0,0,199,0,47,0,209,0,0,0,186,0,50,0,163,0,39,0,175,0,55,0,1,0,134,0,80,0,178,0,19,0,104,0,79,0,212,0,205,0,0,0,140,0,0,0,191,0,151,0,0,0,52,0,128,0,133,0,0,0,0,0,48,0,156,0,79,0,137,0,98,0,0,0,12,0,106,0,0,0,139,0,92,0,16,0,103,0,0,0,246,0,123,0,247,0,151,0,0,0,134,0,62,0,79,0,0,0,0,0,25,0,166,0,117,0,54,0,8,0,0,0,83,0,202,0,167,0,225,0,0,0,100,0,129,0,93,0,151,0,61,0,44,0,182,0,218,0,238,0,80,0,191,0,18,0,0,0,0,0,56,0,0,0,136,0,27,0,21,0,68,0,0,0,205,0,4,0,61,0,200,0,224,0,239,0,204,0,128,0,127,0,112,0,0,0,6,0,153,0,166,0,24,0,120,0,246,0,128,0,213,0,237,0,154,0,194,0,225,0,200,0,139,0,185,0,201,0,48,0,245,0,125,0,0,0,0,0,0,0,58,0,161,0,85,0,243,0,118,0,0,0,130,0,4,0,0,0,193,0,0,0,191,0,37,0,0,0,255,0,57,0,146,0,0,0,151,0,173,0,7,0,0,0,110,0,175,0,0,0,36,0,0,0,9,0,246,0,233,0,0,0,94,0,109,0,0,0,128,0,5,0,0,0,0,0,11,0,14,0,85,0,198,0,0,0,32,0,143,0,69,0,75,0,25,0,69,0,156,0,137,0,225,0,153,0,0,0,132,0,0,0,67,0,16,0,155,0,12,0,72,0,241,0,134,0,163,0,50,0,123,0,54,0,91,0,18,0,0,0,178,0,228,0,104,0,0,0,26,0,152,0,198,0,232,0,50,0,130,0,0,0,0,0,172,0,0,0,242,0,10,0,0,0,0,0,25,0,136,0,66,0,246,0,150,0,97,0,125,0,235,0,15,0,220,0,14,0,230,0,66,0,52,0,17,0,203,0,21,0,52,0,94,0,30,0,0,0,38,0,228,0,162,0,0,0,114,0,85,0,0,0,176,0,49,0,232,0,140,0,34,0,83,0,221,0,67,0,0,0,30,0,37,0,0,0,11,0,84,0,57,0,0,0,136,0,45,0,155,0,1,0,211,0,0,0,69,0,15,0,68,0,0,0,211,0,173,0,201,0,0,0,66,0,185,0,114,0,212,0,24,0,74,0,18,0,217,0,0,0,29,0,0,0,0,0,121,0,215,0,249,0,217,0,128,0,16,0,199,0,0,0,188,0,139,0,142,0,39,0,176,0,65,0,159,0,152,0,91,0,68,0,0,0,176,0,6,0,61,0,163,0,197,0,11,0,239,0,133,0,86,0,138,0,0,0,41,0,99,0,120,0,0,0,238,0,132,0,136,0,42,0,0,0,0,0,184,0,155,0,14,0,111,0,211,0,53,0,33,0,0,0,36,0,0,0,0,0,0,0,0,0,141,0,124,0,0,0,0,0,68,0,15,0,248,0,143,0,204,0,143,0,129,0,94,0,111,0,18,0,123,0,228,0,109,0,235,0,7,0,72,0,41,0,112,0,164,0,74,0,54,0,0,0,165,0,0,0,37,0,0,0,124,0,0,0,220,0,96,0,208,0,0,0,183,0,133,0,0,0,248,0,175,0,6,0,222,0,43,0,7,0,0,0,0,0,244,0,97,0,253,0,69,0,130,0,234,0,0,0,63,0,181,0,34,0,71,0,173,0,64,0,0,0,0,0,169,0,5,0,249,0,224,0,224,0,248,0,254,0,0,0,61,0,166,0,30,0,254,0,51,0,56,0,39,0,52,0,143,0,0,0,61,0,9,0,168,0,69,0,187,0,91,0,38,0,105,0,0,0,218,0,0,0,116,0,219,0,179,0,97,0,158,0,118,0,76,0,0,0,149,0,6,0,0,0,60,0,62,0,169,0,134,0,170,0,0,0,66,0,205,0,156,0,44,0,108,0,37,0,88,0,180,0,104,0,167,0,16,0,2,0,127,0,156,0,92,0,0,0,255,0,220,0,0,0,72,0,157,0,132,0,0,0,191,0,77,0,130,0,0,0,29,0,171,0,112,0,110,0,84,0,65,0,0,0,251,0,165,0,69,0,41,0,0,0,210,0,189,0,0,0,57,0,181,0,83,0,123,0,0,0,221,0,200,0,77,0,52,0,205,0,181,0,50,0,145,0,108,0,76,0,164,0,6,0,165,0,0,0,27,0,56,0,77,0,8,0,0,0,130,0,157,0,8,0,159,0,186,0,11,0,238,0,212,0,179,0,188,0,0,0,91,0,221,0,60,0,0,0,172,0,60,0,205,0,68,0,91,0,172,0,193,0,216,0,40,0,169,0,81,0,242,0,244,0,214,0,0,0,114,0,218,0,243,0,208,0,14,0,97,0,208,0,242,0,0,0,0,0,167,0,87,0,185,0,248,0,44,0,236,0,168,0,0,0,33,0,244,0,0,0,0,0,184,0,225,0,228,0,20,0,0,0,66,0,211,0,115,0,206,0,15,0,61,0,118,0,56,0,18,0,16,0,139,0,227,0,0,0,0,0,82,0,0,0,72,0,231,0,48,0,205,0,143,0,178,0,221,0,217,0,201,0,104,0,240,0,72,0,20,0,70,0,0,0,241,0,206,0,102,0);
signal scenario_full  : scenario_type := (104,31,114,31,114,30,114,29,236,31,177,31,109,31,7,31,255,31,127,31,10,31,156,31,161,31,232,31,31,31,37,31,128,31,234,31,18,31,18,30,102,31,54,31,54,30,34,31,19,31,186,31,186,30,129,31,130,31,103,31,131,31,177,31,144,31,51,31,217,31,19,31,19,30,242,31,122,31,196,31,165,31,157,31,140,31,78,31,89,31,89,30,7,31,179,31,248,31,33,31,206,31,206,30,180,31,250,31,66,31,66,30,66,29,167,31,167,30,167,29,207,31,207,30,34,31,110,31,218,31,218,31,14,31,14,30,14,29,219,31,219,30,100,31,188,31,188,30,210,31,110,31,182,31,75,31,146,31,146,30,146,29,146,28,159,31,135,31,83,31,83,30,240,31,250,31,113,31,92,31,56,31,107,31,107,30,107,31,246,31,100,31,100,30,100,29,156,31,5,31,153,31,248,31,181,31,181,30,179,31,69,31,127,31,160,31,244,31,244,30,203,31,37,31,198,31,49,31,89,31,143,31,74,31,183,31,56,31,56,30,173,31,244,31,244,30,230,31,229,31,214,31,233,31,78,31,167,31,203,31,64,31,64,30,142,31,139,31,220,31,220,30,167,31,23,31,39,31,39,30,38,31,179,31,179,30,227,31,90,31,182,31,64,31,122,31,104,31,178,31,178,30,103,31,103,30,83,31,122,31,165,31,80,31,239,31,216,31,100,31,206,31,97,31,240,31,172,31,231,31,6,31,6,30,34,31,34,30,34,29,218,31,163,31,163,30,131,31,131,30,249,31,56,31,56,30,10,31,64,31,142,31,11,31,129,31,77,31,63,31,111,31,110,31,110,30,249,31,100,31,139,31,204,31,209,31,209,30,251,31,79,31,103,31,82,31,82,30,171,31,203,31,99,31,84,31,217,31,13,31,66,31,89,31,201,31,162,31,184,31,230,31,45,31,116,31,1,31,166,31,61,31,103,31,239,31,239,30,173,31,198,31,158,31,158,30,173,31,178,31,152,31,219,31,78,31,178,31,249,31,151,31,151,30,53,31,6,31,16,31,99,31,214,31,214,30,85,31,85,30,130,31,130,30,199,31,47,31,209,31,209,30,186,31,50,31,163,31,39,31,175,31,55,31,1,31,134,31,80,31,178,31,19,31,104,31,79,31,212,31,205,31,205,30,140,31,140,30,191,31,151,31,151,30,52,31,128,31,133,31,133,30,133,29,48,31,156,31,79,31,137,31,98,31,98,30,12,31,106,31,106,30,139,31,92,31,16,31,103,31,103,30,246,31,123,31,247,31,151,31,151,30,134,31,62,31,79,31,79,30,79,29,25,31,166,31,117,31,54,31,8,31,8,30,83,31,202,31,167,31,225,31,225,30,100,31,129,31,93,31,151,31,61,31,44,31,182,31,218,31,238,31,80,31,191,31,18,31,18,30,18,29,56,31,56,30,136,31,27,31,21,31,68,31,68,30,205,31,4,31,61,31,200,31,224,31,239,31,204,31,128,31,127,31,112,31,112,30,6,31,153,31,166,31,24,31,120,31,246,31,128,31,213,31,237,31,154,31,194,31,225,31,200,31,139,31,185,31,201,31,48,31,245,31,125,31,125,30,125,29,125,28,58,31,161,31,85,31,243,31,118,31,118,30,130,31,4,31,4,30,193,31,193,30,191,31,37,31,37,30,255,31,57,31,146,31,146,30,151,31,173,31,7,31,7,30,110,31,175,31,175,30,36,31,36,30,9,31,246,31,233,31,233,30,94,31,109,31,109,30,128,31,5,31,5,30,5,29,11,31,14,31,85,31,198,31,198,30,32,31,143,31,69,31,75,31,25,31,69,31,156,31,137,31,225,31,153,31,153,30,132,31,132,30,67,31,16,31,155,31,12,31,72,31,241,31,134,31,163,31,50,31,123,31,54,31,91,31,18,31,18,30,178,31,228,31,104,31,104,30,26,31,152,31,198,31,232,31,50,31,130,31,130,30,130,29,172,31,172,30,242,31,10,31,10,30,10,29,25,31,136,31,66,31,246,31,150,31,97,31,125,31,235,31,15,31,220,31,14,31,230,31,66,31,52,31,17,31,203,31,21,31,52,31,94,31,30,31,30,30,38,31,228,31,162,31,162,30,114,31,85,31,85,30,176,31,49,31,232,31,140,31,34,31,83,31,221,31,67,31,67,30,30,31,37,31,37,30,11,31,84,31,57,31,57,30,136,31,45,31,155,31,1,31,211,31,211,30,69,31,15,31,68,31,68,30,211,31,173,31,201,31,201,30,66,31,185,31,114,31,212,31,24,31,74,31,18,31,217,31,217,30,29,31,29,30,29,29,121,31,215,31,249,31,217,31,128,31,16,31,199,31,199,30,188,31,139,31,142,31,39,31,176,31,65,31,159,31,152,31,91,31,68,31,68,30,176,31,6,31,61,31,163,31,197,31,11,31,239,31,133,31,86,31,138,31,138,30,41,31,99,31,120,31,120,30,238,31,132,31,136,31,42,31,42,30,42,29,184,31,155,31,14,31,111,31,211,31,53,31,33,31,33,30,36,31,36,30,36,29,36,28,36,27,141,31,124,31,124,30,124,29,68,31,15,31,248,31,143,31,204,31,143,31,129,31,94,31,111,31,18,31,123,31,228,31,109,31,235,31,7,31,72,31,41,31,112,31,164,31,74,31,54,31,54,30,165,31,165,30,37,31,37,30,124,31,124,30,220,31,96,31,208,31,208,30,183,31,133,31,133,30,248,31,175,31,6,31,222,31,43,31,7,31,7,30,7,29,244,31,97,31,253,31,69,31,130,31,234,31,234,30,63,31,181,31,34,31,71,31,173,31,64,31,64,30,64,29,169,31,5,31,249,31,224,31,224,31,248,31,254,31,254,30,61,31,166,31,30,31,254,31,51,31,56,31,39,31,52,31,143,31,143,30,61,31,9,31,168,31,69,31,187,31,91,31,38,31,105,31,105,30,218,31,218,30,116,31,219,31,179,31,97,31,158,31,118,31,76,31,76,30,149,31,6,31,6,30,60,31,62,31,169,31,134,31,170,31,170,30,66,31,205,31,156,31,44,31,108,31,37,31,88,31,180,31,104,31,167,31,16,31,2,31,127,31,156,31,92,31,92,30,255,31,220,31,220,30,72,31,157,31,132,31,132,30,191,31,77,31,130,31,130,30,29,31,171,31,112,31,110,31,84,31,65,31,65,30,251,31,165,31,69,31,41,31,41,30,210,31,189,31,189,30,57,31,181,31,83,31,123,31,123,30,221,31,200,31,77,31,52,31,205,31,181,31,50,31,145,31,108,31,76,31,164,31,6,31,165,31,165,30,27,31,56,31,77,31,8,31,8,30,130,31,157,31,8,31,159,31,186,31,11,31,238,31,212,31,179,31,188,31,188,30,91,31,221,31,60,31,60,30,172,31,60,31,205,31,68,31,91,31,172,31,193,31,216,31,40,31,169,31,81,31,242,31,244,31,214,31,214,30,114,31,218,31,243,31,208,31,14,31,97,31,208,31,242,31,242,30,242,29,167,31,87,31,185,31,248,31,44,31,236,31,168,31,168,30,33,31,244,31,244,30,244,29,184,31,225,31,228,31,20,31,20,30,66,31,211,31,115,31,206,31,15,31,61,31,118,31,56,31,18,31,16,31,139,31,227,31,227,30,227,29,82,31,82,30,72,31,231,31,48,31,205,31,143,31,178,31,221,31,217,31,201,31,104,31,240,31,72,31,20,31,70,31,70,30,241,31,206,31,102,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
