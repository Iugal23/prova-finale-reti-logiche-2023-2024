-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_748 is
end project_tb_748;

architecture project_tb_arch_748 of project_tb_748 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 183;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (158,0,28,0,0,0,27,0,180,0,1,0,247,0,109,0,112,0,86,0,0,0,106,0,158,0,39,0,3,0,94,0,245,0,0,0,21,0,149,0,24,0,32,0,92,0,74,0,136,0,93,0,104,0,28,0,117,0,155,0,24,0,218,0,0,0,22,0,61,0,177,0,188,0,205,0,210,0,95,0,148,0,50,0,120,0,128,0,239,0,255,0,240,0,21,0,66,0,22,0,0,0,0,0,150,0,168,0,130,0,0,0,63,0,120,0,203,0,0,0,249,0,0,0,6,0,188,0,211,0,0,0,75,0,5,0,61,0,240,0,47,0,0,0,229,0,167,0,216,0,237,0,89,0,0,0,0,0,174,0,0,0,10,0,70,0,246,0,145,0,49,0,42,0,0,0,42,0,74,0,250,0,105,0,134,0,93,0,103,0,79,0,223,0,0,0,154,0,0,0,113,0,129,0,227,0,87,0,0,0,62,0,119,0,7,0,15,0,3,0,45,0,224,0,84,0,163,0,13,0,0,0,166,0,7,0,166,0,74,0,103,0,152,0,28,0,0,0,97,0,221,0,153,0,106,0,188,0,44,0,225,0,46,0,90,0,0,0,0,0,25,0,119,0,0,0,161,0,39,0,17,0,0,0,119,0,86,0,132,0,22,0,23,0,3,0,176,0,145,0,36,0,99,0,253,0,244,0,14,0,250,0,156,0,24,0,0,0,229,0,156,0,108,0,153,0,0,0,99,0,0,0,0,0,39,0,221,0,1,0,224,0,149,0,20,0,177,0,133,0,0,0,215,0,170,0,175,0,26,0,0,0,169,0,255,0);
signal scenario_full  : scenario_type := (158,31,28,31,28,30,27,31,180,31,1,31,247,31,109,31,112,31,86,31,86,30,106,31,158,31,39,31,3,31,94,31,245,31,245,30,21,31,149,31,24,31,32,31,92,31,74,31,136,31,93,31,104,31,28,31,117,31,155,31,24,31,218,31,218,30,22,31,61,31,177,31,188,31,205,31,210,31,95,31,148,31,50,31,120,31,128,31,239,31,255,31,240,31,21,31,66,31,22,31,22,30,22,29,150,31,168,31,130,31,130,30,63,31,120,31,203,31,203,30,249,31,249,30,6,31,188,31,211,31,211,30,75,31,5,31,61,31,240,31,47,31,47,30,229,31,167,31,216,31,237,31,89,31,89,30,89,29,174,31,174,30,10,31,70,31,246,31,145,31,49,31,42,31,42,30,42,31,74,31,250,31,105,31,134,31,93,31,103,31,79,31,223,31,223,30,154,31,154,30,113,31,129,31,227,31,87,31,87,30,62,31,119,31,7,31,15,31,3,31,45,31,224,31,84,31,163,31,13,31,13,30,166,31,7,31,166,31,74,31,103,31,152,31,28,31,28,30,97,31,221,31,153,31,106,31,188,31,44,31,225,31,46,31,90,31,90,30,90,29,25,31,119,31,119,30,161,31,39,31,17,31,17,30,119,31,86,31,132,31,22,31,23,31,3,31,176,31,145,31,36,31,99,31,253,31,244,31,14,31,250,31,156,31,24,31,24,30,229,31,156,31,108,31,153,31,153,30,99,31,99,30,99,29,39,31,221,31,1,31,224,31,149,31,20,31,177,31,133,31,133,30,215,31,170,31,175,31,26,31,26,30,169,31,255,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
