-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 688;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (145,0,7,0,0,0,241,0,95,0,172,0,86,0,0,0,78,0,129,0,66,0,88,0,52,0,39,0,0,0,98,0,226,0,28,0,0,0,49,0,0,0,108,0,75,0,140,0,164,0,9,0,19,0,105,0,67,0,0,0,0,0,76,0,172,0,126,0,216,0,26,0,0,0,55,0,97,0,246,0,0,0,197,0,89,0,144,0,84,0,253,0,171,0,0,0,226,0,154,0,93,0,252,0,67,0,9,0,117,0,220,0,65,0,213,0,50,0,0,0,109,0,228,0,125,0,191,0,224,0,178,0,98,0,154,0,40,0,251,0,0,0,251,0,0,0,105,0,0,0,183,0,91,0,172,0,0,0,142,0,30,0,0,0,126,0,228,0,142,0,0,0,72,0,238,0,4,0,27,0,113,0,59,0,66,0,140,0,194,0,179,0,47,0,0,0,175,0,29,0,231,0,147,0,83,0,157,0,104,0,238,0,16,0,121,0,0,0,0,0,82,0,52,0,93,0,21,0,3,0,0,0,118,0,83,0,30,0,171,0,100,0,212,0,108,0,178,0,0,0,78,0,206,0,100,0,226,0,62,0,149,0,253,0,93,0,4,0,146,0,139,0,50,0,206,0,0,0,111,0,21,0,200,0,5,0,0,0,89,0,191,0,39,0,139,0,19,0,199,0,0,0,239,0,74,0,0,0,200,0,179,0,0,0,124,0,96,0,148,0,0,0,86,0,0,0,0,0,0,0,237,0,0,0,109,0,0,0,13,0,13,0,242,0,85,0,220,0,0,0,0,0,0,0,16,0,216,0,107,0,221,0,246,0,157,0,2,0,157,0,22,0,96,0,88,0,94,0,225,0,115,0,171,0,248,0,85,0,136,0,0,0,248,0,2,0,129,0,248,0,201,0,91,0,13,0,0,0,178,0,35,0,48,0,216,0,178,0,213,0,117,0,12,0,210,0,130,0,219,0,111,0,1,0,167,0,98,0,83,0,72,0,172,0,0,0,83,0,98,0,85,0,218,0,250,0,219,0,118,0,6,0,226,0,100,0,26,0,53,0,158,0,198,0,78,0,109,0,73,0,0,0,10,0,0,0,45,0,231,0,64,0,12,0,65,0,147,0,0,0,0,0,0,0,196,0,0,0,83,0,112,0,23,0,44,0,31,0,0,0,16,0,38,0,3,0,238,0,100,0,159,0,0,0,146,0,216,0,22,0,137,0,0,0,111,0,161,0,89,0,196,0,98,0,0,0,16,0,0,0,15,0,255,0,197,0,204,0,0,0,0,0,77,0,0,0,180,0,13,0,10,0,105,0,120,0,228,0,88,0,69,0,53,0,18,0,199,0,220,0,81,0,71,0,169,0,9,0,21,0,80,0,45,0,25,0,2,0,0,0,186,0,0,0,115,0,139,0,126,0,166,0,0,0,0,0,0,0,92,0,232,0,110,0,134,0,217,0,59,0,20,0,0,0,70,0,218,0,0,0,4,0,14,0,152,0,57,0,228,0,0,0,14,0,49,0,0,0,12,0,242,0,155,0,0,0,0,0,0,0,211,0,155,0,0,0,39,0,222,0,7,0,55,0,0,0,34,0,0,0,182,0,62,0,223,0,66,0,190,0,122,0,202,0,0,0,41,0,33,0,112,0,0,0,0,0,27,0,211,0,86,0,0,0,156,0,64,0,144,0,86,0,0,0,115,0,248,0,191,0,0,0,78,0,0,0,138,0,0,0,132,0,0,0,0,0,174,0,55,0,39,0,111,0,0,0,85,0,0,0,60,0,50,0,182,0,0,0,249,0,91,0,0,0,143,0,252,0,254,0,0,0,181,0,210,0,0,0,240,0,155,0,100,0,0,0,0,0,217,0,244,0,110,0,120,0,45,0,48,0,241,0,117,0,155,0,0,0,0,0,0,0,0,0,233,0,252,0,47,0,74,0,0,0,149,0,68,0,136,0,0,0,0,0,19,0,105,0,102,0,0,0,0,0,93,0,199,0,228,0,45,0,231,0,0,0,0,0,4,0,0,0,38,0,183,0,0,0,136,0,47,0,0,0,199,0,0,0,0,0,154,0,28,0,137,0,143,0,252,0,196,0,216,0,0,0,100,0,212,0,204,0,251,0,160,0,40,0,72,0,132,0,133,0,104,0,173,0,0,0,163,0,231,0,25,0,0,0,145,0,15,0,15,0,228,0,231,0,251,0,0,0,175,0,83,0,158,0,49,0,34,0,43,0,202,0,143,0,25,0,216,0,0,0,165,0,210,0,60,0,0,0,71,0,123,0,125,0,109,0,83,0,226,0,43,0,96,0,76,0,147,0,222,0,0,0,130,0,0,0,13,0,184,0,38,0,42,0,243,0,131,0,0,0,0,0,16,0,0,0,13,0,181,0,96,0,6,0,181,0,13,0,62,0,88,0,44,0,172,0,104,0,0,0,81,0,0,0,0,0,55,0,0,0,51,0,0,0,64,0,132,0,118,0,0,0,151,0,0,0,31,0,0,0,179,0,24,0,150,0,35,0,30,0,245,0,0,0,0,0,63,0,0,0,0,0,49,0,57,0,171,0,72,0,193,0,216,0,177,0,66,0,80,0,0,0,40,0,42,0,147,0,30,0,0,0,105,0,0,0,0,0,95,0,35,0,134,0,152,0,148,0,58,0,36,0,11,0,243,0,129,0,12,0,86,0,191,0,91,0,254,0,218,0,65,0,139,0,0,0,238,0,61,0,16,0,0,0,0,0,106,0,127,0,240,0,128,0,217,0,50,0,202,0,0,0,90,0,15,0,0,0,208,0,199,0,157,0,39,0,0,0,201,0,17,0,20,0,98,0,0,0,63,0,154,0,235,0,71,0,66,0,0,0,97,0,220,0,0,0,0,0,0,0,59,0,233,0,204,0,72,0,153,0,234,0,233,0,148,0,151,0,18,0,0,0,186,0,220,0,4,0,10,0,49,0,0,0,0,0,3,0,251,0,89,0,20,0,92,0,76,0,227,0,37,0,17,0,0,0,13,0,138,0,75,0,87,0,18,0,119,0,85,0,199,0,109,0,122,0,0,0,17,0,252,0,50,0,221,0,0,0,52,0,217,0);
signal scenario_full  : scenario_type := (145,31,7,31,7,30,241,31,95,31,172,31,86,31,86,30,78,31,129,31,66,31,88,31,52,31,39,31,39,30,98,31,226,31,28,31,28,30,49,31,49,30,108,31,75,31,140,31,164,31,9,31,19,31,105,31,67,31,67,30,67,29,76,31,172,31,126,31,216,31,26,31,26,30,55,31,97,31,246,31,246,30,197,31,89,31,144,31,84,31,253,31,171,31,171,30,226,31,154,31,93,31,252,31,67,31,9,31,117,31,220,31,65,31,213,31,50,31,50,30,109,31,228,31,125,31,191,31,224,31,178,31,98,31,154,31,40,31,251,31,251,30,251,31,251,30,105,31,105,30,183,31,91,31,172,31,172,30,142,31,30,31,30,30,126,31,228,31,142,31,142,30,72,31,238,31,4,31,27,31,113,31,59,31,66,31,140,31,194,31,179,31,47,31,47,30,175,31,29,31,231,31,147,31,83,31,157,31,104,31,238,31,16,31,121,31,121,30,121,29,82,31,52,31,93,31,21,31,3,31,3,30,118,31,83,31,30,31,171,31,100,31,212,31,108,31,178,31,178,30,78,31,206,31,100,31,226,31,62,31,149,31,253,31,93,31,4,31,146,31,139,31,50,31,206,31,206,30,111,31,21,31,200,31,5,31,5,30,89,31,191,31,39,31,139,31,19,31,199,31,199,30,239,31,74,31,74,30,200,31,179,31,179,30,124,31,96,31,148,31,148,30,86,31,86,30,86,29,86,28,237,31,237,30,109,31,109,30,13,31,13,31,242,31,85,31,220,31,220,30,220,29,220,28,16,31,216,31,107,31,221,31,246,31,157,31,2,31,157,31,22,31,96,31,88,31,94,31,225,31,115,31,171,31,248,31,85,31,136,31,136,30,248,31,2,31,129,31,248,31,201,31,91,31,13,31,13,30,178,31,35,31,48,31,216,31,178,31,213,31,117,31,12,31,210,31,130,31,219,31,111,31,1,31,167,31,98,31,83,31,72,31,172,31,172,30,83,31,98,31,85,31,218,31,250,31,219,31,118,31,6,31,226,31,100,31,26,31,53,31,158,31,198,31,78,31,109,31,73,31,73,30,10,31,10,30,45,31,231,31,64,31,12,31,65,31,147,31,147,30,147,29,147,28,196,31,196,30,83,31,112,31,23,31,44,31,31,31,31,30,16,31,38,31,3,31,238,31,100,31,159,31,159,30,146,31,216,31,22,31,137,31,137,30,111,31,161,31,89,31,196,31,98,31,98,30,16,31,16,30,15,31,255,31,197,31,204,31,204,30,204,29,77,31,77,30,180,31,13,31,10,31,105,31,120,31,228,31,88,31,69,31,53,31,18,31,199,31,220,31,81,31,71,31,169,31,9,31,21,31,80,31,45,31,25,31,2,31,2,30,186,31,186,30,115,31,139,31,126,31,166,31,166,30,166,29,166,28,92,31,232,31,110,31,134,31,217,31,59,31,20,31,20,30,70,31,218,31,218,30,4,31,14,31,152,31,57,31,228,31,228,30,14,31,49,31,49,30,12,31,242,31,155,31,155,30,155,29,155,28,211,31,155,31,155,30,39,31,222,31,7,31,55,31,55,30,34,31,34,30,182,31,62,31,223,31,66,31,190,31,122,31,202,31,202,30,41,31,33,31,112,31,112,30,112,29,27,31,211,31,86,31,86,30,156,31,64,31,144,31,86,31,86,30,115,31,248,31,191,31,191,30,78,31,78,30,138,31,138,30,132,31,132,30,132,29,174,31,55,31,39,31,111,31,111,30,85,31,85,30,60,31,50,31,182,31,182,30,249,31,91,31,91,30,143,31,252,31,254,31,254,30,181,31,210,31,210,30,240,31,155,31,100,31,100,30,100,29,217,31,244,31,110,31,120,31,45,31,48,31,241,31,117,31,155,31,155,30,155,29,155,28,155,27,233,31,252,31,47,31,74,31,74,30,149,31,68,31,136,31,136,30,136,29,19,31,105,31,102,31,102,30,102,29,93,31,199,31,228,31,45,31,231,31,231,30,231,29,4,31,4,30,38,31,183,31,183,30,136,31,47,31,47,30,199,31,199,30,199,29,154,31,28,31,137,31,143,31,252,31,196,31,216,31,216,30,100,31,212,31,204,31,251,31,160,31,40,31,72,31,132,31,133,31,104,31,173,31,173,30,163,31,231,31,25,31,25,30,145,31,15,31,15,31,228,31,231,31,251,31,251,30,175,31,83,31,158,31,49,31,34,31,43,31,202,31,143,31,25,31,216,31,216,30,165,31,210,31,60,31,60,30,71,31,123,31,125,31,109,31,83,31,226,31,43,31,96,31,76,31,147,31,222,31,222,30,130,31,130,30,13,31,184,31,38,31,42,31,243,31,131,31,131,30,131,29,16,31,16,30,13,31,181,31,96,31,6,31,181,31,13,31,62,31,88,31,44,31,172,31,104,31,104,30,81,31,81,30,81,29,55,31,55,30,51,31,51,30,64,31,132,31,118,31,118,30,151,31,151,30,31,31,31,30,179,31,24,31,150,31,35,31,30,31,245,31,245,30,245,29,63,31,63,30,63,29,49,31,57,31,171,31,72,31,193,31,216,31,177,31,66,31,80,31,80,30,40,31,42,31,147,31,30,31,30,30,105,31,105,30,105,29,95,31,35,31,134,31,152,31,148,31,58,31,36,31,11,31,243,31,129,31,12,31,86,31,191,31,91,31,254,31,218,31,65,31,139,31,139,30,238,31,61,31,16,31,16,30,16,29,106,31,127,31,240,31,128,31,217,31,50,31,202,31,202,30,90,31,15,31,15,30,208,31,199,31,157,31,39,31,39,30,201,31,17,31,20,31,98,31,98,30,63,31,154,31,235,31,71,31,66,31,66,30,97,31,220,31,220,30,220,29,220,28,59,31,233,31,204,31,72,31,153,31,234,31,233,31,148,31,151,31,18,31,18,30,186,31,220,31,4,31,10,31,49,31,49,30,49,29,3,31,251,31,89,31,20,31,92,31,76,31,227,31,37,31,17,31,17,30,13,31,138,31,75,31,87,31,18,31,119,31,85,31,199,31,109,31,122,31,122,30,17,31,252,31,50,31,221,31,221,30,52,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
