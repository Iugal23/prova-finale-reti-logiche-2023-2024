-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 714;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (208,0,97,0,76,0,207,0,229,0,238,0,211,0,77,0,83,0,0,0,0,0,21,0,0,0,207,0,140,0,136,0,107,0,212,0,104,0,208,0,213,0,4,0,46,0,125,0,55,0,65,0,123,0,217,0,109,0,95,0,64,0,130,0,253,0,0,0,162,0,223,0,145,0,77,0,117,0,0,0,94,0,84,0,144,0,50,0,196,0,143,0,116,0,91,0,150,0,0,0,0,0,205,0,0,0,29,0,0,0,223,0,0,0,158,0,131,0,114,0,114,0,238,0,101,0,134,0,220,0,0,0,28,0,140,0,0,0,0,0,82,0,204,0,118,0,212,0,100,0,215,0,82,0,34,0,176,0,23,0,77,0,0,0,44,0,235,0,97,0,185,0,169,0,9,0,255,0,28,0,200,0,37,0,0,0,70,0,163,0,80,0,0,0,176,0,111,0,203,0,37,0,106,0,0,0,4,0,4,0,0,0,66,0,0,0,248,0,11,0,245,0,181,0,211,0,147,0,241,0,0,0,191,0,0,0,159,0,12,0,134,0,0,0,194,0,0,0,0,0,181,0,0,0,217,0,108,0,152,0,250,0,159,0,32,0,222,0,34,0,255,0,50,0,237,0,169,0,56,0,172,0,30,0,240,0,42,0,159,0,39,0,0,0,246,0,0,0,246,0,53,0,63,0,0,0,153,0,240,0,0,0,120,0,0,0,192,0,227,0,0,0,79,0,197,0,78,0,144,0,37,0,90,0,164,0,60,0,34,0,64,0,197,0,88,0,198,0,187,0,111,0,177,0,112,0,75,0,58,0,62,0,0,0,92,0,229,0,63,0,0,0,194,0,0,0,149,0,248,0,39,0,78,0,101,0,199,0,110,0,181,0,178,0,85,0,110,0,153,0,0,0,0,0,149,0,192,0,92,0,72,0,113,0,0,0,23,0,177,0,84,0,228,0,4,0,174,0,204,0,0,0,215,0,238,0,137,0,0,0,44,0,201,0,0,0,56,0,255,0,212,0,37,0,0,0,0,0,190,0,50,0,146,0,0,0,0,0,183,0,0,0,8,0,183,0,0,0,241,0,27,0,244,0,88,0,102,0,94,0,54,0,0,0,110,0,0,0,162,0,6,0,21,0,54,0,127,0,61,0,0,0,99,0,185,0,12,0,22,0,3,0,205,0,0,0,194,0,149,0,207,0,222,0,219,0,57,0,110,0,16,0,196,0,12,0,0,0,84,0,0,0,0,0,0,0,172,0,175,0,0,0,43,0,235,0,102,0,117,0,156,0,105,0,95,0,14,0,96,0,0,0,132,0,228,0,67,0,74,0,250,0,180,0,206,0,45,0,102,0,0,0,10,0,117,0,28,0,0,0,110,0,0,0,0,0,0,0,0,0,163,0,221,0,180,0,0,0,224,0,0,0,0,0,0,0,75,0,172,0,99,0,114,0,130,0,0,0,140,0,0,0,129,0,163,0,106,0,137,0,0,0,0,0,184,0,108,0,71,0,71,0,0,0,0,0,0,0,66,0,115,0,201,0,79,0,66,0,196,0,241,0,216,0,168,0,81,0,158,0,217,0,151,0,27,0,0,0,2,0,99,0,189,0,140,0,199,0,221,0,164,0,7,0,232,0,156,0,0,0,0,0,86,0,177,0,84,0,219,0,0,0,36,0,205,0,48,0,0,0,0,0,124,0,75,0,80,0,23,0,38,0,222,0,0,0,0,0,226,0,109,0,19,0,3,0,42,0,66,0,248,0,39,0,0,0,0,0,73,0,46,0,17,0,0,0,95,0,88,0,0,0,0,0,234,0,0,0,239,0,194,0,21,0,138,0,100,0,1,0,116,0,0,0,82,0,133,0,0,0,241,0,109,0,225,0,147,0,156,0,45,0,243,0,61,0,91,0,24,0,164,0,94,0,0,0,0,0,156,0,200,0,0,0,165,0,130,0,81,0,24,0,127,0,79,0,53,0,59,0,112,0,71,0,110,0,126,0,113,0,215,0,224,0,64,0,90,0,40,0,3,0,123,0,241,0,0,0,35,0,243,0,172,0,236,0,139,0,236,0,191,0,221,0,212,0,197,0,51,0,233,0,38,0,0,0,151,0,169,0,254,0,22,0,28,0,208,0,99,0,244,0,0,0,0,0,184,0,132,0,0,0,200,0,224,0,166,0,0,0,182,0,215,0,108,0,158,0,193,0,164,0,173,0,234,0,255,0,23,0,242,0,130,0,245,0,0,0,175,0,0,0,213,0,172,0,154,0,153,0,133,0,133,0,108,0,0,0,240,0,227,0,0,0,39,0,202,0,129,0,80,0,186,0,0,0,46,0,0,0,72,0,82,0,0,0,0,0,0,0,254,0,155,0,0,0,0,0,0,0,61,0,0,0,85,0,147,0,195,0,132,0,0,0,221,0,13,0,219,0,104,0,12,0,3,0,36,0,184,0,84,0,0,0,0,0,0,0,183,0,35,0,32,0,0,0,71,0,92,0,99,0,68,0,66,0,94,0,31,0,0,0,79,0,84,0,35,0,239,0,201,0,230,0,0,0,62,0,246,0,5,0,41,0,38,0,141,0,178,0,70,0,191,0,253,0,72,0,169,0,0,0,183,0,0,0,85,0,126,0,0,0,72,0,42,0,0,0,0,0,0,0,0,0,156,0,109,0,162,0,140,0,195,0,4,0,71,0,253,0,178,0,0,0,141,0,85,0,146,0,212,0,253,0,0,0,236,0,116,0,68,0,74,0,0,0,216,0,247,0,0,0,197,0,135,0,154,0,223,0,0,0,145,0,167,0,16,0,236,0,216,0,0,0,254,0,47,0,161,0,251,0,178,0,174,0,89,0,34,0,69,0,216,0,140,0,68,0,0,0,0,0,231,0,166,0,184,0,0,0,0,0,213,0,244,0,218,0,0,0,96,0,159,0,58,0,14,0,0,0,167,0,0,0,54,0,0,0,85,0,0,0,223,0,101,0,82,0,131,0,125,0,169,0,0,0,86,0,0,0,223,0,169,0,224,0,161,0,89,0,77,0,100,0,0,0,0,0,58,0,13,0,226,0,239,0,110,0,47,0,137,0,160,0,0,0,0,0,53,0,129,0,157,0,5,0,0,0,200,0,159,0,212,0,0,0,0,0,2,0,106,0,0,0,78,0,6,0,52,0,0,0,184,0,134,0,0,0,89,0,115,0,191,0,112,0,13,0);
signal scenario_full  : scenario_type := (208,31,97,31,76,31,207,31,229,31,238,31,211,31,77,31,83,31,83,30,83,29,21,31,21,30,207,31,140,31,136,31,107,31,212,31,104,31,208,31,213,31,4,31,46,31,125,31,55,31,65,31,123,31,217,31,109,31,95,31,64,31,130,31,253,31,253,30,162,31,223,31,145,31,77,31,117,31,117,30,94,31,84,31,144,31,50,31,196,31,143,31,116,31,91,31,150,31,150,30,150,29,205,31,205,30,29,31,29,30,223,31,223,30,158,31,131,31,114,31,114,31,238,31,101,31,134,31,220,31,220,30,28,31,140,31,140,30,140,29,82,31,204,31,118,31,212,31,100,31,215,31,82,31,34,31,176,31,23,31,77,31,77,30,44,31,235,31,97,31,185,31,169,31,9,31,255,31,28,31,200,31,37,31,37,30,70,31,163,31,80,31,80,30,176,31,111,31,203,31,37,31,106,31,106,30,4,31,4,31,4,30,66,31,66,30,248,31,11,31,245,31,181,31,211,31,147,31,241,31,241,30,191,31,191,30,159,31,12,31,134,31,134,30,194,31,194,30,194,29,181,31,181,30,217,31,108,31,152,31,250,31,159,31,32,31,222,31,34,31,255,31,50,31,237,31,169,31,56,31,172,31,30,31,240,31,42,31,159,31,39,31,39,30,246,31,246,30,246,31,53,31,63,31,63,30,153,31,240,31,240,30,120,31,120,30,192,31,227,31,227,30,79,31,197,31,78,31,144,31,37,31,90,31,164,31,60,31,34,31,64,31,197,31,88,31,198,31,187,31,111,31,177,31,112,31,75,31,58,31,62,31,62,30,92,31,229,31,63,31,63,30,194,31,194,30,149,31,248,31,39,31,78,31,101,31,199,31,110,31,181,31,178,31,85,31,110,31,153,31,153,30,153,29,149,31,192,31,92,31,72,31,113,31,113,30,23,31,177,31,84,31,228,31,4,31,174,31,204,31,204,30,215,31,238,31,137,31,137,30,44,31,201,31,201,30,56,31,255,31,212,31,37,31,37,30,37,29,190,31,50,31,146,31,146,30,146,29,183,31,183,30,8,31,183,31,183,30,241,31,27,31,244,31,88,31,102,31,94,31,54,31,54,30,110,31,110,30,162,31,6,31,21,31,54,31,127,31,61,31,61,30,99,31,185,31,12,31,22,31,3,31,205,31,205,30,194,31,149,31,207,31,222,31,219,31,57,31,110,31,16,31,196,31,12,31,12,30,84,31,84,30,84,29,84,28,172,31,175,31,175,30,43,31,235,31,102,31,117,31,156,31,105,31,95,31,14,31,96,31,96,30,132,31,228,31,67,31,74,31,250,31,180,31,206,31,45,31,102,31,102,30,10,31,117,31,28,31,28,30,110,31,110,30,110,29,110,28,110,27,163,31,221,31,180,31,180,30,224,31,224,30,224,29,224,28,75,31,172,31,99,31,114,31,130,31,130,30,140,31,140,30,129,31,163,31,106,31,137,31,137,30,137,29,184,31,108,31,71,31,71,31,71,30,71,29,71,28,66,31,115,31,201,31,79,31,66,31,196,31,241,31,216,31,168,31,81,31,158,31,217,31,151,31,27,31,27,30,2,31,99,31,189,31,140,31,199,31,221,31,164,31,7,31,232,31,156,31,156,30,156,29,86,31,177,31,84,31,219,31,219,30,36,31,205,31,48,31,48,30,48,29,124,31,75,31,80,31,23,31,38,31,222,31,222,30,222,29,226,31,109,31,19,31,3,31,42,31,66,31,248,31,39,31,39,30,39,29,73,31,46,31,17,31,17,30,95,31,88,31,88,30,88,29,234,31,234,30,239,31,194,31,21,31,138,31,100,31,1,31,116,31,116,30,82,31,133,31,133,30,241,31,109,31,225,31,147,31,156,31,45,31,243,31,61,31,91,31,24,31,164,31,94,31,94,30,94,29,156,31,200,31,200,30,165,31,130,31,81,31,24,31,127,31,79,31,53,31,59,31,112,31,71,31,110,31,126,31,113,31,215,31,224,31,64,31,90,31,40,31,3,31,123,31,241,31,241,30,35,31,243,31,172,31,236,31,139,31,236,31,191,31,221,31,212,31,197,31,51,31,233,31,38,31,38,30,151,31,169,31,254,31,22,31,28,31,208,31,99,31,244,31,244,30,244,29,184,31,132,31,132,30,200,31,224,31,166,31,166,30,182,31,215,31,108,31,158,31,193,31,164,31,173,31,234,31,255,31,23,31,242,31,130,31,245,31,245,30,175,31,175,30,213,31,172,31,154,31,153,31,133,31,133,31,108,31,108,30,240,31,227,31,227,30,39,31,202,31,129,31,80,31,186,31,186,30,46,31,46,30,72,31,82,31,82,30,82,29,82,28,254,31,155,31,155,30,155,29,155,28,61,31,61,30,85,31,147,31,195,31,132,31,132,30,221,31,13,31,219,31,104,31,12,31,3,31,36,31,184,31,84,31,84,30,84,29,84,28,183,31,35,31,32,31,32,30,71,31,92,31,99,31,68,31,66,31,94,31,31,31,31,30,79,31,84,31,35,31,239,31,201,31,230,31,230,30,62,31,246,31,5,31,41,31,38,31,141,31,178,31,70,31,191,31,253,31,72,31,169,31,169,30,183,31,183,30,85,31,126,31,126,30,72,31,42,31,42,30,42,29,42,28,42,27,156,31,109,31,162,31,140,31,195,31,4,31,71,31,253,31,178,31,178,30,141,31,85,31,146,31,212,31,253,31,253,30,236,31,116,31,68,31,74,31,74,30,216,31,247,31,247,30,197,31,135,31,154,31,223,31,223,30,145,31,167,31,16,31,236,31,216,31,216,30,254,31,47,31,161,31,251,31,178,31,174,31,89,31,34,31,69,31,216,31,140,31,68,31,68,30,68,29,231,31,166,31,184,31,184,30,184,29,213,31,244,31,218,31,218,30,96,31,159,31,58,31,14,31,14,30,167,31,167,30,54,31,54,30,85,31,85,30,223,31,101,31,82,31,131,31,125,31,169,31,169,30,86,31,86,30,223,31,169,31,224,31,161,31,89,31,77,31,100,31,100,30,100,29,58,31,13,31,226,31,239,31,110,31,47,31,137,31,160,31,160,30,160,29,53,31,129,31,157,31,5,31,5,30,200,31,159,31,212,31,212,30,212,29,2,31,106,31,106,30,78,31,6,31,52,31,52,30,184,31,134,31,134,30,89,31,115,31,191,31,112,31,13,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
