-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_8 is
end project_tb_8;

architecture project_tb_arch_8 of project_tb_8 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1004;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (86,0,0,0,83,0,107,0,0,0,11,0,34,0,117,0,185,0,171,0,65,0,28,0,0,0,0,0,0,0,0,0,0,0,72,0,131,0,164,0,193,0,0,0,22,0,184,0,199,0,138,0,169,0,90,0,129,0,109,0,29,0,119,0,251,0,31,0,54,0,138,0,115,0,88,0,0,0,227,0,0,0,204,0,63,0,225,0,15,0,149,0,0,0,220,0,206,0,63,0,146,0,24,0,222,0,142,0,128,0,222,0,191,0,0,0,0,0,79,0,166,0,65,0,226,0,149,0,121,0,182,0,127,0,210,0,61,0,123,0,0,0,138,0,223,0,233,0,237,0,0,0,59,0,218,0,83,0,68,0,106,0,0,0,249,0,247,0,17,0,80,0,98,0,105,0,157,0,187,0,17,0,83,0,55,0,170,0,208,0,78,0,227,0,111,0,168,0,150,0,31,0,125,0,73,0,0,0,62,0,146,0,0,0,139,0,0,0,174,0,62,0,0,0,79,0,0,0,211,0,0,0,200,0,174,0,0,0,13,0,115,0,0,0,0,0,12,0,228,0,126,0,208,0,150,0,0,0,158,0,132,0,158,0,0,0,161,0,223,0,15,0,195,0,228,0,77,0,0,0,0,0,0,0,0,0,65,0,24,0,220,0,119,0,0,0,44,0,0,0,227,0,180,0,79,0,0,0,89,0,111,0,0,0,121,0,146,0,179,0,92,0,16,0,240,0,0,0,70,0,121,0,0,0,193,0,0,0,193,0,237,0,243,0,16,0,78,0,236,0,222,0,63,0,76,0,107,0,227,0,0,0,183,0,57,0,215,0,57,0,9,0,0,0,197,0,214,0,0,0,0,0,197,0,229,0,0,0,222,0,255,0,7,0,66,0,96,0,134,0,29,0,0,0,18,0,163,0,88,0,74,0,196,0,16,0,10,0,1,0,184,0,215,0,29,0,11,0,186,0,60,0,34,0,144,0,217,0,45,0,0,0,131,0,253,0,0,0,199,0,180,0,76,0,0,0,0,0,114,0,231,0,0,0,0,0,0,0,201,0,225,0,168,0,190,0,19,0,105,0,28,0,85,0,99,0,0,0,170,0,13,0,28,0,0,0,45,0,207,0,238,0,0,0,254,0,232,0,0,0,7,0,207,0,3,0,115,0,0,0,224,0,223,0,153,0,53,0,181,0,165,0,0,0,141,0,44,0,0,0,11,0,110,0,126,0,83,0,242,0,102,0,0,0,170,0,164,0,0,0,96,0,58,0,129,0,248,0,0,0,0,0,107,0,123,0,160,0,70,0,241,0,0,0,3,0,11,0,249,0,171,0,97,0,3,0,214,0,220,0,43,0,167,0,180,0,0,0,112,0,23,0,53,0,187,0,155,0,45,0,26,0,161,0,78,0,151,0,0,0,209,0,168,0,248,0,0,0,79,0,28,0,0,0,213,0,143,0,2,0,217,0,184,0,106,0,41,0,158,0,70,0,53,0,5,0,0,0,249,0,197,0,180,0,239,0,78,0,155,0,0,0,5,0,0,0,0,0,181,0,55,0,0,0,55,0,162,0,226,0,138,0,0,0,18,0,0,0,4,0,172,0,66,0,0,0,173,0,68,0,0,0,70,0,0,0,244,0,211,0,126,0,1,0,144,0,77,0,0,0,104,0,13,0,218,0,76,0,96,0,214,0,164,0,80,0,249,0,0,0,0,0,227,0,114,0,217,0,75,0,104,0,0,0,110,0,79,0,48,0,151,0,0,0,0,0,131,0,3,0,210,0,218,0,57,0,54,0,170,0,0,0,251,0,166,0,213,0,12,0,8,0,55,0,105,0,77,0,149,0,123,0,0,0,74,0,201,0,203,0,73,0,176,0,28,0,0,0,0,0,180,0,124,0,176,0,189,0,84,0,6,0,237,0,65,0,2,0,75,0,26,0,219,0,220,0,133,0,159,0,134,0,236,0,165,0,71,0,71,0,71,0,0,0,0,0,99,0,0,0,0,0,191,0,0,0,181,0,217,0,58,0,252,0,119,0,80,0,127,0,0,0,21,0,95,0,117,0,184,0,10,0,0,0,88,0,0,0,228,0,203,0,93,0,222,0,0,0,0,0,0,0,0,0,37,0,251,0,222,0,0,0,74,0,158,0,139,0,66,0,0,0,116,0,181,0,171,0,219,0,48,0,191,0,72,0,17,0,182,0,47,0,78,0,175,0,64,0,49,0,0,0,191,0,235,0,12,0,182,0,164,0,0,0,57,0,9,0,11,0,99,0,135,0,0,0,211,0,34,0,0,0,250,0,0,0,0,0,116,0,188,0,126,0,196,0,0,0,121,0,193,0,0,0,92,0,244,0,107,0,106,0,109,0,233,0,0,0,178,0,131,0,80,0,134,0,27,0,50,0,0,0,133,0,230,0,73,0,156,0,55,0,37,0,132,0,0,0,226,0,91,0,65,0,0,0,44,0,221,0,163,0,22,0,53,0,140,0,138,0,162,0,174,0,144,0,0,0,218,0,66,0,52,0,248,0,144,0,208,0,0,0,32,0,0,0,220,0,41,0,107,0,31,0,20,0,184,0,28,0,155,0,8,0,220,0,161,0,0,0,195,0,157,0,38,0,124,0,32,0,121,0,143,0,195,0,102,0,199,0,196,0,252,0,0,0,0,0,212,0,105,0,101,0,112,0,132,0,223,0,121,0,0,0,131,0,133,0,71,0,106,0,254,0,85,0,0,0,181,0,4,0,218,0,0,0,221,0,63,0,53,0,40,0,0,0,68,0,253,0,57,0,0,0,12,0,42,0,0,0,179,0,228,0,0,0,236,0,5,0,179,0,7,0,0,0,132,0,237,0,246,0,90,0,111,0,22,0,188,0,154,0,2,0,0,0,185,0,0,0,88,0,29,0,28,0,108,0,182,0,185,0,182,0,0,0,0,0,42,0,65,0,212,0,233,0,102,0,128,0,204,0,0,0,135,0,191,0,103,0,0,0,0,0,94,0,46,0,0,0,138,0,116,0,124,0,0,0,53,0,0,0,80,0,0,0,169,0,0,0,0,0,32,0,108,0,0,0,47,0,0,0,0,0,0,0,33,0,53,0,174,0,93,0,24,0,81,0,0,0,223,0,13,0,230,0,95,0,143,0,57,0,150,0,92,0,173,0,93,0,241,0,172,0,7,0,192,0,22,0,229,0,4,0,194,0,0,0,46,0,0,0,240,0,32,0,29,0,188,0,12,0,11,0,43,0,249,0,86,0,117,0,227,0,0,0,0,0,0,0,152,0,194,0,247,0,142,0,36,0,35,0,185,0,0,0,0,0,130,0,0,0,0,0,0,0,0,0,206,0,216,0,216,0,173,0,22,0,0,0,69,0,126,0,0,0,134,0,26,0,51,0,0,0,97,0,208,0,246,0,105,0,167,0,0,0,52,0,88,0,188,0,137,0,150,0,14,0,206,0,176,0,146,0,200,0,0,0,153,0,246,0,0,0,204,0,240,0,116,0,0,0,82,0,199,0,182,0,243,0,6,0,4,0,177,0,78,0,15,0,72,0,87,0,47,0,243,0,50,0,89,0,122,0,133,0,45,0,1,0,0,0,0,0,100,0,62,0,11,0,188,0,116,0,0,0,53,0,26,0,0,0,245,0,151,0,96,0,123,0,0,0,107,0,79,0,108,0,211,0,248,0,168,0,112,0,5,0,195,0,246,0,30,0,0,0,0,0,0,0,217,0,230,0,72,0,0,0,12,0,0,0,148,0,174,0,135,0,236,0,185,0,107,0,140,0,0,0,255,0,31,0,173,0,126,0,53,0,124,0,99,0,252,0,54,0,0,0,123,0,170,0,0,0,55,0,246,0,114,0,0,0,105,0,163,0,207,0,47,0,190,0,86,0,19,0,70,0,203,0,204,0,151,0,86,0,232,0,25,0,15,0,162,0,236,0,0,0,70,0,229,0,57,0,0,0,247,0,0,0,222,0,213,0,0,0,197,0,84,0,56,0,144,0,91,0,165,0,140,0,21,0,145,0,168,0,154,0,8,0,49,0,13,0,56,0,0,0,162,0,16,0,0,0,28,0,0,0,0,0,205,0,0,0,235,0,251,0,203,0,142,0,21,0,222,0,76,0,233,0,188,0,220,0,0,0,233,0,248,0,0,0,0,0,199,0,73,0,230,0,142,0,216,0,44,0,39,0,75,0,0,0,211,0,148,0,95,0,110,0,0,0,248,0,69,0,93,0,21,0,66,0,35,0,62,0,70,0,48,0,73,0,174,0,94,0,136,0,214,0,0,0,134,0,0,0,70,0,83,0,178,0,234,0,92,0,213,0,227,0,37,0,232,0,194,0,0,0,0,0,149,0,92,0,0,0,0,0,82,0,12,0,133,0,206,0,0,0,252,0,18,0,0,0,151,0,116,0,0,0,119,0,49,0,97,0,179,0,158,0,42,0,165,0,0,0,151,0,187,0,0,0,138,0,173,0,41,0,97,0,29,0,166,0,0,0,0,0);
signal scenario_full  : scenario_type := (86,31,86,30,83,31,107,31,107,30,11,31,34,31,117,31,185,31,171,31,65,31,28,31,28,30,28,29,28,28,28,27,28,26,72,31,131,31,164,31,193,31,193,30,22,31,184,31,199,31,138,31,169,31,90,31,129,31,109,31,29,31,119,31,251,31,31,31,54,31,138,31,115,31,88,31,88,30,227,31,227,30,204,31,63,31,225,31,15,31,149,31,149,30,220,31,206,31,63,31,146,31,24,31,222,31,142,31,128,31,222,31,191,31,191,30,191,29,79,31,166,31,65,31,226,31,149,31,121,31,182,31,127,31,210,31,61,31,123,31,123,30,138,31,223,31,233,31,237,31,237,30,59,31,218,31,83,31,68,31,106,31,106,30,249,31,247,31,17,31,80,31,98,31,105,31,157,31,187,31,17,31,83,31,55,31,170,31,208,31,78,31,227,31,111,31,168,31,150,31,31,31,125,31,73,31,73,30,62,31,146,31,146,30,139,31,139,30,174,31,62,31,62,30,79,31,79,30,211,31,211,30,200,31,174,31,174,30,13,31,115,31,115,30,115,29,12,31,228,31,126,31,208,31,150,31,150,30,158,31,132,31,158,31,158,30,161,31,223,31,15,31,195,31,228,31,77,31,77,30,77,29,77,28,77,27,65,31,24,31,220,31,119,31,119,30,44,31,44,30,227,31,180,31,79,31,79,30,89,31,111,31,111,30,121,31,146,31,179,31,92,31,16,31,240,31,240,30,70,31,121,31,121,30,193,31,193,30,193,31,237,31,243,31,16,31,78,31,236,31,222,31,63,31,76,31,107,31,227,31,227,30,183,31,57,31,215,31,57,31,9,31,9,30,197,31,214,31,214,30,214,29,197,31,229,31,229,30,222,31,255,31,7,31,66,31,96,31,134,31,29,31,29,30,18,31,163,31,88,31,74,31,196,31,16,31,10,31,1,31,184,31,215,31,29,31,11,31,186,31,60,31,34,31,144,31,217,31,45,31,45,30,131,31,253,31,253,30,199,31,180,31,76,31,76,30,76,29,114,31,231,31,231,30,231,29,231,28,201,31,225,31,168,31,190,31,19,31,105,31,28,31,85,31,99,31,99,30,170,31,13,31,28,31,28,30,45,31,207,31,238,31,238,30,254,31,232,31,232,30,7,31,207,31,3,31,115,31,115,30,224,31,223,31,153,31,53,31,181,31,165,31,165,30,141,31,44,31,44,30,11,31,110,31,126,31,83,31,242,31,102,31,102,30,170,31,164,31,164,30,96,31,58,31,129,31,248,31,248,30,248,29,107,31,123,31,160,31,70,31,241,31,241,30,3,31,11,31,249,31,171,31,97,31,3,31,214,31,220,31,43,31,167,31,180,31,180,30,112,31,23,31,53,31,187,31,155,31,45,31,26,31,161,31,78,31,151,31,151,30,209,31,168,31,248,31,248,30,79,31,28,31,28,30,213,31,143,31,2,31,217,31,184,31,106,31,41,31,158,31,70,31,53,31,5,31,5,30,249,31,197,31,180,31,239,31,78,31,155,31,155,30,5,31,5,30,5,29,181,31,55,31,55,30,55,31,162,31,226,31,138,31,138,30,18,31,18,30,4,31,172,31,66,31,66,30,173,31,68,31,68,30,70,31,70,30,244,31,211,31,126,31,1,31,144,31,77,31,77,30,104,31,13,31,218,31,76,31,96,31,214,31,164,31,80,31,249,31,249,30,249,29,227,31,114,31,217,31,75,31,104,31,104,30,110,31,79,31,48,31,151,31,151,30,151,29,131,31,3,31,210,31,218,31,57,31,54,31,170,31,170,30,251,31,166,31,213,31,12,31,8,31,55,31,105,31,77,31,149,31,123,31,123,30,74,31,201,31,203,31,73,31,176,31,28,31,28,30,28,29,180,31,124,31,176,31,189,31,84,31,6,31,237,31,65,31,2,31,75,31,26,31,219,31,220,31,133,31,159,31,134,31,236,31,165,31,71,31,71,31,71,31,71,30,71,29,99,31,99,30,99,29,191,31,191,30,181,31,217,31,58,31,252,31,119,31,80,31,127,31,127,30,21,31,95,31,117,31,184,31,10,31,10,30,88,31,88,30,228,31,203,31,93,31,222,31,222,30,222,29,222,28,222,27,37,31,251,31,222,31,222,30,74,31,158,31,139,31,66,31,66,30,116,31,181,31,171,31,219,31,48,31,191,31,72,31,17,31,182,31,47,31,78,31,175,31,64,31,49,31,49,30,191,31,235,31,12,31,182,31,164,31,164,30,57,31,9,31,11,31,99,31,135,31,135,30,211,31,34,31,34,30,250,31,250,30,250,29,116,31,188,31,126,31,196,31,196,30,121,31,193,31,193,30,92,31,244,31,107,31,106,31,109,31,233,31,233,30,178,31,131,31,80,31,134,31,27,31,50,31,50,30,133,31,230,31,73,31,156,31,55,31,37,31,132,31,132,30,226,31,91,31,65,31,65,30,44,31,221,31,163,31,22,31,53,31,140,31,138,31,162,31,174,31,144,31,144,30,218,31,66,31,52,31,248,31,144,31,208,31,208,30,32,31,32,30,220,31,41,31,107,31,31,31,20,31,184,31,28,31,155,31,8,31,220,31,161,31,161,30,195,31,157,31,38,31,124,31,32,31,121,31,143,31,195,31,102,31,199,31,196,31,252,31,252,30,252,29,212,31,105,31,101,31,112,31,132,31,223,31,121,31,121,30,131,31,133,31,71,31,106,31,254,31,85,31,85,30,181,31,4,31,218,31,218,30,221,31,63,31,53,31,40,31,40,30,68,31,253,31,57,31,57,30,12,31,42,31,42,30,179,31,228,31,228,30,236,31,5,31,179,31,7,31,7,30,132,31,237,31,246,31,90,31,111,31,22,31,188,31,154,31,2,31,2,30,185,31,185,30,88,31,29,31,28,31,108,31,182,31,185,31,182,31,182,30,182,29,42,31,65,31,212,31,233,31,102,31,128,31,204,31,204,30,135,31,191,31,103,31,103,30,103,29,94,31,46,31,46,30,138,31,116,31,124,31,124,30,53,31,53,30,80,31,80,30,169,31,169,30,169,29,32,31,108,31,108,30,47,31,47,30,47,29,47,28,33,31,53,31,174,31,93,31,24,31,81,31,81,30,223,31,13,31,230,31,95,31,143,31,57,31,150,31,92,31,173,31,93,31,241,31,172,31,7,31,192,31,22,31,229,31,4,31,194,31,194,30,46,31,46,30,240,31,32,31,29,31,188,31,12,31,11,31,43,31,249,31,86,31,117,31,227,31,227,30,227,29,227,28,152,31,194,31,247,31,142,31,36,31,35,31,185,31,185,30,185,29,130,31,130,30,130,29,130,28,130,27,206,31,216,31,216,31,173,31,22,31,22,30,69,31,126,31,126,30,134,31,26,31,51,31,51,30,97,31,208,31,246,31,105,31,167,31,167,30,52,31,88,31,188,31,137,31,150,31,14,31,206,31,176,31,146,31,200,31,200,30,153,31,246,31,246,30,204,31,240,31,116,31,116,30,82,31,199,31,182,31,243,31,6,31,4,31,177,31,78,31,15,31,72,31,87,31,47,31,243,31,50,31,89,31,122,31,133,31,45,31,1,31,1,30,1,29,100,31,62,31,11,31,188,31,116,31,116,30,53,31,26,31,26,30,245,31,151,31,96,31,123,31,123,30,107,31,79,31,108,31,211,31,248,31,168,31,112,31,5,31,195,31,246,31,30,31,30,30,30,29,30,28,217,31,230,31,72,31,72,30,12,31,12,30,148,31,174,31,135,31,236,31,185,31,107,31,140,31,140,30,255,31,31,31,173,31,126,31,53,31,124,31,99,31,252,31,54,31,54,30,123,31,170,31,170,30,55,31,246,31,114,31,114,30,105,31,163,31,207,31,47,31,190,31,86,31,19,31,70,31,203,31,204,31,151,31,86,31,232,31,25,31,15,31,162,31,236,31,236,30,70,31,229,31,57,31,57,30,247,31,247,30,222,31,213,31,213,30,197,31,84,31,56,31,144,31,91,31,165,31,140,31,21,31,145,31,168,31,154,31,8,31,49,31,13,31,56,31,56,30,162,31,16,31,16,30,28,31,28,30,28,29,205,31,205,30,235,31,251,31,203,31,142,31,21,31,222,31,76,31,233,31,188,31,220,31,220,30,233,31,248,31,248,30,248,29,199,31,73,31,230,31,142,31,216,31,44,31,39,31,75,31,75,30,211,31,148,31,95,31,110,31,110,30,248,31,69,31,93,31,21,31,66,31,35,31,62,31,70,31,48,31,73,31,174,31,94,31,136,31,214,31,214,30,134,31,134,30,70,31,83,31,178,31,234,31,92,31,213,31,227,31,37,31,232,31,194,31,194,30,194,29,149,31,92,31,92,30,92,29,82,31,12,31,133,31,206,31,206,30,252,31,18,31,18,30,151,31,116,31,116,30,119,31,49,31,97,31,179,31,158,31,42,31,165,31,165,30,151,31,187,31,187,30,138,31,173,31,41,31,97,31,29,31,166,31,166,30,166,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
