-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 570;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,0,0,0,0,212,0,211,0,252,0,19,0,0,0,9,0,198,0,96,0,55,0,27,0,250,0,183,0,66,0,150,0,155,0,207,0,78,0,0,0,214,0,0,0,0,0,22,0,28,0,132,0,141,0,0,0,0,0,173,0,0,0,149,0,6,0,0,0,159,0,231,0,55,0,0,0,129,0,122,0,0,0,7,0,69,0,0,0,55,0,6,0,122,0,0,0,71,0,22,0,30,0,0,0,156,0,7,0,40,0,57,0,227,0,110,0,58,0,0,0,144,0,156,0,190,0,134,0,168,0,120,0,97,0,0,0,64,0,201,0,244,0,125,0,233,0,47,0,143,0,119,0,243,0,223,0,198,0,27,0,71,0,30,0,163,0,173,0,11,0,221,0,91,0,95,0,161,0,167,0,77,0,0,0,1,0,231,0,49,0,2,0,13,0,92,0,0,0,103,0,184,0,0,0,64,0,0,0,184,0,255,0,207,0,0,0,0,0,221,0,105,0,199,0,207,0,235,0,135,0,203,0,0,0,78,0,155,0,70,0,168,0,254,0,0,0,0,0,103,0,70,0,53,0,0,0,211,0,62,0,240,0,131,0,76,0,40,0,175,0,0,0,168,0,19,0,206,0,156,0,0,0,189,0,0,0,225,0,89,0,89,0,144,0,191,0,193,0,102,0,0,0,0,0,115,0,45,0,250,0,0,0,183,0,195,0,4,0,176,0,158,0,229,0,242,0,48,0,233,0,208,0,103,0,0,0,218,0,23,0,172,0,184,0,166,0,0,0,96,0,199,0,172,0,145,0,70,0,0,0,190,0,0,0,189,0,218,0,31,0,0,0,153,0,61,0,220,0,232,0,103,0,153,0,158,0,0,0,100,0,47,0,25,0,37,0,0,0,221,0,0,0,133,0,80,0,155,0,129,0,148,0,63,0,137,0,0,0,137,0,231,0,191,0,17,0,87,0,0,0,193,0,243,0,60,0,0,0,239,0,249,0,2,0,17,0,156,0,0,0,26,0,0,0,198,0,36,0,0,0,0,0,8,0,0,0,190,0,167,0,229,0,73,0,165,0,133,0,88,0,0,0,1,0,67,0,46,0,160,0,241,0,161,0,69,0,128,0,217,0,169,0,20,0,0,0,11,0,72,0,17,0,160,0,1,0,0,0,22,0,217,0,3,0,253,0,9,0,218,0,164,0,0,0,237,0,131,0,0,0,149,0,0,0,0,0,194,0,11,0,150,0,0,0,176,0,83,0,6,0,232,0,101,0,6,0,234,0,0,0,180,0,172,0,245,0,186,0,82,0,84,0,169,0,146,0,142,0,134,0,49,0,227,0,231,0,255,0,196,0,126,0,21,0,88,0,84,0,118,0,97,0,109,0,93,0,242,0,72,0,40,0,127,0,192,0,139,0,106,0,54,0,34,0,184,0,120,0,139,0,191,0,0,0,112,0,174,0,0,0,178,0,250,0,25,0,141,0,154,0,200,0,0,0,26,0,241,0,26,0,0,0,9,0,194,0,108,0,0,0,0,0,137,0,186,0,0,0,16,0,21,0,217,0,127,0,101,0,167,0,202,0,62,0,200,0,169,0,21,0,147,0,0,0,196,0,43,0,249,0,253,0,162,0,207,0,255,0,193,0,17,0,224,0,10,0,0,0,0,0,90,0,40,0,26,0,178,0,106,0,0,0,37,0,184,0,139,0,205,0,217,0,64,0,48,0,0,0,11,0,245,0,188,0,203,0,198,0,195,0,241,0,0,0,223,0,0,0,251,0,241,0,63,0,214,0,27,0,141,0,72,0,0,0,185,0,0,0,187,0,167,0,0,0,72,0,0,0,157,0,246,0,74,0,165,0,121,0,51,0,23,0,0,0,0,0,126,0,0,0,0,0,6,0,151,0,0,0,0,0,149,0,150,0,103,0,107,0,0,0,184,0,68,0,0,0,181,0,215,0,87,0,147,0,117,0,161,0,0,0,0,0,214,0,127,0,60,0,95,0,208,0,195,0,115,0,93,0,0,0,242,0,143,0,0,0,217,0,20,0,0,0,0,0,48,0,112,0,201,0,8,0,225,0,237,0,233,0,0,0,0,0,0,0,187,0,50,0,45,0,195,0,108,0,144,0,0,0,95,0,30,0,128,0,161,0,201,0,34,0,0,0,105,0,151,0,93,0,0,0,33,0,176,0,105,0,149,0,28,0,0,0,145,0,231,0,70,0,46,0,120,0,195,0,0,0,159,0,247,0,0,0,127,0,35,0,93,0,136,0,203,0,0,0,22,0,41,0,93,0,84,0,71,0,231,0,193,0,80,0,0,0,156,0,195,0,130,0,4,0,31,0,98,0,210,0,215,0,0,0,244,0,129,0,0,0,0,0,181,0,142,0,115,0,236,0,52,0,104,0,239,0,148,0,0,0,40,0,0,0,205,0,245,0,17,0,0,0,42,0,72,0,153,0,0,0,217,0,12,0,148,0,235,0,84,0,0,0,52,0,233,0,211,0,155,0,104,0,134,0,48,0,232,0,233,0,207,0,29,0,59,0,102,0,143,0,171,0);
signal scenario_full  : scenario_type := (35,31,35,30,35,29,212,31,211,31,252,31,19,31,19,30,9,31,198,31,96,31,55,31,27,31,250,31,183,31,66,31,150,31,155,31,207,31,78,31,78,30,214,31,214,30,214,29,22,31,28,31,132,31,141,31,141,30,141,29,173,31,173,30,149,31,6,31,6,30,159,31,231,31,55,31,55,30,129,31,122,31,122,30,7,31,69,31,69,30,55,31,6,31,122,31,122,30,71,31,22,31,30,31,30,30,156,31,7,31,40,31,57,31,227,31,110,31,58,31,58,30,144,31,156,31,190,31,134,31,168,31,120,31,97,31,97,30,64,31,201,31,244,31,125,31,233,31,47,31,143,31,119,31,243,31,223,31,198,31,27,31,71,31,30,31,163,31,173,31,11,31,221,31,91,31,95,31,161,31,167,31,77,31,77,30,1,31,231,31,49,31,2,31,13,31,92,31,92,30,103,31,184,31,184,30,64,31,64,30,184,31,255,31,207,31,207,30,207,29,221,31,105,31,199,31,207,31,235,31,135,31,203,31,203,30,78,31,155,31,70,31,168,31,254,31,254,30,254,29,103,31,70,31,53,31,53,30,211,31,62,31,240,31,131,31,76,31,40,31,175,31,175,30,168,31,19,31,206,31,156,31,156,30,189,31,189,30,225,31,89,31,89,31,144,31,191,31,193,31,102,31,102,30,102,29,115,31,45,31,250,31,250,30,183,31,195,31,4,31,176,31,158,31,229,31,242,31,48,31,233,31,208,31,103,31,103,30,218,31,23,31,172,31,184,31,166,31,166,30,96,31,199,31,172,31,145,31,70,31,70,30,190,31,190,30,189,31,218,31,31,31,31,30,153,31,61,31,220,31,232,31,103,31,153,31,158,31,158,30,100,31,47,31,25,31,37,31,37,30,221,31,221,30,133,31,80,31,155,31,129,31,148,31,63,31,137,31,137,30,137,31,231,31,191,31,17,31,87,31,87,30,193,31,243,31,60,31,60,30,239,31,249,31,2,31,17,31,156,31,156,30,26,31,26,30,198,31,36,31,36,30,36,29,8,31,8,30,190,31,167,31,229,31,73,31,165,31,133,31,88,31,88,30,1,31,67,31,46,31,160,31,241,31,161,31,69,31,128,31,217,31,169,31,20,31,20,30,11,31,72,31,17,31,160,31,1,31,1,30,22,31,217,31,3,31,253,31,9,31,218,31,164,31,164,30,237,31,131,31,131,30,149,31,149,30,149,29,194,31,11,31,150,31,150,30,176,31,83,31,6,31,232,31,101,31,6,31,234,31,234,30,180,31,172,31,245,31,186,31,82,31,84,31,169,31,146,31,142,31,134,31,49,31,227,31,231,31,255,31,196,31,126,31,21,31,88,31,84,31,118,31,97,31,109,31,93,31,242,31,72,31,40,31,127,31,192,31,139,31,106,31,54,31,34,31,184,31,120,31,139,31,191,31,191,30,112,31,174,31,174,30,178,31,250,31,25,31,141,31,154,31,200,31,200,30,26,31,241,31,26,31,26,30,9,31,194,31,108,31,108,30,108,29,137,31,186,31,186,30,16,31,21,31,217,31,127,31,101,31,167,31,202,31,62,31,200,31,169,31,21,31,147,31,147,30,196,31,43,31,249,31,253,31,162,31,207,31,255,31,193,31,17,31,224,31,10,31,10,30,10,29,90,31,40,31,26,31,178,31,106,31,106,30,37,31,184,31,139,31,205,31,217,31,64,31,48,31,48,30,11,31,245,31,188,31,203,31,198,31,195,31,241,31,241,30,223,31,223,30,251,31,241,31,63,31,214,31,27,31,141,31,72,31,72,30,185,31,185,30,187,31,167,31,167,30,72,31,72,30,157,31,246,31,74,31,165,31,121,31,51,31,23,31,23,30,23,29,126,31,126,30,126,29,6,31,151,31,151,30,151,29,149,31,150,31,103,31,107,31,107,30,184,31,68,31,68,30,181,31,215,31,87,31,147,31,117,31,161,31,161,30,161,29,214,31,127,31,60,31,95,31,208,31,195,31,115,31,93,31,93,30,242,31,143,31,143,30,217,31,20,31,20,30,20,29,48,31,112,31,201,31,8,31,225,31,237,31,233,31,233,30,233,29,233,28,187,31,50,31,45,31,195,31,108,31,144,31,144,30,95,31,30,31,128,31,161,31,201,31,34,31,34,30,105,31,151,31,93,31,93,30,33,31,176,31,105,31,149,31,28,31,28,30,145,31,231,31,70,31,46,31,120,31,195,31,195,30,159,31,247,31,247,30,127,31,35,31,93,31,136,31,203,31,203,30,22,31,41,31,93,31,84,31,71,31,231,31,193,31,80,31,80,30,156,31,195,31,130,31,4,31,31,31,98,31,210,31,215,31,215,30,244,31,129,31,129,30,129,29,181,31,142,31,115,31,236,31,52,31,104,31,239,31,148,31,148,30,40,31,40,30,205,31,245,31,17,31,17,30,42,31,72,31,153,31,153,30,217,31,12,31,148,31,235,31,84,31,84,30,52,31,233,31,211,31,155,31,104,31,134,31,48,31,232,31,233,31,207,31,29,31,59,31,102,31,143,31,171,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
