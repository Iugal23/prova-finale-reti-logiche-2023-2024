-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 258;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,233,0,0,0,43,0,94,0,69,0,0,0,219,0,215,0,0,0,241,0,38,0,5,0,213,0,0,0,38,0,115,0,87,0,36,0,90,0,119,0,49,0,7,0,0,0,158,0,82,0,54,0,0,0,4,0,133,0,245,0,45,0,0,0,0,0,49,0,16,0,124,0,209,0,0,0,169,0,21,0,120,0,109,0,45,0,180,0,168,0,32,0,254,0,47,0,187,0,81,0,182,0,0,0,194,0,1,0,199,0,148,0,254,0,219,0,0,0,14,0,158,0,0,0,237,0,0,0,110,0,153,0,0,0,193,0,199,0,55,0,4,0,246,0,0,0,245,0,229,0,190,0,190,0,235,0,163,0,196,0,0,0,0,0,0,0,233,0,178,0,114,0,0,0,124,0,73,0,80,0,109,0,0,0,168,0,126,0,52,0,0,0,0,0,101,0,0,0,39,0,0,0,228,0,185,0,0,0,92,0,191,0,114,0,253,0,112,0,85,0,136,0,209,0,171,0,0,0,147,0,0,0,54,0,87,0,115,0,124,0,0,0,0,0,11,0,45,0,42,0,0,0,31,0,140,0,88,0,67,0,179,0,145,0,99,0,0,0,0,0,0,0,171,0,194,0,196,0,67,0,246,0,0,0,181,0,151,0,231,0,137,0,183,0,0,0,249,0,73,0,48,0,0,0,49,0,110,0,65,0,225,0,195,0,98,0,232,0,228,0,38,0,149,0,0,0,23,0,231,0,0,0,208,0,0,0,70,0,114,0,72,0,200,0,213,0,231,0,0,0,0,0,165,0,104,0,0,0,233,0,182,0,137,0,9,0,198,0,228,0,240,0,112,0,28,0,162,0,98,0,3,0,172,0,0,0,213,0,175,0,251,0,27,0,0,0,141,0,0,0,17,0,156,0,0,0,38,0,172,0,135,0,164,0,0,0,115,0,0,0,13,0,0,0,0,0,48,0,239,0,240,0,37,0,0,0,203,0,204,0,149,0,117,0,21,0,212,0,132,0,230,0,241,0,215,0,215,0,203,0,30,0,104,0,202,0,17,0,119,0,108,0,107,0,183,0,95,0,0,0,224,0,0,0,51,0,61,0,130,0,49,0,170,0,40,0,188,0,0,0,3,0,71,0,166,0,25,0,85,0,61,0,166,0);
signal scenario_full  : scenario_type := (149,31,233,31,233,30,43,31,94,31,69,31,69,30,219,31,215,31,215,30,241,31,38,31,5,31,213,31,213,30,38,31,115,31,87,31,36,31,90,31,119,31,49,31,7,31,7,30,158,31,82,31,54,31,54,30,4,31,133,31,245,31,45,31,45,30,45,29,49,31,16,31,124,31,209,31,209,30,169,31,21,31,120,31,109,31,45,31,180,31,168,31,32,31,254,31,47,31,187,31,81,31,182,31,182,30,194,31,1,31,199,31,148,31,254,31,219,31,219,30,14,31,158,31,158,30,237,31,237,30,110,31,153,31,153,30,193,31,199,31,55,31,4,31,246,31,246,30,245,31,229,31,190,31,190,31,235,31,163,31,196,31,196,30,196,29,196,28,233,31,178,31,114,31,114,30,124,31,73,31,80,31,109,31,109,30,168,31,126,31,52,31,52,30,52,29,101,31,101,30,39,31,39,30,228,31,185,31,185,30,92,31,191,31,114,31,253,31,112,31,85,31,136,31,209,31,171,31,171,30,147,31,147,30,54,31,87,31,115,31,124,31,124,30,124,29,11,31,45,31,42,31,42,30,31,31,140,31,88,31,67,31,179,31,145,31,99,31,99,30,99,29,99,28,171,31,194,31,196,31,67,31,246,31,246,30,181,31,151,31,231,31,137,31,183,31,183,30,249,31,73,31,48,31,48,30,49,31,110,31,65,31,225,31,195,31,98,31,232,31,228,31,38,31,149,31,149,30,23,31,231,31,231,30,208,31,208,30,70,31,114,31,72,31,200,31,213,31,231,31,231,30,231,29,165,31,104,31,104,30,233,31,182,31,137,31,9,31,198,31,228,31,240,31,112,31,28,31,162,31,98,31,3,31,172,31,172,30,213,31,175,31,251,31,27,31,27,30,141,31,141,30,17,31,156,31,156,30,38,31,172,31,135,31,164,31,164,30,115,31,115,30,13,31,13,30,13,29,48,31,239,31,240,31,37,31,37,30,203,31,204,31,149,31,117,31,21,31,212,31,132,31,230,31,241,31,215,31,215,31,203,31,30,31,104,31,202,31,17,31,119,31,108,31,107,31,183,31,95,31,95,30,224,31,224,30,51,31,61,31,130,31,49,31,170,31,40,31,188,31,188,30,3,31,71,31,166,31,25,31,85,31,61,31,166,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
