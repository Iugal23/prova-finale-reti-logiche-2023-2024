-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 649;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,162,0,6,0,144,0,252,0,79,0,0,0,50,0,0,0,76,0,35,0,215,0,186,0,228,0,245,0,187,0,8,0,254,0,116,0,0,0,117,0,164,0,123,0,11,0,127,0,31,0,78,0,61,0,225,0,252,0,229,0,103,0,223,0,0,0,0,0,116,0,0,0,0,0,108,0,110,0,0,0,16,0,86,0,7,0,232,0,0,0,0,0,186,0,236,0,212,0,11,0,0,0,239,0,0,0,236,0,189,0,0,0,68,0,50,0,221,0,248,0,181,0,222,0,3,0,208,0,224,0,0,0,54,0,95,0,245,0,64,0,0,0,0,0,22,0,0,0,254,0,107,0,0,0,188,0,0,0,246,0,161,0,205,0,217,0,53,0,38,0,235,0,63,0,148,0,137,0,185,0,21,0,10,0,213,0,28,0,69,0,207,0,67,0,222,0,199,0,0,0,248,0,205,0,146,0,26,0,0,0,0,0,0,0,0,0,66,0,50,0,227,0,96,0,196,0,87,0,102,0,0,0,65,0,0,0,120,0,0,0,107,0,129,0,145,0,154,0,215,0,253,0,0,0,50,0,29,0,171,0,23,0,108,0,0,0,212,0,209,0,198,0,135,0,225,0,194,0,103,0,181,0,15,0,0,0,149,0,94,0,66,0,71,0,176,0,57,0,39,0,0,0,68,0,235,0,45,0,136,0,66,0,86,0,168,0,0,0,172,0,180,0,87,0,191,0,7,0,68,0,0,0,0,0,233,0,152,0,86,0,169,0,11,0,87,0,40,0,197,0,65,0,104,0,63,0,99,0,0,0,128,0,0,0,91,0,189,0,246,0,239,0,194,0,115,0,96,0,25,0,187,0,222,0,0,0,210,0,160,0,83,0,140,0,234,0,0,0,148,0,218,0,203,0,13,0,53,0,59,0,46,0,195,0,112,0,51,0,24,0,251,0,40,0,200,0,198,0,218,0,39,0,22,0,162,0,49,0,32,0,129,0,33,0,40,0,4,0,50,0,0,0,30,0,250,0,0,0,0,0,0,0,202,0,0,0,0,0,212,0,172,0,235,0,231,0,179,0,0,0,50,0,86,0,80,0,44,0,0,0,54,0,0,0,97,0,20,0,144,0,161,0,31,0,51,0,56,0,0,0,45,0,148,0,0,0,0,0,92,0,68,0,251,0,252,0,189,0,226,0,179,0,0,0,120,0,153,0,0,0,106,0,9,0,66,0,28,0,110,0,0,0,165,0,0,0,1,0,67,0,0,0,154,0,200,0,238,0,0,0,48,0,238,0,0,0,215,0,0,0,0,0,116,0,249,0,0,0,86,0,171,0,150,0,128,0,7,0,238,0,77,0,105,0,0,0,101,0,236,0,190,0,11,0,98,0,154,0,0,0,23,0,10,0,173,0,139,0,240,0,54,0,238,0,0,0,252,0,217,0,124,0,244,0,45,0,137,0,191,0,125,0,241,0,215,0,215,0,0,0,0,0,253,0,70,0,15,0,14,0,145,0,254,0,0,0,0,0,90,0,242,0,0,0,21,0,108,0,41,0,40,0,179,0,162,0,17,0,0,0,230,0,209,0,189,0,0,0,143,0,205,0,23,0,204,0,201,0,180,0,27,0,39,0,243,0,69,0,7,0,0,0,226,0,140,0,144,0,112,0,200,0,160,0,173,0,0,0,244,0,10,0,86,0,0,0,69,0,73,0,26,0,90,0,108,0,224,0,162,0,116,0,197,0,133,0,56,0,170,0,90,0,245,0,123,0,170,0,105,0,197,0,0,0,85,0,229,0,0,0,0,0,11,0,162,0,110,0,136,0,187,0,0,0,253,0,0,0,0,0,77,0,72,0,182,0,94,0,0,0,51,0,107,0,0,0,233,0,52,0,154,0,223,0,0,0,0,0,19,0,210,0,0,0,116,0,0,0,0,0,255,0,249,0,121,0,0,0,0,0,185,0,116,0,171,0,224,0,39,0,235,0,23,0,89,0,68,0,155,0,112,0,0,0,0,0,176,0,30,0,198,0,15,0,107,0,30,0,17,0,34,0,206,0,173,0,0,0,104,0,0,0,250,0,120,0,156,0,82,0,108,0,129,0,1,0,222,0,0,0,158,0,0,0,0,0,0,0,177,0,145,0,237,0,0,0,24,0,66,0,209,0,74,0,49,0,104,0,46,0,222,0,196,0,192,0,205,0,214,0,0,0,0,0,176,0,25,0,121,0,6,0,99,0,84,0,10,0,118,0,172,0,182,0,148,0,173,0,64,0,140,0,26,0,87,0,245,0,206,0,0,0,54,0,1,0,61,0,196,0,30,0,234,0,25,0,0,0,227,0,122,0,118,0,170,0,109,0,52,0,75,0,0,0,128,0,6,0,0,0,244,0,0,0,46,0,55,0,0,0,78,0,208,0,49,0,156,0,40,0,232,0,176,0,253,0,139,0,80,0,61,0,138,0,249,0,101,0,71,0,251,0,254,0,2,0,119,0,130,0,13,0,5,0,0,0,107,0,75,0,0,0,111,0,0,0,4,0,126,0,3,0,0,0,9,0,47,0,206,0,86,0,197,0,4,0,25,0,116,0,50,0,0,0,61,0,10,0,11,0,0,0,46,0,107,0,215,0,156,0,182,0,0,0,122,0,249,0,157,0,7,0,0,0,68,0,98,0,116,0,234,0,0,0,0,0,162,0,35,0,216,0,142,0,231,0,95,0,46,0,19,0,202,0,0,0,0,0,0,0,61,0,253,0,163,0,185,0,67,0,63,0,103,0,227,0,118,0,215,0,0,0,192,0,253,0,123,0,94,0,26,0,0,0,0,0,0,0,32,0,238,0,200,0,12,0,70,0,203,0,225,0,118,0,198,0,36,0,196,0,212,0,59,0,191,0,0,0,171,0,49,0,197,0,245,0);
signal scenario_full  : scenario_type := (35,31,162,31,6,31,144,31,252,31,79,31,79,30,50,31,50,30,76,31,35,31,215,31,186,31,228,31,245,31,187,31,8,31,254,31,116,31,116,30,117,31,164,31,123,31,11,31,127,31,31,31,78,31,61,31,225,31,252,31,229,31,103,31,223,31,223,30,223,29,116,31,116,30,116,29,108,31,110,31,110,30,16,31,86,31,7,31,232,31,232,30,232,29,186,31,236,31,212,31,11,31,11,30,239,31,239,30,236,31,189,31,189,30,68,31,50,31,221,31,248,31,181,31,222,31,3,31,208,31,224,31,224,30,54,31,95,31,245,31,64,31,64,30,64,29,22,31,22,30,254,31,107,31,107,30,188,31,188,30,246,31,161,31,205,31,217,31,53,31,38,31,235,31,63,31,148,31,137,31,185,31,21,31,10,31,213,31,28,31,69,31,207,31,67,31,222,31,199,31,199,30,248,31,205,31,146,31,26,31,26,30,26,29,26,28,26,27,66,31,50,31,227,31,96,31,196,31,87,31,102,31,102,30,65,31,65,30,120,31,120,30,107,31,129,31,145,31,154,31,215,31,253,31,253,30,50,31,29,31,171,31,23,31,108,31,108,30,212,31,209,31,198,31,135,31,225,31,194,31,103,31,181,31,15,31,15,30,149,31,94,31,66,31,71,31,176,31,57,31,39,31,39,30,68,31,235,31,45,31,136,31,66,31,86,31,168,31,168,30,172,31,180,31,87,31,191,31,7,31,68,31,68,30,68,29,233,31,152,31,86,31,169,31,11,31,87,31,40,31,197,31,65,31,104,31,63,31,99,31,99,30,128,31,128,30,91,31,189,31,246,31,239,31,194,31,115,31,96,31,25,31,187,31,222,31,222,30,210,31,160,31,83,31,140,31,234,31,234,30,148,31,218,31,203,31,13,31,53,31,59,31,46,31,195,31,112,31,51,31,24,31,251,31,40,31,200,31,198,31,218,31,39,31,22,31,162,31,49,31,32,31,129,31,33,31,40,31,4,31,50,31,50,30,30,31,250,31,250,30,250,29,250,28,202,31,202,30,202,29,212,31,172,31,235,31,231,31,179,31,179,30,50,31,86,31,80,31,44,31,44,30,54,31,54,30,97,31,20,31,144,31,161,31,31,31,51,31,56,31,56,30,45,31,148,31,148,30,148,29,92,31,68,31,251,31,252,31,189,31,226,31,179,31,179,30,120,31,153,31,153,30,106,31,9,31,66,31,28,31,110,31,110,30,165,31,165,30,1,31,67,31,67,30,154,31,200,31,238,31,238,30,48,31,238,31,238,30,215,31,215,30,215,29,116,31,249,31,249,30,86,31,171,31,150,31,128,31,7,31,238,31,77,31,105,31,105,30,101,31,236,31,190,31,11,31,98,31,154,31,154,30,23,31,10,31,173,31,139,31,240,31,54,31,238,31,238,30,252,31,217,31,124,31,244,31,45,31,137,31,191,31,125,31,241,31,215,31,215,31,215,30,215,29,253,31,70,31,15,31,14,31,145,31,254,31,254,30,254,29,90,31,242,31,242,30,21,31,108,31,41,31,40,31,179,31,162,31,17,31,17,30,230,31,209,31,189,31,189,30,143,31,205,31,23,31,204,31,201,31,180,31,27,31,39,31,243,31,69,31,7,31,7,30,226,31,140,31,144,31,112,31,200,31,160,31,173,31,173,30,244,31,10,31,86,31,86,30,69,31,73,31,26,31,90,31,108,31,224,31,162,31,116,31,197,31,133,31,56,31,170,31,90,31,245,31,123,31,170,31,105,31,197,31,197,30,85,31,229,31,229,30,229,29,11,31,162,31,110,31,136,31,187,31,187,30,253,31,253,30,253,29,77,31,72,31,182,31,94,31,94,30,51,31,107,31,107,30,233,31,52,31,154,31,223,31,223,30,223,29,19,31,210,31,210,30,116,31,116,30,116,29,255,31,249,31,121,31,121,30,121,29,185,31,116,31,171,31,224,31,39,31,235,31,23,31,89,31,68,31,155,31,112,31,112,30,112,29,176,31,30,31,198,31,15,31,107,31,30,31,17,31,34,31,206,31,173,31,173,30,104,31,104,30,250,31,120,31,156,31,82,31,108,31,129,31,1,31,222,31,222,30,158,31,158,30,158,29,158,28,177,31,145,31,237,31,237,30,24,31,66,31,209,31,74,31,49,31,104,31,46,31,222,31,196,31,192,31,205,31,214,31,214,30,214,29,176,31,25,31,121,31,6,31,99,31,84,31,10,31,118,31,172,31,182,31,148,31,173,31,64,31,140,31,26,31,87,31,245,31,206,31,206,30,54,31,1,31,61,31,196,31,30,31,234,31,25,31,25,30,227,31,122,31,118,31,170,31,109,31,52,31,75,31,75,30,128,31,6,31,6,30,244,31,244,30,46,31,55,31,55,30,78,31,208,31,49,31,156,31,40,31,232,31,176,31,253,31,139,31,80,31,61,31,138,31,249,31,101,31,71,31,251,31,254,31,2,31,119,31,130,31,13,31,5,31,5,30,107,31,75,31,75,30,111,31,111,30,4,31,126,31,3,31,3,30,9,31,47,31,206,31,86,31,197,31,4,31,25,31,116,31,50,31,50,30,61,31,10,31,11,31,11,30,46,31,107,31,215,31,156,31,182,31,182,30,122,31,249,31,157,31,7,31,7,30,68,31,98,31,116,31,234,31,234,30,234,29,162,31,35,31,216,31,142,31,231,31,95,31,46,31,19,31,202,31,202,30,202,29,202,28,61,31,253,31,163,31,185,31,67,31,63,31,103,31,227,31,118,31,215,31,215,30,192,31,253,31,123,31,94,31,26,31,26,30,26,29,26,28,32,31,238,31,200,31,12,31,70,31,203,31,225,31,118,31,198,31,36,31,196,31,212,31,59,31,191,31,191,30,171,31,49,31,197,31,245,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
