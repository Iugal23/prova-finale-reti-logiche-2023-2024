-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 559;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (2,0,0,0,64,0,111,0,0,0,68,0,131,0,176,0,208,0,13,0,10,0,0,0,123,0,85,0,96,0,0,0,136,0,0,0,93,0,26,0,213,0,127,0,104,0,195,0,89,0,165,0,0,0,219,0,245,0,0,0,133,0,27,0,196,0,142,0,137,0,79,0,32,0,52,0,69,0,206,0,0,0,181,0,0,0,248,0,240,0,0,0,0,0,92,0,131,0,141,0,0,0,150,0,134,0,79,0,0,0,0,0,0,0,176,0,0,0,76,0,19,0,179,0,191,0,249,0,0,0,18,0,42,0,184,0,248,0,116,0,177,0,149,0,128,0,10,0,226,0,0,0,58,0,72,0,0,0,149,0,101,0,149,0,225,0,134,0,95,0,104,0,231,0,202,0,0,0,0,0,86,0,251,0,243,0,215,0,162,0,135,0,203,0,136,0,137,0,165,0,157,0,0,0,144,0,93,0,105,0,165,0,95,0,156,0,0,0,86,0,40,0,185,0,230,0,57,0,35,0,0,0,238,0,0,0,0,0,140,0,150,0,15,0,126,0,170,0,125,0,19,0,11,0,16,0,0,0,100,0,0,0,176,0,11,0,54,0,0,0,160,0,230,0,83,0,149,0,207,0,187,0,190,0,226,0,27,0,68,0,64,0,168,0,112,0,0,0,164,0,156,0,71,0,0,0,63,0,69,0,116,0,162,0,193,0,134,0,0,0,151,0,95,0,193,0,108,0,149,0,163,0,237,0,250,0,0,0,75,0,90,0,196,0,37,0,0,0,60,0,225,0,205,0,83,0,35,0,41,0,72,0,43,0,227,0,0,0,147,0,37,0,5,0,164,0,188,0,0,0,0,0,214,0,145,0,81,0,0,0,0,0,28,0,0,0,0,0,0,0,204,0,248,0,253,0,130,0,241,0,81,0,236,0,166,0,0,0,142,0,253,0,232,0,2,0,117,0,21,0,0,0,181,0,25,0,0,0,112,0,129,0,0,0,173,0,58,0,130,0,243,0,75,0,255,0,231,0,0,0,101,0,182,0,27,0,7,0,197,0,141,0,0,0,40,0,105,0,204,0,15,0,172,0,187,0,3,0,28,0,206,0,64,0,41,0,175,0,21,0,132,0,90,0,139,0,192,0,90,0,217,0,86,0,220,0,242,0,131,0,0,0,134,0,92,0,0,0,156,0,248,0,138,0,52,0,71,0,50,0,46,0,0,0,95,0,167,0,0,0,0,0,0,0,161,0,0,0,0,0,233,0,14,0,128,0,0,0,15,0,61,0,194,0,169,0,237,0,96,0,0,0,15,0,126,0,33,0,247,0,0,0,0,0,251,0,68,0,133,0,187,0,0,0,0,0,243,0,0,0,0,0,204,0,54,0,0,0,14,0,0,0,0,0,206,0,128,0,19,0,167,0,0,0,153,0,47,0,189,0,95,0,125,0,19,0,13,0,38,0,22,0,0,0,204,0,52,0,0,0,0,0,139,0,39,0,230,0,64,0,131,0,0,0,117,0,115,0,89,0,142,0,97,0,175,0,78,0,120,0,96,0,217,0,158,0,205,0,31,0,0,0,0,0,0,0,114,0,0,0,246,0,104,0,223,0,235,0,229,0,57,0,0,0,117,0,58,0,160,0,123,0,168,0,27,0,26,0,105,0,243,0,0,0,0,0,0,0,63,0,80,0,205,0,101,0,123,0,74,0,142,0,0,0,15,0,137,0,86,0,136,0,133,0,11,0,140,0,0,0,34,0,234,0,148,0,211,0,122,0,0,0,0,0,235,0,184,0,207,0,207,0,132,0,175,0,124,0,237,0,0,0,52,0,230,0,181,0,73,0,0,0,64,0,186,0,204,0,0,0,80,0,87,0,73,0,145,0,124,0,186,0,12,0,5,0,0,0,248,0,212,0,120,0,180,0,140,0,183,0,105,0,120,0,73,0,122,0,200,0,217,0,219,0,84,0,36,0,24,0,251,0,67,0,0,0,75,0,13,0,0,0,16,0,145,0,213,0,125,0,57,0,233,0,0,0,129,0,5,0,126,0,64,0,10,0,175,0,0,0,3,0,226,0,70,0,81,0,0,0,0,0,175,0,220,0,134,0,112,0,155,0,0,0,193,0,246,0,78,0,203,0,117,0,208,0,22,0,232,0,194,0,0,0,65,0,234,0,38,0,111,0,227,0,255,0,250,0,0,0,234,0,44,0,0,0,237,0,0,0,254,0,0,0,51,0,0,0,94,0,0,0,62,0,255,0,39,0,106,0,0,0,175,0,53,0,169,0,102,0,206,0,39,0,0,0,0,0,252,0,212,0,187,0,14,0,218,0,0,0,82,0,100,0,85,0,231,0,113,0,5,0,143,0,67,0,88,0,239,0,120,0,46,0,151,0,0,0,159,0,149,0,0,0,34,0,111,0,239,0,147,0,3,0,130,0,33,0,145,0,4,0,165,0,0,0,144,0,248,0,0,0,127,0,167,0,70,0,239,0,122,0,29,0,0,0,191,0);
signal scenario_full  : scenario_type := (2,31,2,30,64,31,111,31,111,30,68,31,131,31,176,31,208,31,13,31,10,31,10,30,123,31,85,31,96,31,96,30,136,31,136,30,93,31,26,31,213,31,127,31,104,31,195,31,89,31,165,31,165,30,219,31,245,31,245,30,133,31,27,31,196,31,142,31,137,31,79,31,32,31,52,31,69,31,206,31,206,30,181,31,181,30,248,31,240,31,240,30,240,29,92,31,131,31,141,31,141,30,150,31,134,31,79,31,79,30,79,29,79,28,176,31,176,30,76,31,19,31,179,31,191,31,249,31,249,30,18,31,42,31,184,31,248,31,116,31,177,31,149,31,128,31,10,31,226,31,226,30,58,31,72,31,72,30,149,31,101,31,149,31,225,31,134,31,95,31,104,31,231,31,202,31,202,30,202,29,86,31,251,31,243,31,215,31,162,31,135,31,203,31,136,31,137,31,165,31,157,31,157,30,144,31,93,31,105,31,165,31,95,31,156,31,156,30,86,31,40,31,185,31,230,31,57,31,35,31,35,30,238,31,238,30,238,29,140,31,150,31,15,31,126,31,170,31,125,31,19,31,11,31,16,31,16,30,100,31,100,30,176,31,11,31,54,31,54,30,160,31,230,31,83,31,149,31,207,31,187,31,190,31,226,31,27,31,68,31,64,31,168,31,112,31,112,30,164,31,156,31,71,31,71,30,63,31,69,31,116,31,162,31,193,31,134,31,134,30,151,31,95,31,193,31,108,31,149,31,163,31,237,31,250,31,250,30,75,31,90,31,196,31,37,31,37,30,60,31,225,31,205,31,83,31,35,31,41,31,72,31,43,31,227,31,227,30,147,31,37,31,5,31,164,31,188,31,188,30,188,29,214,31,145,31,81,31,81,30,81,29,28,31,28,30,28,29,28,28,204,31,248,31,253,31,130,31,241,31,81,31,236,31,166,31,166,30,142,31,253,31,232,31,2,31,117,31,21,31,21,30,181,31,25,31,25,30,112,31,129,31,129,30,173,31,58,31,130,31,243,31,75,31,255,31,231,31,231,30,101,31,182,31,27,31,7,31,197,31,141,31,141,30,40,31,105,31,204,31,15,31,172,31,187,31,3,31,28,31,206,31,64,31,41,31,175,31,21,31,132,31,90,31,139,31,192,31,90,31,217,31,86,31,220,31,242,31,131,31,131,30,134,31,92,31,92,30,156,31,248,31,138,31,52,31,71,31,50,31,46,31,46,30,95,31,167,31,167,30,167,29,167,28,161,31,161,30,161,29,233,31,14,31,128,31,128,30,15,31,61,31,194,31,169,31,237,31,96,31,96,30,15,31,126,31,33,31,247,31,247,30,247,29,251,31,68,31,133,31,187,31,187,30,187,29,243,31,243,30,243,29,204,31,54,31,54,30,14,31,14,30,14,29,206,31,128,31,19,31,167,31,167,30,153,31,47,31,189,31,95,31,125,31,19,31,13,31,38,31,22,31,22,30,204,31,52,31,52,30,52,29,139,31,39,31,230,31,64,31,131,31,131,30,117,31,115,31,89,31,142,31,97,31,175,31,78,31,120,31,96,31,217,31,158,31,205,31,31,31,31,30,31,29,31,28,114,31,114,30,246,31,104,31,223,31,235,31,229,31,57,31,57,30,117,31,58,31,160,31,123,31,168,31,27,31,26,31,105,31,243,31,243,30,243,29,243,28,63,31,80,31,205,31,101,31,123,31,74,31,142,31,142,30,15,31,137,31,86,31,136,31,133,31,11,31,140,31,140,30,34,31,234,31,148,31,211,31,122,31,122,30,122,29,235,31,184,31,207,31,207,31,132,31,175,31,124,31,237,31,237,30,52,31,230,31,181,31,73,31,73,30,64,31,186,31,204,31,204,30,80,31,87,31,73,31,145,31,124,31,186,31,12,31,5,31,5,30,248,31,212,31,120,31,180,31,140,31,183,31,105,31,120,31,73,31,122,31,200,31,217,31,219,31,84,31,36,31,24,31,251,31,67,31,67,30,75,31,13,31,13,30,16,31,145,31,213,31,125,31,57,31,233,31,233,30,129,31,5,31,126,31,64,31,10,31,175,31,175,30,3,31,226,31,70,31,81,31,81,30,81,29,175,31,220,31,134,31,112,31,155,31,155,30,193,31,246,31,78,31,203,31,117,31,208,31,22,31,232,31,194,31,194,30,65,31,234,31,38,31,111,31,227,31,255,31,250,31,250,30,234,31,44,31,44,30,237,31,237,30,254,31,254,30,51,31,51,30,94,31,94,30,62,31,255,31,39,31,106,31,106,30,175,31,53,31,169,31,102,31,206,31,39,31,39,30,39,29,252,31,212,31,187,31,14,31,218,31,218,30,82,31,100,31,85,31,231,31,113,31,5,31,143,31,67,31,88,31,239,31,120,31,46,31,151,31,151,30,159,31,149,31,149,30,34,31,111,31,239,31,147,31,3,31,130,31,33,31,145,31,4,31,165,31,165,30,144,31,248,31,248,30,127,31,167,31,70,31,239,31,122,31,29,31,29,30,191,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
