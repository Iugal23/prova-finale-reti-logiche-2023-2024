-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_323 is
end project_tb_323;

architecture project_tb_arch_323 of project_tb_323 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 859;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,167,0,140,0,218,0,60,0,66,0,40,0,75,0,25,0,130,0,0,0,53,0,141,0,0,0,170,0,22,0,0,0,46,0,93,0,0,0,138,0,121,0,198,0,10,0,118,0,35,0,221,0,0,0,142,0,0,0,22,0,0,0,21,0,246,0,197,0,154,0,253,0,25,0,191,0,247,0,46,0,73,0,210,0,0,0,200,0,0,0,84,0,106,0,179,0,215,0,186,0,0,0,249,0,172,0,33,0,42,0,4,0,179,0,76,0,169,0,29,0,135,0,0,0,241,0,91,0,248,0,164,0,194,0,212,0,0,0,153,0,0,0,198,0,74,0,57,0,94,0,177,0,165,0,73,0,152,0,225,0,6,0,223,0,147,0,62,0,179,0,181,0,0,0,20,0,55,0,33,0,67,0,226,0,0,0,0,0,216,0,115,0,0,0,0,0,172,0,196,0,98,0,0,0,41,0,209,0,130,0,104,0,147,0,17,0,165,0,41,0,151,0,184,0,19,0,163,0,97,0,0,0,191,0,0,0,66,0,36,0,159,0,147,0,233,0,103,0,0,0,42,0,0,0,168,0,139,0,208,0,66,0,0,0,45,0,146,0,132,0,122,0,243,0,115,0,249,0,38,0,143,0,0,0,0,0,118,0,106,0,193,0,122,0,17,0,82,0,251,0,2,0,19,0,0,0,95,0,229,0,53,0,247,0,0,0,63,0,116,0,94,0,17,0,45,0,130,0,219,0,67,0,220,0,16,0,188,0,85,0,62,0,31,0,161,0,0,0,13,0,31,0,0,0,3,0,179,0,242,0,250,0,13,0,0,0,0,0,54,0,111,0,0,0,84,0,21,0,155,0,122,0,47,0,167,0,143,0,0,0,92,0,58,0,104,0,222,0,69,0,140,0,201,0,148,0,40,0,109,0,0,0,186,0,225,0,59,0,211,0,0,0,194,0,45,0,141,0,0,0,97,0,212,0,223,0,0,0,113,0,7,0,124,0,203,0,226,0,110,0,147,0,147,0,177,0,228,0,190,0,0,0,178,0,225,0,0,0,224,0,209,0,0,0,180,0,0,0,142,0,144,0,103,0,52,0,84,0,215,0,244,0,216,0,219,0,164,0,61,0,0,0,223,0,104,0,40,0,163,0,4,0,69,0,0,0,0,0,136,0,253,0,0,0,62,0,111,0,0,0,192,0,113,0,95,0,0,0,159,0,0,0,130,0,89,0,10,0,201,0,25,0,159,0,0,0,101,0,61,0,0,0,0,0,0,0,2,0,0,0,92,0,97,0,32,0,213,0,0,0,40,0,233,0,210,0,114,0,31,0,20,0,216,0,84,0,113,0,241,0,51,0,185,0,139,0,217,0,0,0,169,0,211,0,83,0,85,0,0,0,202,0,234,0,167,0,0,0,34,0,85,0,63,0,19,0,152,0,28,0,0,0,105,0,0,0,103,0,109,0,85,0,115,0,0,0,145,0,83,0,76,0,42,0,27,0,41,0,223,0,0,0,174,0,173,0,151,0,116,0,148,0,214,0,209,0,123,0,87,0,167,0,167,0,184,0,0,0,135,0,66,0,210,0,168,0,20,0,226,0,0,0,44,0,36,0,235,0,19,0,192,0,0,0,211,0,201,0,231,0,95,0,0,0,0,0,51,0,0,0,0,0,89,0,133,0,68,0,39,0,116,0,59,0,31,0,19,0,0,0,0,0,45,0,0,0,0,0,49,0,113,0,123,0,21,0,213,0,33,0,140,0,24,0,25,0,25,0,173,0,50,0,47,0,27,0,16,0,98,0,0,0,142,0,253,0,50,0,113,0,158,0,115,0,19,0,89,0,249,0,56,0,81,0,0,0,58,0,122,0,3,0,52,0,16,0,16,0,0,0,114,0,254,0,55,0,175,0,186,0,3,0,62,0,0,0,53,0,0,0,121,0,197,0,0,0,129,0,95,0,208,0,173,0,0,0,129,0,8,0,96,0,86,0,0,0,171,0,212,0,48,0,0,0,32,0,158,0,0,0,60,0,48,0,235,0,0,0,217,0,162,0,0,0,193,0,244,0,39,0,188,0,6,0,249,0,206,0,0,0,44,0,148,0,114,0,15,0,195,0,0,0,252,0,51,0,101,0,85,0,5,0,211,0,33,0,209,0,0,0,19,0,0,0,85,0,45,0,95,0,242,0,43,0,0,0,180,0,63,0,168,0,195,0,0,0,133,0,182,0,247,0,36,0,154,0,251,0,181,0,0,0,124,0,0,0,90,0,231,0,240,0,0,0,0,0,198,0,232,0,129,0,36,0,0,0,226,0,227,0,0,0,23,0,249,0,187,0,159,0,0,0,140,0,201,0,0,0,0,0,229,0,248,0,169,0,0,0,30,0,173,0,205,0,186,0,252,0,67,0,224,0,34,0,222,0,95,0,254,0,180,0,216,0,240,0,0,0,71,0,32,0,202,0,162,0,52,0,211,0,100,0,65,0,59,0,0,0,208,0,204,0,253,0,0,0,246,0,133,0,0,0,122,0,200,0,154,0,159,0,155,0,60,0,154,0,240,0,2,0,145,0,170,0,243,0,0,0,127,0,213,0,239,0,223,0,228,0,0,0,41,0,180,0,160,0,70,0,106,0,160,0,215,0,191,0,0,0,86,0,147,0,116,0,125,0,154,0,0,0,43,0,183,0,166,0,161,0,0,0,0,0,0,0,24,0,75,0,171,0,245,0,101,0,41,0,11,0,196,0,173,0,0,0,0,0,0,0,231,0,150,0,0,0,164,0,254,0,175,0,81,0,139,0,252,0,12,0,132,0,241,0,185,0,111,0,125,0,157,0,143,0,56,0,22,0,235,0,229,0,74,0,0,0,245,0,97,0,198,0,155,0,20,0,0,0,0,0,217,0,0,0,199,0,214,0,98,0,0,0,106,0,236,0,27,0,148,0,0,0,254,0,0,0,190,0,0,0,22,0,49,0,60,0,95,0,105,0,106,0,232,0,0,0,152,0,242,0,250,0,0,0,252,0,254,0,35,0,207,0,0,0,0,0,102,0,150,0,100,0,11,0,17,0,213,0,0,0,0,0,53,0,127,0,243,0,147,0,0,0,0,0,14,0,44,0,144,0,34,0,111,0,65,0,0,0,136,0,70,0,203,0,117,0,179,0,18,0,204,0,235,0,0,0,235,0,51,0,49,0,132,0,6,0,145,0,223,0,175,0,235,0,118,0,178,0,0,0,0,0,226,0,175,0,176,0,129,0,183,0,164,0,117,0,52,0,157,0,0,0,63,0,73,0,0,0,171,0,31,0,56,0,0,0,227,0,128,0,34,0,149,0,0,0,109,0,0,0,0,0,69,0,140,0,95,0,62,0,8,0,124,0,100,0,152,0,106,0,162,0,0,0,177,0,106,0,115,0,186,0,105,0,34,0,99,0,222,0,151,0,241,0,56,0,25,0,88,0,142,0,131,0,178,0,145,0,166,0,25,0,136,0,142,0,101,0,126,0,13,0,215,0,0,0,118,0,208,0,166,0,90,0,211,0,222,0,0,0,22,0,254,0,253,0,6,0,88,0,58,0,0,0,64,0,0,0,83,0,11,0,0,0,166,0,74,0,53,0,127,0,110,0,236,0,109,0,45,0,0,0,135,0,109,0,45,0,67,0,164,0,252,0,116,0,196,0,31,0,153,0,68,0,194,0,115,0,187,0,0,0,0,0,95,0,248,0,41,0,223,0,57,0,122,0,204,0,163,0,76,0,192,0,108,0,0,0,36,0,35,0,215,0,100,0,0,0,153,0,158,0,50,0,162,0,192,0,22,0,151,0,13,0,0,0,120,0,206,0,188,0,37,0,42,0,30,0);
signal scenario_full  : scenario_type := (0,0,167,31,140,31,218,31,60,31,66,31,40,31,75,31,25,31,130,31,130,30,53,31,141,31,141,30,170,31,22,31,22,30,46,31,93,31,93,30,138,31,121,31,198,31,10,31,118,31,35,31,221,31,221,30,142,31,142,30,22,31,22,30,21,31,246,31,197,31,154,31,253,31,25,31,191,31,247,31,46,31,73,31,210,31,210,30,200,31,200,30,84,31,106,31,179,31,215,31,186,31,186,30,249,31,172,31,33,31,42,31,4,31,179,31,76,31,169,31,29,31,135,31,135,30,241,31,91,31,248,31,164,31,194,31,212,31,212,30,153,31,153,30,198,31,74,31,57,31,94,31,177,31,165,31,73,31,152,31,225,31,6,31,223,31,147,31,62,31,179,31,181,31,181,30,20,31,55,31,33,31,67,31,226,31,226,30,226,29,216,31,115,31,115,30,115,29,172,31,196,31,98,31,98,30,41,31,209,31,130,31,104,31,147,31,17,31,165,31,41,31,151,31,184,31,19,31,163,31,97,31,97,30,191,31,191,30,66,31,36,31,159,31,147,31,233,31,103,31,103,30,42,31,42,30,168,31,139,31,208,31,66,31,66,30,45,31,146,31,132,31,122,31,243,31,115,31,249,31,38,31,143,31,143,30,143,29,118,31,106,31,193,31,122,31,17,31,82,31,251,31,2,31,19,31,19,30,95,31,229,31,53,31,247,31,247,30,63,31,116,31,94,31,17,31,45,31,130,31,219,31,67,31,220,31,16,31,188,31,85,31,62,31,31,31,161,31,161,30,13,31,31,31,31,30,3,31,179,31,242,31,250,31,13,31,13,30,13,29,54,31,111,31,111,30,84,31,21,31,155,31,122,31,47,31,167,31,143,31,143,30,92,31,58,31,104,31,222,31,69,31,140,31,201,31,148,31,40,31,109,31,109,30,186,31,225,31,59,31,211,31,211,30,194,31,45,31,141,31,141,30,97,31,212,31,223,31,223,30,113,31,7,31,124,31,203,31,226,31,110,31,147,31,147,31,177,31,228,31,190,31,190,30,178,31,225,31,225,30,224,31,209,31,209,30,180,31,180,30,142,31,144,31,103,31,52,31,84,31,215,31,244,31,216,31,219,31,164,31,61,31,61,30,223,31,104,31,40,31,163,31,4,31,69,31,69,30,69,29,136,31,253,31,253,30,62,31,111,31,111,30,192,31,113,31,95,31,95,30,159,31,159,30,130,31,89,31,10,31,201,31,25,31,159,31,159,30,101,31,61,31,61,30,61,29,61,28,2,31,2,30,92,31,97,31,32,31,213,31,213,30,40,31,233,31,210,31,114,31,31,31,20,31,216,31,84,31,113,31,241,31,51,31,185,31,139,31,217,31,217,30,169,31,211,31,83,31,85,31,85,30,202,31,234,31,167,31,167,30,34,31,85,31,63,31,19,31,152,31,28,31,28,30,105,31,105,30,103,31,109,31,85,31,115,31,115,30,145,31,83,31,76,31,42,31,27,31,41,31,223,31,223,30,174,31,173,31,151,31,116,31,148,31,214,31,209,31,123,31,87,31,167,31,167,31,184,31,184,30,135,31,66,31,210,31,168,31,20,31,226,31,226,30,44,31,36,31,235,31,19,31,192,31,192,30,211,31,201,31,231,31,95,31,95,30,95,29,51,31,51,30,51,29,89,31,133,31,68,31,39,31,116,31,59,31,31,31,19,31,19,30,19,29,45,31,45,30,45,29,49,31,113,31,123,31,21,31,213,31,33,31,140,31,24,31,25,31,25,31,173,31,50,31,47,31,27,31,16,31,98,31,98,30,142,31,253,31,50,31,113,31,158,31,115,31,19,31,89,31,249,31,56,31,81,31,81,30,58,31,122,31,3,31,52,31,16,31,16,31,16,30,114,31,254,31,55,31,175,31,186,31,3,31,62,31,62,30,53,31,53,30,121,31,197,31,197,30,129,31,95,31,208,31,173,31,173,30,129,31,8,31,96,31,86,31,86,30,171,31,212,31,48,31,48,30,32,31,158,31,158,30,60,31,48,31,235,31,235,30,217,31,162,31,162,30,193,31,244,31,39,31,188,31,6,31,249,31,206,31,206,30,44,31,148,31,114,31,15,31,195,31,195,30,252,31,51,31,101,31,85,31,5,31,211,31,33,31,209,31,209,30,19,31,19,30,85,31,45,31,95,31,242,31,43,31,43,30,180,31,63,31,168,31,195,31,195,30,133,31,182,31,247,31,36,31,154,31,251,31,181,31,181,30,124,31,124,30,90,31,231,31,240,31,240,30,240,29,198,31,232,31,129,31,36,31,36,30,226,31,227,31,227,30,23,31,249,31,187,31,159,31,159,30,140,31,201,31,201,30,201,29,229,31,248,31,169,31,169,30,30,31,173,31,205,31,186,31,252,31,67,31,224,31,34,31,222,31,95,31,254,31,180,31,216,31,240,31,240,30,71,31,32,31,202,31,162,31,52,31,211,31,100,31,65,31,59,31,59,30,208,31,204,31,253,31,253,30,246,31,133,31,133,30,122,31,200,31,154,31,159,31,155,31,60,31,154,31,240,31,2,31,145,31,170,31,243,31,243,30,127,31,213,31,239,31,223,31,228,31,228,30,41,31,180,31,160,31,70,31,106,31,160,31,215,31,191,31,191,30,86,31,147,31,116,31,125,31,154,31,154,30,43,31,183,31,166,31,161,31,161,30,161,29,161,28,24,31,75,31,171,31,245,31,101,31,41,31,11,31,196,31,173,31,173,30,173,29,173,28,231,31,150,31,150,30,164,31,254,31,175,31,81,31,139,31,252,31,12,31,132,31,241,31,185,31,111,31,125,31,157,31,143,31,56,31,22,31,235,31,229,31,74,31,74,30,245,31,97,31,198,31,155,31,20,31,20,30,20,29,217,31,217,30,199,31,214,31,98,31,98,30,106,31,236,31,27,31,148,31,148,30,254,31,254,30,190,31,190,30,22,31,49,31,60,31,95,31,105,31,106,31,232,31,232,30,152,31,242,31,250,31,250,30,252,31,254,31,35,31,207,31,207,30,207,29,102,31,150,31,100,31,11,31,17,31,213,31,213,30,213,29,53,31,127,31,243,31,147,31,147,30,147,29,14,31,44,31,144,31,34,31,111,31,65,31,65,30,136,31,70,31,203,31,117,31,179,31,18,31,204,31,235,31,235,30,235,31,51,31,49,31,132,31,6,31,145,31,223,31,175,31,235,31,118,31,178,31,178,30,178,29,226,31,175,31,176,31,129,31,183,31,164,31,117,31,52,31,157,31,157,30,63,31,73,31,73,30,171,31,31,31,56,31,56,30,227,31,128,31,34,31,149,31,149,30,109,31,109,30,109,29,69,31,140,31,95,31,62,31,8,31,124,31,100,31,152,31,106,31,162,31,162,30,177,31,106,31,115,31,186,31,105,31,34,31,99,31,222,31,151,31,241,31,56,31,25,31,88,31,142,31,131,31,178,31,145,31,166,31,25,31,136,31,142,31,101,31,126,31,13,31,215,31,215,30,118,31,208,31,166,31,90,31,211,31,222,31,222,30,22,31,254,31,253,31,6,31,88,31,58,31,58,30,64,31,64,30,83,31,11,31,11,30,166,31,74,31,53,31,127,31,110,31,236,31,109,31,45,31,45,30,135,31,109,31,45,31,67,31,164,31,252,31,116,31,196,31,31,31,153,31,68,31,194,31,115,31,187,31,187,30,187,29,95,31,248,31,41,31,223,31,57,31,122,31,204,31,163,31,76,31,192,31,108,31,108,30,36,31,35,31,215,31,100,31,100,30,153,31,158,31,50,31,162,31,192,31,22,31,151,31,13,31,13,30,120,31,206,31,188,31,37,31,42,31,30,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
