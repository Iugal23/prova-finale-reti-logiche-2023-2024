-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_983 is
end project_tb_983;

architecture project_tb_arch_983 of project_tb_983 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 715;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,108,0,177,0,16,0,0,0,21,0,185,0,149,0,44,0,89,0,75,0,231,0,27,0,209,0,181,0,251,0,82,0,40,0,11,0,198,0,79,0,0,0,178,0,94,0,239,0,183,0,58,0,133,0,0,0,0,0,55,0,173,0,245,0,63,0,240,0,216,0,210,0,60,0,149,0,129,0,147,0,118,0,0,0,193,0,53,0,75,0,211,0,199,0,119,0,195,0,104,0,163,0,239,0,0,0,0,0,167,0,14,0,248,0,24,0,87,0,17,0,42,0,135,0,0,0,252,0,77,0,197,0,0,0,3,0,0,0,84,0,198,0,191,0,0,0,0,0,138,0,170,0,210,0,209,0,128,0,39,0,0,0,229,0,0,0,11,0,100,0,127,0,95,0,174,0,108,0,191,0,138,0,47,0,100,0,203,0,44,0,28,0,36,0,0,0,0,0,0,0,249,0,0,0,0,0,153,0,0,0,251,0,131,0,253,0,181,0,235,0,199,0,0,0,0,0,114,0,88,0,115,0,154,0,120,0,161,0,177,0,0,0,159,0,0,0,6,0,189,0,155,0,105,0,203,0,0,0,131,0,154,0,173,0,196,0,181,0,0,0,172,0,138,0,44,0,61,0,0,0,67,0,0,0,243,0,230,0,23,0,250,0,209,0,0,0,123,0,114,0,106,0,48,0,195,0,0,0,30,0,245,0,113,0,175,0,27,0,48,0,203,0,29,0,221,0,227,0,82,0,0,0,0,0,0,0,170,0,77,0,0,0,202,0,0,0,51,0,202,0,231,0,153,0,185,0,76,0,0,0,203,0,58,0,146,0,63,0,114,0,171,0,0,0,131,0,55,0,0,0,165,0,26,0,150,0,197,0,18,0,86,0,216,0,52,0,187,0,209,0,106,0,76,0,23,0,76,0,88,0,0,0,153,0,212,0,112,0,135,0,62,0,12,0,182,0,34,0,57,0,0,0,206,0,182,0,1,0,80,0,91,0,176,0,0,0,23,0,89,0,246,0,0,0,56,0,25,0,150,0,213,0,43,0,0,0,66,0,187,0,198,0,249,0,52,0,95,0,78,0,66,0,110,0,0,0,0,0,86,0,184,0,0,0,0,0,0,0,172,0,88,0,170,0,215,0,44,0,0,0,67,0,0,0,41,0,127,0,241,0,32,0,0,0,0,0,41,0,166,0,92,0,202,0,217,0,137,0,55,0,0,0,0,0,11,0,231,0,0,0,42,0,101,0,41,0,0,0,250,0,93,0,150,0,250,0,7,0,37,0,9,0,123,0,250,0,0,0,3,0,211,0,61,0,247,0,135,0,49,0,0,0,100,0,23,0,243,0,95,0,92,0,55,0,253,0,85,0,20,0,173,0,244,0,45,0,83,0,156,0,174,0,0,0,109,0,0,0,200,0,55,0,179,0,238,0,179,0,254,0,175,0,55,0,131,0,0,0,17,0,212,0,223,0,0,0,218,0,240,0,149,0,62,0,25,0,0,0,0,0,134,0,239,0,143,0,66,0,153,0,125,0,208,0,36,0,51,0,153,0,94,0,61,0,123,0,216,0,194,0,0,0,0,0,24,0,4,0,20,0,0,0,0,0,33,0,236,0,170,0,85,0,141,0,113,0,1,0,7,0,133,0,20,0,27,0,229,0,239,0,19,0,183,0,1,0,0,0,0,0,29,0,76,0,59,0,7,0,168,0,0,0,75,0,0,0,82,0,105,0,59,0,211,0,87,0,50,0,0,0,0,0,227,0,0,0,200,0,44,0,76,0,103,0,188,0,0,0,68,0,0,0,134,0,0,0,0,0,194,0,191,0,73,0,161,0,49,0,237,0,245,0,36,0,52,0,44,0,179,0,40,0,228,0,81,0,211,0,163,0,133,0,0,0,0,0,50,0,254,0,200,0,159,0,176,0,126,0,39,0,102,0,169,0,162,0,146,0,196,0,160,0,42,0,165,0,162,0,242,0,163,0,95,0,65,0,228,0,32,0,0,0,82,0,148,0,211,0,234,0,0,0,36,0,24,0,254,0,203,0,95,0,199,0,62,0,200,0,183,0,209,0,8,0,242,0,0,0,54,0,213,0,104,0,123,0,168,0,0,0,233,0,239,0,182,0,115,0,0,0,88,0,172,0,37,0,99,0,0,0,75,0,0,0,0,0,47,0,0,0,42,0,88,0,26,0,251,0,246,0,249,0,53,0,0,0,107,0,51,0,89,0,2,0,179,0,210,0,33,0,84,0,0,0,117,0,0,0,197,0,0,0,154,0,168,0,147,0,144,0,60,0,52,0,23,0,254,0,151,0,145,0,0,0,183,0,175,0,219,0,0,0,50,0,0,0,130,0,94,0,249,0,75,0,0,0,184,0,96,0,67,0,0,0,77,0,96,0,236,0,113,0,0,0,153,0,4,0,0,0,96,0,250,0,57,0,128,0,204,0,254,0,244,0,199,0,238,0,179,0,243,0,249,0,168,0,235,0,126,0,243,0,196,0,89,0,132,0,148,0,0,0,192,0,113,0,0,0,244,0,176,0,109,0,39,0,150,0,0,0,102,0,68,0,151,0,254,0,179,0,148,0,45,0,60,0,0,0,27,0,0,0,241,0,0,0,144,0,205,0,219,0,0,0,0,0,0,0,54,0,252,0,167,0,116,0,254,0,61,0,151,0,22,0,82,0,2,0,0,0,87,0,245,0,189,0,199,0,252,0,30,0,106,0,218,0,0,0,0,0,45,0,0,0,207,0,108,0,4,0,252,0,195,0,73,0,0,0,209,0,135,0,103,0,12,0,183,0,97,0,0,0,229,0,62,0,148,0,1,0,60,0,28,0,0,0,99,0,237,0,241,0,218,0,234,0,28,0,190,0,174,0,51,0,0,0,81,0,91,0,242,0,0,0,0,0,52,0,154,0,10,0,0,0,10,0,4,0,220,0,43,0,0,0,41,0,0,0,220,0,85,0,7,0,173,0,72,0,0,0,107,0,64,0,184,0,60,0,132,0,35,0,106,0,72,0,248,0,0,0,142,0,118,0,81,0,119,0,0,0,2,0,22,0,89,0,110,0,210,0,103,0,76,0,107,0,105,0,185,0,189,0,166,0,151,0,109,0,64,0,108,0,86,0,194,0,164,0,148,0,217,0,0,0,54,0,0,0,208,0,92,0,254,0,87,0,108,0,101,0,42,0,114,0,85,0,191,0);
signal scenario_full  : scenario_type := (0,0,108,31,177,31,16,31,16,30,21,31,185,31,149,31,44,31,89,31,75,31,231,31,27,31,209,31,181,31,251,31,82,31,40,31,11,31,198,31,79,31,79,30,178,31,94,31,239,31,183,31,58,31,133,31,133,30,133,29,55,31,173,31,245,31,63,31,240,31,216,31,210,31,60,31,149,31,129,31,147,31,118,31,118,30,193,31,53,31,75,31,211,31,199,31,119,31,195,31,104,31,163,31,239,31,239,30,239,29,167,31,14,31,248,31,24,31,87,31,17,31,42,31,135,31,135,30,252,31,77,31,197,31,197,30,3,31,3,30,84,31,198,31,191,31,191,30,191,29,138,31,170,31,210,31,209,31,128,31,39,31,39,30,229,31,229,30,11,31,100,31,127,31,95,31,174,31,108,31,191,31,138,31,47,31,100,31,203,31,44,31,28,31,36,31,36,30,36,29,36,28,249,31,249,30,249,29,153,31,153,30,251,31,131,31,253,31,181,31,235,31,199,31,199,30,199,29,114,31,88,31,115,31,154,31,120,31,161,31,177,31,177,30,159,31,159,30,6,31,189,31,155,31,105,31,203,31,203,30,131,31,154,31,173,31,196,31,181,31,181,30,172,31,138,31,44,31,61,31,61,30,67,31,67,30,243,31,230,31,23,31,250,31,209,31,209,30,123,31,114,31,106,31,48,31,195,31,195,30,30,31,245,31,113,31,175,31,27,31,48,31,203,31,29,31,221,31,227,31,82,31,82,30,82,29,82,28,170,31,77,31,77,30,202,31,202,30,51,31,202,31,231,31,153,31,185,31,76,31,76,30,203,31,58,31,146,31,63,31,114,31,171,31,171,30,131,31,55,31,55,30,165,31,26,31,150,31,197,31,18,31,86,31,216,31,52,31,187,31,209,31,106,31,76,31,23,31,76,31,88,31,88,30,153,31,212,31,112,31,135,31,62,31,12,31,182,31,34,31,57,31,57,30,206,31,182,31,1,31,80,31,91,31,176,31,176,30,23,31,89,31,246,31,246,30,56,31,25,31,150,31,213,31,43,31,43,30,66,31,187,31,198,31,249,31,52,31,95,31,78,31,66,31,110,31,110,30,110,29,86,31,184,31,184,30,184,29,184,28,172,31,88,31,170,31,215,31,44,31,44,30,67,31,67,30,41,31,127,31,241,31,32,31,32,30,32,29,41,31,166,31,92,31,202,31,217,31,137,31,55,31,55,30,55,29,11,31,231,31,231,30,42,31,101,31,41,31,41,30,250,31,93,31,150,31,250,31,7,31,37,31,9,31,123,31,250,31,250,30,3,31,211,31,61,31,247,31,135,31,49,31,49,30,100,31,23,31,243,31,95,31,92,31,55,31,253,31,85,31,20,31,173,31,244,31,45,31,83,31,156,31,174,31,174,30,109,31,109,30,200,31,55,31,179,31,238,31,179,31,254,31,175,31,55,31,131,31,131,30,17,31,212,31,223,31,223,30,218,31,240,31,149,31,62,31,25,31,25,30,25,29,134,31,239,31,143,31,66,31,153,31,125,31,208,31,36,31,51,31,153,31,94,31,61,31,123,31,216,31,194,31,194,30,194,29,24,31,4,31,20,31,20,30,20,29,33,31,236,31,170,31,85,31,141,31,113,31,1,31,7,31,133,31,20,31,27,31,229,31,239,31,19,31,183,31,1,31,1,30,1,29,29,31,76,31,59,31,7,31,168,31,168,30,75,31,75,30,82,31,105,31,59,31,211,31,87,31,50,31,50,30,50,29,227,31,227,30,200,31,44,31,76,31,103,31,188,31,188,30,68,31,68,30,134,31,134,30,134,29,194,31,191,31,73,31,161,31,49,31,237,31,245,31,36,31,52,31,44,31,179,31,40,31,228,31,81,31,211,31,163,31,133,31,133,30,133,29,50,31,254,31,200,31,159,31,176,31,126,31,39,31,102,31,169,31,162,31,146,31,196,31,160,31,42,31,165,31,162,31,242,31,163,31,95,31,65,31,228,31,32,31,32,30,82,31,148,31,211,31,234,31,234,30,36,31,24,31,254,31,203,31,95,31,199,31,62,31,200,31,183,31,209,31,8,31,242,31,242,30,54,31,213,31,104,31,123,31,168,31,168,30,233,31,239,31,182,31,115,31,115,30,88,31,172,31,37,31,99,31,99,30,75,31,75,30,75,29,47,31,47,30,42,31,88,31,26,31,251,31,246,31,249,31,53,31,53,30,107,31,51,31,89,31,2,31,179,31,210,31,33,31,84,31,84,30,117,31,117,30,197,31,197,30,154,31,168,31,147,31,144,31,60,31,52,31,23,31,254,31,151,31,145,31,145,30,183,31,175,31,219,31,219,30,50,31,50,30,130,31,94,31,249,31,75,31,75,30,184,31,96,31,67,31,67,30,77,31,96,31,236,31,113,31,113,30,153,31,4,31,4,30,96,31,250,31,57,31,128,31,204,31,254,31,244,31,199,31,238,31,179,31,243,31,249,31,168,31,235,31,126,31,243,31,196,31,89,31,132,31,148,31,148,30,192,31,113,31,113,30,244,31,176,31,109,31,39,31,150,31,150,30,102,31,68,31,151,31,254,31,179,31,148,31,45,31,60,31,60,30,27,31,27,30,241,31,241,30,144,31,205,31,219,31,219,30,219,29,219,28,54,31,252,31,167,31,116,31,254,31,61,31,151,31,22,31,82,31,2,31,2,30,87,31,245,31,189,31,199,31,252,31,30,31,106,31,218,31,218,30,218,29,45,31,45,30,207,31,108,31,4,31,252,31,195,31,73,31,73,30,209,31,135,31,103,31,12,31,183,31,97,31,97,30,229,31,62,31,148,31,1,31,60,31,28,31,28,30,99,31,237,31,241,31,218,31,234,31,28,31,190,31,174,31,51,31,51,30,81,31,91,31,242,31,242,30,242,29,52,31,154,31,10,31,10,30,10,31,4,31,220,31,43,31,43,30,41,31,41,30,220,31,85,31,7,31,173,31,72,31,72,30,107,31,64,31,184,31,60,31,132,31,35,31,106,31,72,31,248,31,248,30,142,31,118,31,81,31,119,31,119,30,2,31,22,31,89,31,110,31,210,31,103,31,76,31,107,31,105,31,185,31,189,31,166,31,151,31,109,31,64,31,108,31,86,31,194,31,164,31,148,31,217,31,217,30,54,31,54,30,208,31,92,31,254,31,87,31,108,31,101,31,42,31,114,31,85,31,191,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
