-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_730 is
end project_tb_730;

architecture project_tb_arch_730 of project_tb_730 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 208;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,1,0,79,0,57,0,60,0,185,0,170,0,90,0,178,0,78,0,0,0,68,0,70,0,52,0,172,0,67,0,40,0,0,0,173,0,67,0,234,0,9,0,52,0,0,0,102,0,77,0,99,0,64,0,60,0,220,0,0,0,176,0,70,0,61,0,0,0,0,0,109,0,138,0,213,0,182,0,0,0,172,0,232,0,180,0,0,0,69,0,19,0,0,0,209,0,115,0,0,0,177,0,204,0,48,0,48,0,0,0,31,0,0,0,48,0,177,0,230,0,144,0,52,0,93,0,60,0,0,0,253,0,227,0,144,0,121,0,107,0,29,0,0,0,0,0,8,0,127,0,30,0,77,0,239,0,62,0,0,0,148,0,245,0,67,0,0,0,49,0,83,0,152,0,6,0,14,0,22,0,25,0,213,0,134,0,247,0,149,0,61,0,116,0,185,0,0,0,60,0,0,0,143,0,20,0,163,0,0,0,0,0,71,0,3,0,123,0,136,0,203,0,164,0,116,0,180,0,79,0,0,0,159,0,0,0,229,0,124,0,90,0,140,0,126,0,234,0,116,0,244,0,80,0,21,0,0,0,0,0,200,0,122,0,5,0,85,0,101,0,133,0,0,0,150,0,219,0,97,0,87,0,210,0,47,0,36,0,164,0,0,0,118,0,179,0,86,0,232,0,213,0,119,0,0,0,70,0,71,0,56,0,43,0,0,0,97,0,64,0,204,0,185,0,0,0,130,0,171,0,203,0,0,0,186,0,0,0,173,0,38,0,36,0,0,0,0,0,0,0,177,0,0,0,8,0,69,0,73,0,230,0,0,0,140,0,85,0,252,0,144,0,47,0,252,0,126,0,74,0,83,0,144,0,0,0,71,0,8,0,54,0,203,0,199,0,0,0,184,0,209,0,0,0,0,0,0,0,3,0,104,0,234,0);
signal scenario_full  : scenario_type := (49,31,1,31,79,31,57,31,60,31,185,31,170,31,90,31,178,31,78,31,78,30,68,31,70,31,52,31,172,31,67,31,40,31,40,30,173,31,67,31,234,31,9,31,52,31,52,30,102,31,77,31,99,31,64,31,60,31,220,31,220,30,176,31,70,31,61,31,61,30,61,29,109,31,138,31,213,31,182,31,182,30,172,31,232,31,180,31,180,30,69,31,19,31,19,30,209,31,115,31,115,30,177,31,204,31,48,31,48,31,48,30,31,31,31,30,48,31,177,31,230,31,144,31,52,31,93,31,60,31,60,30,253,31,227,31,144,31,121,31,107,31,29,31,29,30,29,29,8,31,127,31,30,31,77,31,239,31,62,31,62,30,148,31,245,31,67,31,67,30,49,31,83,31,152,31,6,31,14,31,22,31,25,31,213,31,134,31,247,31,149,31,61,31,116,31,185,31,185,30,60,31,60,30,143,31,20,31,163,31,163,30,163,29,71,31,3,31,123,31,136,31,203,31,164,31,116,31,180,31,79,31,79,30,159,31,159,30,229,31,124,31,90,31,140,31,126,31,234,31,116,31,244,31,80,31,21,31,21,30,21,29,200,31,122,31,5,31,85,31,101,31,133,31,133,30,150,31,219,31,97,31,87,31,210,31,47,31,36,31,164,31,164,30,118,31,179,31,86,31,232,31,213,31,119,31,119,30,70,31,71,31,56,31,43,31,43,30,97,31,64,31,204,31,185,31,185,30,130,31,171,31,203,31,203,30,186,31,186,30,173,31,38,31,36,31,36,30,36,29,36,28,177,31,177,30,8,31,69,31,73,31,230,31,230,30,140,31,85,31,252,31,144,31,47,31,252,31,126,31,74,31,83,31,144,31,144,30,71,31,8,31,54,31,203,31,199,31,199,30,184,31,209,31,209,30,209,29,209,28,3,31,104,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
