-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_798 is
end project_tb_798;

architecture project_tb_arch_798 of project_tb_798 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 778;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,254,0,102,0,245,0,242,0,3,0,83,0,145,0,188,0,114,0,111,0,150,0,0,0,148,0,151,0,186,0,0,0,170,0,36,0,197,0,120,0,240,0,0,0,154,0,116,0,194,0,53,0,10,0,0,0,193,0,159,0,4,0,0,0,132,0,158,0,188,0,97,0,130,0,0,0,12,0,0,0,0,0,58,0,0,0,53,0,0,0,60,0,0,0,201,0,26,0,30,0,0,0,111,0,0,0,35,0,207,0,140,0,132,0,0,0,188,0,0,0,0,0,174,0,46,0,116,0,223,0,94,0,152,0,0,0,68,0,232,0,107,0,142,0,38,0,169,0,215,0,250,0,0,0,183,0,0,0,49,0,0,0,197,0,89,0,90,0,43,0,252,0,43,0,90,0,36,0,187,0,224,0,236,0,177,0,159,0,66,0,202,0,0,0,228,0,113,0,0,0,0,0,156,0,63,0,58,0,210,0,167,0,144,0,133,0,241,0,82,0,0,0,149,0,89,0,0,0,0,0,0,0,0,0,64,0,0,0,0,0,0,0,118,0,182,0,174,0,137,0,0,0,60,0,59,0,0,0,0,0,46,0,76,0,62,0,16,0,51,0,190,0,0,0,99,0,161,0,165,0,24,0,93,0,0,0,0,0,126,0,138,0,59,0,163,0,43,0,248,0,107,0,74,0,14,0,187,0,177,0,3,0,0,0,49,0,0,0,8,0,107,0,0,0,0,0,6,0,23,0,216,0,103,0,205,0,224,0,29,0,115,0,0,0,28,0,253,0,123,0,0,0,37,0,246,0,152,0,186,0,54,0,0,0,215,0,33,0,7,0,37,0,0,0,226,0,216,0,4,0,224,0,198,0,168,0,0,0,253,0,225,0,13,0,164,0,165,0,203,0,1,0,99,0,152,0,0,0,103,0,134,0,0,0,199,0,0,0,154,0,0,0,153,0,177,0,0,0,236,0,210,0,226,0,0,0,30,0,68,0,43,0,62,0,176,0,192,0,184,0,119,0,0,0,87,0,57,0,41,0,15,0,101,0,95,0,94,0,198,0,186,0,0,0,106,0,82,0,0,0,0,0,11,0,45,0,164,0,67,0,153,0,100,0,0,0,148,0,195,0,90,0,111,0,22,0,119,0,201,0,23,0,91,0,252,0,185,0,0,0,135,0,64,0,115,0,179,0,38,0,114,0,0,0,79,0,64,0,102,0,147,0,144,0,49,0,220,0,205,0,0,0,199,0,67,0,108,0,0,0,54,0,46,0,42,0,83,0,192,0,0,0,219,0,205,0,0,0,67,0,144,0,80,0,204,0,223,0,0,0,224,0,159,0,0,0,7,0,107,0,166,0,100,0,115,0,103,0,156,0,69,0,253,0,76,0,2,0,216,0,210,0,243,0,229,0,57,0,64,0,229,0,147,0,3,0,92,0,191,0,98,0,88,0,64,0,179,0,236,0,38,0,206,0,0,0,167,0,5,0,0,0,203,0,208,0,0,0,191,0,44,0,245,0,90,0,0,0,0,0,0,0,0,0,0,0,194,0,202,0,164,0,66,0,130,0,63,0,9,0,31,0,221,0,0,0,182,0,113,0,0,0,59,0,13,0,73,0,35,0,21,0,108,0,145,0,51,0,209,0,96,0,39,0,116,0,154,0,88,0,148,0,253,0,187,0,227,0,58,0,211,0,136,0,178,0,0,0,126,0,0,0,212,0,0,0,183,0,18,0,63,0,0,0,14,0,212,0,0,0,214,0,242,0,65,0,239,0,34,0,72,0,122,0,0,0,93,0,151,0,111,0,166,0,48,0,0,0,164,0,129,0,118,0,203,0,240,0,114,0,0,0,0,0,69,0,7,0,85,0,39,0,90,0,18,0,85,0,137,0,0,0,172,0,46,0,146,0,189,0,43,0,124,0,12,0,0,0,33,0,210,0,230,0,204,0,127,0,21,0,140,0,168,0,39,0,166,0,16,0,146,0,0,0,0,0,13,0,79,0,0,0,14,0,0,0,225,0,116,0,134,0,0,0,0,0,0,0,64,0,192,0,182,0,73,0,65,0,3,0,0,0,153,0,34,0,0,0,23,0,3,0,17,0,101,0,211,0,11,0,165,0,156,0,50,0,0,0,225,0,81,0,245,0,90,0,64,0,20,0,0,0,134,0,83,0,0,0,242,0,52,0,159,0,113,0,0,0,170,0,0,0,0,0,37,0,195,0,168,0,120,0,28,0,186,0,0,0,97,0,198,0,213,0,253,0,0,0,18,0,20,0,79,0,76,0,246,0,241,0,143,0,169,0,179,0,0,0,157,0,59,0,248,0,10,0,158,0,242,0,185,0,228,0,213,0,202,0,129,0,0,0,99,0,243,0,77,0,0,0,24,0,0,0,207,0,235,0,41,0,138,0,186,0,141,0,119,0,113,0,17,0,118,0,86,0,151,0,56,0,19,0,233,0,37,0,233,0,52,0,0,0,239,0,109,0,200,0,86,0,46,0,175,0,115,0,87,0,25,0,85,0,202,0,69,0,0,0,225,0,0,0,221,0,248,0,27,0,217,0,0,0,220,0,253,0,155,0,0,0,152,0,184,0,127,0,17,0,39,0,0,0,215,0,223,0,59,0,101,0,62,0,0,0,0,0,67,0,114,0,100,0,148,0,99,0,0,0,247,0,101,0,138,0,147,0,173,0,17,0,189,0,2,0,0,0,255,0,88,0,86,0,60,0,0,0,12,0,94,0,141,0,0,0,0,0,89,0,0,0,0,0,0,0,0,0,99,0,60,0,91,0,65,0,150,0,0,0,29,0,9,0,147,0,225,0,0,0,60,0,197,0,0,0,174,0,19,0,0,0,64,0,182,0,13,0,65,0,0,0,95,0,192,0,160,0,151,0,36,0,2,0,76,0,175,0,48,0,0,0,219,0,191,0,85,0,227,0,128,0,153,0,236,0,17,0,134,0,48,0,253,0,21,0,0,0,193,0,0,0,180,0,67,0,154,0,23,0,145,0,137,0,250,0,0,0,113,0,237,0,166,0,230,0,12,0,121,0,227,0,102,0,0,0,247,0,0,0,177,0,143,0,85,0,168,0,40,0,211,0,0,0,81,0,0,0,116,0,0,0,22,0,28,0,234,0,176,0,7,0,184,0,197,0,0,0,0,0,195,0,121,0,175,0,142,0,118,0,125,0,109,0,48,0,0,0,163,0,0,0,0,0,97,0,7,0,82,0,197,0,241,0,47,0,100,0,0,0,66,0,138,0,77,0,205,0,29,0,252,0,219,0,154,0,167,0,201,0,128,0,225,0,0,0,203,0,86,0,244,0,108,0,136,0,250,0,0,0,0,0,152,0,0,0,0,0,0,0,0,0,216,0,143,0,54,0,17,0,222,0,17,0,145,0,65,0,134,0,159,0,0,0,201,0,0,0,0,0,38,0,0,0,53,0,239,0,244,0,213,0,69,0,242,0,174,0,122,0,72,0,14,0,238,0);
signal scenario_full  : scenario_type := (232,31,254,31,102,31,245,31,242,31,3,31,83,31,145,31,188,31,114,31,111,31,150,31,150,30,148,31,151,31,186,31,186,30,170,31,36,31,197,31,120,31,240,31,240,30,154,31,116,31,194,31,53,31,10,31,10,30,193,31,159,31,4,31,4,30,132,31,158,31,188,31,97,31,130,31,130,30,12,31,12,30,12,29,58,31,58,30,53,31,53,30,60,31,60,30,201,31,26,31,30,31,30,30,111,31,111,30,35,31,207,31,140,31,132,31,132,30,188,31,188,30,188,29,174,31,46,31,116,31,223,31,94,31,152,31,152,30,68,31,232,31,107,31,142,31,38,31,169,31,215,31,250,31,250,30,183,31,183,30,49,31,49,30,197,31,89,31,90,31,43,31,252,31,43,31,90,31,36,31,187,31,224,31,236,31,177,31,159,31,66,31,202,31,202,30,228,31,113,31,113,30,113,29,156,31,63,31,58,31,210,31,167,31,144,31,133,31,241,31,82,31,82,30,149,31,89,31,89,30,89,29,89,28,89,27,64,31,64,30,64,29,64,28,118,31,182,31,174,31,137,31,137,30,60,31,59,31,59,30,59,29,46,31,76,31,62,31,16,31,51,31,190,31,190,30,99,31,161,31,165,31,24,31,93,31,93,30,93,29,126,31,138,31,59,31,163,31,43,31,248,31,107,31,74,31,14,31,187,31,177,31,3,31,3,30,49,31,49,30,8,31,107,31,107,30,107,29,6,31,23,31,216,31,103,31,205,31,224,31,29,31,115,31,115,30,28,31,253,31,123,31,123,30,37,31,246,31,152,31,186,31,54,31,54,30,215,31,33,31,7,31,37,31,37,30,226,31,216,31,4,31,224,31,198,31,168,31,168,30,253,31,225,31,13,31,164,31,165,31,203,31,1,31,99,31,152,31,152,30,103,31,134,31,134,30,199,31,199,30,154,31,154,30,153,31,177,31,177,30,236,31,210,31,226,31,226,30,30,31,68,31,43,31,62,31,176,31,192,31,184,31,119,31,119,30,87,31,57,31,41,31,15,31,101,31,95,31,94,31,198,31,186,31,186,30,106,31,82,31,82,30,82,29,11,31,45,31,164,31,67,31,153,31,100,31,100,30,148,31,195,31,90,31,111,31,22,31,119,31,201,31,23,31,91,31,252,31,185,31,185,30,135,31,64,31,115,31,179,31,38,31,114,31,114,30,79,31,64,31,102,31,147,31,144,31,49,31,220,31,205,31,205,30,199,31,67,31,108,31,108,30,54,31,46,31,42,31,83,31,192,31,192,30,219,31,205,31,205,30,67,31,144,31,80,31,204,31,223,31,223,30,224,31,159,31,159,30,7,31,107,31,166,31,100,31,115,31,103,31,156,31,69,31,253,31,76,31,2,31,216,31,210,31,243,31,229,31,57,31,64,31,229,31,147,31,3,31,92,31,191,31,98,31,88,31,64,31,179,31,236,31,38,31,206,31,206,30,167,31,5,31,5,30,203,31,208,31,208,30,191,31,44,31,245,31,90,31,90,30,90,29,90,28,90,27,90,26,194,31,202,31,164,31,66,31,130,31,63,31,9,31,31,31,221,31,221,30,182,31,113,31,113,30,59,31,13,31,73,31,35,31,21,31,108,31,145,31,51,31,209,31,96,31,39,31,116,31,154,31,88,31,148,31,253,31,187,31,227,31,58,31,211,31,136,31,178,31,178,30,126,31,126,30,212,31,212,30,183,31,18,31,63,31,63,30,14,31,212,31,212,30,214,31,242,31,65,31,239,31,34,31,72,31,122,31,122,30,93,31,151,31,111,31,166,31,48,31,48,30,164,31,129,31,118,31,203,31,240,31,114,31,114,30,114,29,69,31,7,31,85,31,39,31,90,31,18,31,85,31,137,31,137,30,172,31,46,31,146,31,189,31,43,31,124,31,12,31,12,30,33,31,210,31,230,31,204,31,127,31,21,31,140,31,168,31,39,31,166,31,16,31,146,31,146,30,146,29,13,31,79,31,79,30,14,31,14,30,225,31,116,31,134,31,134,30,134,29,134,28,64,31,192,31,182,31,73,31,65,31,3,31,3,30,153,31,34,31,34,30,23,31,3,31,17,31,101,31,211,31,11,31,165,31,156,31,50,31,50,30,225,31,81,31,245,31,90,31,64,31,20,31,20,30,134,31,83,31,83,30,242,31,52,31,159,31,113,31,113,30,170,31,170,30,170,29,37,31,195,31,168,31,120,31,28,31,186,31,186,30,97,31,198,31,213,31,253,31,253,30,18,31,20,31,79,31,76,31,246,31,241,31,143,31,169,31,179,31,179,30,157,31,59,31,248,31,10,31,158,31,242,31,185,31,228,31,213,31,202,31,129,31,129,30,99,31,243,31,77,31,77,30,24,31,24,30,207,31,235,31,41,31,138,31,186,31,141,31,119,31,113,31,17,31,118,31,86,31,151,31,56,31,19,31,233,31,37,31,233,31,52,31,52,30,239,31,109,31,200,31,86,31,46,31,175,31,115,31,87,31,25,31,85,31,202,31,69,31,69,30,225,31,225,30,221,31,248,31,27,31,217,31,217,30,220,31,253,31,155,31,155,30,152,31,184,31,127,31,17,31,39,31,39,30,215,31,223,31,59,31,101,31,62,31,62,30,62,29,67,31,114,31,100,31,148,31,99,31,99,30,247,31,101,31,138,31,147,31,173,31,17,31,189,31,2,31,2,30,255,31,88,31,86,31,60,31,60,30,12,31,94,31,141,31,141,30,141,29,89,31,89,30,89,29,89,28,89,27,99,31,60,31,91,31,65,31,150,31,150,30,29,31,9,31,147,31,225,31,225,30,60,31,197,31,197,30,174,31,19,31,19,30,64,31,182,31,13,31,65,31,65,30,95,31,192,31,160,31,151,31,36,31,2,31,76,31,175,31,48,31,48,30,219,31,191,31,85,31,227,31,128,31,153,31,236,31,17,31,134,31,48,31,253,31,21,31,21,30,193,31,193,30,180,31,67,31,154,31,23,31,145,31,137,31,250,31,250,30,113,31,237,31,166,31,230,31,12,31,121,31,227,31,102,31,102,30,247,31,247,30,177,31,143,31,85,31,168,31,40,31,211,31,211,30,81,31,81,30,116,31,116,30,22,31,28,31,234,31,176,31,7,31,184,31,197,31,197,30,197,29,195,31,121,31,175,31,142,31,118,31,125,31,109,31,48,31,48,30,163,31,163,30,163,29,97,31,7,31,82,31,197,31,241,31,47,31,100,31,100,30,66,31,138,31,77,31,205,31,29,31,252,31,219,31,154,31,167,31,201,31,128,31,225,31,225,30,203,31,86,31,244,31,108,31,136,31,250,31,250,30,250,29,152,31,152,30,152,29,152,28,152,27,216,31,143,31,54,31,17,31,222,31,17,31,145,31,65,31,134,31,159,31,159,30,201,31,201,30,201,29,38,31,38,30,53,31,239,31,244,31,213,31,69,31,242,31,174,31,122,31,72,31,14,31,238,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
