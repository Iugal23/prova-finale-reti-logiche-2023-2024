-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 912;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (131,0,0,0,55,0,68,0,82,0,109,0,63,0,188,0,195,0,212,0,159,0,0,0,0,0,52,0,0,0,16,0,0,0,91,0,243,0,0,0,0,0,250,0,149,0,215,0,0,0,226,0,11,0,233,0,196,0,0,0,68,0,0,0,96,0,242,0,0,0,24,0,19,0,53,0,103,0,138,0,247,0,0,0,0,0,227,0,0,0,248,0,0,0,0,0,49,0,74,0,24,0,98,0,0,0,27,0,125,0,247,0,141,0,17,0,59,0,7,0,152,0,0,0,0,0,61,0,15,0,247,0,89,0,202,0,105,0,119,0,0,0,10,0,183,0,108,0,98,0,136,0,14,0,1,0,64,0,144,0,163,0,181,0,220,0,26,0,13,0,191,0,249,0,157,0,165,0,146,0,125,0,91,0,137,0,25,0,229,0,0,0,154,0,0,0,0,0,181,0,0,0,127,0,60,0,0,0,216,0,0,0,0,0,22,0,248,0,166,0,28,0,0,0,166,0,41,0,152,0,107,0,158,0,12,0,0,0,0,0,114,0,217,0,154,0,101,0,90,0,0,0,178,0,106,0,8,0,104,0,195,0,43,0,31,0,243,0,147,0,152,0,231,0,197,0,207,0,234,0,0,0,170,0,58,0,0,0,18,0,5,0,101,0,0,0,25,0,221,0,0,0,7,0,19,0,0,0,61,0,78,0,27,0,179,0,0,0,248,0,110,0,79,0,122,0,46,0,35,0,214,0,0,0,0,0,203,0,127,0,246,0,219,0,3,0,123,0,0,0,0,0,0,0,190,0,162,0,161,0,0,0,0,0,65,0,102,0,189,0,32,0,0,0,166,0,45,0,129,0,230,0,34,0,88,0,181,0,104,0,52,0,237,0,0,0,46,0,172,0,98,0,0,0,89,0,194,0,218,0,243,0,0,0,0,0,105,0,53,0,206,0,0,0,42,0,85,0,124,0,87,0,90,0,137,0,208,0,0,0,0,0,98,0,163,0,240,0,249,0,183,0,212,0,146,0,80,0,0,0,75,0,81,0,71,0,17,0,125,0,38,0,0,0,220,0,63,0,0,0,211,0,84,0,124,0,59,0,0,0,0,0,0,0,77,0,198,0,94,0,66,0,45,0,89,0,172,0,153,0,20,0,83,0,217,0,255,0,52,0,0,0,0,0,95,0,69,0,17,0,137,0,226,0,44,0,0,0,26,0,57,0,223,0,178,0,166,0,150,0,166,0,0,0,46,0,50,0,0,0,20,0,0,0,229,0,0,0,211,0,223,0,1,0,0,0,3,0,0,0,231,0,172,0,0,0,72,0,157,0,243,0,16,0,171,0,202,0,217,0,64,0,18,0,0,0,252,0,153,0,173,0,234,0,2,0,163,0,0,0,1,0,126,0,25,0,243,0,220,0,192,0,0,0,0,0,192,0,118,0,142,0,10,0,243,0,174,0,71,0,94,0,144,0,0,0,88,0,23,0,106,0,238,0,178,0,78,0,145,0,55,0,236,0,88,0,37,0,197,0,80,0,27,0,4,0,137,0,8,0,66,0,0,0,210,0,189,0,108,0,0,0,65,0,27,0,90,0,95,0,141,0,136,0,0,0,148,0,189,0,214,0,74,0,0,0,41,0,202,0,100,0,100,0,0,0,0,0,187,0,134,0,0,0,63,0,95,0,115,0,172,0,217,0,37,0,245,0,245,0,0,0,0,0,158,0,247,0,0,0,167,0,245,0,178,0,132,0,159,0,116,0,227,0,205,0,0,0,149,0,86,0,148,0,218,0,28,0,217,0,166,0,237,0,208,0,0,0,144,0,95,0,10,0,0,0,57,0,3,0,237,0,236,0,121,0,92,0,66,0,0,0,105,0,146,0,17,0,69,0,0,0,0,0,0,0,175,0,189,0,226,0,4,0,0,0,0,0,109,0,170,0,71,0,214,0,113,0,223,0,60,0,22,0,241,0,73,0,137,0,137,0,220,0,0,0,35,0,93,0,122,0,185,0,181,0,145,0,127,0,0,0,223,0,58,0,92,0,105,0,0,0,82,0,239,0,251,0,0,0,0,0,207,0,24,0,167,0,130,0,172,0,0,0,199,0,0,0,11,0,160,0,84,0,0,0,114,0,66,0,251,0,158,0,170,0,145,0,70,0,174,0,143,0,237,0,78,0,27,0,118,0,0,0,0,0,151,0,0,0,0,0,39,0,0,0,130,0,141,0,0,0,0,0,133,0,0,0,239,0,134,0,0,0,0,0,11,0,121,0,209,0,0,0,41,0,106,0,138,0,204,0,175,0,166,0,23,0,143,0,160,0,82,0,227,0,0,0,115,0,0,0,157,0,0,0,181,0,64,0,58,0,0,0,201,0,0,0,103,0,26,0,107,0,118,0,0,0,121,0,157,0,81,0,37,0,216,0,57,0,0,0,249,0,8,0,0,0,92,0,192,0,95,0,7,0,0,0,192,0,201,0,243,0,202,0,242,0,0,0,0,0,110,0,213,0,51,0,129,0,199,0,0,0,37,0,9,0,116,0,0,0,53,0,110,0,196,0,144,0,0,0,234,0,50,0,63,0,0,0,150,0,82,0,126,0,196,0,0,0,149,0,0,0,87,0,0,0,125,0,203,0,117,0,12,0,86,0,2,0,103,0,0,0,125,0,102,0,209,0,190,0,18,0,181,0,0,0,163,0,104,0,87,0,173,0,43,0,0,0,87,0,150,0,0,0,58,0,171,0,96,0,0,0,122,0,0,0,67,0,85,0,64,0,190,0,161,0,24,0,105,0,68,0,64,0,179,0,163,0,0,0,41,0,92,0,9,0,0,0,0,0,75,0,223,0,149,0,255,0,100,0,163,0,70,0,50,0,48,0,254,0,0,0,241,0,0,0,227,0,0,0,158,0,132,0,142,0,0,0,172,0,84,0,61,0,196,0,0,0,0,0,144,0,255,0,0,0,152,0,0,0,29,0,56,0,138,0,123,0,0,0,11,0,83,0,11,0,183,0,57,0,9,0,162,0,240,0,33,0,88,0,0,0,221,0,201,0,206,0,65,0,26,0,119,0,216,0,82,0,240,0,166,0,127,0,99,0,114,0,83,0,186,0,140,0,22,0,76,0,131,0,84,0,113,0,131,0,81,0,231,0,134,0,113,0,109,0,142,0,0,0,47,0,43,0,56,0,215,0,35,0,106,0,250,0,118,0,210,0,0,0,75,0,184,0,112,0,207,0,156,0,88,0,78,0,0,0,0,0,93,0,19,0,0,0,177,0,0,0,169,0,24,0,0,0,0,0,0,0,97,0,0,0,0,0,151,0,0,0,0,0,159,0,234,0,220,0,114,0,129,0,97,0,150,0,149,0,78,0,0,0,209,0,119,0,239,0,0,0,29,0,124,0,0,0,167,0,231,0,188,0,0,0,185,0,0,0,31,0,216,0,0,0,224,0,0,0,7,0,199,0,60,0,88,0,63,0,0,0,0,0,0,0,109,0,206,0,0,0,0,0,167,0,207,0,160,0,12,0,65,0,14,0,233,0,0,0,252,0,17,0,196,0,28,0,159,0,0,0,146,0,151,0,3,0,36,0,181,0,254,0,178,0,137,0,133,0,31,0,146,0,224,0,98,0,182,0,56,0,232,0,169,0,0,0,0,0,80,0,21,0,88,0,0,0,232,0,34,0,220,0,250,0,41,0,112,0,222,0,11,0,128,0,124,0,103,0,111,0,254,0,35,0,59,0,0,0,199,0,19,0,30,0,133,0,114,0,36,0,207,0,189,0,0,0,238,0,86,0,62,0,101,0,138,0,150,0,197,0,0,0,53,0,112,0,126,0,88,0,26,0,255,0,15,0,40,0,0,0,159,0,116,0,84,0,0,0,246,0,0,0,88,0,0,0,0,0,0,0,0,0,87,0,254,0,42,0,0,0,4,0,120,0,194,0,238,0,10,0,0,0,0,0,248,0,69,0,170,0,183,0,155,0,0,0,212,0,0,0,251,0,87,0,90,0,220,0,0,0,75,0,239,0,77,0,132,0,140,0,0,0,71,0,128,0,30,0,151,0,134,0,240,0,145,0,0,0,0,0,41,0,226,0);
signal scenario_full  : scenario_type := (131,31,131,30,55,31,68,31,82,31,109,31,63,31,188,31,195,31,212,31,159,31,159,30,159,29,52,31,52,30,16,31,16,30,91,31,243,31,243,30,243,29,250,31,149,31,215,31,215,30,226,31,11,31,233,31,196,31,196,30,68,31,68,30,96,31,242,31,242,30,24,31,19,31,53,31,103,31,138,31,247,31,247,30,247,29,227,31,227,30,248,31,248,30,248,29,49,31,74,31,24,31,98,31,98,30,27,31,125,31,247,31,141,31,17,31,59,31,7,31,152,31,152,30,152,29,61,31,15,31,247,31,89,31,202,31,105,31,119,31,119,30,10,31,183,31,108,31,98,31,136,31,14,31,1,31,64,31,144,31,163,31,181,31,220,31,26,31,13,31,191,31,249,31,157,31,165,31,146,31,125,31,91,31,137,31,25,31,229,31,229,30,154,31,154,30,154,29,181,31,181,30,127,31,60,31,60,30,216,31,216,30,216,29,22,31,248,31,166,31,28,31,28,30,166,31,41,31,152,31,107,31,158,31,12,31,12,30,12,29,114,31,217,31,154,31,101,31,90,31,90,30,178,31,106,31,8,31,104,31,195,31,43,31,31,31,243,31,147,31,152,31,231,31,197,31,207,31,234,31,234,30,170,31,58,31,58,30,18,31,5,31,101,31,101,30,25,31,221,31,221,30,7,31,19,31,19,30,61,31,78,31,27,31,179,31,179,30,248,31,110,31,79,31,122,31,46,31,35,31,214,31,214,30,214,29,203,31,127,31,246,31,219,31,3,31,123,31,123,30,123,29,123,28,190,31,162,31,161,31,161,30,161,29,65,31,102,31,189,31,32,31,32,30,166,31,45,31,129,31,230,31,34,31,88,31,181,31,104,31,52,31,237,31,237,30,46,31,172,31,98,31,98,30,89,31,194,31,218,31,243,31,243,30,243,29,105,31,53,31,206,31,206,30,42,31,85,31,124,31,87,31,90,31,137,31,208,31,208,30,208,29,98,31,163,31,240,31,249,31,183,31,212,31,146,31,80,31,80,30,75,31,81,31,71,31,17,31,125,31,38,31,38,30,220,31,63,31,63,30,211,31,84,31,124,31,59,31,59,30,59,29,59,28,77,31,198,31,94,31,66,31,45,31,89,31,172,31,153,31,20,31,83,31,217,31,255,31,52,31,52,30,52,29,95,31,69,31,17,31,137,31,226,31,44,31,44,30,26,31,57,31,223,31,178,31,166,31,150,31,166,31,166,30,46,31,50,31,50,30,20,31,20,30,229,31,229,30,211,31,223,31,1,31,1,30,3,31,3,30,231,31,172,31,172,30,72,31,157,31,243,31,16,31,171,31,202,31,217,31,64,31,18,31,18,30,252,31,153,31,173,31,234,31,2,31,163,31,163,30,1,31,126,31,25,31,243,31,220,31,192,31,192,30,192,29,192,31,118,31,142,31,10,31,243,31,174,31,71,31,94,31,144,31,144,30,88,31,23,31,106,31,238,31,178,31,78,31,145,31,55,31,236,31,88,31,37,31,197,31,80,31,27,31,4,31,137,31,8,31,66,31,66,30,210,31,189,31,108,31,108,30,65,31,27,31,90,31,95,31,141,31,136,31,136,30,148,31,189,31,214,31,74,31,74,30,41,31,202,31,100,31,100,31,100,30,100,29,187,31,134,31,134,30,63,31,95,31,115,31,172,31,217,31,37,31,245,31,245,31,245,30,245,29,158,31,247,31,247,30,167,31,245,31,178,31,132,31,159,31,116,31,227,31,205,31,205,30,149,31,86,31,148,31,218,31,28,31,217,31,166,31,237,31,208,31,208,30,144,31,95,31,10,31,10,30,57,31,3,31,237,31,236,31,121,31,92,31,66,31,66,30,105,31,146,31,17,31,69,31,69,30,69,29,69,28,175,31,189,31,226,31,4,31,4,30,4,29,109,31,170,31,71,31,214,31,113,31,223,31,60,31,22,31,241,31,73,31,137,31,137,31,220,31,220,30,35,31,93,31,122,31,185,31,181,31,145,31,127,31,127,30,223,31,58,31,92,31,105,31,105,30,82,31,239,31,251,31,251,30,251,29,207,31,24,31,167,31,130,31,172,31,172,30,199,31,199,30,11,31,160,31,84,31,84,30,114,31,66,31,251,31,158,31,170,31,145,31,70,31,174,31,143,31,237,31,78,31,27,31,118,31,118,30,118,29,151,31,151,30,151,29,39,31,39,30,130,31,141,31,141,30,141,29,133,31,133,30,239,31,134,31,134,30,134,29,11,31,121,31,209,31,209,30,41,31,106,31,138,31,204,31,175,31,166,31,23,31,143,31,160,31,82,31,227,31,227,30,115,31,115,30,157,31,157,30,181,31,64,31,58,31,58,30,201,31,201,30,103,31,26,31,107,31,118,31,118,30,121,31,157,31,81,31,37,31,216,31,57,31,57,30,249,31,8,31,8,30,92,31,192,31,95,31,7,31,7,30,192,31,201,31,243,31,202,31,242,31,242,30,242,29,110,31,213,31,51,31,129,31,199,31,199,30,37,31,9,31,116,31,116,30,53,31,110,31,196,31,144,31,144,30,234,31,50,31,63,31,63,30,150,31,82,31,126,31,196,31,196,30,149,31,149,30,87,31,87,30,125,31,203,31,117,31,12,31,86,31,2,31,103,31,103,30,125,31,102,31,209,31,190,31,18,31,181,31,181,30,163,31,104,31,87,31,173,31,43,31,43,30,87,31,150,31,150,30,58,31,171,31,96,31,96,30,122,31,122,30,67,31,85,31,64,31,190,31,161,31,24,31,105,31,68,31,64,31,179,31,163,31,163,30,41,31,92,31,9,31,9,30,9,29,75,31,223,31,149,31,255,31,100,31,163,31,70,31,50,31,48,31,254,31,254,30,241,31,241,30,227,31,227,30,158,31,132,31,142,31,142,30,172,31,84,31,61,31,196,31,196,30,196,29,144,31,255,31,255,30,152,31,152,30,29,31,56,31,138,31,123,31,123,30,11,31,83,31,11,31,183,31,57,31,9,31,162,31,240,31,33,31,88,31,88,30,221,31,201,31,206,31,65,31,26,31,119,31,216,31,82,31,240,31,166,31,127,31,99,31,114,31,83,31,186,31,140,31,22,31,76,31,131,31,84,31,113,31,131,31,81,31,231,31,134,31,113,31,109,31,142,31,142,30,47,31,43,31,56,31,215,31,35,31,106,31,250,31,118,31,210,31,210,30,75,31,184,31,112,31,207,31,156,31,88,31,78,31,78,30,78,29,93,31,19,31,19,30,177,31,177,30,169,31,24,31,24,30,24,29,24,28,97,31,97,30,97,29,151,31,151,30,151,29,159,31,234,31,220,31,114,31,129,31,97,31,150,31,149,31,78,31,78,30,209,31,119,31,239,31,239,30,29,31,124,31,124,30,167,31,231,31,188,31,188,30,185,31,185,30,31,31,216,31,216,30,224,31,224,30,7,31,199,31,60,31,88,31,63,31,63,30,63,29,63,28,109,31,206,31,206,30,206,29,167,31,207,31,160,31,12,31,65,31,14,31,233,31,233,30,252,31,17,31,196,31,28,31,159,31,159,30,146,31,151,31,3,31,36,31,181,31,254,31,178,31,137,31,133,31,31,31,146,31,224,31,98,31,182,31,56,31,232,31,169,31,169,30,169,29,80,31,21,31,88,31,88,30,232,31,34,31,220,31,250,31,41,31,112,31,222,31,11,31,128,31,124,31,103,31,111,31,254,31,35,31,59,31,59,30,199,31,19,31,30,31,133,31,114,31,36,31,207,31,189,31,189,30,238,31,86,31,62,31,101,31,138,31,150,31,197,31,197,30,53,31,112,31,126,31,88,31,26,31,255,31,15,31,40,31,40,30,159,31,116,31,84,31,84,30,246,31,246,30,88,31,88,30,88,29,88,28,88,27,87,31,254,31,42,31,42,30,4,31,120,31,194,31,238,31,10,31,10,30,10,29,248,31,69,31,170,31,183,31,155,31,155,30,212,31,212,30,251,31,87,31,90,31,220,31,220,30,75,31,239,31,77,31,132,31,140,31,140,30,71,31,128,31,30,31,151,31,134,31,240,31,145,31,145,30,145,29,41,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
