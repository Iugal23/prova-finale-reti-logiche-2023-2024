-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_392 is
end project_tb_392;

architecture project_tb_arch_392 of project_tb_392 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 929;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (187,0,21,0,142,0,40,0,192,0,3,0,134,0,4,0,0,0,0,0,0,0,0,0,138,0,208,0,53,0,162,0,223,0,80,0,247,0,0,0,210,0,0,0,39,0,188,0,0,0,6,0,209,0,60,0,37,0,81,0,241,0,192,0,183,0,24,0,0,0,128,0,52,0,0,0,229,0,0,0,115,0,159,0,48,0,166,0,240,0,200,0,104,0,117,0,31,0,121,0,184,0,214,0,37,0,0,0,22,0,241,0,147,0,174,0,168,0,0,0,246,0,113,0,71,0,0,0,120,0,53,0,184,0,23,0,156,0,95,0,147,0,154,0,78,0,255,0,192,0,78,0,71,0,108,0,127,0,60,0,242,0,124,0,19,0,0,0,222,0,53,0,0,0,0,0,0,0,147,0,0,0,252,0,183,0,179,0,0,0,60,0,197,0,0,0,0,0,28,0,208,0,86,0,73,0,0,0,233,0,154,0,42,0,26,0,160,0,69,0,148,0,0,0,196,0,97,0,145,0,141,0,50,0,0,0,122,0,172,0,212,0,52,0,0,0,37,0,14,0,0,0,244,0,0,0,20,0,0,0,0,0,157,0,201,0,0,0,82,0,202,0,127,0,36,0,28,0,169,0,161,0,122,0,234,0,151,0,149,0,146,0,252,0,0,0,64,0,90,0,215,0,94,0,195,0,0,0,15,0,89,0,7,0,217,0,93,0,0,0,147,0,220,0,75,0,201,0,105,0,197,0,0,0,144,0,94,0,179,0,236,0,196,0,96,0,0,0,30,0,134,0,231,0,0,0,0,0,0,0,50,0,224,0,64,0,209,0,255,0,73,0,0,0,90,0,11,0,169,0,0,0,231,0,142,0,134,0,103,0,0,0,0,0,227,0,107,0,174,0,111,0,197,0,105,0,172,0,145,0,83,0,200,0,25,0,153,0,61,0,137,0,101,0,124,0,149,0,109,0,124,0,130,0,51,0,14,0,75,0,177,0,64,0,200,0,0,0,82,0,221,0,154,0,156,0,165,0,106,0,106,0,106,0,9,0,56,0,70,0,0,0,152,0,9,0,184,0,179,0,72,0,117,0,177,0,11,0,0,0,45,0,20,0,182,0,227,0,134,0,119,0,161,0,215,0,38,0,0,0,238,0,92,0,0,0,0,0,0,0,248,0,0,0,16,0,191,0,194,0,124,0,0,0,18,0,130,0,251,0,160,0,81,0,0,0,31,0,251,0,46,0,230,0,0,0,129,0,0,0,6,0,194,0,0,0,0,0,177,0,151,0,0,0,235,0,74,0,14,0,182,0,154,0,23,0,0,0,65,0,109,0,251,0,34,0,0,0,186,0,0,0,211,0,182,0,65,0,178,0,0,0,91,0,187,0,48,0,35,0,55,0,53,0,0,0,114,0,3,0,245,0,86,0,174,0,0,0,93,0,221,0,72,0,96,0,122,0,77,0,98,0,0,0,1,0,105,0,83,0,5,0,0,0,96,0,105,0,193,0,0,0,211,0,128,0,149,0,140,0,125,0,0,0,170,0,249,0,141,0,0,0,136,0,43,0,0,0,135,0,128,0,107,0,181,0,168,0,104,0,107,0,169,0,121,0,182,0,147,0,192,0,32,0,66,0,193,0,227,0,167,0,0,0,198,0,143,0,0,0,50,0,0,0,45,0,107,0,192,0,127,0,170,0,84,0,0,0,103,0,210,0,0,0,221,0,55,0,115,0,246,0,180,0,97,0,0,0,35,0,0,0,0,0,62,0,31,0,28,0,247,0,193,0,139,0,0,0,0,0,221,0,40,0,229,0,212,0,64,0,134,0,44,0,0,0,0,0,69,0,0,0,235,0,121,0,253,0,138,0,122,0,156,0,33,0,52,0,0,0,0,0,91,0,33,0,111,0,0,0,242,0,0,0,235,0,0,0,48,0,143,0,3,0,0,0,0,0,138,0,222,0,0,0,241,0,122,0,123,0,50,0,101,0,66,0,0,0,2,0,56,0,132,0,239,0,0,0,134,0,0,0,0,0,117,0,227,0,0,0,33,0,148,0,213,0,31,0,91,0,251,0,0,0,187,0,0,0,229,0,0,0,200,0,74,0,202,0,82,0,0,0,49,0,175,0,102,0,28,0,103,0,170,0,34,0,172,0,0,0,132,0,206,0,250,0,47,0,135,0,72,0,0,0,174,0,0,0,0,0,0,0,118,0,0,0,125,0,42,0,117,0,60,0,0,0,170,0,155,0,204,0,186,0,92,0,239,0,181,0,164,0,34,0,249,0,60,0,61,0,0,0,104,0,125,0,219,0,183,0,132,0,225,0,22,0,93,0,79,0,35,0,199,0,201,0,0,0,70,0,246,0,0,0,213,0,106,0,111,0,4,0,80,0,42,0,112,0,0,0,46,0,0,0,0,0,220,0,0,0,0,0,174,0,29,0,212,0,132,0,0,0,222,0,0,0,40,0,127,0,24,0,73,0,18,0,59,0,146,0,194,0,42,0,214,0,160,0,172,0,215,0,200,0,142,0,228,0,199,0,47,0,0,0,0,0,153,0,108,0,90,0,130,0,46,0,246,0,180,0,97,0,0,0,4,0,0,0,165,0,68,0,101,0,131,0,0,0,14,0,26,0,117,0,225,0,232,0,186,0,90,0,231,0,19,0,131,0,219,0,0,0,67,0,43,0,191,0,79,0,111,0,137,0,143,0,237,0,118,0,216,0,176,0,243,0,122,0,204,0,0,0,2,0,236,0,138,0,57,0,148,0,0,0,142,0,243,0,193,0,0,0,160,0,0,0,217,0,215,0,155,0,0,0,0,0,244,0,190,0,140,0,26,0,26,0,64,0,204,0,0,0,0,0,231,0,29,0,124,0,210,0,135,0,22,0,86,0,0,0,60,0,182,0,176,0,0,0,85,0,29,0,223,0,159,0,0,0,121,0,23,0,198,0,87,0,0,0,0,0,200,0,0,0,0,0,123,0,4,0,42,0,0,0,116,0,147,0,101,0,0,0,172,0,0,0,18,0,36,0,4,0,129,0,176,0,0,0,176,0,230,0,96,0,166,0,114,0,0,0,244,0,47,0,11,0,28,0,0,0,43,0,119,0,0,0,138,0,0,0,134,0,237,0,96,0,0,0,51,0,222,0,4,0,204,0,198,0,182,0,231,0,0,0,91,0,71,0,41,0,137,0,172,0,138,0,0,0,110,0,130,0,208,0,147,0,189,0,12,0,0,0,0,0,150,0,131,0,189,0,158,0,234,0,58,0,252,0,77,0,151,0,109,0,195,0,0,0,198,0,94,0,199,0,122,0,187,0,176,0,0,0,94,0,0,0,10,0,15,0,203,0,0,0,163,0,240,0,0,0,32,0,57,0,0,0,0,0,212,0,176,0,0,0,0,0,212,0,125,0,0,0,209,0,33,0,240,0,246,0,130,0,245,0,209,0,5,0,102,0,39,0,186,0,10,0,196,0,68,0,87,0,253,0,237,0,0,0,0,0,0,0,255,0,83,0,147,0,16,0,0,0,0,0,212,0,87,0,130,0,202,0,122,0,171,0,198,0,0,0,218,0,0,0,193,0,0,0,106,0,0,0,55,0,177,0,106,0,0,0,0,0,216,0,142,0,253,0,228,0,121,0,207,0,119,0,72,0,200,0,172,0,164,0,0,0,111,0,63,0,0,0,114,0,12,0,0,0,147,0,11,0,163,0,187,0,114,0,29,0,5,0,215,0,118,0,141,0,54,0,217,0,112,0,246,0,147,0,93,0,244,0,95,0,87,0,26,0,169,0,129,0,3,0,44,0,0,0,0,0,2,0,211,0,187,0,199,0,78,0,0,0,0,0,133,0,0,0,0,0,229,0,0,0,134,0,0,0,4,0,136,0,173,0,24,0,51,0,56,0,237,0,156,0,2,0,169,0,183,0,0,0,0,0,112,0,114,0,77,0,228,0,23,0,25,0,62,0,95,0,102,0,34,0,154,0,44,0,13,0,0,0,60,0,180,0,0,0,0,0,23,0,116,0,99,0,210,0,0,0,46,0,44,0,215,0,192,0,232,0,65,0,250,0,8,0,133,0,0,0,21,0,244,0,83,0,59,0,0,0,45,0,65,0,132,0,82,0,210,0,201,0,7,0,198,0,0,0,38,0,52,0,122,0,0,0,87,0);
signal scenario_full  : scenario_type := (187,31,21,31,142,31,40,31,192,31,3,31,134,31,4,31,4,30,4,29,4,28,4,27,138,31,208,31,53,31,162,31,223,31,80,31,247,31,247,30,210,31,210,30,39,31,188,31,188,30,6,31,209,31,60,31,37,31,81,31,241,31,192,31,183,31,24,31,24,30,128,31,52,31,52,30,229,31,229,30,115,31,159,31,48,31,166,31,240,31,200,31,104,31,117,31,31,31,121,31,184,31,214,31,37,31,37,30,22,31,241,31,147,31,174,31,168,31,168,30,246,31,113,31,71,31,71,30,120,31,53,31,184,31,23,31,156,31,95,31,147,31,154,31,78,31,255,31,192,31,78,31,71,31,108,31,127,31,60,31,242,31,124,31,19,31,19,30,222,31,53,31,53,30,53,29,53,28,147,31,147,30,252,31,183,31,179,31,179,30,60,31,197,31,197,30,197,29,28,31,208,31,86,31,73,31,73,30,233,31,154,31,42,31,26,31,160,31,69,31,148,31,148,30,196,31,97,31,145,31,141,31,50,31,50,30,122,31,172,31,212,31,52,31,52,30,37,31,14,31,14,30,244,31,244,30,20,31,20,30,20,29,157,31,201,31,201,30,82,31,202,31,127,31,36,31,28,31,169,31,161,31,122,31,234,31,151,31,149,31,146,31,252,31,252,30,64,31,90,31,215,31,94,31,195,31,195,30,15,31,89,31,7,31,217,31,93,31,93,30,147,31,220,31,75,31,201,31,105,31,197,31,197,30,144,31,94,31,179,31,236,31,196,31,96,31,96,30,30,31,134,31,231,31,231,30,231,29,231,28,50,31,224,31,64,31,209,31,255,31,73,31,73,30,90,31,11,31,169,31,169,30,231,31,142,31,134,31,103,31,103,30,103,29,227,31,107,31,174,31,111,31,197,31,105,31,172,31,145,31,83,31,200,31,25,31,153,31,61,31,137,31,101,31,124,31,149,31,109,31,124,31,130,31,51,31,14,31,75,31,177,31,64,31,200,31,200,30,82,31,221,31,154,31,156,31,165,31,106,31,106,31,106,31,9,31,56,31,70,31,70,30,152,31,9,31,184,31,179,31,72,31,117,31,177,31,11,31,11,30,45,31,20,31,182,31,227,31,134,31,119,31,161,31,215,31,38,31,38,30,238,31,92,31,92,30,92,29,92,28,248,31,248,30,16,31,191,31,194,31,124,31,124,30,18,31,130,31,251,31,160,31,81,31,81,30,31,31,251,31,46,31,230,31,230,30,129,31,129,30,6,31,194,31,194,30,194,29,177,31,151,31,151,30,235,31,74,31,14,31,182,31,154,31,23,31,23,30,65,31,109,31,251,31,34,31,34,30,186,31,186,30,211,31,182,31,65,31,178,31,178,30,91,31,187,31,48,31,35,31,55,31,53,31,53,30,114,31,3,31,245,31,86,31,174,31,174,30,93,31,221,31,72,31,96,31,122,31,77,31,98,31,98,30,1,31,105,31,83,31,5,31,5,30,96,31,105,31,193,31,193,30,211,31,128,31,149,31,140,31,125,31,125,30,170,31,249,31,141,31,141,30,136,31,43,31,43,30,135,31,128,31,107,31,181,31,168,31,104,31,107,31,169,31,121,31,182,31,147,31,192,31,32,31,66,31,193,31,227,31,167,31,167,30,198,31,143,31,143,30,50,31,50,30,45,31,107,31,192,31,127,31,170,31,84,31,84,30,103,31,210,31,210,30,221,31,55,31,115,31,246,31,180,31,97,31,97,30,35,31,35,30,35,29,62,31,31,31,28,31,247,31,193,31,139,31,139,30,139,29,221,31,40,31,229,31,212,31,64,31,134,31,44,31,44,30,44,29,69,31,69,30,235,31,121,31,253,31,138,31,122,31,156,31,33,31,52,31,52,30,52,29,91,31,33,31,111,31,111,30,242,31,242,30,235,31,235,30,48,31,143,31,3,31,3,30,3,29,138,31,222,31,222,30,241,31,122,31,123,31,50,31,101,31,66,31,66,30,2,31,56,31,132,31,239,31,239,30,134,31,134,30,134,29,117,31,227,31,227,30,33,31,148,31,213,31,31,31,91,31,251,31,251,30,187,31,187,30,229,31,229,30,200,31,74,31,202,31,82,31,82,30,49,31,175,31,102,31,28,31,103,31,170,31,34,31,172,31,172,30,132,31,206,31,250,31,47,31,135,31,72,31,72,30,174,31,174,30,174,29,174,28,118,31,118,30,125,31,42,31,117,31,60,31,60,30,170,31,155,31,204,31,186,31,92,31,239,31,181,31,164,31,34,31,249,31,60,31,61,31,61,30,104,31,125,31,219,31,183,31,132,31,225,31,22,31,93,31,79,31,35,31,199,31,201,31,201,30,70,31,246,31,246,30,213,31,106,31,111,31,4,31,80,31,42,31,112,31,112,30,46,31,46,30,46,29,220,31,220,30,220,29,174,31,29,31,212,31,132,31,132,30,222,31,222,30,40,31,127,31,24,31,73,31,18,31,59,31,146,31,194,31,42,31,214,31,160,31,172,31,215,31,200,31,142,31,228,31,199,31,47,31,47,30,47,29,153,31,108,31,90,31,130,31,46,31,246,31,180,31,97,31,97,30,4,31,4,30,165,31,68,31,101,31,131,31,131,30,14,31,26,31,117,31,225,31,232,31,186,31,90,31,231,31,19,31,131,31,219,31,219,30,67,31,43,31,191,31,79,31,111,31,137,31,143,31,237,31,118,31,216,31,176,31,243,31,122,31,204,31,204,30,2,31,236,31,138,31,57,31,148,31,148,30,142,31,243,31,193,31,193,30,160,31,160,30,217,31,215,31,155,31,155,30,155,29,244,31,190,31,140,31,26,31,26,31,64,31,204,31,204,30,204,29,231,31,29,31,124,31,210,31,135,31,22,31,86,31,86,30,60,31,182,31,176,31,176,30,85,31,29,31,223,31,159,31,159,30,121,31,23,31,198,31,87,31,87,30,87,29,200,31,200,30,200,29,123,31,4,31,42,31,42,30,116,31,147,31,101,31,101,30,172,31,172,30,18,31,36,31,4,31,129,31,176,31,176,30,176,31,230,31,96,31,166,31,114,31,114,30,244,31,47,31,11,31,28,31,28,30,43,31,119,31,119,30,138,31,138,30,134,31,237,31,96,31,96,30,51,31,222,31,4,31,204,31,198,31,182,31,231,31,231,30,91,31,71,31,41,31,137,31,172,31,138,31,138,30,110,31,130,31,208,31,147,31,189,31,12,31,12,30,12,29,150,31,131,31,189,31,158,31,234,31,58,31,252,31,77,31,151,31,109,31,195,31,195,30,198,31,94,31,199,31,122,31,187,31,176,31,176,30,94,31,94,30,10,31,15,31,203,31,203,30,163,31,240,31,240,30,32,31,57,31,57,30,57,29,212,31,176,31,176,30,176,29,212,31,125,31,125,30,209,31,33,31,240,31,246,31,130,31,245,31,209,31,5,31,102,31,39,31,186,31,10,31,196,31,68,31,87,31,253,31,237,31,237,30,237,29,237,28,255,31,83,31,147,31,16,31,16,30,16,29,212,31,87,31,130,31,202,31,122,31,171,31,198,31,198,30,218,31,218,30,193,31,193,30,106,31,106,30,55,31,177,31,106,31,106,30,106,29,216,31,142,31,253,31,228,31,121,31,207,31,119,31,72,31,200,31,172,31,164,31,164,30,111,31,63,31,63,30,114,31,12,31,12,30,147,31,11,31,163,31,187,31,114,31,29,31,5,31,215,31,118,31,141,31,54,31,217,31,112,31,246,31,147,31,93,31,244,31,95,31,87,31,26,31,169,31,129,31,3,31,44,31,44,30,44,29,2,31,211,31,187,31,199,31,78,31,78,30,78,29,133,31,133,30,133,29,229,31,229,30,134,31,134,30,4,31,136,31,173,31,24,31,51,31,56,31,237,31,156,31,2,31,169,31,183,31,183,30,183,29,112,31,114,31,77,31,228,31,23,31,25,31,62,31,95,31,102,31,34,31,154,31,44,31,13,31,13,30,60,31,180,31,180,30,180,29,23,31,116,31,99,31,210,31,210,30,46,31,44,31,215,31,192,31,232,31,65,31,250,31,8,31,133,31,133,30,21,31,244,31,83,31,59,31,59,30,45,31,65,31,132,31,82,31,210,31,201,31,7,31,198,31,198,30,38,31,52,31,122,31,122,30,87,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
