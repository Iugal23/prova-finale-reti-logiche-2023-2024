-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_663 is
end project_tb_663;

architecture project_tb_arch_663 of project_tb_663 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 492;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (198,0,235,0,32,0,0,0,0,0,88,0,29,0,92,0,207,0,0,0,161,0,99,0,153,0,69,0,230,0,0,0,202,0,156,0,243,0,254,0,76,0,108,0,90,0,227,0,87,0,128,0,213,0,42,0,71,0,99,0,17,0,2,0,107,0,100,0,156,0,125,0,0,0,31,0,90,0,76,0,242,0,180,0,62,0,0,0,0,0,154,0,163,0,217,0,48,0,202,0,178,0,235,0,161,0,105,0,156,0,228,0,0,0,0,0,217,0,0,0,149,0,18,0,0,0,0,0,0,0,199,0,246,0,45,0,162,0,117,0,0,0,0,0,243,0,188,0,71,0,0,0,102,0,237,0,0,0,0,0,62,0,27,0,94,0,41,0,0,0,0,0,79,0,54,0,234,0,222,0,0,0,119,0,237,0,95,0,2,0,178,0,33,0,0,0,135,0,0,0,0,0,33,0,70,0,235,0,0,0,19,0,88,0,84,0,0,0,211,0,48,0,0,0,0,0,17,0,15,0,5,0,0,0,0,0,24,0,101,0,232,0,146,0,0,0,219,0,0,0,103,0,170,0,139,0,9,0,0,0,0,0,0,0,27,0,189,0,0,0,183,0,0,0,116,0,145,0,161,0,0,0,18,0,0,0,219,0,254,0,149,0,142,0,29,0,221,0,126,0,46,0,249,0,237,0,179,0,182,0,100,0,0,0,0,0,0,0,186,0,88,0,0,0,23,0,100,0,43,0,242,0,0,0,0,0,0,0,0,0,188,0,18,0,144,0,0,0,2,0,198,0,0,0,0,0,37,0,214,0,162,0,47,0,147,0,243,0,67,0,9,0,231,0,236,0,203,0,45,0,250,0,0,0,200,0,105,0,165,0,183,0,124,0,152,0,52,0,113,0,148,0,244,0,140,0,0,0,0,0,0,0,15,0,179,0,0,0,29,0,106,0,0,0,195,0,176,0,52,0,168,0,0,0,139,0,121,0,120,0,103,0,115,0,220,0,157,0,191,0,14,0,44,0,75,0,12,0,210,0,207,0,61,0,163,0,184,0,0,0,0,0,215,0,231,0,208,0,165,0,185,0,130,0,8,0,0,0,149,0,46,0,108,0,0,0,123,0,245,0,110,0,0,0,156,0,0,0,79,0,52,0,153,0,0,0,116,0,143,0,209,0,181,0,171,0,203,0,213,0,162,0,26,0,50,0,13,0,207,0,86,0,96,0,205,0,193,0,207,0,21,0,0,0,0,0,0,0,0,0,37,0,254,0,194,0,138,0,45,0,211,0,140,0,198,0,188,0,0,0,0,0,0,0,24,0,170,0,95,0,151,0,211,0,211,0,177,0,48,0,184,0,145,0,162,0,52,0,95,0,0,0,51,0,0,0,227,0,209,0,0,0,111,0,74,0,142,0,238,0,150,0,0,0,0,0,7,0,0,0,191,0,0,0,202,0,153,0,70,0,70,0,33,0,240,0,0,0,0,0,167,0,24,0,42,0,20,0,219,0,8,0,108,0,143,0,216,0,176,0,109,0,174,0,193,0,0,0,147,0,38,0,0,0,55,0,0,0,0,0,203,0,174,0,0,0,78,0,248,0,37,0,10,0,215,0,0,0,237,0,0,0,243,0,83,0,0,0,0,0,137,0,85,0,240,0,157,0,0,0,84,0,215,0,0,0,179,0,133,0,233,0,9,0,0,0,106,0,0,0,39,0,20,0,174,0,0,0,61,0,104,0,71,0,20,0,78,0,23,0,199,0,205,0,87,0,2,0,161,0,39,0,200,0,190,0,168,0,104,0,0,0,159,0,0,0,148,0,213,0,154,0,233,0,186,0,254,0,114,0,198,0,116,0,0,0,0,0,26,0,31,0,197,0,74,0,134,0,65,0,20,0,95,0,3,0,49,0,10,0,122,0,205,0,0,0,242,0,218,0,140,0,130,0,95,0,217,0,180,0,94,0,227,0,237,0,0,0,160,0,235,0,101,0,0,0,136,0,255,0,110,0,46,0,54,0,242,0,51,0,175,0,86,0,209,0,0,0,0,0,66,0,87,0,54,0,131,0,0,0,237,0,248,0,0,0,253,0,0,0,147,0,21,0,120,0,222,0,0,0,197,0,0,0,249,0,0,0,95,0,0,0,15,0,0,0,69,0,0,0,159,0,87,0,35,0,111,0,0,0,163,0,118,0,3,0,0,0,225,0,91,0,75,0);
signal scenario_full  : scenario_type := (198,31,235,31,32,31,32,30,32,29,88,31,29,31,92,31,207,31,207,30,161,31,99,31,153,31,69,31,230,31,230,30,202,31,156,31,243,31,254,31,76,31,108,31,90,31,227,31,87,31,128,31,213,31,42,31,71,31,99,31,17,31,2,31,107,31,100,31,156,31,125,31,125,30,31,31,90,31,76,31,242,31,180,31,62,31,62,30,62,29,154,31,163,31,217,31,48,31,202,31,178,31,235,31,161,31,105,31,156,31,228,31,228,30,228,29,217,31,217,30,149,31,18,31,18,30,18,29,18,28,199,31,246,31,45,31,162,31,117,31,117,30,117,29,243,31,188,31,71,31,71,30,102,31,237,31,237,30,237,29,62,31,27,31,94,31,41,31,41,30,41,29,79,31,54,31,234,31,222,31,222,30,119,31,237,31,95,31,2,31,178,31,33,31,33,30,135,31,135,30,135,29,33,31,70,31,235,31,235,30,19,31,88,31,84,31,84,30,211,31,48,31,48,30,48,29,17,31,15,31,5,31,5,30,5,29,24,31,101,31,232,31,146,31,146,30,219,31,219,30,103,31,170,31,139,31,9,31,9,30,9,29,9,28,27,31,189,31,189,30,183,31,183,30,116,31,145,31,161,31,161,30,18,31,18,30,219,31,254,31,149,31,142,31,29,31,221,31,126,31,46,31,249,31,237,31,179,31,182,31,100,31,100,30,100,29,100,28,186,31,88,31,88,30,23,31,100,31,43,31,242,31,242,30,242,29,242,28,242,27,188,31,18,31,144,31,144,30,2,31,198,31,198,30,198,29,37,31,214,31,162,31,47,31,147,31,243,31,67,31,9,31,231,31,236,31,203,31,45,31,250,31,250,30,200,31,105,31,165,31,183,31,124,31,152,31,52,31,113,31,148,31,244,31,140,31,140,30,140,29,140,28,15,31,179,31,179,30,29,31,106,31,106,30,195,31,176,31,52,31,168,31,168,30,139,31,121,31,120,31,103,31,115,31,220,31,157,31,191,31,14,31,44,31,75,31,12,31,210,31,207,31,61,31,163,31,184,31,184,30,184,29,215,31,231,31,208,31,165,31,185,31,130,31,8,31,8,30,149,31,46,31,108,31,108,30,123,31,245,31,110,31,110,30,156,31,156,30,79,31,52,31,153,31,153,30,116,31,143,31,209,31,181,31,171,31,203,31,213,31,162,31,26,31,50,31,13,31,207,31,86,31,96,31,205,31,193,31,207,31,21,31,21,30,21,29,21,28,21,27,37,31,254,31,194,31,138,31,45,31,211,31,140,31,198,31,188,31,188,30,188,29,188,28,24,31,170,31,95,31,151,31,211,31,211,31,177,31,48,31,184,31,145,31,162,31,52,31,95,31,95,30,51,31,51,30,227,31,209,31,209,30,111,31,74,31,142,31,238,31,150,31,150,30,150,29,7,31,7,30,191,31,191,30,202,31,153,31,70,31,70,31,33,31,240,31,240,30,240,29,167,31,24,31,42,31,20,31,219,31,8,31,108,31,143,31,216,31,176,31,109,31,174,31,193,31,193,30,147,31,38,31,38,30,55,31,55,30,55,29,203,31,174,31,174,30,78,31,248,31,37,31,10,31,215,31,215,30,237,31,237,30,243,31,83,31,83,30,83,29,137,31,85,31,240,31,157,31,157,30,84,31,215,31,215,30,179,31,133,31,233,31,9,31,9,30,106,31,106,30,39,31,20,31,174,31,174,30,61,31,104,31,71,31,20,31,78,31,23,31,199,31,205,31,87,31,2,31,161,31,39,31,200,31,190,31,168,31,104,31,104,30,159,31,159,30,148,31,213,31,154,31,233,31,186,31,254,31,114,31,198,31,116,31,116,30,116,29,26,31,31,31,197,31,74,31,134,31,65,31,20,31,95,31,3,31,49,31,10,31,122,31,205,31,205,30,242,31,218,31,140,31,130,31,95,31,217,31,180,31,94,31,227,31,237,31,237,30,160,31,235,31,101,31,101,30,136,31,255,31,110,31,46,31,54,31,242,31,51,31,175,31,86,31,209,31,209,30,209,29,66,31,87,31,54,31,131,31,131,30,237,31,248,31,248,30,253,31,253,30,147,31,21,31,120,31,222,31,222,30,197,31,197,30,249,31,249,30,95,31,95,30,15,31,15,30,69,31,69,30,159,31,87,31,35,31,111,31,111,30,163,31,118,31,3,31,3,30,225,31,91,31,75,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
