-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 762;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (235,0,93,0,213,0,227,0,140,0,36,0,219,0,23,0,148,0,14,0,0,0,211,0,0,0,21,0,10,0,159,0,152,0,80,0,218,0,112,0,107,0,224,0,95,0,0,0,76,0,50,0,0,0,44,0,28,0,0,0,226,0,134,0,0,0,144,0,14,0,148,0,175,0,55,0,0,0,219,0,18,0,0,0,97,0,232,0,12,0,154,0,82,0,107,0,155,0,20,0,94,0,210,0,0,0,244,0,0,0,116,0,35,0,203,0,101,0,0,0,207,0,0,0,144,0,220,0,0,0,10,0,95,0,186,0,168,0,0,0,57,0,0,0,0,0,0,0,16,0,216,0,102,0,115,0,97,0,46,0,206,0,0,0,0,0,196,0,97,0,140,0,37,0,172,0,44,0,100,0,64,0,65,0,0,0,0,0,0,0,213,0,34,0,84,0,96,0,81,0,11,0,99,0,194,0,0,0,81,0,0,0,0,0,201,0,0,0,0,0,82,0,205,0,252,0,180,0,96,0,76,0,121,0,133,0,0,0,206,0,80,0,0,0,0,0,0,0,76,0,38,0,186,0,152,0,18,0,220,0,89,0,130,0,173,0,153,0,98,0,86,0,192,0,108,0,178,0,0,0,251,0,157,0,154,0,0,0,0,0,86,0,118,0,0,0,0,0,226,0,0,0,47,0,28,0,73,0,0,0,61,0,204,0,104,0,0,0,55,0,214,0,98,0,0,0,126,0,0,0,237,0,74,0,79,0,112,0,0,0,8,0,212,0,8,0,0,0,30,0,233,0,177,0,84,0,62,0,63,0,177,0,166,0,73,0,0,0,74,0,122,0,202,0,144,0,0,0,0,0,0,0,162,0,50,0,164,0,231,0,0,0,34,0,193,0,238,0,50,0,180,0,215,0,218,0,0,0,24,0,0,0,103,0,0,0,0,0,250,0,0,0,198,0,37,0,106,0,165,0,0,0,125,0,161,0,37,0,43,0,44,0,14,0,61,0,23,0,58,0,0,0,252,0,253,0,34,0,0,0,0,0,185,0,8,0,0,0,47,0,34,0,216,0,60,0,218,0,0,0,10,0,199,0,136,0,158,0,0,0,56,0,87,0,71,0,95,0,107,0,216,0,92,0,127,0,171,0,0,0,154,0,35,0,0,0,83,0,122,0,64,0,161,0,83,0,86,0,75,0,93,0,0,0,252,0,0,0,89,0,64,0,0,0,0,0,81,0,111,0,23,0,170,0,61,0,31,0,5,0,191,0,96,0,45,0,149,0,0,0,0,0,0,0,211,0,125,0,0,0,252,0,57,0,60,0,0,0,119,0,207,0,2,0,0,0,71,0,84,0,198,0,215,0,173,0,188,0,194,0,0,0,119,0,210,0,183,0,0,0,25,0,28,0,0,0,194,0,0,0,90,0,64,0,0,0,29,0,37,0,0,0,218,0,177,0,199,0,212,0,24,0,168,0,128,0,26,0,100,0,73,0,231,0,0,0,97,0,59,0,0,0,2,0,0,0,0,0,0,0,120,0,54,0,76,0,7,0,151,0,76,0,197,0,143,0,0,0,213,0,103,0,149,0,36,0,205,0,125,0,0,0,0,0,179,0,0,0,132,0,49,0,88,0,134,0,240,0,16,0,0,0,0,0,187,0,54,0,212,0,188,0,75,0,217,0,87,0,194,0,38,0,31,0,0,0,219,0,40,0,22,0,152,0,17,0,65,0,229,0,32,0,79,0,95,0,112,0,161,0,102,0,208,0,185,0,167,0,0,0,207,0,39,0,71,0,196,0,0,0,0,0,0,0,144,0,0,0,96,0,11,0,225,0,0,0,203,0,104,0,97,0,40,0,160,0,22,0,195,0,0,0,154,0,72,0,250,0,249,0,190,0,0,0,178,0,231,0,30,0,49,0,185,0,0,0,0,0,193,0,39,0,10,0,14,0,183,0,36,0,186,0,224,0,161,0,0,0,57,0,246,0,206,0,0,0,0,0,30,0,57,0,0,0,78,0,104,0,113,0,79,0,87,0,120,0,125,0,0,0,91,0,239,0,194,0,0,0,125,0,142,0,218,0,166,0,48,0,186,0,71,0,25,0,0,0,102,0,204,0,95,0,215,0,64,0,17,0,103,0,250,0,204,0,209,0,253,0,19,0,73,0,218,0,0,0,163,0,0,0,0,0,195,0,165,0,72,0,80,0,72,0,73,0,161,0,172,0,126,0,160,0,191,0,176,0,222,0,102,0,32,0,90,0,148,0,138,0,0,0,255,0,135,0,120,0,163,0,33,0,214,0,209,0,160,0,76,0,240,0,0,0,32,0,35,0,200,0,40,0,146,0,108,0,0,0,60,0,0,0,195,0,10,0,58,0,238,0,56,0,84,0,149,0,250,0,11,0,190,0,120,0,208,0,182,0,121,0,0,0,236,0,201,0,12,0,186,0,0,0,204,0,170,0,80,0,164,0,253,0,25,0,172,0,58,0,94,0,235,0,142,0,255,0,216,0,0,0,152,0,32,0,19,0,20,0,244,0,0,0,158,0,219,0,76,0,163,0,0,0,0,0,0,0,208,0,214,0,0,0,0,0,98,0,167,0,109,0,3,0,89,0,112,0,0,0,0,0,100,0,236,0,22,0,172,0,106,0,0,0,155,0,182,0,148,0,86,0,172,0,39,0,57,0,154,0,114,0,131,0,0,0,10,0,0,0,0,0,137,0,235,0,176,0,154,0,0,0,97,0,119,0,131,0,39,0,182,0,0,0,217,0,134,0,188,0,0,0,23,0,0,0,235,0,145,0,97,0,1,0,135,0,0,0,207,0,113,0,10,0,175,0,148,0,47,0,41,0,49,0,0,0,255,0,0,0,221,0,36,0,208,0,198,0,98,0,31,0,0,0,181,0,40,0,4,0,85,0,149,0,134,0,204,0,192,0,34,0,185,0,202,0,147,0,171,0,141,0,0,0,5,0,46,0,143,0,7,0,243,0,250,0,101,0,1,0,97,0,0,0,179,0,0,0,141,0,254,0,164,0,226,0,58,0,222,0,0,0,0,0,20,0,0,0,0,0,186,0,0,0,250,0,75,0,91,0,0,0,208,0,0,0,121,0,113,0,152,0,0,0,169,0,0,0,0,0,143,0,181,0,0,0,229,0,0,0,0,0,169,0,0,0,0,0,132,0,0,0,112,0,145,0,186,0,124,0,34,0,93,0,83,0,218,0,46,0,143,0,174,0,0,0,196,0,111,0,214,0,205,0,85,0,6,0,0,0,0,0,195,0,26,0,105,0,0,0,0,0,37,0,79,0,65,0,206,0,187,0,165,0,101,0,159,0,129,0,114,0,211,0,17,0,53,0,144,0,0,0,158,0,90,0,0,0,240,0,138,0,66,0,26,0,124,0,36,0,144,0,164,0,102,0,23,0);
signal scenario_full  : scenario_type := (235,31,93,31,213,31,227,31,140,31,36,31,219,31,23,31,148,31,14,31,14,30,211,31,211,30,21,31,10,31,159,31,152,31,80,31,218,31,112,31,107,31,224,31,95,31,95,30,76,31,50,31,50,30,44,31,28,31,28,30,226,31,134,31,134,30,144,31,14,31,148,31,175,31,55,31,55,30,219,31,18,31,18,30,97,31,232,31,12,31,154,31,82,31,107,31,155,31,20,31,94,31,210,31,210,30,244,31,244,30,116,31,35,31,203,31,101,31,101,30,207,31,207,30,144,31,220,31,220,30,10,31,95,31,186,31,168,31,168,30,57,31,57,30,57,29,57,28,16,31,216,31,102,31,115,31,97,31,46,31,206,31,206,30,206,29,196,31,97,31,140,31,37,31,172,31,44,31,100,31,64,31,65,31,65,30,65,29,65,28,213,31,34,31,84,31,96,31,81,31,11,31,99,31,194,31,194,30,81,31,81,30,81,29,201,31,201,30,201,29,82,31,205,31,252,31,180,31,96,31,76,31,121,31,133,31,133,30,206,31,80,31,80,30,80,29,80,28,76,31,38,31,186,31,152,31,18,31,220,31,89,31,130,31,173,31,153,31,98,31,86,31,192,31,108,31,178,31,178,30,251,31,157,31,154,31,154,30,154,29,86,31,118,31,118,30,118,29,226,31,226,30,47,31,28,31,73,31,73,30,61,31,204,31,104,31,104,30,55,31,214,31,98,31,98,30,126,31,126,30,237,31,74,31,79,31,112,31,112,30,8,31,212,31,8,31,8,30,30,31,233,31,177,31,84,31,62,31,63,31,177,31,166,31,73,31,73,30,74,31,122,31,202,31,144,31,144,30,144,29,144,28,162,31,50,31,164,31,231,31,231,30,34,31,193,31,238,31,50,31,180,31,215,31,218,31,218,30,24,31,24,30,103,31,103,30,103,29,250,31,250,30,198,31,37,31,106,31,165,31,165,30,125,31,161,31,37,31,43,31,44,31,14,31,61,31,23,31,58,31,58,30,252,31,253,31,34,31,34,30,34,29,185,31,8,31,8,30,47,31,34,31,216,31,60,31,218,31,218,30,10,31,199,31,136,31,158,31,158,30,56,31,87,31,71,31,95,31,107,31,216,31,92,31,127,31,171,31,171,30,154,31,35,31,35,30,83,31,122,31,64,31,161,31,83,31,86,31,75,31,93,31,93,30,252,31,252,30,89,31,64,31,64,30,64,29,81,31,111,31,23,31,170,31,61,31,31,31,5,31,191,31,96,31,45,31,149,31,149,30,149,29,149,28,211,31,125,31,125,30,252,31,57,31,60,31,60,30,119,31,207,31,2,31,2,30,71,31,84,31,198,31,215,31,173,31,188,31,194,31,194,30,119,31,210,31,183,31,183,30,25,31,28,31,28,30,194,31,194,30,90,31,64,31,64,30,29,31,37,31,37,30,218,31,177,31,199,31,212,31,24,31,168,31,128,31,26,31,100,31,73,31,231,31,231,30,97,31,59,31,59,30,2,31,2,30,2,29,2,28,120,31,54,31,76,31,7,31,151,31,76,31,197,31,143,31,143,30,213,31,103,31,149,31,36,31,205,31,125,31,125,30,125,29,179,31,179,30,132,31,49,31,88,31,134,31,240,31,16,31,16,30,16,29,187,31,54,31,212,31,188,31,75,31,217,31,87,31,194,31,38,31,31,31,31,30,219,31,40,31,22,31,152,31,17,31,65,31,229,31,32,31,79,31,95,31,112,31,161,31,102,31,208,31,185,31,167,31,167,30,207,31,39,31,71,31,196,31,196,30,196,29,196,28,144,31,144,30,96,31,11,31,225,31,225,30,203,31,104,31,97,31,40,31,160,31,22,31,195,31,195,30,154,31,72,31,250,31,249,31,190,31,190,30,178,31,231,31,30,31,49,31,185,31,185,30,185,29,193,31,39,31,10,31,14,31,183,31,36,31,186,31,224,31,161,31,161,30,57,31,246,31,206,31,206,30,206,29,30,31,57,31,57,30,78,31,104,31,113,31,79,31,87,31,120,31,125,31,125,30,91,31,239,31,194,31,194,30,125,31,142,31,218,31,166,31,48,31,186,31,71,31,25,31,25,30,102,31,204,31,95,31,215,31,64,31,17,31,103,31,250,31,204,31,209,31,253,31,19,31,73,31,218,31,218,30,163,31,163,30,163,29,195,31,165,31,72,31,80,31,72,31,73,31,161,31,172,31,126,31,160,31,191,31,176,31,222,31,102,31,32,31,90,31,148,31,138,31,138,30,255,31,135,31,120,31,163,31,33,31,214,31,209,31,160,31,76,31,240,31,240,30,32,31,35,31,200,31,40,31,146,31,108,31,108,30,60,31,60,30,195,31,10,31,58,31,238,31,56,31,84,31,149,31,250,31,11,31,190,31,120,31,208,31,182,31,121,31,121,30,236,31,201,31,12,31,186,31,186,30,204,31,170,31,80,31,164,31,253,31,25,31,172,31,58,31,94,31,235,31,142,31,255,31,216,31,216,30,152,31,32,31,19,31,20,31,244,31,244,30,158,31,219,31,76,31,163,31,163,30,163,29,163,28,208,31,214,31,214,30,214,29,98,31,167,31,109,31,3,31,89,31,112,31,112,30,112,29,100,31,236,31,22,31,172,31,106,31,106,30,155,31,182,31,148,31,86,31,172,31,39,31,57,31,154,31,114,31,131,31,131,30,10,31,10,30,10,29,137,31,235,31,176,31,154,31,154,30,97,31,119,31,131,31,39,31,182,31,182,30,217,31,134,31,188,31,188,30,23,31,23,30,235,31,145,31,97,31,1,31,135,31,135,30,207,31,113,31,10,31,175,31,148,31,47,31,41,31,49,31,49,30,255,31,255,30,221,31,36,31,208,31,198,31,98,31,31,31,31,30,181,31,40,31,4,31,85,31,149,31,134,31,204,31,192,31,34,31,185,31,202,31,147,31,171,31,141,31,141,30,5,31,46,31,143,31,7,31,243,31,250,31,101,31,1,31,97,31,97,30,179,31,179,30,141,31,254,31,164,31,226,31,58,31,222,31,222,30,222,29,20,31,20,30,20,29,186,31,186,30,250,31,75,31,91,31,91,30,208,31,208,30,121,31,113,31,152,31,152,30,169,31,169,30,169,29,143,31,181,31,181,30,229,31,229,30,229,29,169,31,169,30,169,29,132,31,132,30,112,31,145,31,186,31,124,31,34,31,93,31,83,31,218,31,46,31,143,31,174,31,174,30,196,31,111,31,214,31,205,31,85,31,6,31,6,30,6,29,195,31,26,31,105,31,105,30,105,29,37,31,79,31,65,31,206,31,187,31,165,31,101,31,159,31,129,31,114,31,211,31,17,31,53,31,144,31,144,30,158,31,90,31,90,30,240,31,138,31,66,31,26,31,124,31,36,31,144,31,164,31,102,31,23,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
