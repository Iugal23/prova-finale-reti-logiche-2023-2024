-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 916;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,31,0,86,0,206,0,0,0,203,0,124,0,122,0,233,0,26,0,229,0,214,0,253,0,227,0,0,0,140,0,152,0,166,0,60,0,218,0,103,0,248,0,0,0,0,0,4,0,153,0,78,0,141,0,216,0,149,0,102,0,98,0,0,0,0,0,179,0,240,0,195,0,0,0,0,0,79,0,113,0,224,0,60,0,254,0,214,0,128,0,83,0,0,0,161,0,118,0,68,0,0,0,57,0,0,0,184,0,108,0,13,0,220,0,95,0,51,0,79,0,181,0,74,0,103,0,149,0,0,0,20,0,24,0,53,0,0,0,186,0,93,0,29,0,0,0,219,0,191,0,253,0,132,0,0,0,73,0,0,0,165,0,0,0,0,0,48,0,116,0,157,0,0,0,108,0,0,0,188,0,31,0,0,0,21,0,68,0,173,0,0,0,115,0,171,0,0,0,90,0,100,0,188,0,0,0,94,0,44,0,57,0,208,0,139,0,0,0,105,0,221,0,13,0,44,0,233,0,219,0,0,0,25,0,210,0,222,0,70,0,59,0,136,0,0,0,0,0,91,0,206,0,0,0,117,0,28,0,214,0,252,0,200,0,232,0,51,0,245,0,166,0,0,0,255,0,192,0,0,0,182,0,147,0,114,0,173,0,223,0,95,0,179,0,44,0,0,0,216,0,234,0,252,0,0,0,86,0,112,0,193,0,0,0,201,0,26,0,0,0,77,0,0,0,79,0,67,0,3,0,0,0,34,0,162,0,95,0,234,0,41,0,110,0,41,0,0,0,0,0,194,0,212,0,162,0,111,0,221,0,55,0,214,0,0,0,239,0,108,0,109,0,216,0,178,0,12,0,63,0,103,0,74,0,0,0,0,0,173,0,109,0,109,0,0,0,0,0,11,0,0,0,222,0,95,0,55,0,190,0,97,0,0,0,10,0,93,0,201,0,65,0,0,0,239,0,103,0,31,0,46,0,150,0,34,0,0,0,14,0,95,0,209,0,102,0,253,0,0,0,47,0,24,0,161,0,139,0,0,0,0,0,215,0,39,0,207,0,82,0,25,0,199,0,0,0,175,0,251,0,93,0,0,0,244,0,185,0,80,0,37,0,184,0,31,0,116,0,120,0,11,0,0,0,105,0,8,0,249,0,28,0,60,0,0,0,5,0,39,0,221,0,224,0,218,0,0,0,193,0,240,0,61,0,124,0,47,0,2,0,152,0,14,0,135,0,4,0,65,0,139,0,24,0,217,0,225,0,186,0,140,0,29,0,171,0,0,0,200,0,102,0,157,0,204,0,107,0,0,0,67,0,0,0,1,0,159,0,0,0,79,0,8,0,191,0,98,0,117,0,0,0,77,0,1,0,168,0,89,0,0,0,176,0,169,0,0,0,0,0,133,0,0,0,10,0,244,0,108,0,0,0,115,0,113,0,101,0,101,0,53,0,34,0,0,0,16,0,0,0,202,0,143,0,177,0,233,0,0,0,215,0,198,0,149,0,95,0,69,0,0,0,102,0,153,0,0,0,0,0,137,0,8,0,67,0,176,0,42,0,0,0,0,0,246,0,68,0,238,0,34,0,212,0,228,0,108,0,202,0,198,0,0,0,166,0,19,0,181,0,62,0,161,0,166,0,174,0,148,0,241,0,20,0,219,0,48,0,0,0,222,0,0,0,10,0,0,0,72,0,114,0,185,0,241,0,242,0,0,0,0,0,187,0,210,0,0,0,150,0,0,0,205,0,0,0,62,0,105,0,0,0,198,0,167,0,127,0,247,0,123,0,0,0,112,0,135,0,0,0,151,0,194,0,25,0,0,0,0,0,238,0,251,0,48,0,0,0,0,0,255,0,78,0,123,0,135,0,0,0,31,0,66,0,0,0,0,0,219,0,98,0,236,0,0,0,79,0,185,0,13,0,143,0,0,0,173,0,74,0,46,0,234,0,147,0,3,0,144,0,94,0,55,0,235,0,116,0,157,0,151,0,47,0,95,0,171,0,145,0,173,0,206,0,0,0,0,0,25,0,0,0,0,0,113,0,203,0,117,0,155,0,89,0,0,0,60,0,238,0,84,0,227,0,227,0,0,0,7,0,187,0,44,0,130,0,94,0,0,0,98,0,61,0,130,0,197,0,0,0,179,0,242,0,178,0,120,0,80,0,45,0,170,0,134,0,164,0,0,0,161,0,179,0,40,0,0,0,28,0,210,0,18,0,0,0,0,0,40,0,20,0,140,0,0,0,0,0,154,0,0,0,134,0,0,0,211,0,169,0,0,0,7,0,67,0,58,0,111,0,0,0,39,0,0,0,253,0,112,0,0,0,210,0,193,0,20,0,237,0,185,0,18,0,0,0,237,0,184,0,48,0,167,0,221,0,59,0,134,0,194,0,133,0,228,0,0,0,39,0,114,0,52,0,214,0,0,0,0,0,244,0,122,0,74,0,86,0,228,0,246,0,17,0,250,0,9,0,0,0,224,0,0,0,233,0,100,0,57,0,160,0,94,0,237,0,66,0,0,0,247,0,70,0,0,0,0,0,158,0,128,0,45,0,166,0,215,0,92,0,19,0,0,0,41,0,21,0,93,0,229,0,206,0,242,0,58,0,135,0,0,0,59,0,221,0,44,0,43,0,0,0,116,0,0,0,60,0,244,0,144,0,0,0,90,0,150,0,199,0,210,0,215,0,202,0,107,0,104,0,51,0,35,0,108,0,0,0,162,0,173,0,210,0,168,0,0,0,210,0,0,0,191,0,76,0,194,0,33,0,113,0,36,0,102,0,89,0,196,0,0,0,213,0,3,0,236,0,0,0,138,0,0,0,136,0,19,0,67,0,185,0,148,0,226,0,0,0,6,0,234,0,74,0,131,0,244,0,92,0,0,0,179,0,92,0,117,0,216,0,238,0,181,0,48,0,52,0,0,0,153,0,202,0,10,0,122,0,235,0,0,0,0,0,241,0,0,0,0,0,78,0,44,0,84,0,182,0,198,0,47,0,230,0,202,0,0,0,191,0,0,0,169,0,100,0,173,0,207,0,0,0,17,0,188,0,250,0,250,0,16,0,191,0,253,0,19,0,74,0,136,0,111,0,110,0,24,0,97,0,157,0,225,0,124,0,176,0,196,0,93,0,74,0,68,0,0,0,0,0,0,0,127,0,0,0,120,0,71,0,0,0,252,0,47,0,207,0,134,0,174,0,0,0,6,0,82,0,62,0,83,0,0,0,59,0,61,0,89,0,0,0,0,0,210,0,106,0,206,0,59,0,225,0,0,0,87,0,59,0,239,0,94,0,112,0,162,0,127,0,250,0,132,0,0,0,98,0,177,0,53,0,37,0,76,0,205,0,12,0,114,0,177,0,0,0,0,0,7,0,31,0,0,0,254,0,0,0,144,0,48,0,0,0,208,0,165,0,0,0,64,0,144,0,0,0,148,0,255,0,110,0,0,0,183,0,225,0,97,0,56,0,9,0,63,0,81,0,0,0,240,0,158,0,24,0,35,0,244,0,208,0,54,0,222,0,66,0,0,0,252,0,88,0,239,0,0,0,58,0,109,0,0,0,0,0,2,0,112,0,192,0,0,0,156,0,156,0,226,0,170,0,105,0,229,0,237,0,25,0,0,0,48,0,147,0,0,0,0,0,28,0,0,0,145,0,204,0,213,0,0,0,156,0,0,0,0,0,231,0,128,0,0,0,136,0,43,0,0,0,248,0,0,0,153,0,244,0,0,0,0,0,0,0,143,0,0,0,0,0,0,0,194,0,176,0,33,0,0,0,105,0,0,0,193,0,45,0,196,0,221,0,166,0,252,0,91,0,215,0,164,0,56,0,107,0,188,0,143,0,205,0,81,0,81,0,4,0,246,0,0,0,208,0,159,0,201,0,28,0,90,0,252,0,169,0,111,0,0,0,0,0,219,0,91,0,176,0,147,0,236,0,0,0,139,0,23,0,23,0,0,0,0,0,244,0,74,0,0,0,240,0,209,0,0,0,134,0,219,0,4,0,50,0,14,0,0,0,95,0,109,0,41,0,237,0,223,0,218,0,212,0,203,0,46,0,90,0,139,0,60,0,0,0,27,0,206,0,0,0,0,0,152,0,0,0,195,0,149,0);
signal scenario_full  : scenario_type := (168,31,31,31,86,31,206,31,206,30,203,31,124,31,122,31,233,31,26,31,229,31,214,31,253,31,227,31,227,30,140,31,152,31,166,31,60,31,218,31,103,31,248,31,248,30,248,29,4,31,153,31,78,31,141,31,216,31,149,31,102,31,98,31,98,30,98,29,179,31,240,31,195,31,195,30,195,29,79,31,113,31,224,31,60,31,254,31,214,31,128,31,83,31,83,30,161,31,118,31,68,31,68,30,57,31,57,30,184,31,108,31,13,31,220,31,95,31,51,31,79,31,181,31,74,31,103,31,149,31,149,30,20,31,24,31,53,31,53,30,186,31,93,31,29,31,29,30,219,31,191,31,253,31,132,31,132,30,73,31,73,30,165,31,165,30,165,29,48,31,116,31,157,31,157,30,108,31,108,30,188,31,31,31,31,30,21,31,68,31,173,31,173,30,115,31,171,31,171,30,90,31,100,31,188,31,188,30,94,31,44,31,57,31,208,31,139,31,139,30,105,31,221,31,13,31,44,31,233,31,219,31,219,30,25,31,210,31,222,31,70,31,59,31,136,31,136,30,136,29,91,31,206,31,206,30,117,31,28,31,214,31,252,31,200,31,232,31,51,31,245,31,166,31,166,30,255,31,192,31,192,30,182,31,147,31,114,31,173,31,223,31,95,31,179,31,44,31,44,30,216,31,234,31,252,31,252,30,86,31,112,31,193,31,193,30,201,31,26,31,26,30,77,31,77,30,79,31,67,31,3,31,3,30,34,31,162,31,95,31,234,31,41,31,110,31,41,31,41,30,41,29,194,31,212,31,162,31,111,31,221,31,55,31,214,31,214,30,239,31,108,31,109,31,216,31,178,31,12,31,63,31,103,31,74,31,74,30,74,29,173,31,109,31,109,31,109,30,109,29,11,31,11,30,222,31,95,31,55,31,190,31,97,31,97,30,10,31,93,31,201,31,65,31,65,30,239,31,103,31,31,31,46,31,150,31,34,31,34,30,14,31,95,31,209,31,102,31,253,31,253,30,47,31,24,31,161,31,139,31,139,30,139,29,215,31,39,31,207,31,82,31,25,31,199,31,199,30,175,31,251,31,93,31,93,30,244,31,185,31,80,31,37,31,184,31,31,31,116,31,120,31,11,31,11,30,105,31,8,31,249,31,28,31,60,31,60,30,5,31,39,31,221,31,224,31,218,31,218,30,193,31,240,31,61,31,124,31,47,31,2,31,152,31,14,31,135,31,4,31,65,31,139,31,24,31,217,31,225,31,186,31,140,31,29,31,171,31,171,30,200,31,102,31,157,31,204,31,107,31,107,30,67,31,67,30,1,31,159,31,159,30,79,31,8,31,191,31,98,31,117,31,117,30,77,31,1,31,168,31,89,31,89,30,176,31,169,31,169,30,169,29,133,31,133,30,10,31,244,31,108,31,108,30,115,31,113,31,101,31,101,31,53,31,34,31,34,30,16,31,16,30,202,31,143,31,177,31,233,31,233,30,215,31,198,31,149,31,95,31,69,31,69,30,102,31,153,31,153,30,153,29,137,31,8,31,67,31,176,31,42,31,42,30,42,29,246,31,68,31,238,31,34,31,212,31,228,31,108,31,202,31,198,31,198,30,166,31,19,31,181,31,62,31,161,31,166,31,174,31,148,31,241,31,20,31,219,31,48,31,48,30,222,31,222,30,10,31,10,30,72,31,114,31,185,31,241,31,242,31,242,30,242,29,187,31,210,31,210,30,150,31,150,30,205,31,205,30,62,31,105,31,105,30,198,31,167,31,127,31,247,31,123,31,123,30,112,31,135,31,135,30,151,31,194,31,25,31,25,30,25,29,238,31,251,31,48,31,48,30,48,29,255,31,78,31,123,31,135,31,135,30,31,31,66,31,66,30,66,29,219,31,98,31,236,31,236,30,79,31,185,31,13,31,143,31,143,30,173,31,74,31,46,31,234,31,147,31,3,31,144,31,94,31,55,31,235,31,116,31,157,31,151,31,47,31,95,31,171,31,145,31,173,31,206,31,206,30,206,29,25,31,25,30,25,29,113,31,203,31,117,31,155,31,89,31,89,30,60,31,238,31,84,31,227,31,227,31,227,30,7,31,187,31,44,31,130,31,94,31,94,30,98,31,61,31,130,31,197,31,197,30,179,31,242,31,178,31,120,31,80,31,45,31,170,31,134,31,164,31,164,30,161,31,179,31,40,31,40,30,28,31,210,31,18,31,18,30,18,29,40,31,20,31,140,31,140,30,140,29,154,31,154,30,134,31,134,30,211,31,169,31,169,30,7,31,67,31,58,31,111,31,111,30,39,31,39,30,253,31,112,31,112,30,210,31,193,31,20,31,237,31,185,31,18,31,18,30,237,31,184,31,48,31,167,31,221,31,59,31,134,31,194,31,133,31,228,31,228,30,39,31,114,31,52,31,214,31,214,30,214,29,244,31,122,31,74,31,86,31,228,31,246,31,17,31,250,31,9,31,9,30,224,31,224,30,233,31,100,31,57,31,160,31,94,31,237,31,66,31,66,30,247,31,70,31,70,30,70,29,158,31,128,31,45,31,166,31,215,31,92,31,19,31,19,30,41,31,21,31,93,31,229,31,206,31,242,31,58,31,135,31,135,30,59,31,221,31,44,31,43,31,43,30,116,31,116,30,60,31,244,31,144,31,144,30,90,31,150,31,199,31,210,31,215,31,202,31,107,31,104,31,51,31,35,31,108,31,108,30,162,31,173,31,210,31,168,31,168,30,210,31,210,30,191,31,76,31,194,31,33,31,113,31,36,31,102,31,89,31,196,31,196,30,213,31,3,31,236,31,236,30,138,31,138,30,136,31,19,31,67,31,185,31,148,31,226,31,226,30,6,31,234,31,74,31,131,31,244,31,92,31,92,30,179,31,92,31,117,31,216,31,238,31,181,31,48,31,52,31,52,30,153,31,202,31,10,31,122,31,235,31,235,30,235,29,241,31,241,30,241,29,78,31,44,31,84,31,182,31,198,31,47,31,230,31,202,31,202,30,191,31,191,30,169,31,100,31,173,31,207,31,207,30,17,31,188,31,250,31,250,31,16,31,191,31,253,31,19,31,74,31,136,31,111,31,110,31,24,31,97,31,157,31,225,31,124,31,176,31,196,31,93,31,74,31,68,31,68,30,68,29,68,28,127,31,127,30,120,31,71,31,71,30,252,31,47,31,207,31,134,31,174,31,174,30,6,31,82,31,62,31,83,31,83,30,59,31,61,31,89,31,89,30,89,29,210,31,106,31,206,31,59,31,225,31,225,30,87,31,59,31,239,31,94,31,112,31,162,31,127,31,250,31,132,31,132,30,98,31,177,31,53,31,37,31,76,31,205,31,12,31,114,31,177,31,177,30,177,29,7,31,31,31,31,30,254,31,254,30,144,31,48,31,48,30,208,31,165,31,165,30,64,31,144,31,144,30,148,31,255,31,110,31,110,30,183,31,225,31,97,31,56,31,9,31,63,31,81,31,81,30,240,31,158,31,24,31,35,31,244,31,208,31,54,31,222,31,66,31,66,30,252,31,88,31,239,31,239,30,58,31,109,31,109,30,109,29,2,31,112,31,192,31,192,30,156,31,156,31,226,31,170,31,105,31,229,31,237,31,25,31,25,30,48,31,147,31,147,30,147,29,28,31,28,30,145,31,204,31,213,31,213,30,156,31,156,30,156,29,231,31,128,31,128,30,136,31,43,31,43,30,248,31,248,30,153,31,244,31,244,30,244,29,244,28,143,31,143,30,143,29,143,28,194,31,176,31,33,31,33,30,105,31,105,30,193,31,45,31,196,31,221,31,166,31,252,31,91,31,215,31,164,31,56,31,107,31,188,31,143,31,205,31,81,31,81,31,4,31,246,31,246,30,208,31,159,31,201,31,28,31,90,31,252,31,169,31,111,31,111,30,111,29,219,31,91,31,176,31,147,31,236,31,236,30,139,31,23,31,23,31,23,30,23,29,244,31,74,31,74,30,240,31,209,31,209,30,134,31,219,31,4,31,50,31,14,31,14,30,95,31,109,31,41,31,237,31,223,31,218,31,212,31,203,31,46,31,90,31,139,31,60,31,60,30,27,31,206,31,206,30,206,29,152,31,152,30,195,31,149,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
