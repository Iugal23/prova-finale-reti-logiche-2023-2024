-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 660;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (14,0,78,0,7,0,237,0,79,0,8,0,173,0,109,0,66,0,106,0,147,0,246,0,203,0,0,0,110,0,206,0,34,0,176,0,49,0,108,0,164,0,0,0,16,0,247,0,193,0,12,0,65,0,50,0,129,0,225,0,0,0,170,0,241,0,194,0,85,0,137,0,16,0,79,0,19,0,1,0,151,0,118,0,165,0,246,0,240,0,146,0,8,0,81,0,0,0,8,0,226,0,0,0,149,0,228,0,210,0,0,0,13,0,201,0,91,0,49,0,43,0,222,0,2,0,240,0,196,0,197,0,130,0,32,0,50,0,209,0,8,0,131,0,0,0,184,0,0,0,243,0,140,0,0,0,0,0,154,0,0,0,248,0,51,0,253,0,0,0,37,0,115,0,255,0,46,0,248,0,40,0,204,0,0,0,73,0,23,0,0,0,133,0,252,0,161,0,0,0,10,0,39,0,196,0,96,0,233,0,0,0,125,0,0,0,78,0,45,0,18,0,0,0,127,0,169,0,189,0,200,0,0,0,44,0,18,0,223,0,179,0,223,0,0,0,80,0,187,0,4,0,0,0,48,0,48,0,111,0,0,0,100,0,0,0,35,0,57,0,0,0,50,0,247,0,58,0,184,0,34,0,11,0,118,0,148,0,128,0,122,0,168,0,0,0,9,0,174,0,27,0,151,0,0,0,196,0,190,0,199,0,0,0,222,0,152,0,91,0,239,0,125,0,171,0,30,0,0,0,26,0,70,0,58,0,229,0,0,0,26,0,16,0,0,0,0,0,121,0,181,0,252,0,62,0,216,0,154,0,123,0,249,0,198,0,247,0,162,0,237,0,38,0,133,0,235,0,113,0,38,0,0,0,36,0,216,0,0,0,241,0,0,0,0,0,25,0,0,0,92,0,149,0,197,0,124,0,16,0,189,0,0,0,15,0,213,0,158,0,118,0,169,0,0,0,12,0,182,0,243,0,26,0,254,0,47,0,0,0,45,0,0,0,134,0,0,0,197,0,147,0,82,0,252,0,0,0,72,0,177,0,115,0,0,0,240,0,137,0,4,0,184,0,217,0,97,0,249,0,0,0,0,0,223,0,184,0,231,0,138,0,122,0,229,0,38,0,172,0,178,0,0,0,11,0,219,0,193,0,234,0,239,0,233,0,175,0,32,0,0,0,151,0,19,0,93,0,131,0,59,0,61,0,0,0,129,0,33,0,109,0,135,0,164,0,109,0,0,0,0,0,73,0,175,0,194,0,68,0,88,0,204,0,249,0,52,0,0,0,184,0,27,0,229,0,24,0,147,0,155,0,0,0,141,0,252,0,0,0,0,0,0,0,198,0,233,0,0,0,0,0,0,0,196,0,203,0,175,0,110,0,209,0,0,0,164,0,214,0,0,0,144,0,0,0,99,0,81,0,0,0,227,0,129,0,0,0,234,0,253,0,92,0,0,0,120,0,0,0,0,0,29,0,0,0,0,0,160,0,190,0,153,0,0,0,0,0,0,0,220,0,0,0,9,0,136,0,146,0,229,0,171,0,0,0,0,0,141,0,6,0,0,0,0,0,0,0,0,0,164,0,0,0,68,0,248,0,0,0,134,0,119,0,65,0,203,0,236,0,0,0,237,0,66,0,0,0,31,0,175,0,175,0,231,0,233,0,18,0,65,0,0,0,219,0,126,0,0,0,0,0,0,0,169,0,171,0,0,0,249,0,0,0,3,0,0,0,187,0,246,0,56,0,0,0,203,0,30,0,197,0,197,0,135,0,245,0,99,0,0,0,231,0,236,0,254,0,52,0,0,0,0,0,38,0,215,0,93,0,22,0,161,0,0,0,0,0,0,0,180,0,88,0,121,0,0,0,130,0,10,0,199,0,0,0,203,0,160,0,194,0,65,0,151,0,135,0,214,0,131,0,49,0,99,0,0,0,63,0,22,0,0,0,0,0,176,0,213,0,23,0,3,0,32,0,212,0,0,0,221,0,174,0,213,0,156,0,214,0,42,0,245,0,203,0,0,0,0,0,135,0,83,0,75,0,42,0,0,0,22,0,40,0,0,0,198,0,213,0,0,0,184,0,0,0,30,0,76,0,203,0,43,0,0,0,165,0,0,0,116,0,190,0,205,0,0,0,0,0,106,0,210,0,139,0,163,0,0,0,0,0,162,0,33,0,25,0,0,0,98,0,81,0,66,0,0,0,212,0,58,0,0,0,9,0,223,0,51,0,48,0,78,0,221,0,252,0,36,0,223,0,188,0,0,0,149,0,0,0,155,0,106,0,0,0,114,0,238,0,183,0,21,0,109,0,0,0,194,0,0,0,0,0,231,0,209,0,235,0,52,0,114,0,58,0,66,0,175,0,82,0,193,0,0,0,70,0,11,0,182,0,33,0,240,0,4,0,0,0,8,0,230,0,69,0,99,0,182,0,134,0,90,0,26,0,9,0,191,0,59,0,140,0,0,0,137,0,29,0,123,0,147,0,0,0,107,0,38,0,0,0,0,0,8,0,241,0,80,0,0,0,137,0,171,0,243,0,0,0,0,0,0,0,92,0,40,0,149,0,103,0,54,0,0,0,242,0,0,0,225,0,201,0,151,0,106,0,181,0,19,0,0,0,126,0,71,0,28,0,124,0,207,0,31,0,202,0,110,0,109,0,0,0,0,0,214,0,44,0,192,0,111,0,25,0,138,0,97,0,228,0,99,0,103,0,0,0,112,0,0,0,128,0,236,0,117,0,143,0,0,0,111,0,100,0,238,0,143,0,15,0,0,0,189,0,162,0,0,0,228,0,101,0,0,0,0,0,215,0,157,0,216,0,218,0,150,0,236,0,2,0,0,0,244,0,194,0,24,0,221,0,251,0,0,0,17,0,50,0,0,0,208,0,38,0,43,0,126,0,134,0,0,0,185,0,148,0,0,0,0,0,116,0,180,0,130,0,251,0,33,0,49,0,109,0,0,0,104,0);
signal scenario_full  : scenario_type := (14,31,78,31,7,31,237,31,79,31,8,31,173,31,109,31,66,31,106,31,147,31,246,31,203,31,203,30,110,31,206,31,34,31,176,31,49,31,108,31,164,31,164,30,16,31,247,31,193,31,12,31,65,31,50,31,129,31,225,31,225,30,170,31,241,31,194,31,85,31,137,31,16,31,79,31,19,31,1,31,151,31,118,31,165,31,246,31,240,31,146,31,8,31,81,31,81,30,8,31,226,31,226,30,149,31,228,31,210,31,210,30,13,31,201,31,91,31,49,31,43,31,222,31,2,31,240,31,196,31,197,31,130,31,32,31,50,31,209,31,8,31,131,31,131,30,184,31,184,30,243,31,140,31,140,30,140,29,154,31,154,30,248,31,51,31,253,31,253,30,37,31,115,31,255,31,46,31,248,31,40,31,204,31,204,30,73,31,23,31,23,30,133,31,252,31,161,31,161,30,10,31,39,31,196,31,96,31,233,31,233,30,125,31,125,30,78,31,45,31,18,31,18,30,127,31,169,31,189,31,200,31,200,30,44,31,18,31,223,31,179,31,223,31,223,30,80,31,187,31,4,31,4,30,48,31,48,31,111,31,111,30,100,31,100,30,35,31,57,31,57,30,50,31,247,31,58,31,184,31,34,31,11,31,118,31,148,31,128,31,122,31,168,31,168,30,9,31,174,31,27,31,151,31,151,30,196,31,190,31,199,31,199,30,222,31,152,31,91,31,239,31,125,31,171,31,30,31,30,30,26,31,70,31,58,31,229,31,229,30,26,31,16,31,16,30,16,29,121,31,181,31,252,31,62,31,216,31,154,31,123,31,249,31,198,31,247,31,162,31,237,31,38,31,133,31,235,31,113,31,38,31,38,30,36,31,216,31,216,30,241,31,241,30,241,29,25,31,25,30,92,31,149,31,197,31,124,31,16,31,189,31,189,30,15,31,213,31,158,31,118,31,169,31,169,30,12,31,182,31,243,31,26,31,254,31,47,31,47,30,45,31,45,30,134,31,134,30,197,31,147,31,82,31,252,31,252,30,72,31,177,31,115,31,115,30,240,31,137,31,4,31,184,31,217,31,97,31,249,31,249,30,249,29,223,31,184,31,231,31,138,31,122,31,229,31,38,31,172,31,178,31,178,30,11,31,219,31,193,31,234,31,239,31,233,31,175,31,32,31,32,30,151,31,19,31,93,31,131,31,59,31,61,31,61,30,129,31,33,31,109,31,135,31,164,31,109,31,109,30,109,29,73,31,175,31,194,31,68,31,88,31,204,31,249,31,52,31,52,30,184,31,27,31,229,31,24,31,147,31,155,31,155,30,141,31,252,31,252,30,252,29,252,28,198,31,233,31,233,30,233,29,233,28,196,31,203,31,175,31,110,31,209,31,209,30,164,31,214,31,214,30,144,31,144,30,99,31,81,31,81,30,227,31,129,31,129,30,234,31,253,31,92,31,92,30,120,31,120,30,120,29,29,31,29,30,29,29,160,31,190,31,153,31,153,30,153,29,153,28,220,31,220,30,9,31,136,31,146,31,229,31,171,31,171,30,171,29,141,31,6,31,6,30,6,29,6,28,6,27,164,31,164,30,68,31,248,31,248,30,134,31,119,31,65,31,203,31,236,31,236,30,237,31,66,31,66,30,31,31,175,31,175,31,231,31,233,31,18,31,65,31,65,30,219,31,126,31,126,30,126,29,126,28,169,31,171,31,171,30,249,31,249,30,3,31,3,30,187,31,246,31,56,31,56,30,203,31,30,31,197,31,197,31,135,31,245,31,99,31,99,30,231,31,236,31,254,31,52,31,52,30,52,29,38,31,215,31,93,31,22,31,161,31,161,30,161,29,161,28,180,31,88,31,121,31,121,30,130,31,10,31,199,31,199,30,203,31,160,31,194,31,65,31,151,31,135,31,214,31,131,31,49,31,99,31,99,30,63,31,22,31,22,30,22,29,176,31,213,31,23,31,3,31,32,31,212,31,212,30,221,31,174,31,213,31,156,31,214,31,42,31,245,31,203,31,203,30,203,29,135,31,83,31,75,31,42,31,42,30,22,31,40,31,40,30,198,31,213,31,213,30,184,31,184,30,30,31,76,31,203,31,43,31,43,30,165,31,165,30,116,31,190,31,205,31,205,30,205,29,106,31,210,31,139,31,163,31,163,30,163,29,162,31,33,31,25,31,25,30,98,31,81,31,66,31,66,30,212,31,58,31,58,30,9,31,223,31,51,31,48,31,78,31,221,31,252,31,36,31,223,31,188,31,188,30,149,31,149,30,155,31,106,31,106,30,114,31,238,31,183,31,21,31,109,31,109,30,194,31,194,30,194,29,231,31,209,31,235,31,52,31,114,31,58,31,66,31,175,31,82,31,193,31,193,30,70,31,11,31,182,31,33,31,240,31,4,31,4,30,8,31,230,31,69,31,99,31,182,31,134,31,90,31,26,31,9,31,191,31,59,31,140,31,140,30,137,31,29,31,123,31,147,31,147,30,107,31,38,31,38,30,38,29,8,31,241,31,80,31,80,30,137,31,171,31,243,31,243,30,243,29,243,28,92,31,40,31,149,31,103,31,54,31,54,30,242,31,242,30,225,31,201,31,151,31,106,31,181,31,19,31,19,30,126,31,71,31,28,31,124,31,207,31,31,31,202,31,110,31,109,31,109,30,109,29,214,31,44,31,192,31,111,31,25,31,138,31,97,31,228,31,99,31,103,31,103,30,112,31,112,30,128,31,236,31,117,31,143,31,143,30,111,31,100,31,238,31,143,31,15,31,15,30,189,31,162,31,162,30,228,31,101,31,101,30,101,29,215,31,157,31,216,31,218,31,150,31,236,31,2,31,2,30,244,31,194,31,24,31,221,31,251,31,251,30,17,31,50,31,50,30,208,31,38,31,43,31,126,31,134,31,134,30,185,31,148,31,148,30,148,29,116,31,180,31,130,31,251,31,33,31,49,31,109,31,109,30,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
