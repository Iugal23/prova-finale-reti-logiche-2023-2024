-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 960;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (200,0,213,0,138,0,64,0,4,0,0,0,175,0,0,0,120,0,0,0,249,0,209,0,243,0,117,0,125,0,0,0,0,0,251,0,98,0,253,0,162,0,207,0,0,0,0,0,0,0,38,0,202,0,253,0,50,0,0,0,141,0,121,0,66,0,2,0,11,0,99,0,0,0,77,0,0,0,23,0,252,0,157,0,73,0,105,0,0,0,121,0,170,0,44,0,150,0,55,0,37,0,188,0,0,0,56,0,0,0,160,0,180,0,229,0,26,0,247,0,92,0,0,0,104,0,38,0,75,0,97,0,93,0,129,0,244,0,0,0,182,0,0,0,93,0,0,0,138,0,0,0,0,0,224,0,0,0,119,0,0,0,198,0,205,0,0,0,231,0,70,0,32,0,0,0,252,0,64,0,125,0,230,0,101,0,154,0,1,0,100,0,48,0,80,0,37,0,32,0,0,0,196,0,15,0,216,0,0,0,238,0,123,0,20,0,185,0,204,0,179,0,242,0,0,0,0,0,160,0,128,0,222,0,219,0,204,0,254,0,29,0,95,0,18,0,0,0,92,0,87,0,50,0,252,0,140,0,249,0,172,0,129,0,231,0,87,0,59,0,113,0,21,0,84,0,119,0,0,0,123,0,195,0,241,0,0,0,0,0,44,0,227,0,219,0,18,0,136,0,160,0,217,0,0,0,130,0,137,0,0,0,18,0,190,0,42,0,90,0,227,0,168,0,80,0,103,0,9,0,138,0,85,0,0,0,41,0,91,0,199,0,180,0,227,0,0,0,7,0,67,0,179,0,8,0,0,0,98,0,243,0,95,0,2,0,187,0,215,0,83,0,81,0,236,0,114,0,191,0,156,0,14,0,0,0,248,0,121,0,234,0,157,0,201,0,177,0,128,0,219,0,0,0,217,0,0,0,36,0,217,0,156,0,0,0,70,0,104,0,143,0,77,0,153,0,0,0,15,0,222,0,202,0,92,0,229,0,136,0,69,0,103,0,41,0,148,0,73,0,56,0,234,0,152,0,93,0,141,0,167,0,0,0,23,0,0,0,193,0,219,0,252,0,0,0,169,0,49,0,6,0,0,0,127,0,228,0,62,0,30,0,221,0,75,0,171,0,139,0,62,0,6,0,0,0,0,0,227,0,111,0,0,0,158,0,160,0,0,0,0,0,59,0,0,0,222,0,241,0,0,0,246,0,119,0,88,0,0,0,251,0,179,0,69,0,15,0,0,0,151,0,43,0,54,0,8,0,91,0,242,0,183,0,0,0,168,0,122,0,179,0,83,0,109,0,117,0,0,0,197,0,19,0,70,0,24,0,25,0,50,0,124,0,65,0,202,0,119,0,203,0,88,0,168,0,81,0,0,0,0,0,222,0,17,0,62,0,100,0,140,0,0,0,0,0,5,0,147,0,0,0,167,0,221,0,219,0,202,0,238,0,199,0,232,0,175,0,176,0,28,0,83,0,215,0,168,0,207,0,0,0,197,0,190,0,178,0,0,0,183,0,115,0,162,0,217,0,0,0,53,0,3,0,0,0,192,0,168,0,158,0,105,0,124,0,185,0,222,0,171,0,113,0,110,0,20,0,0,0,2,0,0,0,156,0,0,0,0,0,192,0,193,0,39,0,0,0,109,0,24,0,14,0,0,0,221,0,0,0,51,0,26,0,217,0,53,0,209,0,0,0,205,0,234,0,198,0,20,0,0,0,0,0,134,0,3,0,158,0,211,0,0,0,44,0,217,0,0,0,28,0,228,0,231,0,74,0,213,0,40,0,0,0,13,0,147,0,96,0,0,0,124,0,0,0,0,0,71,0,0,0,135,0,249,0,20,0,140,0,86,0,21,0,130,0,227,0,190,0,49,0,60,0,0,0,40,0,0,0,165,0,166,0,207,0,42,0,0,0,0,0,189,0,65,0,227,0,72,0,168,0,129,0,0,0,251,0,1,0,157,0,252,0,63,0,207,0,243,0,21,0,239,0,0,0,59,0,196,0,182,0,57,0,0,0,80,0,0,0,33,0,167,0,157,0,14,0,123,0,250,0,0,0,0,0,57,0,52,0,25,0,16,0,161,0,50,0,143,0,224,0,122,0,143,0,88,0,53,0,0,0,190,0,109,0,154,0,160,0,99,0,172,0,200,0,203,0,50,0,193,0,179,0,251,0,201,0,19,0,33,0,75,0,0,0,0,0,86,0,124,0,224,0,142,0,217,0,187,0,171,0,253,0,197,0,216,0,240,0,217,0,118,0,30,0,134,0,49,0,0,0,35,0,100,0,96,0,109,0,111,0,200,0,122,0,60,0,68,0,0,0,122,0,216,0,54,0,148,0,0,0,142,0,0,0,0,0,0,0,159,0,137,0,124,0,26,0,187,0,12,0,152,0,154,0,0,0,0,0,150,0,0,0,0,0,103,0,49,0,233,0,0,0,78,0,0,0,105,0,150,0,68,0,222,0,0,0,3,0,30,0,139,0,199,0,123,0,219,0,0,0,154,0,0,0,214,0,177,0,42,0,0,0,116,0,222,0,59,0,24,0,0,0,193,0,242,0,60,0,215,0,52,0,206,0,115,0,0,0,239,0,14,0,229,0,0,0,42,0,232,0,15,0,113,0,92,0,0,0,153,0,188,0,225,0,227,0,120,0,50,0,116,0,126,0,62,0,55,0,114,0,43,0,4,0,102,0,134,0,39,0,128,0,204,0,179,0,0,0,0,0,25,0,38,0,130,0,0,0,61,0,112,0,0,0,170,0,0,0,61,0,230,0,77,0,195,0,171,0,16,0,242,0,0,0,11,0,177,0,102,0,24,0,13,0,0,0,251,0,221,0,161,0,0,0,71,0,202,0,95,0,95,0,74,0,35,0,84,0,0,0,40,0,232,0,253,0,0,0,60,0,97,0,0,0,234,0,93,0,111,0,181,0,0,0,184,0,166,0,0,0,0,0,33,0,22,0,0,0,106,0,58,0,151,0,0,0,0,0,101,0,95,0,226,0,253,0,0,0,211,0,129,0,0,0,224,0,0,0,162,0,117,0,220,0,162,0,245,0,106,0,6,0,220,0,183,0,83,0,0,0,165,0,101,0,149,0,190,0,244,0,169,0,0,0,145,0,26,0,0,0,73,0,101,0,0,0,235,0,155,0,119,0,0,0,25,0,178,0,225,0,253,0,38,0,106,0,236,0,0,0,214,0,0,0,205,0,33,0,135,0,30,0,0,0,24,0,169,0,101,0,23,0,192,0,126,0,207,0,0,0,157,0,25,0,22,0,194,0,0,0,245,0,124,0,33,0,172,0,167,0,95,0,102,0,15,0,161,0,51,0,202,0,86,0,254,0,244,0,0,0,161,0,148,0,73,0,0,0,235,0,92,0,98,0,0,0,0,0,0,0,157,0,0,0,157,0,250,0,0,0,6,0,180,0,0,0,0,0,112,0,212,0,184,0,241,0,0,0,1,0,253,0,24,0,175,0,37,0,0,0,132,0,0,0,0,0,42,0,0,0,0,0,138,0,111,0,193,0,238,0,83,0,0,0,178,0,75,0,0,0,56,0,0,0,220,0,193,0,96,0,91,0,125,0,0,0,158,0,0,0,0,0,229,0,0,0,187,0,105,0,0,0,243,0,156,0,0,0,1,0,48,0,239,0,67,0,225,0,82,0,165,0,167,0,99,0,43,0,98,0,252,0,176,0,138,0,0,0,104,0,26,0,0,0,118,0,29,0,123,0,28,0,187,0,0,0,134,0,0,0,27,0,226,0,0,0,116,0,179,0,78,0,0,0,62,0,0,0,106,0,14,0,197,0,160,0,0,0,236,0,195,0,0,0,120,0,0,0,166,0,142,0,80,0,178,0,0,0,0,0,0,0,0,0,221,0,33,0,177,0,168,0,221,0,0,0,0,0,246,0,171,0,81,0,198,0,189,0,11,0,72,0,127,0,0,0,65,0,0,0,0,0,193,0,142,0,0,0,202,0,80,0,164,0,154,0,7,0,93,0,4,0,29,0,231,0,21,0,53,0,195,0,13,0,56,0,217,0,188,0,55,0,247,0,96,0,155,0,39,0,180,0,220,0,2,0,98,0,119,0,241,0,74,0,161,0,88,0,175,0,0,0,138,0,5,0,76,0,120,0,44,0,219,0,21,0,0,0,152,0,40,0,0,0,183,0,61,0,51,0,0,0,0,0,0,0,0,0,20,0,94,0,198,0,20,0,231,0,233,0,210,0,11,0,136,0,17,0,188,0,74,0,160,0,218,0,9,0,45,0,11,0,21,0,1,0,150,0,14,0,102,0,180,0,0,0,0,0);
signal scenario_full  : scenario_type := (200,31,213,31,138,31,64,31,4,31,4,30,175,31,175,30,120,31,120,30,249,31,209,31,243,31,117,31,125,31,125,30,125,29,251,31,98,31,253,31,162,31,207,31,207,30,207,29,207,28,38,31,202,31,253,31,50,31,50,30,141,31,121,31,66,31,2,31,11,31,99,31,99,30,77,31,77,30,23,31,252,31,157,31,73,31,105,31,105,30,121,31,170,31,44,31,150,31,55,31,37,31,188,31,188,30,56,31,56,30,160,31,180,31,229,31,26,31,247,31,92,31,92,30,104,31,38,31,75,31,97,31,93,31,129,31,244,31,244,30,182,31,182,30,93,31,93,30,138,31,138,30,138,29,224,31,224,30,119,31,119,30,198,31,205,31,205,30,231,31,70,31,32,31,32,30,252,31,64,31,125,31,230,31,101,31,154,31,1,31,100,31,48,31,80,31,37,31,32,31,32,30,196,31,15,31,216,31,216,30,238,31,123,31,20,31,185,31,204,31,179,31,242,31,242,30,242,29,160,31,128,31,222,31,219,31,204,31,254,31,29,31,95,31,18,31,18,30,92,31,87,31,50,31,252,31,140,31,249,31,172,31,129,31,231,31,87,31,59,31,113,31,21,31,84,31,119,31,119,30,123,31,195,31,241,31,241,30,241,29,44,31,227,31,219,31,18,31,136,31,160,31,217,31,217,30,130,31,137,31,137,30,18,31,190,31,42,31,90,31,227,31,168,31,80,31,103,31,9,31,138,31,85,31,85,30,41,31,91,31,199,31,180,31,227,31,227,30,7,31,67,31,179,31,8,31,8,30,98,31,243,31,95,31,2,31,187,31,215,31,83,31,81,31,236,31,114,31,191,31,156,31,14,31,14,30,248,31,121,31,234,31,157,31,201,31,177,31,128,31,219,31,219,30,217,31,217,30,36,31,217,31,156,31,156,30,70,31,104,31,143,31,77,31,153,31,153,30,15,31,222,31,202,31,92,31,229,31,136,31,69,31,103,31,41,31,148,31,73,31,56,31,234,31,152,31,93,31,141,31,167,31,167,30,23,31,23,30,193,31,219,31,252,31,252,30,169,31,49,31,6,31,6,30,127,31,228,31,62,31,30,31,221,31,75,31,171,31,139,31,62,31,6,31,6,30,6,29,227,31,111,31,111,30,158,31,160,31,160,30,160,29,59,31,59,30,222,31,241,31,241,30,246,31,119,31,88,31,88,30,251,31,179,31,69,31,15,31,15,30,151,31,43,31,54,31,8,31,91,31,242,31,183,31,183,30,168,31,122,31,179,31,83,31,109,31,117,31,117,30,197,31,19,31,70,31,24,31,25,31,50,31,124,31,65,31,202,31,119,31,203,31,88,31,168,31,81,31,81,30,81,29,222,31,17,31,62,31,100,31,140,31,140,30,140,29,5,31,147,31,147,30,167,31,221,31,219,31,202,31,238,31,199,31,232,31,175,31,176,31,28,31,83,31,215,31,168,31,207,31,207,30,197,31,190,31,178,31,178,30,183,31,115,31,162,31,217,31,217,30,53,31,3,31,3,30,192,31,168,31,158,31,105,31,124,31,185,31,222,31,171,31,113,31,110,31,20,31,20,30,2,31,2,30,156,31,156,30,156,29,192,31,193,31,39,31,39,30,109,31,24,31,14,31,14,30,221,31,221,30,51,31,26,31,217,31,53,31,209,31,209,30,205,31,234,31,198,31,20,31,20,30,20,29,134,31,3,31,158,31,211,31,211,30,44,31,217,31,217,30,28,31,228,31,231,31,74,31,213,31,40,31,40,30,13,31,147,31,96,31,96,30,124,31,124,30,124,29,71,31,71,30,135,31,249,31,20,31,140,31,86,31,21,31,130,31,227,31,190,31,49,31,60,31,60,30,40,31,40,30,165,31,166,31,207,31,42,31,42,30,42,29,189,31,65,31,227,31,72,31,168,31,129,31,129,30,251,31,1,31,157,31,252,31,63,31,207,31,243,31,21,31,239,31,239,30,59,31,196,31,182,31,57,31,57,30,80,31,80,30,33,31,167,31,157,31,14,31,123,31,250,31,250,30,250,29,57,31,52,31,25,31,16,31,161,31,50,31,143,31,224,31,122,31,143,31,88,31,53,31,53,30,190,31,109,31,154,31,160,31,99,31,172,31,200,31,203,31,50,31,193,31,179,31,251,31,201,31,19,31,33,31,75,31,75,30,75,29,86,31,124,31,224,31,142,31,217,31,187,31,171,31,253,31,197,31,216,31,240,31,217,31,118,31,30,31,134,31,49,31,49,30,35,31,100,31,96,31,109,31,111,31,200,31,122,31,60,31,68,31,68,30,122,31,216,31,54,31,148,31,148,30,142,31,142,30,142,29,142,28,159,31,137,31,124,31,26,31,187,31,12,31,152,31,154,31,154,30,154,29,150,31,150,30,150,29,103,31,49,31,233,31,233,30,78,31,78,30,105,31,150,31,68,31,222,31,222,30,3,31,30,31,139,31,199,31,123,31,219,31,219,30,154,31,154,30,214,31,177,31,42,31,42,30,116,31,222,31,59,31,24,31,24,30,193,31,242,31,60,31,215,31,52,31,206,31,115,31,115,30,239,31,14,31,229,31,229,30,42,31,232,31,15,31,113,31,92,31,92,30,153,31,188,31,225,31,227,31,120,31,50,31,116,31,126,31,62,31,55,31,114,31,43,31,4,31,102,31,134,31,39,31,128,31,204,31,179,31,179,30,179,29,25,31,38,31,130,31,130,30,61,31,112,31,112,30,170,31,170,30,61,31,230,31,77,31,195,31,171,31,16,31,242,31,242,30,11,31,177,31,102,31,24,31,13,31,13,30,251,31,221,31,161,31,161,30,71,31,202,31,95,31,95,31,74,31,35,31,84,31,84,30,40,31,232,31,253,31,253,30,60,31,97,31,97,30,234,31,93,31,111,31,181,31,181,30,184,31,166,31,166,30,166,29,33,31,22,31,22,30,106,31,58,31,151,31,151,30,151,29,101,31,95,31,226,31,253,31,253,30,211,31,129,31,129,30,224,31,224,30,162,31,117,31,220,31,162,31,245,31,106,31,6,31,220,31,183,31,83,31,83,30,165,31,101,31,149,31,190,31,244,31,169,31,169,30,145,31,26,31,26,30,73,31,101,31,101,30,235,31,155,31,119,31,119,30,25,31,178,31,225,31,253,31,38,31,106,31,236,31,236,30,214,31,214,30,205,31,33,31,135,31,30,31,30,30,24,31,169,31,101,31,23,31,192,31,126,31,207,31,207,30,157,31,25,31,22,31,194,31,194,30,245,31,124,31,33,31,172,31,167,31,95,31,102,31,15,31,161,31,51,31,202,31,86,31,254,31,244,31,244,30,161,31,148,31,73,31,73,30,235,31,92,31,98,31,98,30,98,29,98,28,157,31,157,30,157,31,250,31,250,30,6,31,180,31,180,30,180,29,112,31,212,31,184,31,241,31,241,30,1,31,253,31,24,31,175,31,37,31,37,30,132,31,132,30,132,29,42,31,42,30,42,29,138,31,111,31,193,31,238,31,83,31,83,30,178,31,75,31,75,30,56,31,56,30,220,31,193,31,96,31,91,31,125,31,125,30,158,31,158,30,158,29,229,31,229,30,187,31,105,31,105,30,243,31,156,31,156,30,1,31,48,31,239,31,67,31,225,31,82,31,165,31,167,31,99,31,43,31,98,31,252,31,176,31,138,31,138,30,104,31,26,31,26,30,118,31,29,31,123,31,28,31,187,31,187,30,134,31,134,30,27,31,226,31,226,30,116,31,179,31,78,31,78,30,62,31,62,30,106,31,14,31,197,31,160,31,160,30,236,31,195,31,195,30,120,31,120,30,166,31,142,31,80,31,178,31,178,30,178,29,178,28,178,27,221,31,33,31,177,31,168,31,221,31,221,30,221,29,246,31,171,31,81,31,198,31,189,31,11,31,72,31,127,31,127,30,65,31,65,30,65,29,193,31,142,31,142,30,202,31,80,31,164,31,154,31,7,31,93,31,4,31,29,31,231,31,21,31,53,31,195,31,13,31,56,31,217,31,188,31,55,31,247,31,96,31,155,31,39,31,180,31,220,31,2,31,98,31,119,31,241,31,74,31,161,31,88,31,175,31,175,30,138,31,5,31,76,31,120,31,44,31,219,31,21,31,21,30,152,31,40,31,40,30,183,31,61,31,51,31,51,30,51,29,51,28,51,27,20,31,94,31,198,31,20,31,231,31,233,31,210,31,11,31,136,31,17,31,188,31,74,31,160,31,218,31,9,31,45,31,11,31,21,31,1,31,150,31,14,31,102,31,180,31,180,30,180,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
