-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 253;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,0,0,0,0,91,0,33,0,60,0,104,0,0,0,0,0,109,0,96,0,183,0,38,0,244,0,20,0,0,0,254,0,143,0,97,0,110,0,248,0,95,0,169,0,0,0,19,0,159,0,68,0,91,0,184,0,0,0,204,0,242,0,109,0,23,0,0,0,192,0,160,0,0,0,5,0,167,0,27,0,147,0,79,0,32,0,245,0,0,0,215,0,0,0,194,0,130,0,207,0,150,0,135,0,0,0,124,0,255,0,77,0,0,0,165,0,128,0,117,0,4,0,196,0,220,0,230,0,223,0,174,0,83,0,18,0,0,0,75,0,183,0,30,0,100,0,31,0,0,0,43,0,195,0,0,0,20,0,84,0,45,0,0,0,116,0,107,0,121,0,25,0,125,0,0,0,137,0,0,0,222,0,137,0,56,0,0,0,57,0,127,0,218,0,6,0,35,0,148,0,0,0,203,0,0,0,255,0,187,0,138,0,138,0,39,0,49,0,49,0,57,0,240,0,138,0,0,0,208,0,237,0,0,0,229,0,117,0,216,0,0,0,220,0,167,0,45,0,8,0,165,0,189,0,0,0,217,0,235,0,0,0,114,0,28,0,96,0,0,0,169,0,42,0,0,0,55,0,163,0,0,0,91,0,1,0,82,0,194,0,6,0,24,0,228,0,232,0,0,0,140,0,96,0,53,0,0,0,129,0,224,0,47,0,19,0,122,0,38,0,239,0,128,0,136,0,0,0,46,0,0,0,247,0,177,0,95,0,245,0,0,0,64,0,66,0,220,0,12,0,0,0,61,0,93,0,146,0,189,0,92,0,119,0,138,0,9,0,21,0,152,0,55,0,44,0,0,0,0,0,229,0,0,0,85,0,0,0,49,0,88,0,59,0,0,0,0,0,162,0,69,0,23,0,175,0,144,0,87,0,178,0,16,0,208,0,0,0,191,0,105,0,16,0,133,0,227,0,85,0,237,0,0,0,39,0,77,0,40,0,0,0,161,0,174,0,186,0,10,0,0,0,250,0,0,0,44,0,97,0,0,0,29,0,242,0,104,0,247,0,34,0,23,0,54,0,0,0,91,0,67,0,0,0,103,0,162,0,0,0,97,0,0,0,79,0,120,0,249,0,153,0,84,0);
signal scenario_full  : scenario_type := (34,31,34,30,34,29,91,31,33,31,60,31,104,31,104,30,104,29,109,31,96,31,183,31,38,31,244,31,20,31,20,30,254,31,143,31,97,31,110,31,248,31,95,31,169,31,169,30,19,31,159,31,68,31,91,31,184,31,184,30,204,31,242,31,109,31,23,31,23,30,192,31,160,31,160,30,5,31,167,31,27,31,147,31,79,31,32,31,245,31,245,30,215,31,215,30,194,31,130,31,207,31,150,31,135,31,135,30,124,31,255,31,77,31,77,30,165,31,128,31,117,31,4,31,196,31,220,31,230,31,223,31,174,31,83,31,18,31,18,30,75,31,183,31,30,31,100,31,31,31,31,30,43,31,195,31,195,30,20,31,84,31,45,31,45,30,116,31,107,31,121,31,25,31,125,31,125,30,137,31,137,30,222,31,137,31,56,31,56,30,57,31,127,31,218,31,6,31,35,31,148,31,148,30,203,31,203,30,255,31,187,31,138,31,138,31,39,31,49,31,49,31,57,31,240,31,138,31,138,30,208,31,237,31,237,30,229,31,117,31,216,31,216,30,220,31,167,31,45,31,8,31,165,31,189,31,189,30,217,31,235,31,235,30,114,31,28,31,96,31,96,30,169,31,42,31,42,30,55,31,163,31,163,30,91,31,1,31,82,31,194,31,6,31,24,31,228,31,232,31,232,30,140,31,96,31,53,31,53,30,129,31,224,31,47,31,19,31,122,31,38,31,239,31,128,31,136,31,136,30,46,31,46,30,247,31,177,31,95,31,245,31,245,30,64,31,66,31,220,31,12,31,12,30,61,31,93,31,146,31,189,31,92,31,119,31,138,31,9,31,21,31,152,31,55,31,44,31,44,30,44,29,229,31,229,30,85,31,85,30,49,31,88,31,59,31,59,30,59,29,162,31,69,31,23,31,175,31,144,31,87,31,178,31,16,31,208,31,208,30,191,31,105,31,16,31,133,31,227,31,85,31,237,31,237,30,39,31,77,31,40,31,40,30,161,31,174,31,186,31,10,31,10,30,250,31,250,30,44,31,97,31,97,30,29,31,242,31,104,31,247,31,34,31,23,31,54,31,54,30,91,31,67,31,67,30,103,31,162,31,162,30,97,31,97,30,79,31,120,31,249,31,153,31,84,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
