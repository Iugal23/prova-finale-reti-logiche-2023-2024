-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_417 is
end project_tb_417;

architecture project_tb_arch_417 of project_tb_417 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 980;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (151,0,0,0,11,0,160,0,209,0,181,0,0,0,129,0,217,0,175,0,223,0,89,0,0,0,112,0,20,0,172,0,196,0,22,0,124,0,14,0,203,0,215,0,15,0,89,0,104,0,194,0,197,0,137,0,156,0,0,0,43,0,134,0,15,0,167,0,0,0,173,0,240,0,0,0,0,0,130,0,242,0,118,0,234,0,117,0,97,0,206,0,0,0,0,0,65,0,35,0,38,0,136,0,125,0,12,0,219,0,224,0,0,0,39,0,0,0,17,0,19,0,190,0,33,0,47,0,186,0,172,0,213,0,242,0,34,0,72,0,124,0,131,0,208,0,0,0,0,0,216,0,23,0,58,0,65,0,0,0,211,0,185,0,210,0,223,0,0,0,173,0,235,0,0,0,190,0,27,0,136,0,195,0,0,0,248,0,5,0,47,0,246,0,0,0,206,0,206,0,0,0,137,0,0,0,0,0,9,0,190,0,98,0,31,0,32,0,161,0,153,0,35,0,68,0,39,0,0,0,44,0,247,0,0,0,112,0,223,0,54,0,192,0,0,0,0,0,110,0,39,0,152,0,0,0,146,0,86,0,127,0,108,0,209,0,148,0,161,0,129,0,0,0,157,0,0,0,44,0,91,0,131,0,233,0,97,0,240,0,11,0,85,0,131,0,87,0,0,0,198,0,185,0,0,0,21,0,35,0,143,0,0,0,80,0,0,0,28,0,0,0,62,0,92,0,201,0,78,0,254,0,0,0,0,0,168,0,37,0,242,0,29,0,0,0,0,0,155,0,180,0,0,0,80,0,189,0,58,0,207,0,111,0,97,0,47,0,250,0,170,0,0,0,0,0,54,0,146,0,0,0,83,0,26,0,140,0,67,0,15,0,240,0,17,0,104,0,0,0,56,0,0,0,26,0,0,0,231,0,202,0,2,0,110,0,134,0,193,0,150,0,240,0,80,0,42,0,0,0,101,0,176,0,156,0,0,0,111,0,0,0,39,0,0,0,226,0,0,0,0,0,142,0,132,0,196,0,12,0,0,0,0,0,31,0,0,0,55,0,134,0,73,0,158,0,81,0,155,0,126,0,0,0,0,0,0,0,73,0,162,0,0,0,213,0,0,0,0,0,171,0,210,0,0,0,0,0,0,0,201,0,0,0,26,0,37,0,120,0,0,0,95,0,71,0,0,0,0,0,200,0,75,0,37,0,55,0,225,0,115,0,9,0,239,0,113,0,159,0,71,0,12,0,26,0,195,0,0,0,120,0,150,0,129,0,222,0,186,0,98,0,25,0,89,0,186,0,59,0,216,0,49,0,26,0,34,0,165,0,171,0,147,0,87,0,125,0,143,0,45,0,89,0,210,0,187,0,69,0,233,0,0,0,38,0,0,0,223,0,97,0,0,0,96,0,26,0,0,0,0,0,153,0,81,0,219,0,0,0,95,0,175,0,0,0,228,0,67,0,0,0,239,0,107,0,195,0,0,0,0,0,56,0,164,0,48,0,39,0,68,0,0,0,177,0,188,0,151,0,101,0,73,0,0,0,147,0,0,0,234,0,70,0,83,0,0,0,0,0,123,0,60,0,148,0,0,0,0,0,0,0,0,0,7,0,92,0,172,0,0,0,0,0,236,0,157,0,0,0,0,0,157,0,142,0,205,0,0,0,196,0,94,0,226,0,158,0,186,0,0,0,213,0,0,0,169,0,161,0,171,0,185,0,21,0,231,0,133,0,56,0,0,0,240,0,0,0,13,0,235,0,8,0,113,0,42,0,5,0,14,0,102,0,0,0,71,0,79,0,26,0,216,0,189,0,122,0,0,0,228,0,202,0,0,0,81,0,81,0,0,0,24,0,168,0,25,0,140,0,0,0,59,0,122,0,0,0,172,0,156,0,0,0,198,0,0,0,9,0,147,0,37,0,224,0,209,0,142,0,74,0,0,0,110,0,241,0,0,0,0,0,54,0,109,0,184,0,91,0,20,0,200,0,212,0,227,0,3,0,70,0,236,0,16,0,7,0,87,0,179,0,89,0,39,0,108,0,201,0,205,0,18,0,156,0,180,0,15,0,210,0,184,0,131,0,240,0,72,0,166,0,27,0,172,0,152,0,28,0,229,0,0,0,0,0,118,0,0,0,170,0,112,0,152,0,84,0,167,0,84,0,0,0,202,0,249,0,244,0,67,0,76,0,216,0,15,0,0,0,126,0,0,0,153,0,175,0,177,0,193,0,0,0,0,0,11,0,77,0,129,0,190,0,52,0,209,0,12,0,11,0,22,0,223,0,0,0,226,0,53,0,0,0,21,0,59,0,194,0,102,0,0,0,0,0,240,0,198,0,190,0,153,0,251,0,64,0,174,0,95,0,227,0,0,0,0,0,198,0,187,0,8,0,221,0,70,0,0,0,55,0,162,0,0,0,251,0,202,0,0,0,13,0,93,0,215,0,0,0,161,0,88,0,37,0,217,0,247,0,119,0,31,0,188,0,30,0,70,0,47,0,0,0,0,0,50,0,0,0,163,0,207,0,162,0,161,0,113,0,98,0,204,0,46,0,0,0,211,0,171,0,1,0,0,0,8,0,0,0,88,0,0,0,243,0,41,0,184,0,0,0,172,0,64,0,223,0,173,0,221,0,92,0,18,0,247,0,210,0,204,0,3,0,199,0,55,0,69,0,0,0,183,0,53,0,36,0,190,0,103,0,247,0,0,0,0,0,0,0,31,0,149,0,133,0,155,0,84,0,212,0,0,0,0,0,8,0,179,0,213,0,134,0,193,0,0,0,12,0,99,0,220,0,0,0,42,0,124,0,0,0,32,0,239,0,210,0,0,0,51,0,224,0,169,0,193,0,0,0,0,0,85,0,0,0,115,0,231,0,0,0,78,0,242,0,138,0,0,0,0,0,251,0,85,0,0,0,245,0,91,0,20,0,3,0,42,0,0,0,41,0,154,0,58,0,93,0,108,0,44,0,39,0,2,0,17,0,0,0,30,0,229,0,69,0,0,0,0,0,246,0,211,0,144,0,100,0,210,0,15,0,60,0,177,0,22,0,170,0,0,0,87,0,164,0,147,0,18,0,100,0,97,0,153,0,62,0,133,0,105,0,216,0,214,0,0,0,166,0,164,0,236,0,239,0,24,0,218,0,0,0,0,0,0,0,35,0,79,0,246,0,142,0,81,0,0,0,141,0,249,0,143,0,95,0,63,0,220,0,242,0,114,0,204,0,225,0,235,0,126,0,0,0,65,0,39,0,62,0,147,0,0,0,53,0,216,0,30,0,0,0,180,0,178,0,106,0,0,0,221,0,79,0,49,0,215,0,32,0,211,0,253,0,59,0,46,0,74,0,202,0,0,0,157,0,240,0,204,0,222,0,67,0,64,0,57,0,25,0,173,0,217,0,44,0,149,0,197,0,210,0,0,0,21,0,199,0,57,0,180,0,29,0,206,0,131,0,68,0,0,0,42,0,26,0,0,0,94,0,0,0,61,0,212,0,65,0,228,0,207,0,3,0,53,0,26,0,191,0,106,0,109,0,215,0,232,0,249,0,162,0,211,0,94,0,214,0,200,0,58,0,140,0,174,0,0,0,254,0,163,0,218,0,2,0,145,0,76,0,8,0,0,0,169,0,119,0,109,0,89,0,183,0,185,0,179,0,238,0,68,0,127,0,4,0,127,0,138,0,0,0,26,0,45,0,34,0,226,0,226,0,255,0,245,0,224,0,167,0,43,0,204,0,26,0,233,0,158,0,250,0,63,0,0,0,160,0,98,0,53,0,161,0,0,0,148,0,138,0,4,0,172,0,100,0,121,0,43,0,102,0,105,0,135,0,0,0,105,0,199,0,37,0,173,0,99,0,165,0,53,0,206,0,68,0,137,0,30,0,144,0,0,0,227,0,209,0,104,0,0,0,144,0,0,0,67,0,145,0,167,0,0,0,0,0,189,0,129,0,83,0,0,0,32,0,88,0,7,0,58,0,148,0,0,0,20,0,0,0,110,0,180,0,127,0,55,0,0,0,57,0,0,0,107,0,180,0,63,0,0,0,87,0,0,0,43,0,99,0,0,0,172,0,0,0,152,0,79,0,13,0,156,0,20,0,158,0,0,0,236,0,0,0,161,0,168,0,207,0,0,0,0,0,226,0,180,0,178,0,189,0,22,0,193,0,239,0,226,0,224,0,0,0,123,0,132,0,42,0,120,0,0,0,169,0,3,0,0,0,32,0,27,0,223,0,110,0,201,0,0,0,0,0,123,0,0,0,249,0,116,0,121,0,211,0,142,0,231,0,0,0,226,0,0,0,0,0,125,0,0,0,181,0,13,0,240,0,61,0,184,0,42,0,228,0,5,0,35,0,131,0,215,0,0,0,0,0,169,0,13,0,14,0,0,0,130,0,120,0);
signal scenario_full  : scenario_type := (151,31,151,30,11,31,160,31,209,31,181,31,181,30,129,31,217,31,175,31,223,31,89,31,89,30,112,31,20,31,172,31,196,31,22,31,124,31,14,31,203,31,215,31,15,31,89,31,104,31,194,31,197,31,137,31,156,31,156,30,43,31,134,31,15,31,167,31,167,30,173,31,240,31,240,30,240,29,130,31,242,31,118,31,234,31,117,31,97,31,206,31,206,30,206,29,65,31,35,31,38,31,136,31,125,31,12,31,219,31,224,31,224,30,39,31,39,30,17,31,19,31,190,31,33,31,47,31,186,31,172,31,213,31,242,31,34,31,72,31,124,31,131,31,208,31,208,30,208,29,216,31,23,31,58,31,65,31,65,30,211,31,185,31,210,31,223,31,223,30,173,31,235,31,235,30,190,31,27,31,136,31,195,31,195,30,248,31,5,31,47,31,246,31,246,30,206,31,206,31,206,30,137,31,137,30,137,29,9,31,190,31,98,31,31,31,32,31,161,31,153,31,35,31,68,31,39,31,39,30,44,31,247,31,247,30,112,31,223,31,54,31,192,31,192,30,192,29,110,31,39,31,152,31,152,30,146,31,86,31,127,31,108,31,209,31,148,31,161,31,129,31,129,30,157,31,157,30,44,31,91,31,131,31,233,31,97,31,240,31,11,31,85,31,131,31,87,31,87,30,198,31,185,31,185,30,21,31,35,31,143,31,143,30,80,31,80,30,28,31,28,30,62,31,92,31,201,31,78,31,254,31,254,30,254,29,168,31,37,31,242,31,29,31,29,30,29,29,155,31,180,31,180,30,80,31,189,31,58,31,207,31,111,31,97,31,47,31,250,31,170,31,170,30,170,29,54,31,146,31,146,30,83,31,26,31,140,31,67,31,15,31,240,31,17,31,104,31,104,30,56,31,56,30,26,31,26,30,231,31,202,31,2,31,110,31,134,31,193,31,150,31,240,31,80,31,42,31,42,30,101,31,176,31,156,31,156,30,111,31,111,30,39,31,39,30,226,31,226,30,226,29,142,31,132,31,196,31,12,31,12,30,12,29,31,31,31,30,55,31,134,31,73,31,158,31,81,31,155,31,126,31,126,30,126,29,126,28,73,31,162,31,162,30,213,31,213,30,213,29,171,31,210,31,210,30,210,29,210,28,201,31,201,30,26,31,37,31,120,31,120,30,95,31,71,31,71,30,71,29,200,31,75,31,37,31,55,31,225,31,115,31,9,31,239,31,113,31,159,31,71,31,12,31,26,31,195,31,195,30,120,31,150,31,129,31,222,31,186,31,98,31,25,31,89,31,186,31,59,31,216,31,49,31,26,31,34,31,165,31,171,31,147,31,87,31,125,31,143,31,45,31,89,31,210,31,187,31,69,31,233,31,233,30,38,31,38,30,223,31,97,31,97,30,96,31,26,31,26,30,26,29,153,31,81,31,219,31,219,30,95,31,175,31,175,30,228,31,67,31,67,30,239,31,107,31,195,31,195,30,195,29,56,31,164,31,48,31,39,31,68,31,68,30,177,31,188,31,151,31,101,31,73,31,73,30,147,31,147,30,234,31,70,31,83,31,83,30,83,29,123,31,60,31,148,31,148,30,148,29,148,28,148,27,7,31,92,31,172,31,172,30,172,29,236,31,157,31,157,30,157,29,157,31,142,31,205,31,205,30,196,31,94,31,226,31,158,31,186,31,186,30,213,31,213,30,169,31,161,31,171,31,185,31,21,31,231,31,133,31,56,31,56,30,240,31,240,30,13,31,235,31,8,31,113,31,42,31,5,31,14,31,102,31,102,30,71,31,79,31,26,31,216,31,189,31,122,31,122,30,228,31,202,31,202,30,81,31,81,31,81,30,24,31,168,31,25,31,140,31,140,30,59,31,122,31,122,30,172,31,156,31,156,30,198,31,198,30,9,31,147,31,37,31,224,31,209,31,142,31,74,31,74,30,110,31,241,31,241,30,241,29,54,31,109,31,184,31,91,31,20,31,200,31,212,31,227,31,3,31,70,31,236,31,16,31,7,31,87,31,179,31,89,31,39,31,108,31,201,31,205,31,18,31,156,31,180,31,15,31,210,31,184,31,131,31,240,31,72,31,166,31,27,31,172,31,152,31,28,31,229,31,229,30,229,29,118,31,118,30,170,31,112,31,152,31,84,31,167,31,84,31,84,30,202,31,249,31,244,31,67,31,76,31,216,31,15,31,15,30,126,31,126,30,153,31,175,31,177,31,193,31,193,30,193,29,11,31,77,31,129,31,190,31,52,31,209,31,12,31,11,31,22,31,223,31,223,30,226,31,53,31,53,30,21,31,59,31,194,31,102,31,102,30,102,29,240,31,198,31,190,31,153,31,251,31,64,31,174,31,95,31,227,31,227,30,227,29,198,31,187,31,8,31,221,31,70,31,70,30,55,31,162,31,162,30,251,31,202,31,202,30,13,31,93,31,215,31,215,30,161,31,88,31,37,31,217,31,247,31,119,31,31,31,188,31,30,31,70,31,47,31,47,30,47,29,50,31,50,30,163,31,207,31,162,31,161,31,113,31,98,31,204,31,46,31,46,30,211,31,171,31,1,31,1,30,8,31,8,30,88,31,88,30,243,31,41,31,184,31,184,30,172,31,64,31,223,31,173,31,221,31,92,31,18,31,247,31,210,31,204,31,3,31,199,31,55,31,69,31,69,30,183,31,53,31,36,31,190,31,103,31,247,31,247,30,247,29,247,28,31,31,149,31,133,31,155,31,84,31,212,31,212,30,212,29,8,31,179,31,213,31,134,31,193,31,193,30,12,31,99,31,220,31,220,30,42,31,124,31,124,30,32,31,239,31,210,31,210,30,51,31,224,31,169,31,193,31,193,30,193,29,85,31,85,30,115,31,231,31,231,30,78,31,242,31,138,31,138,30,138,29,251,31,85,31,85,30,245,31,91,31,20,31,3,31,42,31,42,30,41,31,154,31,58,31,93,31,108,31,44,31,39,31,2,31,17,31,17,30,30,31,229,31,69,31,69,30,69,29,246,31,211,31,144,31,100,31,210,31,15,31,60,31,177,31,22,31,170,31,170,30,87,31,164,31,147,31,18,31,100,31,97,31,153,31,62,31,133,31,105,31,216,31,214,31,214,30,166,31,164,31,236,31,239,31,24,31,218,31,218,30,218,29,218,28,35,31,79,31,246,31,142,31,81,31,81,30,141,31,249,31,143,31,95,31,63,31,220,31,242,31,114,31,204,31,225,31,235,31,126,31,126,30,65,31,39,31,62,31,147,31,147,30,53,31,216,31,30,31,30,30,180,31,178,31,106,31,106,30,221,31,79,31,49,31,215,31,32,31,211,31,253,31,59,31,46,31,74,31,202,31,202,30,157,31,240,31,204,31,222,31,67,31,64,31,57,31,25,31,173,31,217,31,44,31,149,31,197,31,210,31,210,30,21,31,199,31,57,31,180,31,29,31,206,31,131,31,68,31,68,30,42,31,26,31,26,30,94,31,94,30,61,31,212,31,65,31,228,31,207,31,3,31,53,31,26,31,191,31,106,31,109,31,215,31,232,31,249,31,162,31,211,31,94,31,214,31,200,31,58,31,140,31,174,31,174,30,254,31,163,31,218,31,2,31,145,31,76,31,8,31,8,30,169,31,119,31,109,31,89,31,183,31,185,31,179,31,238,31,68,31,127,31,4,31,127,31,138,31,138,30,26,31,45,31,34,31,226,31,226,31,255,31,245,31,224,31,167,31,43,31,204,31,26,31,233,31,158,31,250,31,63,31,63,30,160,31,98,31,53,31,161,31,161,30,148,31,138,31,4,31,172,31,100,31,121,31,43,31,102,31,105,31,135,31,135,30,105,31,199,31,37,31,173,31,99,31,165,31,53,31,206,31,68,31,137,31,30,31,144,31,144,30,227,31,209,31,104,31,104,30,144,31,144,30,67,31,145,31,167,31,167,30,167,29,189,31,129,31,83,31,83,30,32,31,88,31,7,31,58,31,148,31,148,30,20,31,20,30,110,31,180,31,127,31,55,31,55,30,57,31,57,30,107,31,180,31,63,31,63,30,87,31,87,30,43,31,99,31,99,30,172,31,172,30,152,31,79,31,13,31,156,31,20,31,158,31,158,30,236,31,236,30,161,31,168,31,207,31,207,30,207,29,226,31,180,31,178,31,189,31,22,31,193,31,239,31,226,31,224,31,224,30,123,31,132,31,42,31,120,31,120,30,169,31,3,31,3,30,32,31,27,31,223,31,110,31,201,31,201,30,201,29,123,31,123,30,249,31,116,31,121,31,211,31,142,31,231,31,231,30,226,31,226,30,226,29,125,31,125,30,181,31,13,31,240,31,61,31,184,31,42,31,228,31,5,31,35,31,131,31,215,31,215,30,215,29,169,31,13,31,14,31,14,30,130,31,120,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
