-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_75 is
end project_tb_75;

architecture project_tb_arch_75 of project_tb_75 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 312;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,219,0,41,0,239,0,0,0,210,0,139,0,95,0,116,0,243,0,255,0,0,0,0,0,137,0,0,0,166,0,28,0,116,0,233,0,223,0,153,0,150,0,117,0,254,0,0,0,112,0,82,0,235,0,13,0,175,0,0,0,147,0,0,0,157,0,0,0,9,0,24,0,248,0,78,0,70,0,12,0,236,0,73,0,0,0,6,0,94,0,135,0,210,0,0,0,119,0,147,0,110,0,142,0,0,0,212,0,248,0,58,0,112,0,0,0,4,0,212,0,0,0,197,0,49,0,0,0,104,0,248,0,97,0,186,0,218,0,214,0,106,0,190,0,103,0,100,0,0,0,84,0,93,0,0,0,35,0,233,0,226,0,105,0,153,0,0,0,29,0,115,0,162,0,60,0,191,0,65,0,195,0,79,0,172,0,55,0,8,0,158,0,190,0,211,0,5,0,200,0,196,0,0,0,81,0,147,0,176,0,4,0,183,0,240,0,3,0,39,0,38,0,50,0,0,0,0,0,56,0,34,0,186,0,0,0,92,0,0,0,178,0,43,0,0,0,46,0,103,0,126,0,99,0,159,0,53,0,53,0,0,0,61,0,156,0,194,0,98,0,221,0,58,0,0,0,209,0,107,0,168,0,60,0,124,0,158,0,166,0,192,0,0,0,195,0,223,0,0,0,86,0,213,0,0,0,76,0,190,0,109,0,0,0,140,0,67,0,0,0,196,0,13,0,115,0,0,0,38,0,104,0,76,0,193,0,27,0,89,0,27,0,100,0,16,0,100,0,0,0,173,0,0,0,221,0,214,0,216,0,228,0,230,0,100,0,0,0,0,0,70,0,0,0,202,0,25,0,0,0,247,0,93,0,204,0,0,0,0,0,172,0,84,0,238,0,61,0,66,0,109,0,0,0,208,0,206,0,110,0,0,0,153,0,195,0,59,0,215,0,133,0,202,0,101,0,0,0,151,0,0,0,0,0,213,0,71,0,177,0,226,0,43,0,136,0,218,0,0,0,35,0,52,0,99,0,27,0,0,0,66,0,34,0,127,0,156,0,235,0,104,0,0,0,69,0,0,0,0,0,0,0,93,0,26,0,118,0,111,0,131,0,125,0,47,0,248,0,13,0,131,0,244,0,4,0,13,0,63,0,200,0,102,0,61,0,146,0,113,0,0,0,95,0,175,0,203,0,0,0,159,0,0,0,69,0,133,0,88,0,214,0,42,0,229,0,226,0,21,0,210,0,180,0,180,0,214,0,0,0,185,0,196,0,23,0,225,0,165,0,0,0,86,0,134,0,95,0,44,0,9,0,23,0,84,0,149,0,0,0,56,0,223,0,249,0,117,0,62,0,18,0,78,0,147,0,57,0,221,0,106,0,93,0,233,0,0,0,248,0,0,0);
signal scenario_full  : scenario_type := (0,0,219,31,41,31,239,31,239,30,210,31,139,31,95,31,116,31,243,31,255,31,255,30,255,29,137,31,137,30,166,31,28,31,116,31,233,31,223,31,153,31,150,31,117,31,254,31,254,30,112,31,82,31,235,31,13,31,175,31,175,30,147,31,147,30,157,31,157,30,9,31,24,31,248,31,78,31,70,31,12,31,236,31,73,31,73,30,6,31,94,31,135,31,210,31,210,30,119,31,147,31,110,31,142,31,142,30,212,31,248,31,58,31,112,31,112,30,4,31,212,31,212,30,197,31,49,31,49,30,104,31,248,31,97,31,186,31,218,31,214,31,106,31,190,31,103,31,100,31,100,30,84,31,93,31,93,30,35,31,233,31,226,31,105,31,153,31,153,30,29,31,115,31,162,31,60,31,191,31,65,31,195,31,79,31,172,31,55,31,8,31,158,31,190,31,211,31,5,31,200,31,196,31,196,30,81,31,147,31,176,31,4,31,183,31,240,31,3,31,39,31,38,31,50,31,50,30,50,29,56,31,34,31,186,31,186,30,92,31,92,30,178,31,43,31,43,30,46,31,103,31,126,31,99,31,159,31,53,31,53,31,53,30,61,31,156,31,194,31,98,31,221,31,58,31,58,30,209,31,107,31,168,31,60,31,124,31,158,31,166,31,192,31,192,30,195,31,223,31,223,30,86,31,213,31,213,30,76,31,190,31,109,31,109,30,140,31,67,31,67,30,196,31,13,31,115,31,115,30,38,31,104,31,76,31,193,31,27,31,89,31,27,31,100,31,16,31,100,31,100,30,173,31,173,30,221,31,214,31,216,31,228,31,230,31,100,31,100,30,100,29,70,31,70,30,202,31,25,31,25,30,247,31,93,31,204,31,204,30,204,29,172,31,84,31,238,31,61,31,66,31,109,31,109,30,208,31,206,31,110,31,110,30,153,31,195,31,59,31,215,31,133,31,202,31,101,31,101,30,151,31,151,30,151,29,213,31,71,31,177,31,226,31,43,31,136,31,218,31,218,30,35,31,52,31,99,31,27,31,27,30,66,31,34,31,127,31,156,31,235,31,104,31,104,30,69,31,69,30,69,29,69,28,93,31,26,31,118,31,111,31,131,31,125,31,47,31,248,31,13,31,131,31,244,31,4,31,13,31,63,31,200,31,102,31,61,31,146,31,113,31,113,30,95,31,175,31,203,31,203,30,159,31,159,30,69,31,133,31,88,31,214,31,42,31,229,31,226,31,21,31,210,31,180,31,180,31,214,31,214,30,185,31,196,31,23,31,225,31,165,31,165,30,86,31,134,31,95,31,44,31,9,31,23,31,84,31,149,31,149,30,56,31,223,31,249,31,117,31,62,31,18,31,78,31,147,31,57,31,221,31,106,31,93,31,233,31,233,30,248,31,248,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
