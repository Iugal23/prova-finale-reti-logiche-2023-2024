-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 294;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (198,0,224,0,150,0,0,0,0,0,246,0,162,0,178,0,226,0,49,0,28,0,0,0,0,0,0,0,158,0,27,0,116,0,186,0,194,0,30,0,208,0,0,0,46,0,0,0,151,0,45,0,0,0,162,0,0,0,6,0,180,0,242,0,45,0,144,0,75,0,240,0,177,0,0,0,7,0,204,0,44,0,29,0,223,0,23,0,120,0,28,0,166,0,37,0,34,0,0,0,3,0,0,0,61,0,188,0,26,0,56,0,81,0,230,0,164,0,28,0,225,0,0,0,41,0,96,0,205,0,77,0,187,0,197,0,91,0,105,0,238,0,31,0,144,0,0,0,205,0,101,0,25,0,198,0,121,0,211,0,23,0,0,0,94,0,197,0,0,0,53,0,188,0,56,0,185,0,14,0,160,0,179,0,129,0,77,0,187,0,126,0,183,0,225,0,201,0,154,0,42,0,184,0,0,0,43,0,49,0,165,0,191,0,154,0,0,0,67,0,211,0,0,0,91,0,117,0,110,0,123,0,0,0,0,0,0,0,127,0,0,0,0,0,3,0,150,0,16,0,103,0,22,0,22,0,24,0,171,0,0,0,20,0,94,0,0,0,178,0,52,0,109,0,97,0,248,0,0,0,194,0,31,0,134,0,28,0,136,0,140,0,77,0,0,0,226,0,83,0,250,0,220,0,85,0,85,0,0,0,0,0,157,0,184,0,124,0,123,0,178,0,0,0,0,0,202,0,63,0,0,0,204,0,215,0,79,0,249,0,182,0,221,0,211,0,0,0,82,0,229,0,165,0,149,0,248,0,54,0,158,0,0,0,232,0,62,0,7,0,85,0,149,0,191,0,167,0,80,0,240,0,5,0,0,0,70,0,194,0,77,0,130,0,0,0,50,0,0,0,53,0,149,0,0,0,67,0,0,0,85,0,0,0,166,0,87,0,66,0,102,0,124,0,96,0,0,0,160,0,0,0,216,0,0,0,40,0,81,0,203,0,27,0,110,0,96,0,141,0,46,0,121,0,144,0,32,0,144,0,0,0,192,0,0,0,138,0,0,0,112,0,186,0,101,0,199,0,82,0,0,0,244,0,246,0,249,0,39,0,19,0,95,0,84,0,237,0,182,0,0,0,55,0,44,0,154,0,136,0,74,0,32,0,126,0,173,0,234,0,13,0,0,0,137,0,0,0,211,0,54,0,56,0,0,0,113,0,187,0,227,0,144,0,244,0,0,0,0,0,0,0,133,0,175,0,0,0,0,0,68,0,0,0,141,0,171,0,24,0,112,0,34,0,187,0,136,0,76,0,206,0,173,0,125,0,125,0);
signal scenario_full  : scenario_type := (198,31,224,31,150,31,150,30,150,29,246,31,162,31,178,31,226,31,49,31,28,31,28,30,28,29,28,28,158,31,27,31,116,31,186,31,194,31,30,31,208,31,208,30,46,31,46,30,151,31,45,31,45,30,162,31,162,30,6,31,180,31,242,31,45,31,144,31,75,31,240,31,177,31,177,30,7,31,204,31,44,31,29,31,223,31,23,31,120,31,28,31,166,31,37,31,34,31,34,30,3,31,3,30,61,31,188,31,26,31,56,31,81,31,230,31,164,31,28,31,225,31,225,30,41,31,96,31,205,31,77,31,187,31,197,31,91,31,105,31,238,31,31,31,144,31,144,30,205,31,101,31,25,31,198,31,121,31,211,31,23,31,23,30,94,31,197,31,197,30,53,31,188,31,56,31,185,31,14,31,160,31,179,31,129,31,77,31,187,31,126,31,183,31,225,31,201,31,154,31,42,31,184,31,184,30,43,31,49,31,165,31,191,31,154,31,154,30,67,31,211,31,211,30,91,31,117,31,110,31,123,31,123,30,123,29,123,28,127,31,127,30,127,29,3,31,150,31,16,31,103,31,22,31,22,31,24,31,171,31,171,30,20,31,94,31,94,30,178,31,52,31,109,31,97,31,248,31,248,30,194,31,31,31,134,31,28,31,136,31,140,31,77,31,77,30,226,31,83,31,250,31,220,31,85,31,85,31,85,30,85,29,157,31,184,31,124,31,123,31,178,31,178,30,178,29,202,31,63,31,63,30,204,31,215,31,79,31,249,31,182,31,221,31,211,31,211,30,82,31,229,31,165,31,149,31,248,31,54,31,158,31,158,30,232,31,62,31,7,31,85,31,149,31,191,31,167,31,80,31,240,31,5,31,5,30,70,31,194,31,77,31,130,31,130,30,50,31,50,30,53,31,149,31,149,30,67,31,67,30,85,31,85,30,166,31,87,31,66,31,102,31,124,31,96,31,96,30,160,31,160,30,216,31,216,30,40,31,81,31,203,31,27,31,110,31,96,31,141,31,46,31,121,31,144,31,32,31,144,31,144,30,192,31,192,30,138,31,138,30,112,31,186,31,101,31,199,31,82,31,82,30,244,31,246,31,249,31,39,31,19,31,95,31,84,31,237,31,182,31,182,30,55,31,44,31,154,31,136,31,74,31,32,31,126,31,173,31,234,31,13,31,13,30,137,31,137,30,211,31,54,31,56,31,56,30,113,31,187,31,227,31,144,31,244,31,244,30,244,29,244,28,133,31,175,31,175,30,175,29,68,31,68,30,141,31,171,31,24,31,112,31,34,31,187,31,136,31,76,31,206,31,173,31,125,31,125,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
