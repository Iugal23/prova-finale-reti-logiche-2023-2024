-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 620;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (52,0,3,0,129,0,142,0,39,0,5,0,228,0,16,0,106,0,19,0,95,0,14,0,87,0,226,0,0,0,185,0,223,0,0,0,182,0,154,0,181,0,117,0,28,0,75,0,0,0,241,0,163,0,119,0,0,0,194,0,18,0,195,0,218,0,238,0,91,0,186,0,140,0,130,0,214,0,145,0,158,0,119,0,155,0,131,0,0,0,110,0,15,0,0,0,0,0,0,0,0,0,187,0,20,0,66,0,0,0,0,0,0,0,218,0,154,0,236,0,0,0,0,0,233,0,0,0,155,0,169,0,0,0,0,0,200,0,0,0,0,0,0,0,213,0,194,0,193,0,26,0,0,0,54,0,40,0,95,0,162,0,154,0,92,0,0,0,8,0,214,0,0,0,238,0,212,0,58,0,58,0,57,0,190,0,25,0,212,0,0,0,72,0,0,0,17,0,27,0,27,0,0,0,123,0,77,0,145,0,0,0,254,0,217,0,117,0,0,0,239,0,120,0,31,0,62,0,198,0,182,0,81,0,0,0,168,0,0,0,147,0,231,0,149,0,90,0,29,0,178,0,0,0,144,0,0,0,74,0,214,0,0,0,113,0,0,0,66,0,21,0,128,0,155,0,61,0,247,0,137,0,42,0,215,0,61,0,232,0,117,0,112,0,234,0,0,0,184,0,178,0,76,0,250,0,0,0,148,0,0,0,0,0,62,0,18,0,211,0,0,0,95,0,237,0,62,0,115,0,79,0,212,0,211,0,0,0,34,0,175,0,191,0,0,0,83,0,191,0,193,0,128,0,231,0,106,0,87,0,89,0,50,0,0,0,0,0,84,0,41,0,140,0,160,0,0,0,175,0,0,0,246,0,0,0,193,0,200,0,2,0,0,0,224,0,0,0,0,0,150,0,230,0,39,0,164,0,62,0,199,0,152,0,229,0,216,0,69,0,236,0,151,0,252,0,123,0,20,0,0,0,232,0,49,0,163,0,0,0,219,0,91,0,13,0,154,0,169,0,5,0,0,0,71,0,0,0,112,0,0,0,0,0,58,0,95,0,137,0,106,0,125,0,166,0,15,0,238,0,26,0,184,0,176,0,0,0,0,0,72,0,205,0,0,0,0,0,252,0,187,0,100,0,193,0,67,0,198,0,181,0,0,0,14,0,69,0,134,0,34,0,105,0,61,0,16,0,26,0,194,0,100,0,199,0,208,0,216,0,242,0,0,0,20,0,196,0,0,0,237,0,104,0,0,0,139,0,0,0,228,0,72,0,129,0,0,0,139,0,178,0,95,0,216,0,172,0,134,0,61,0,34,0,166,0,132,0,199,0,121,0,56,0,30,0,252,0,70,0,0,0,63,0,28,0,0,0,131,0,0,0,70,0,182,0,230,0,159,0,0,0,95,0,136,0,202,0,0,0,45,0,219,0,156,0,170,0,94,0,201,0,0,0,28,0,120,0,0,0,0,0,41,0,254,0,176,0,79,0,231,0,0,0,105,0,0,0,166,0,114,0,60,0,28,0,0,0,85,0,87,0,130,0,213,0,245,0,0,0,20,0,184,0,169,0,95,0,200,0,246,0,0,0,13,0,166,0,20,0,0,0,2,0,0,0,0,0,186,0,147,0,199,0,247,0,129,0,26,0,127,0,155,0,3,0,191,0,0,0,0,0,37,0,52,0,8,0,18,0,215,0,204,0,106,0,0,0,116,0,115,0,0,0,0,0,68,0,3,0,178,0,21,0,102,0,131,0,181,0,0,0,0,0,5,0,0,0,72,0,55,0,75,0,55,0,95,0,71,0,0,0,31,0,30,0,181,0,50,0,0,0,12,0,198,0,225,0,111,0,207,0,245,0,0,0,8,0,191,0,16,0,140,0,0,0,138,0,22,0,149,0,187,0,96,0,240,0,164,0,159,0,0,0,145,0,0,0,251,0,0,0,35,0,223,0,240,0,0,0,0,0,140,0,188,0,238,0,183,0,248,0,231,0,32,0,163,0,0,0,185,0,0,0,31,0,26,0,59,0,106,0,99,0,235,0,202,0,98,0,92,0,157,0,236,0,152,0,0,0,81,0,204,0,157,0,26,0,0,0,67,0,195,0,211,0,69,0,41,0,0,0,40,0,177,0,76,0,38,0,121,0,235,0,96,0,82,0,0,0,233,0,104,0,67,0,151,0,116,0,222,0,0,0,0,0,252,0,64,0,201,0,0,0,194,0,0,0,62,0,0,0,69,0,0,0,245,0,91,0,0,0,7,0,184,0,0,0,58,0,189,0,0,0,0,0,43,0,48,0,218,0,0,0,172,0,215,0,0,0,21,0,88,0,0,0,162,0,188,0,210,0,91,0,0,0,54,0,110,0,89,0,86,0,39,0,0,0,10,0,251,0,57,0,227,0,51,0,183,0,198,0,249,0,141,0,129,0,141,0,5,0,182,0,80,0,103,0,144,0,123,0,90,0,221,0,17,0,200,0,82,0,0,0,0,0,0,0,85,0,212,0,186,0,183,0,71,0,151,0,246,0,144,0,34,0,0,0,237,0,206,0,226,0,0,0,0,0,0,0,0,0,0,0,227,0,7,0,44,0,97,0,71,0,227,0,176,0,46,0,237,0,0,0,64,0,197,0,0,0,0,0,252,0,221,0,0,0,69,0,0,0,177,0,0,0,212,0,18,0,101,0,124,0,230,0,0,0,54,0,98,0,246,0,239,0,117,0,0,0,216,0,127,0,110,0,0,0,161,0,234,0,15,0,112,0,15,0,0,0,0,0,161,0,103,0,138,0,0,0);
signal scenario_full  : scenario_type := (52,31,3,31,129,31,142,31,39,31,5,31,228,31,16,31,106,31,19,31,95,31,14,31,87,31,226,31,226,30,185,31,223,31,223,30,182,31,154,31,181,31,117,31,28,31,75,31,75,30,241,31,163,31,119,31,119,30,194,31,18,31,195,31,218,31,238,31,91,31,186,31,140,31,130,31,214,31,145,31,158,31,119,31,155,31,131,31,131,30,110,31,15,31,15,30,15,29,15,28,15,27,187,31,20,31,66,31,66,30,66,29,66,28,218,31,154,31,236,31,236,30,236,29,233,31,233,30,155,31,169,31,169,30,169,29,200,31,200,30,200,29,200,28,213,31,194,31,193,31,26,31,26,30,54,31,40,31,95,31,162,31,154,31,92,31,92,30,8,31,214,31,214,30,238,31,212,31,58,31,58,31,57,31,190,31,25,31,212,31,212,30,72,31,72,30,17,31,27,31,27,31,27,30,123,31,77,31,145,31,145,30,254,31,217,31,117,31,117,30,239,31,120,31,31,31,62,31,198,31,182,31,81,31,81,30,168,31,168,30,147,31,231,31,149,31,90,31,29,31,178,31,178,30,144,31,144,30,74,31,214,31,214,30,113,31,113,30,66,31,21,31,128,31,155,31,61,31,247,31,137,31,42,31,215,31,61,31,232,31,117,31,112,31,234,31,234,30,184,31,178,31,76,31,250,31,250,30,148,31,148,30,148,29,62,31,18,31,211,31,211,30,95,31,237,31,62,31,115,31,79,31,212,31,211,31,211,30,34,31,175,31,191,31,191,30,83,31,191,31,193,31,128,31,231,31,106,31,87,31,89,31,50,31,50,30,50,29,84,31,41,31,140,31,160,31,160,30,175,31,175,30,246,31,246,30,193,31,200,31,2,31,2,30,224,31,224,30,224,29,150,31,230,31,39,31,164,31,62,31,199,31,152,31,229,31,216,31,69,31,236,31,151,31,252,31,123,31,20,31,20,30,232,31,49,31,163,31,163,30,219,31,91,31,13,31,154,31,169,31,5,31,5,30,71,31,71,30,112,31,112,30,112,29,58,31,95,31,137,31,106,31,125,31,166,31,15,31,238,31,26,31,184,31,176,31,176,30,176,29,72,31,205,31,205,30,205,29,252,31,187,31,100,31,193,31,67,31,198,31,181,31,181,30,14,31,69,31,134,31,34,31,105,31,61,31,16,31,26,31,194,31,100,31,199,31,208,31,216,31,242,31,242,30,20,31,196,31,196,30,237,31,104,31,104,30,139,31,139,30,228,31,72,31,129,31,129,30,139,31,178,31,95,31,216,31,172,31,134,31,61,31,34,31,166,31,132,31,199,31,121,31,56,31,30,31,252,31,70,31,70,30,63,31,28,31,28,30,131,31,131,30,70,31,182,31,230,31,159,31,159,30,95,31,136,31,202,31,202,30,45,31,219,31,156,31,170,31,94,31,201,31,201,30,28,31,120,31,120,30,120,29,41,31,254,31,176,31,79,31,231,31,231,30,105,31,105,30,166,31,114,31,60,31,28,31,28,30,85,31,87,31,130,31,213,31,245,31,245,30,20,31,184,31,169,31,95,31,200,31,246,31,246,30,13,31,166,31,20,31,20,30,2,31,2,30,2,29,186,31,147,31,199,31,247,31,129,31,26,31,127,31,155,31,3,31,191,31,191,30,191,29,37,31,52,31,8,31,18,31,215,31,204,31,106,31,106,30,116,31,115,31,115,30,115,29,68,31,3,31,178,31,21,31,102,31,131,31,181,31,181,30,181,29,5,31,5,30,72,31,55,31,75,31,55,31,95,31,71,31,71,30,31,31,30,31,181,31,50,31,50,30,12,31,198,31,225,31,111,31,207,31,245,31,245,30,8,31,191,31,16,31,140,31,140,30,138,31,22,31,149,31,187,31,96,31,240,31,164,31,159,31,159,30,145,31,145,30,251,31,251,30,35,31,223,31,240,31,240,30,240,29,140,31,188,31,238,31,183,31,248,31,231,31,32,31,163,31,163,30,185,31,185,30,31,31,26,31,59,31,106,31,99,31,235,31,202,31,98,31,92,31,157,31,236,31,152,31,152,30,81,31,204,31,157,31,26,31,26,30,67,31,195,31,211,31,69,31,41,31,41,30,40,31,177,31,76,31,38,31,121,31,235,31,96,31,82,31,82,30,233,31,104,31,67,31,151,31,116,31,222,31,222,30,222,29,252,31,64,31,201,31,201,30,194,31,194,30,62,31,62,30,69,31,69,30,245,31,91,31,91,30,7,31,184,31,184,30,58,31,189,31,189,30,189,29,43,31,48,31,218,31,218,30,172,31,215,31,215,30,21,31,88,31,88,30,162,31,188,31,210,31,91,31,91,30,54,31,110,31,89,31,86,31,39,31,39,30,10,31,251,31,57,31,227,31,51,31,183,31,198,31,249,31,141,31,129,31,141,31,5,31,182,31,80,31,103,31,144,31,123,31,90,31,221,31,17,31,200,31,82,31,82,30,82,29,82,28,85,31,212,31,186,31,183,31,71,31,151,31,246,31,144,31,34,31,34,30,237,31,206,31,226,31,226,30,226,29,226,28,226,27,226,26,227,31,7,31,44,31,97,31,71,31,227,31,176,31,46,31,237,31,237,30,64,31,197,31,197,30,197,29,252,31,221,31,221,30,69,31,69,30,177,31,177,30,212,31,18,31,101,31,124,31,230,31,230,30,54,31,98,31,246,31,239,31,117,31,117,30,216,31,127,31,110,31,110,30,161,31,234,31,15,31,112,31,15,31,15,30,15,29,161,31,103,31,138,31,138,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
