-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_882 is
end project_tb_882;

architecture project_tb_arch_882 of project_tb_882 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 668;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (119,0,133,0,31,0,246,0,38,0,117,0,76,0,94,0,64,0,19,0,0,0,180,0,92,0,183,0,176,0,147,0,154,0,121,0,247,0,221,0,185,0,152,0,0,0,255,0,228,0,0,0,202,0,75,0,157,0,0,0,17,0,0,0,60,0,0,0,76,0,100,0,224,0,95,0,201,0,98,0,85,0,0,0,245,0,184,0,11,0,33,0,51,0,0,0,0,0,165,0,53,0,64,0,0,0,0,0,210,0,74,0,41,0,142,0,162,0,201,0,0,0,208,0,0,0,82,0,156,0,181,0,216,0,0,0,240,0,38,0,162,0,0,0,174,0,150,0,108,0,0,0,166,0,60,0,197,0,5,0,167,0,250,0,199,0,53,0,198,0,75,0,237,0,64,0,65,0,219,0,55,0,114,0,0,0,0,0,172,0,32,0,193,0,35,0,53,0,117,0,92,0,17,0,179,0,0,0,220,0,222,0,228,0,0,0,42,0,11,0,202,0,0,0,223,0,218,0,102,0,74,0,0,0,3,0,117,0,26,0,0,0,25,0,0,0,18,0,28,0,0,0,14,0,232,0,249,0,108,0,0,0,0,0,236,0,50,0,0,0,184,0,155,0,120,0,180,0,211,0,0,0,0,0,0,0,149,0,76,0,83,0,248,0,74,0,0,0,0,0,250,0,0,0,125,0,0,0,177,0,244,0,212,0,238,0,189,0,99,0,0,0,0,0,0,0,164,0,254,0,110,0,122,0,141,0,68,0,91,0,0,0,0,0,0,0,14,0,0,0,3,0,0,0,0,0,136,0,133,0,221,0,0,0,56,0,120,0,0,0,0,0,0,0,138,0,0,0,120,0,76,0,0,0,92,0,253,0,191,0,188,0,0,0,50,0,221,0,107,0,57,0,149,0,91,0,243,0,0,0,0,0,59,0,180,0,0,0,15,0,7,0,0,0,225,0,210,0,227,0,185,0,178,0,0,0,0,0,0,0,168,0,101,0,0,0,0,0,0,0,0,0,0,0,174,0,212,0,115,0,247,0,133,0,0,0,248,0,44,0,201,0,55,0,233,0,112,0,24,0,148,0,231,0,221,0,0,0,214,0,55,0,0,0,113,0,72,0,0,0,223,0,231,0,119,0,0,0,111,0,0,0,152,0,0,0,151,0,72,0,76,0,236,0,244,0,12,0,94,0,28,0,135,0,0,0,250,0,33,0,7,0,177,0,86,0,141,0,71,0,116,0,10,0,98,0,216,0,69,0,0,0,0,0,50,0,82,0,0,0,168,0,196,0,0,0,126,0,0,0,49,0,124,0,163,0,114,0,69,0,41,0,56,0,79,0,216,0,255,0,190,0,16,0,72,0,0,0,111,0,176,0,4,0,6,0,0,0,7,0,0,0,182,0,65,0,86,0,252,0,69,0,114,0,221,0,128,0,148,0,83,0,2,0,0,0,108,0,79,0,185,0,156,0,78,0,208,0,153,0,5,0,243,0,0,0,64,0,11,0,108,0,0,0,0,0,142,0,104,0,86,0,156,0,116,0,155,0,114,0,188,0,8,0,249,0,74,0,41,0,34,0,196,0,198,0,244,0,232,0,0,0,0,0,245,0,0,0,244,0,144,0,136,0,224,0,151,0,210,0,252,0,123,0,0,0,54,0,54,0,242,0,44,0,37,0,66,0,33,0,34,0,65,0,221,0,199,0,175,0,43,0,175,0,187,0,0,0,33,0,122,0,224,0,82,0,191,0,197,0,142,0,0,0,144,0,16,0,185,0,165,0,64,0,0,0,170,0,114,0,126,0,56,0,31,0,200,0,87,0,0,0,91,0,30,0,4,0,194,0,77,0,221,0,165,0,0,0,253,0,198,0,120,0,243,0,104,0,189,0,40,0,200,0,103,0,141,0,0,0,80,0,220,0,6,0,68,0,207,0,125,0,153,0,142,0,181,0,7,0,193,0,0,0,188,0,0,0,78,0,41,0,162,0,49,0,133,0,0,0,122,0,0,0,247,0,124,0,122,0,219,0,18,0,0,0,180,0,251,0,89,0,222,0,149,0,139,0,92,0,139,0,0,0,33,0,76,0,237,0,238,0,44,0,95,0,27,0,0,0,63,0,0,0,116,0,0,0,0,0,193,0,90,0,0,0,221,0,0,0,220,0,246,0,108,0,145,0,188,0,143,0,21,0,30,0,252,0,143,0,251,0,104,0,143,0,119,0,90,0,0,0,0,0,45,0,243,0,88,0,0,0,33,0,219,0,0,0,222,0,93,0,0,0,86,0,161,0,0,0,20,0,138,0,47,0,0,0,199,0,231,0,50,0,52,0,0,0,0,0,104,0,0,0,22,0,107,0,0,0,240,0,139,0,0,0,45,0,121,0,176,0,11,0,0,0,0,0,30,0,0,0,124,0,177,0,240,0,0,0,6,0,38,0,0,0,53,0,0,0,175,0,248,0,187,0,234,0,236,0,102,0,42,0,0,0,0,0,226,0,215,0,32,0,117,0,217,0,251,0,47,0,131,0,223,0,127,0,46,0,65,0,96,0,130,0,168,0,0,0,203,0,31,0,132,0,0,0,137,0,13,0,159,0,114,0,189,0,49,0,203,0,185,0,250,0,255,0,111,0,0,0,59,0,11,0,53,0,39,0,0,0,64,0,217,0,29,0,84,0,109,0,56,0,0,0,157,0,106,0,239,0,34,0,12,0,96,0,0,0,158,0,49,0,0,0,238,0,128,0,195,0,0,0,71,0,0,0,0,0,190,0,0,0,158,0,0,0,141,0,104,0,150,0,200,0,0,0,225,0,0,0,40,0,128,0,102,0,105,0,245,0,102,0,190,0,249,0,0,0,214,0,176,0,203,0,64,0,66,0,252,0,93,0,12,0,98,0,62,0,183,0,175,0,213,0,227,0,186,0,201,0,247,0,0,0,203,0,91,0,0,0,0,0,0,0,85,0,201,0,0,0,32,0,0,0,0,0,176,0,0,0,75,0,209,0);
signal scenario_full  : scenario_type := (119,31,133,31,31,31,246,31,38,31,117,31,76,31,94,31,64,31,19,31,19,30,180,31,92,31,183,31,176,31,147,31,154,31,121,31,247,31,221,31,185,31,152,31,152,30,255,31,228,31,228,30,202,31,75,31,157,31,157,30,17,31,17,30,60,31,60,30,76,31,100,31,224,31,95,31,201,31,98,31,85,31,85,30,245,31,184,31,11,31,33,31,51,31,51,30,51,29,165,31,53,31,64,31,64,30,64,29,210,31,74,31,41,31,142,31,162,31,201,31,201,30,208,31,208,30,82,31,156,31,181,31,216,31,216,30,240,31,38,31,162,31,162,30,174,31,150,31,108,31,108,30,166,31,60,31,197,31,5,31,167,31,250,31,199,31,53,31,198,31,75,31,237,31,64,31,65,31,219,31,55,31,114,31,114,30,114,29,172,31,32,31,193,31,35,31,53,31,117,31,92,31,17,31,179,31,179,30,220,31,222,31,228,31,228,30,42,31,11,31,202,31,202,30,223,31,218,31,102,31,74,31,74,30,3,31,117,31,26,31,26,30,25,31,25,30,18,31,28,31,28,30,14,31,232,31,249,31,108,31,108,30,108,29,236,31,50,31,50,30,184,31,155,31,120,31,180,31,211,31,211,30,211,29,211,28,149,31,76,31,83,31,248,31,74,31,74,30,74,29,250,31,250,30,125,31,125,30,177,31,244,31,212,31,238,31,189,31,99,31,99,30,99,29,99,28,164,31,254,31,110,31,122,31,141,31,68,31,91,31,91,30,91,29,91,28,14,31,14,30,3,31,3,30,3,29,136,31,133,31,221,31,221,30,56,31,120,31,120,30,120,29,120,28,138,31,138,30,120,31,76,31,76,30,92,31,253,31,191,31,188,31,188,30,50,31,221,31,107,31,57,31,149,31,91,31,243,31,243,30,243,29,59,31,180,31,180,30,15,31,7,31,7,30,225,31,210,31,227,31,185,31,178,31,178,30,178,29,178,28,168,31,101,31,101,30,101,29,101,28,101,27,101,26,174,31,212,31,115,31,247,31,133,31,133,30,248,31,44,31,201,31,55,31,233,31,112,31,24,31,148,31,231,31,221,31,221,30,214,31,55,31,55,30,113,31,72,31,72,30,223,31,231,31,119,31,119,30,111,31,111,30,152,31,152,30,151,31,72,31,76,31,236,31,244,31,12,31,94,31,28,31,135,31,135,30,250,31,33,31,7,31,177,31,86,31,141,31,71,31,116,31,10,31,98,31,216,31,69,31,69,30,69,29,50,31,82,31,82,30,168,31,196,31,196,30,126,31,126,30,49,31,124,31,163,31,114,31,69,31,41,31,56,31,79,31,216,31,255,31,190,31,16,31,72,31,72,30,111,31,176,31,4,31,6,31,6,30,7,31,7,30,182,31,65,31,86,31,252,31,69,31,114,31,221,31,128,31,148,31,83,31,2,31,2,30,108,31,79,31,185,31,156,31,78,31,208,31,153,31,5,31,243,31,243,30,64,31,11,31,108,31,108,30,108,29,142,31,104,31,86,31,156,31,116,31,155,31,114,31,188,31,8,31,249,31,74,31,41,31,34,31,196,31,198,31,244,31,232,31,232,30,232,29,245,31,245,30,244,31,144,31,136,31,224,31,151,31,210,31,252,31,123,31,123,30,54,31,54,31,242,31,44,31,37,31,66,31,33,31,34,31,65,31,221,31,199,31,175,31,43,31,175,31,187,31,187,30,33,31,122,31,224,31,82,31,191,31,197,31,142,31,142,30,144,31,16,31,185,31,165,31,64,31,64,30,170,31,114,31,126,31,56,31,31,31,200,31,87,31,87,30,91,31,30,31,4,31,194,31,77,31,221,31,165,31,165,30,253,31,198,31,120,31,243,31,104,31,189,31,40,31,200,31,103,31,141,31,141,30,80,31,220,31,6,31,68,31,207,31,125,31,153,31,142,31,181,31,7,31,193,31,193,30,188,31,188,30,78,31,41,31,162,31,49,31,133,31,133,30,122,31,122,30,247,31,124,31,122,31,219,31,18,31,18,30,180,31,251,31,89,31,222,31,149,31,139,31,92,31,139,31,139,30,33,31,76,31,237,31,238,31,44,31,95,31,27,31,27,30,63,31,63,30,116,31,116,30,116,29,193,31,90,31,90,30,221,31,221,30,220,31,246,31,108,31,145,31,188,31,143,31,21,31,30,31,252,31,143,31,251,31,104,31,143,31,119,31,90,31,90,30,90,29,45,31,243,31,88,31,88,30,33,31,219,31,219,30,222,31,93,31,93,30,86,31,161,31,161,30,20,31,138,31,47,31,47,30,199,31,231,31,50,31,52,31,52,30,52,29,104,31,104,30,22,31,107,31,107,30,240,31,139,31,139,30,45,31,121,31,176,31,11,31,11,30,11,29,30,31,30,30,124,31,177,31,240,31,240,30,6,31,38,31,38,30,53,31,53,30,175,31,248,31,187,31,234,31,236,31,102,31,42,31,42,30,42,29,226,31,215,31,32,31,117,31,217,31,251,31,47,31,131,31,223,31,127,31,46,31,65,31,96,31,130,31,168,31,168,30,203,31,31,31,132,31,132,30,137,31,13,31,159,31,114,31,189,31,49,31,203,31,185,31,250,31,255,31,111,31,111,30,59,31,11,31,53,31,39,31,39,30,64,31,217,31,29,31,84,31,109,31,56,31,56,30,157,31,106,31,239,31,34,31,12,31,96,31,96,30,158,31,49,31,49,30,238,31,128,31,195,31,195,30,71,31,71,30,71,29,190,31,190,30,158,31,158,30,141,31,104,31,150,31,200,31,200,30,225,31,225,30,40,31,128,31,102,31,105,31,245,31,102,31,190,31,249,31,249,30,214,31,176,31,203,31,64,31,66,31,252,31,93,31,12,31,98,31,62,31,183,31,175,31,213,31,227,31,186,31,201,31,247,31,247,30,203,31,91,31,91,30,91,29,91,28,85,31,201,31,201,30,32,31,32,30,32,29,176,31,176,30,75,31,209,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
