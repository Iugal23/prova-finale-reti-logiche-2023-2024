-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_432 is
end project_tb_432;

architecture project_tb_arch_432 of project_tb_432 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 350;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (160,0,255,0,156,0,53,0,251,0,0,0,125,0,104,0,60,0,89,0,0,0,232,0,218,0,242,0,0,0,68,0,0,0,36,0,141,0,189,0,50,0,69,0,165,0,65,0,6,0,143,0,81,0,4,0,219,0,238,0,37,0,109,0,225,0,0,0,0,0,0,0,230,0,243,0,0,0,59,0,110,0,237,0,173,0,5,0,54,0,43,0,124,0,16,0,169,0,231,0,223,0,0,0,119,0,16,0,251,0,103,0,121,0,176,0,243,0,0,0,8,0,101,0,33,0,43,0,34,0,225,0,192,0,54,0,80,0,203,0,164,0,169,0,188,0,73,0,83,0,126,0,183,0,79,0,46,0,0,0,44,0,0,0,96,0,19,0,0,0,111,0,125,0,0,0,2,0,41,0,0,0,42,0,19,0,129,0,168,0,33,0,129,0,243,0,13,0,246,0,102,0,43,0,0,0,129,0,119,0,236,0,18,0,1,0,205,0,75,0,61,0,15,0,247,0,202,0,55,0,0,0,210,0,61,0,0,0,164,0,77,0,0,0,142,0,237,0,0,0,186,0,125,0,0,0,89,0,229,0,69,0,51,0,134,0,0,0,121,0,76,0,4,0,206,0,73,0,19,0,112,0,0,0,148,0,219,0,28,0,194,0,113,0,0,0,10,0,0,0,50,0,188,0,0,0,156,0,109,0,179,0,107,0,198,0,187,0,44,0,0,0,195,0,217,0,214,0,0,0,45,0,133,0,0,0,31,0,0,0,60,0,24,0,222,0,75,0,173,0,0,0,118,0,116,0,0,0,231,0,195,0,195,0,176,0,3,0,83,0,0,0,117,0,33,0,0,0,26,0,36,0,32,0,164,0,73,0,50,0,173,0,143,0,132,0,140,0,226,0,72,0,151,0,0,0,226,0,210,0,0,0,250,0,0,0,0,0,32,0,230,0,0,0,89,0,0,0,0,0,131,0,0,0,159,0,206,0,201,0,0,0,88,0,229,0,0,0,231,0,23,0,152,0,0,0,54,0,0,0,0,0,42,0,0,0,70,0,123,0,233,0,79,0,230,0,206,0,229,0,125,0,159,0,0,0,32,0,233,0,0,0,221,0,242,0,2,0,5,0,0,0,229,0,0,0,187,0,239,0,201,0,0,0,86,0,198,0,0,0,143,0,85,0,112,0,87,0,0,0,224,0,227,0,59,0,74,0,150,0,160,0,0,0,87,0,30,0,172,0,0,0,128,0,223,0,118,0,28,0,114,0,103,0,234,0,6,0,194,0,44,0,75,0,0,0,26,0,221,0,165,0,175,0,0,0,128,0,86,0,0,0,179,0,237,0,0,0,0,0,111,0,198,0,0,0,7,0,154,0,2,0,0,0,24,0,103,0,193,0,69,0,64,0,209,0,0,0,225,0,227,0,171,0,119,0,199,0,168,0,203,0,0,0,0,0,147,0,233,0,27,0,227,0,0,0,48,0,0,0,56,0,160,0,184,0,78,0,114,0,149,0,240,0,180,0,0,0,0,0,176,0,0,0,109,0,85,0,0,0,4,0,24,0,139,0,148,0,162,0);
signal scenario_full  : scenario_type := (160,31,255,31,156,31,53,31,251,31,251,30,125,31,104,31,60,31,89,31,89,30,232,31,218,31,242,31,242,30,68,31,68,30,36,31,141,31,189,31,50,31,69,31,165,31,65,31,6,31,143,31,81,31,4,31,219,31,238,31,37,31,109,31,225,31,225,30,225,29,225,28,230,31,243,31,243,30,59,31,110,31,237,31,173,31,5,31,54,31,43,31,124,31,16,31,169,31,231,31,223,31,223,30,119,31,16,31,251,31,103,31,121,31,176,31,243,31,243,30,8,31,101,31,33,31,43,31,34,31,225,31,192,31,54,31,80,31,203,31,164,31,169,31,188,31,73,31,83,31,126,31,183,31,79,31,46,31,46,30,44,31,44,30,96,31,19,31,19,30,111,31,125,31,125,30,2,31,41,31,41,30,42,31,19,31,129,31,168,31,33,31,129,31,243,31,13,31,246,31,102,31,43,31,43,30,129,31,119,31,236,31,18,31,1,31,205,31,75,31,61,31,15,31,247,31,202,31,55,31,55,30,210,31,61,31,61,30,164,31,77,31,77,30,142,31,237,31,237,30,186,31,125,31,125,30,89,31,229,31,69,31,51,31,134,31,134,30,121,31,76,31,4,31,206,31,73,31,19,31,112,31,112,30,148,31,219,31,28,31,194,31,113,31,113,30,10,31,10,30,50,31,188,31,188,30,156,31,109,31,179,31,107,31,198,31,187,31,44,31,44,30,195,31,217,31,214,31,214,30,45,31,133,31,133,30,31,31,31,30,60,31,24,31,222,31,75,31,173,31,173,30,118,31,116,31,116,30,231,31,195,31,195,31,176,31,3,31,83,31,83,30,117,31,33,31,33,30,26,31,36,31,32,31,164,31,73,31,50,31,173,31,143,31,132,31,140,31,226,31,72,31,151,31,151,30,226,31,210,31,210,30,250,31,250,30,250,29,32,31,230,31,230,30,89,31,89,30,89,29,131,31,131,30,159,31,206,31,201,31,201,30,88,31,229,31,229,30,231,31,23,31,152,31,152,30,54,31,54,30,54,29,42,31,42,30,70,31,123,31,233,31,79,31,230,31,206,31,229,31,125,31,159,31,159,30,32,31,233,31,233,30,221,31,242,31,2,31,5,31,5,30,229,31,229,30,187,31,239,31,201,31,201,30,86,31,198,31,198,30,143,31,85,31,112,31,87,31,87,30,224,31,227,31,59,31,74,31,150,31,160,31,160,30,87,31,30,31,172,31,172,30,128,31,223,31,118,31,28,31,114,31,103,31,234,31,6,31,194,31,44,31,75,31,75,30,26,31,221,31,165,31,175,31,175,30,128,31,86,31,86,30,179,31,237,31,237,30,237,29,111,31,198,31,198,30,7,31,154,31,2,31,2,30,24,31,103,31,193,31,69,31,64,31,209,31,209,30,225,31,227,31,171,31,119,31,199,31,168,31,203,31,203,30,203,29,147,31,233,31,27,31,227,31,227,30,48,31,48,30,56,31,160,31,184,31,78,31,114,31,149,31,240,31,180,31,180,30,180,29,176,31,176,30,109,31,85,31,85,30,4,31,24,31,139,31,148,31,162,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
