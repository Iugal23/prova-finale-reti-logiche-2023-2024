-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 957;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (23,0,0,0,238,0,146,0,46,0,131,0,200,0,104,0,96,0,0,0,85,0,144,0,0,0,82,0,0,0,207,0,0,0,0,0,43,0,226,0,140,0,239,0,0,0,137,0,1,0,57,0,76,0,245,0,2,0,217,0,0,0,26,0,38,0,0,0,0,0,212,0,157,0,189,0,0,0,69,0,192,0,10,0,0,0,42,0,122,0,219,0,93,0,213,0,130,0,4,0,125,0,0,0,163,0,79,0,142,0,0,0,230,0,0,0,60,0,170,0,233,0,65,0,186,0,61,0,79,0,175,0,23,0,29,0,239,0,0,0,0,0,25,0,119,0,60,0,214,0,10,0,102,0,0,0,0,0,173,0,230,0,0,0,90,0,172,0,175,0,179,0,251,0,169,0,245,0,152,0,186,0,20,0,135,0,0,0,119,0,195,0,128,0,209,0,0,0,0,0,241,0,0,0,133,0,72,0,2,0,0,0,0,0,118,0,218,0,116,0,181,0,255,0,43,0,7,0,0,0,0,0,126,0,168,0,92,0,234,0,209,0,196,0,16,0,74,0,232,0,91,0,142,0,0,0,44,0,0,0,111,0,0,0,123,0,91,0,57,0,0,0,154,0,0,0,135,0,13,0,42,0,173,0,0,0,112,0,86,0,136,0,52,0,178,0,3,0,53,0,159,0,0,0,150,0,167,0,119,0,2,0,143,0,253,0,125,0,47,0,44,0,106,0,19,0,85,0,199,0,237,0,45,0,246,0,131,0,132,0,0,0,83,0,3,0,162,0,66,0,201,0,0,0,0,0,78,0,94,0,0,0,88,0,53,0,0,0,17,0,12,0,53,0,61,0,94,0,173,0,89,0,255,0,247,0,0,0,209,0,157,0,117,0,251,0,0,0,214,0,229,0,140,0,149,0,0,0,184,0,90,0,224,0,71,0,155,0,132,0,0,0,0,0,222,0,67,0,0,0,0,0,0,0,238,0,78,0,13,0,115,0,212,0,142,0,229,0,0,0,187,0,0,0,0,0,162,0,47,0,0,0,112,0,59,0,0,0,152,0,99,0,3,0,213,0,252,0,58,0,246,0,119,0,84,0,196,0,18,0,0,0,144,0,0,0,0,0,131,0,14,0,9,0,0,0,0,0,39,0,241,0,251,0,242,0,0,0,4,0,158,0,221,0,8,0,107,0,88,0,2,0,0,0,0,0,133,0,0,0,38,0,0,0,234,0,48,0,143,0,24,0,64,0,95,0,98,0,0,0,121,0,79,0,46,0,22,0,64,0,137,0,0,0,70,0,76,0,185,0,109,0,58,0,113,0,59,0,0,0,66,0,131,0,141,0,71,0,51,0,213,0,42,0,183,0,9,0,0,0,66,0,10,0,188,0,101,0,83,0,36,0,178,0,149,0,52,0,211,0,95,0,255,0,202,0,149,0,126,0,28,0,217,0,243,0,0,0,117,0,18,0,0,0,49,0,172,0,206,0,23,0,58,0,0,0,61,0,27,0,231,0,53,0,2,0,69,0,0,0,20,0,253,0,72,0,151,0,159,0,81,0,0,0,221,0,0,0,54,0,236,0,136,0,238,0,0,0,246,0,49,0,48,0,0,0,0,0,6,0,188,0,14,0,0,0,128,0,183,0,205,0,36,0,13,0,164,0,129,0,187,0,191,0,116,0,0,0,0,0,115,0,65,0,129,0,124,0,222,0,75,0,77,0,34,0,28,0,232,0,157,0,11,0,215,0,168,0,165,0,0,0,10,0,0,0,91,0,41,0,0,0,189,0,98,0,191,0,135,0,2,0,251,0,230,0,79,0,218,0,196,0,89,0,204,0,0,0,255,0,2,0,164,0,0,0,45,0,127,0,122,0,0,0,105,0,235,0,0,0,93,0,48,0,99,0,167,0,0,0,41,0,230,0,134,0,212,0,199,0,0,0,64,0,236,0,85,0,243,0,188,0,71,0,212,0,99,0,64,0,194,0,56,0,28,0,0,0,50,0,0,0,224,0,239,0,113,0,151,0,129,0,0,0,162,0,0,0,66,0,202,0,0,0,125,0,80,0,12,0,175,0,109,0,231,0,189,0,222,0,56,0,0,0,0,0,117,0,0,0,0,0,0,0,234,0,0,0,0,0,105,0,59,0,235,0,0,0,122,0,0,0,53,0,0,0,0,0,116,0,106,0,0,0,215,0,0,0,157,0,63,0,0,0,61,0,147,0,44,0,200,0,244,0,0,0,35,0,140,0,0,0,0,0,13,0,101,0,64,0,34,0,169,0,68,0,164,0,189,0,62,0,37,0,248,0,222,0,149,0,0,0,116,0,114,0,0,0,0,0,41,0,157,0,220,0,65,0,82,0,222,0,166,0,149,0,17,0,0,0,200,0,147,0,0,0,249,0,106,0,0,0,174,0,0,0,61,0,248,0,40,0,254,0,0,0,72,0,13,0,141,0,4,0,104,0,169,0,204,0,224,0,177,0,16,0,207,0,102,0,45,0,19,0,180,0,0,0,0,0,25,0,250,0,138,0,0,0,66,0,94,0,0,0,0,0,241,0,0,0,16,0,24,0,154,0,2,0,70,0,138,0,123,0,214,0,166,0,130,0,88,0,181,0,153,0,118,0,175,0,63,0,0,0,252,0,123,0,166,0,0,0,0,0,85,0,144,0,79,0,0,0,0,0,26,0,0,0,0,0,73,0,120,0,217,0,45,0,0,0,89,0,107,0,0,0,65,0,0,0,160,0,73,0,200,0,47,0,149,0,181,0,1,0,70,0,0,0,5,0,0,0,0,0,245,0,101,0,53,0,26,0,197,0,128,0,0,0,148,0,190,0,201,0,0,0,70,0,108,0,0,0,46,0,0,0,204,0,180,0,94,0,0,0,140,0,0,0,2,0,55,0,77,0,0,0,44,0,3,0,125,0,90,0,0,0,87,0,170,0,0,0,18,0,0,0,95,0,77,0,124,0,203,0,3,0,186,0,0,0,177,0,143,0,71,0,127,0,0,0,132,0,232,0,253,0,149,0,194,0,171,0,85,0,160,0,251,0,150,0,141,0,91,0,53,0,30,0,0,0,132,0,194,0,114,0,24,0,74,0,75,0,139,0,189,0,255,0,0,0,47,0,154,0,125,0,147,0,237,0,60,0,110,0,21,0,151,0,0,0,107,0,172,0,69,0,224,0,185,0,13,0,175,0,175,0,121,0,102,0,244,0,211,0,0,0,90,0,21,0,0,0,56,0,187,0,164,0,161,0,53,0,135,0,0,0,0,0,86,0,170,0,26,0,0,0,6,0,240,0,226,0,190,0,80,0,0,0,96,0,244,0,234,0,0,0,94,0,0,0,170,0,0,0,73,0,115,0,111,0,101,0,186,0,0,0,161,0,122,0,85,0,237,0,173,0,250,0,82,0,62,0,76,0,0,0,0,0,0,0,249,0,0,0,46,0,0,0,6,0,0,0,81,0,116,0,113,0,0,0,0,0,131,0,64,0,91,0,194,0,124,0,0,0,220,0,236,0,247,0,253,0,79,0,130,0,66,0,220,0,253,0,0,0,77,0,0,0,0,0,116,0,240,0,194,0,114,0,57,0,0,0,28,0,3,0,82,0,135,0,231,0,213,0,0,0,0,0,0,0,5,0,136,0,0,0,186,0,237,0,203,0,108,0,0,0,97,0,42,0,132,0,202,0,229,0,10,0,109,0,0,0,182,0,110,0,56,0,118,0,215,0,214,0,96,0,65,0,233,0,139,0,0,0,130,0,144,0,137,0,7,0,157,0,5,0,32,0,89,0,86,0,0,0,13,0,177,0,8,0,0,0,61,0,183,0,0,0,157,0,0,0,89,0,9,0,196,0,115,0,32,0,49,0,0,0,158,0,4,0,228,0,0,0,0,0,169,0,235,0,0,0,0,0,0,0,0,0,0,0,59,0,148,0,148,0,165,0,64,0,152,0,0,0,0,0,232,0,182,0,0,0,46,0,2,0,32,0,47,0,209,0,93,0,0,0,0,0,121,0,188,0,249,0,131,0,142,0,77,0,0,0,214,0,122,0,6,0,23,0,42,0,160,0,220,0,87,0,39,0,253,0,229,0,170,0,6,0,69,0,157,0,107,0,65,0,214,0,124,0,61,0,172,0,0,0,0,0,174,0,0,0,0,0,0,0,77,0,180,0,0,0,192,0,164,0,210,0,114,0,250,0,158,0,0,0,38,0,91,0,0,0,235,0,20,0,177,0,59,0,202,0,171,0,115,0,0,0,157,0,36,0,213,0,48,0,142,0,0,0,233,0,0,0);
signal scenario_full  : scenario_type := (23,31,23,30,238,31,146,31,46,31,131,31,200,31,104,31,96,31,96,30,85,31,144,31,144,30,82,31,82,30,207,31,207,30,207,29,43,31,226,31,140,31,239,31,239,30,137,31,1,31,57,31,76,31,245,31,2,31,217,31,217,30,26,31,38,31,38,30,38,29,212,31,157,31,189,31,189,30,69,31,192,31,10,31,10,30,42,31,122,31,219,31,93,31,213,31,130,31,4,31,125,31,125,30,163,31,79,31,142,31,142,30,230,31,230,30,60,31,170,31,233,31,65,31,186,31,61,31,79,31,175,31,23,31,29,31,239,31,239,30,239,29,25,31,119,31,60,31,214,31,10,31,102,31,102,30,102,29,173,31,230,31,230,30,90,31,172,31,175,31,179,31,251,31,169,31,245,31,152,31,186,31,20,31,135,31,135,30,119,31,195,31,128,31,209,31,209,30,209,29,241,31,241,30,133,31,72,31,2,31,2,30,2,29,118,31,218,31,116,31,181,31,255,31,43,31,7,31,7,30,7,29,126,31,168,31,92,31,234,31,209,31,196,31,16,31,74,31,232,31,91,31,142,31,142,30,44,31,44,30,111,31,111,30,123,31,91,31,57,31,57,30,154,31,154,30,135,31,13,31,42,31,173,31,173,30,112,31,86,31,136,31,52,31,178,31,3,31,53,31,159,31,159,30,150,31,167,31,119,31,2,31,143,31,253,31,125,31,47,31,44,31,106,31,19,31,85,31,199,31,237,31,45,31,246,31,131,31,132,31,132,30,83,31,3,31,162,31,66,31,201,31,201,30,201,29,78,31,94,31,94,30,88,31,53,31,53,30,17,31,12,31,53,31,61,31,94,31,173,31,89,31,255,31,247,31,247,30,209,31,157,31,117,31,251,31,251,30,214,31,229,31,140,31,149,31,149,30,184,31,90,31,224,31,71,31,155,31,132,31,132,30,132,29,222,31,67,31,67,30,67,29,67,28,238,31,78,31,13,31,115,31,212,31,142,31,229,31,229,30,187,31,187,30,187,29,162,31,47,31,47,30,112,31,59,31,59,30,152,31,99,31,3,31,213,31,252,31,58,31,246,31,119,31,84,31,196,31,18,31,18,30,144,31,144,30,144,29,131,31,14,31,9,31,9,30,9,29,39,31,241,31,251,31,242,31,242,30,4,31,158,31,221,31,8,31,107,31,88,31,2,31,2,30,2,29,133,31,133,30,38,31,38,30,234,31,48,31,143,31,24,31,64,31,95,31,98,31,98,30,121,31,79,31,46,31,22,31,64,31,137,31,137,30,70,31,76,31,185,31,109,31,58,31,113,31,59,31,59,30,66,31,131,31,141,31,71,31,51,31,213,31,42,31,183,31,9,31,9,30,66,31,10,31,188,31,101,31,83,31,36,31,178,31,149,31,52,31,211,31,95,31,255,31,202,31,149,31,126,31,28,31,217,31,243,31,243,30,117,31,18,31,18,30,49,31,172,31,206,31,23,31,58,31,58,30,61,31,27,31,231,31,53,31,2,31,69,31,69,30,20,31,253,31,72,31,151,31,159,31,81,31,81,30,221,31,221,30,54,31,236,31,136,31,238,31,238,30,246,31,49,31,48,31,48,30,48,29,6,31,188,31,14,31,14,30,128,31,183,31,205,31,36,31,13,31,164,31,129,31,187,31,191,31,116,31,116,30,116,29,115,31,65,31,129,31,124,31,222,31,75,31,77,31,34,31,28,31,232,31,157,31,11,31,215,31,168,31,165,31,165,30,10,31,10,30,91,31,41,31,41,30,189,31,98,31,191,31,135,31,2,31,251,31,230,31,79,31,218,31,196,31,89,31,204,31,204,30,255,31,2,31,164,31,164,30,45,31,127,31,122,31,122,30,105,31,235,31,235,30,93,31,48,31,99,31,167,31,167,30,41,31,230,31,134,31,212,31,199,31,199,30,64,31,236,31,85,31,243,31,188,31,71,31,212,31,99,31,64,31,194,31,56,31,28,31,28,30,50,31,50,30,224,31,239,31,113,31,151,31,129,31,129,30,162,31,162,30,66,31,202,31,202,30,125,31,80,31,12,31,175,31,109,31,231,31,189,31,222,31,56,31,56,30,56,29,117,31,117,30,117,29,117,28,234,31,234,30,234,29,105,31,59,31,235,31,235,30,122,31,122,30,53,31,53,30,53,29,116,31,106,31,106,30,215,31,215,30,157,31,63,31,63,30,61,31,147,31,44,31,200,31,244,31,244,30,35,31,140,31,140,30,140,29,13,31,101,31,64,31,34,31,169,31,68,31,164,31,189,31,62,31,37,31,248,31,222,31,149,31,149,30,116,31,114,31,114,30,114,29,41,31,157,31,220,31,65,31,82,31,222,31,166,31,149,31,17,31,17,30,200,31,147,31,147,30,249,31,106,31,106,30,174,31,174,30,61,31,248,31,40,31,254,31,254,30,72,31,13,31,141,31,4,31,104,31,169,31,204,31,224,31,177,31,16,31,207,31,102,31,45,31,19,31,180,31,180,30,180,29,25,31,250,31,138,31,138,30,66,31,94,31,94,30,94,29,241,31,241,30,16,31,24,31,154,31,2,31,70,31,138,31,123,31,214,31,166,31,130,31,88,31,181,31,153,31,118,31,175,31,63,31,63,30,252,31,123,31,166,31,166,30,166,29,85,31,144,31,79,31,79,30,79,29,26,31,26,30,26,29,73,31,120,31,217,31,45,31,45,30,89,31,107,31,107,30,65,31,65,30,160,31,73,31,200,31,47,31,149,31,181,31,1,31,70,31,70,30,5,31,5,30,5,29,245,31,101,31,53,31,26,31,197,31,128,31,128,30,148,31,190,31,201,31,201,30,70,31,108,31,108,30,46,31,46,30,204,31,180,31,94,31,94,30,140,31,140,30,2,31,55,31,77,31,77,30,44,31,3,31,125,31,90,31,90,30,87,31,170,31,170,30,18,31,18,30,95,31,77,31,124,31,203,31,3,31,186,31,186,30,177,31,143,31,71,31,127,31,127,30,132,31,232,31,253,31,149,31,194,31,171,31,85,31,160,31,251,31,150,31,141,31,91,31,53,31,30,31,30,30,132,31,194,31,114,31,24,31,74,31,75,31,139,31,189,31,255,31,255,30,47,31,154,31,125,31,147,31,237,31,60,31,110,31,21,31,151,31,151,30,107,31,172,31,69,31,224,31,185,31,13,31,175,31,175,31,121,31,102,31,244,31,211,31,211,30,90,31,21,31,21,30,56,31,187,31,164,31,161,31,53,31,135,31,135,30,135,29,86,31,170,31,26,31,26,30,6,31,240,31,226,31,190,31,80,31,80,30,96,31,244,31,234,31,234,30,94,31,94,30,170,31,170,30,73,31,115,31,111,31,101,31,186,31,186,30,161,31,122,31,85,31,237,31,173,31,250,31,82,31,62,31,76,31,76,30,76,29,76,28,249,31,249,30,46,31,46,30,6,31,6,30,81,31,116,31,113,31,113,30,113,29,131,31,64,31,91,31,194,31,124,31,124,30,220,31,236,31,247,31,253,31,79,31,130,31,66,31,220,31,253,31,253,30,77,31,77,30,77,29,116,31,240,31,194,31,114,31,57,31,57,30,28,31,3,31,82,31,135,31,231,31,213,31,213,30,213,29,213,28,5,31,136,31,136,30,186,31,237,31,203,31,108,31,108,30,97,31,42,31,132,31,202,31,229,31,10,31,109,31,109,30,182,31,110,31,56,31,118,31,215,31,214,31,96,31,65,31,233,31,139,31,139,30,130,31,144,31,137,31,7,31,157,31,5,31,32,31,89,31,86,31,86,30,13,31,177,31,8,31,8,30,61,31,183,31,183,30,157,31,157,30,89,31,9,31,196,31,115,31,32,31,49,31,49,30,158,31,4,31,228,31,228,30,228,29,169,31,235,31,235,30,235,29,235,28,235,27,235,26,59,31,148,31,148,31,165,31,64,31,152,31,152,30,152,29,232,31,182,31,182,30,46,31,2,31,32,31,47,31,209,31,93,31,93,30,93,29,121,31,188,31,249,31,131,31,142,31,77,31,77,30,214,31,122,31,6,31,23,31,42,31,160,31,220,31,87,31,39,31,253,31,229,31,170,31,6,31,69,31,157,31,107,31,65,31,214,31,124,31,61,31,172,31,172,30,172,29,174,31,174,30,174,29,174,28,77,31,180,31,180,30,192,31,164,31,210,31,114,31,250,31,158,31,158,30,38,31,91,31,91,30,235,31,20,31,177,31,59,31,202,31,171,31,115,31,115,30,157,31,36,31,213,31,48,31,142,31,142,30,233,31,233,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
