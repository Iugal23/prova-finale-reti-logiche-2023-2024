-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_721 is
end project_tb_721;

architecture project_tb_arch_721 of project_tb_721 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 185;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (251,0,0,0,15,0,10,0,152,0,200,0,129,0,15,0,243,0,1,0,134,0,78,0,0,0,195,0,223,0,72,0,185,0,215,0,155,0,158,0,39,0,63,0,0,0,43,0,0,0,173,0,111,0,60,0,41,0,150,0,223,0,138,0,47,0,1,0,41,0,228,0,87,0,248,0,98,0,0,0,222,0,0,0,227,0,76,0,119,0,174,0,125,0,0,0,0,0,251,0,130,0,181,0,0,0,224,0,33,0,160,0,191,0,90,0,190,0,145,0,0,0,108,0,0,0,37,0,126,0,75,0,247,0,178,0,112,0,12,0,20,0,119,0,201,0,3,0,103,0,47,0,0,0,83,0,0,0,129,0,253,0,63,0,73,0,206,0,134,0,16,0,16,0,45,0,47,0,28,0,0,0,67,0,116,0,127,0,255,0,169,0,56,0,121,0,0,0,0,0,0,0,178,0,0,0,136,0,114,0,201,0,143,0,0,0,113,0,0,0,0,0,41,0,2,0,127,0,252,0,250,0,0,0,0,0,203,0,0,0,59,0,98,0,0,0,13,0,135,0,0,0,9,0,0,0,38,0,110,0,90,0,94,0,63,0,66,0,125,0,92,0,0,0,0,0,0,0,126,0,47,0,181,0,0,0,128,0,156,0,187,0,159,0,73,0,13,0,79,0,6,0,168,0,149,0,0,0,142,0,72,0,101,0,78,0,0,0,60,0,134,0,121,0,114,0,215,0,0,0,16,0,150,0,25,0,96,0,110,0,197,0,0,0,157,0,100,0,126,0,111,0,0,0,72,0,3,0,166,0,215,0,0,0,0,0,0,0,148,0);
signal scenario_full  : scenario_type := (251,31,251,30,15,31,10,31,152,31,200,31,129,31,15,31,243,31,1,31,134,31,78,31,78,30,195,31,223,31,72,31,185,31,215,31,155,31,158,31,39,31,63,31,63,30,43,31,43,30,173,31,111,31,60,31,41,31,150,31,223,31,138,31,47,31,1,31,41,31,228,31,87,31,248,31,98,31,98,30,222,31,222,30,227,31,76,31,119,31,174,31,125,31,125,30,125,29,251,31,130,31,181,31,181,30,224,31,33,31,160,31,191,31,90,31,190,31,145,31,145,30,108,31,108,30,37,31,126,31,75,31,247,31,178,31,112,31,12,31,20,31,119,31,201,31,3,31,103,31,47,31,47,30,83,31,83,30,129,31,253,31,63,31,73,31,206,31,134,31,16,31,16,31,45,31,47,31,28,31,28,30,67,31,116,31,127,31,255,31,169,31,56,31,121,31,121,30,121,29,121,28,178,31,178,30,136,31,114,31,201,31,143,31,143,30,113,31,113,30,113,29,41,31,2,31,127,31,252,31,250,31,250,30,250,29,203,31,203,30,59,31,98,31,98,30,13,31,135,31,135,30,9,31,9,30,38,31,110,31,90,31,94,31,63,31,66,31,125,31,92,31,92,30,92,29,92,28,126,31,47,31,181,31,181,30,128,31,156,31,187,31,159,31,73,31,13,31,79,31,6,31,168,31,149,31,149,30,142,31,72,31,101,31,78,31,78,30,60,31,134,31,121,31,114,31,215,31,215,30,16,31,150,31,25,31,96,31,110,31,197,31,197,30,157,31,100,31,126,31,111,31,111,30,72,31,3,31,166,31,215,31,215,30,215,29,215,28,148,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
