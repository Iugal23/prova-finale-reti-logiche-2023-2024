-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 753;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (74,0,247,0,106,0,28,0,165,0,253,0,116,0,0,0,0,0,217,0,48,0,164,0,243,0,131,0,0,0,76,0,135,0,98,0,136,0,118,0,52,0,173,0,31,0,2,0,53,0,136,0,4,0,136,0,62,0,107,0,38,0,93,0,0,0,152,0,0,0,243,0,88,0,112,0,125,0,54,0,14,0,165,0,214,0,63,0,5,0,8,0,248,0,114,0,141,0,31,0,51,0,184,0,19,0,30,0,213,0,0,0,236,0,0,0,28,0,136,0,30,0,246,0,38,0,214,0,235,0,68,0,191,0,155,0,121,0,0,0,243,0,85,0,209,0,187,0,0,0,109,0,21,0,90,0,0,0,25,0,10,0,0,0,127,0,176,0,125,0,179,0,199,0,235,0,179,0,0,0,254,0,164,0,185,0,0,0,92,0,0,0,86,0,137,0,209,0,37,0,189,0,213,0,91,0,192,0,78,0,113,0,182,0,136,0,35,0,0,0,152,0,67,0,7,0,78,0,84,0,117,0,211,0,184,0,0,0,169,0,207,0,220,0,0,0,48,0,188,0,0,0,122,0,171,0,239,0,0,0,0,0,0,0,0,0,224,0,110,0,113,0,48,0,138,0,144,0,0,0,0,0,58,0,66,0,0,0,0,0,44,0,0,0,103,0,20,0,174,0,95,0,0,0,185,0,140,0,108,0,152,0,0,0,117,0,189,0,124,0,207,0,118,0,211,0,214,0,69,0,122,0,88,0,0,0,0,0,0,0,69,0,0,0,255,0,204,0,179,0,68,0,216,0,0,0,63,0,99,0,101,0,61,0,72,0,240,0,174,0,249,0,83,0,74,0,105,0,198,0,254,0,227,0,219,0,15,0,0,0,0,0,236,0,192,0,177,0,0,0,50,0,0,0,228,0,23,0,241,0,80,0,54,0,0,0,0,0,7,0,0,0,155,0,23,0,227,0,176,0,188,0,113,0,122,0,204,0,44,0,0,0,184,0,23,0,64,0,0,0,63,0,122,0,76,0,124,0,1,0,81,0,38,0,0,0,0,0,237,0,71,0,0,0,115,0,63,0,3,0,174,0,132,0,98,0,66,0,86,0,0,0,84,0,27,0,6,0,81,0,0,0,46,0,233,0,231,0,0,0,86,0,57,0,0,0,239,0,88,0,26,0,21,0,79,0,108,0,0,0,0,0,148,0,2,0,0,0,116,0,238,0,220,0,192,0,20,0,131,0,14,0,87,0,227,0,19,0,21,0,187,0,146,0,223,0,162,0,83,0,120,0,61,0,63,0,202,0,50,0,0,0,51,0,172,0,55,0,0,0,163,0,50,0,114,0,99,0,52,0,140,0,251,0,235,0,21,0,41,0,69,0,202,0,42,0,42,0,240,0,213,0,0,0,2,0,200,0,109,0,53,0,33,0,205,0,124,0,0,0,75,0,104,0,0,0,137,0,16,0,18,0,165,0,186,0,0,0,148,0,200,0,0,0,131,0,225,0,0,0,7,0,0,0,0,0,0,0,0,0,155,0,96,0,137,0,54,0,146,0,195,0,0,0,0,0,24,0,62,0,7,0,184,0,166,0,158,0,13,0,124,0,103,0,56,0,199,0,149,0,38,0,55,0,31,0,55,0,0,0,236,0,86,0,148,0,52,0,180,0,72,0,6,0,92,0,136,0,0,0,207,0,150,0,0,0,239,0,24,0,35,0,215,0,86,0,199,0,25,0,46,0,168,0,0,0,96,0,164,0,0,0,196,0,115,0,116,0,126,0,107,0,174,0,0,0,0,0,18,0,107,0,0,0,88,0,0,0,147,0,12,0,239,0,0,0,30,0,136,0,109,0,0,0,63,0,164,0,33,0,254,0,113,0,140,0,237,0,191,0,234,0,151,0,0,0,104,0,118,0,0,0,154,0,0,0,230,0,18,0,69,0,124,0,53,0,236,0,249,0,0,0,232,0,93,0,34,0,134,0,114,0,0,0,0,0,72,0,75,0,0,0,217,0,160,0,38,0,29,0,125,0,131,0,112,0,196,0,62,0,142,0,0,0,6,0,27,0,86,0,129,0,0,0,10,0,205,0,0,0,51,0,12,0,7,0,212,0,162,0,119,0,22,0,49,0,164,0,172,0,0,0,194,0,181,0,65,0,38,0,249,0,46,0,172,0,222,0,140,0,192,0,219,0,71,0,87,0,0,0,225,0,86,0,242,0,128,0,122,0,197,0,64,0,101,0,235,0,2,0,191,0,0,0,225,0,80,0,59,0,135,0,107,0,214,0,246,0,131,0,213,0,147,0,0,0,210,0,150,0,228,0,121,0,115,0,118,0,86,0,0,0,66,0,241,0,200,0,87,0,18,0,81,0,44,0,158,0,14,0,131,0,132,0,0,0,177,0,125,0,88,0,128,0,243,0,148,0,143,0,0,0,47,0,0,0,92,0,26,0,212,0,0,0,159,0,0,0,0,0,239,0,66,0,35,0,244,0,13,0,32,0,104,0,68,0,106,0,219,0,0,0,0,0,170,0,0,0,0,0,29,0,0,0,92,0,76,0,11,0,55,0,42,0,0,0,144,0,200,0,245,0,0,0,82,0,185,0,0,0,56,0,8,0,154,0,235,0,0,0,145,0,184,0,60,0,181,0,148,0,0,0,244,0,125,0,236,0,59,0,184,0,227,0,39,0,0,0,44,0,0,0,160,0,211,0,0,0,202,0,0,0,155,0,93,0,0,0,92,0,161,0,90,0,197,0,7,0,72,0,161,0,0,0,0,0,141,0,153,0,128,0,36,0,0,0,0,0,105,0,0,0,11,0,252,0,53,0,82,0,73,0,217,0,64,0,151,0,47,0,242,0,111,0,36,0,222,0,61,0,17,0,68,0,110,0,80,0,183,0,139,0,227,0,125,0,179,0,42,0,14,0,0,0,0,0,156,0,0,0,91,0,52,0,200,0,187,0,202,0,69,0,44,0,0,0,76,0,188,0,120,0,229,0,148,0,82,0,185,0,118,0,127,0,68,0,157,0,0,0,75,0,0,0,0,0,0,0,0,0,128,0,23,0,0,0,62,0,18,0,56,0,0,0,116,0,39,0,101,0,176,0,147,0,0,0,79,0,229,0,0,0,247,0,223,0,8,0,0,0,161,0,175,0,229,0,224,0,253,0,197,0,39,0,0,0,109,0,0,0,51,0,159,0,98,0,76,0,13,0,45,0,0,0,19,0,0,0,116,0,187,0,57,0,0,0,68,0,133,0,0,0,0,0,165,0,176,0,151,0,11,0,0,0,37,0,59,0,143,0,10,0,49,0,162,0,67,0,68,0,137,0,2,0,231,0,90,0,3,0,109,0,172,0,146,0,51,0,137,0,63,0,0,0,39,0);
signal scenario_full  : scenario_type := (74,31,247,31,106,31,28,31,165,31,253,31,116,31,116,30,116,29,217,31,48,31,164,31,243,31,131,31,131,30,76,31,135,31,98,31,136,31,118,31,52,31,173,31,31,31,2,31,53,31,136,31,4,31,136,31,62,31,107,31,38,31,93,31,93,30,152,31,152,30,243,31,88,31,112,31,125,31,54,31,14,31,165,31,214,31,63,31,5,31,8,31,248,31,114,31,141,31,31,31,51,31,184,31,19,31,30,31,213,31,213,30,236,31,236,30,28,31,136,31,30,31,246,31,38,31,214,31,235,31,68,31,191,31,155,31,121,31,121,30,243,31,85,31,209,31,187,31,187,30,109,31,21,31,90,31,90,30,25,31,10,31,10,30,127,31,176,31,125,31,179,31,199,31,235,31,179,31,179,30,254,31,164,31,185,31,185,30,92,31,92,30,86,31,137,31,209,31,37,31,189,31,213,31,91,31,192,31,78,31,113,31,182,31,136,31,35,31,35,30,152,31,67,31,7,31,78,31,84,31,117,31,211,31,184,31,184,30,169,31,207,31,220,31,220,30,48,31,188,31,188,30,122,31,171,31,239,31,239,30,239,29,239,28,239,27,224,31,110,31,113,31,48,31,138,31,144,31,144,30,144,29,58,31,66,31,66,30,66,29,44,31,44,30,103,31,20,31,174,31,95,31,95,30,185,31,140,31,108,31,152,31,152,30,117,31,189,31,124,31,207,31,118,31,211,31,214,31,69,31,122,31,88,31,88,30,88,29,88,28,69,31,69,30,255,31,204,31,179,31,68,31,216,31,216,30,63,31,99,31,101,31,61,31,72,31,240,31,174,31,249,31,83,31,74,31,105,31,198,31,254,31,227,31,219,31,15,31,15,30,15,29,236,31,192,31,177,31,177,30,50,31,50,30,228,31,23,31,241,31,80,31,54,31,54,30,54,29,7,31,7,30,155,31,23,31,227,31,176,31,188,31,113,31,122,31,204,31,44,31,44,30,184,31,23,31,64,31,64,30,63,31,122,31,76,31,124,31,1,31,81,31,38,31,38,30,38,29,237,31,71,31,71,30,115,31,63,31,3,31,174,31,132,31,98,31,66,31,86,31,86,30,84,31,27,31,6,31,81,31,81,30,46,31,233,31,231,31,231,30,86,31,57,31,57,30,239,31,88,31,26,31,21,31,79,31,108,31,108,30,108,29,148,31,2,31,2,30,116,31,238,31,220,31,192,31,20,31,131,31,14,31,87,31,227,31,19,31,21,31,187,31,146,31,223,31,162,31,83,31,120,31,61,31,63,31,202,31,50,31,50,30,51,31,172,31,55,31,55,30,163,31,50,31,114,31,99,31,52,31,140,31,251,31,235,31,21,31,41,31,69,31,202,31,42,31,42,31,240,31,213,31,213,30,2,31,200,31,109,31,53,31,33,31,205,31,124,31,124,30,75,31,104,31,104,30,137,31,16,31,18,31,165,31,186,31,186,30,148,31,200,31,200,30,131,31,225,31,225,30,7,31,7,30,7,29,7,28,7,27,155,31,96,31,137,31,54,31,146,31,195,31,195,30,195,29,24,31,62,31,7,31,184,31,166,31,158,31,13,31,124,31,103,31,56,31,199,31,149,31,38,31,55,31,31,31,55,31,55,30,236,31,86,31,148,31,52,31,180,31,72,31,6,31,92,31,136,31,136,30,207,31,150,31,150,30,239,31,24,31,35,31,215,31,86,31,199,31,25,31,46,31,168,31,168,30,96,31,164,31,164,30,196,31,115,31,116,31,126,31,107,31,174,31,174,30,174,29,18,31,107,31,107,30,88,31,88,30,147,31,12,31,239,31,239,30,30,31,136,31,109,31,109,30,63,31,164,31,33,31,254,31,113,31,140,31,237,31,191,31,234,31,151,31,151,30,104,31,118,31,118,30,154,31,154,30,230,31,18,31,69,31,124,31,53,31,236,31,249,31,249,30,232,31,93,31,34,31,134,31,114,31,114,30,114,29,72,31,75,31,75,30,217,31,160,31,38,31,29,31,125,31,131,31,112,31,196,31,62,31,142,31,142,30,6,31,27,31,86,31,129,31,129,30,10,31,205,31,205,30,51,31,12,31,7,31,212,31,162,31,119,31,22,31,49,31,164,31,172,31,172,30,194,31,181,31,65,31,38,31,249,31,46,31,172,31,222,31,140,31,192,31,219,31,71,31,87,31,87,30,225,31,86,31,242,31,128,31,122,31,197,31,64,31,101,31,235,31,2,31,191,31,191,30,225,31,80,31,59,31,135,31,107,31,214,31,246,31,131,31,213,31,147,31,147,30,210,31,150,31,228,31,121,31,115,31,118,31,86,31,86,30,66,31,241,31,200,31,87,31,18,31,81,31,44,31,158,31,14,31,131,31,132,31,132,30,177,31,125,31,88,31,128,31,243,31,148,31,143,31,143,30,47,31,47,30,92,31,26,31,212,31,212,30,159,31,159,30,159,29,239,31,66,31,35,31,244,31,13,31,32,31,104,31,68,31,106,31,219,31,219,30,219,29,170,31,170,30,170,29,29,31,29,30,92,31,76,31,11,31,55,31,42,31,42,30,144,31,200,31,245,31,245,30,82,31,185,31,185,30,56,31,8,31,154,31,235,31,235,30,145,31,184,31,60,31,181,31,148,31,148,30,244,31,125,31,236,31,59,31,184,31,227,31,39,31,39,30,44,31,44,30,160,31,211,31,211,30,202,31,202,30,155,31,93,31,93,30,92,31,161,31,90,31,197,31,7,31,72,31,161,31,161,30,161,29,141,31,153,31,128,31,36,31,36,30,36,29,105,31,105,30,11,31,252,31,53,31,82,31,73,31,217,31,64,31,151,31,47,31,242,31,111,31,36,31,222,31,61,31,17,31,68,31,110,31,80,31,183,31,139,31,227,31,125,31,179,31,42,31,14,31,14,30,14,29,156,31,156,30,91,31,52,31,200,31,187,31,202,31,69,31,44,31,44,30,76,31,188,31,120,31,229,31,148,31,82,31,185,31,118,31,127,31,68,31,157,31,157,30,75,31,75,30,75,29,75,28,75,27,128,31,23,31,23,30,62,31,18,31,56,31,56,30,116,31,39,31,101,31,176,31,147,31,147,30,79,31,229,31,229,30,247,31,223,31,8,31,8,30,161,31,175,31,229,31,224,31,253,31,197,31,39,31,39,30,109,31,109,30,51,31,159,31,98,31,76,31,13,31,45,31,45,30,19,31,19,30,116,31,187,31,57,31,57,30,68,31,133,31,133,30,133,29,165,31,176,31,151,31,11,31,11,30,37,31,59,31,143,31,10,31,49,31,162,31,67,31,68,31,137,31,2,31,231,31,90,31,3,31,109,31,172,31,146,31,51,31,137,31,63,31,63,30,39,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
