-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_672 is
end project_tb_672;

architecture project_tb_arch_672 of project_tb_672 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 647;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (15,0,13,0,166,0,69,0,125,0,164,0,122,0,215,0,110,0,223,0,0,0,124,0,238,0,37,0,0,0,50,0,23,0,102,0,244,0,94,0,198,0,0,0,105,0,208,0,0,0,223,0,0,0,170,0,126,0,25,0,130,0,4,0,103,0,0,0,234,0,201,0,0,0,21,0,134,0,39,0,1,0,186,0,193,0,179,0,27,0,225,0,54,0,108,0,151,0,0,0,84,0,52,0,81,0,46,0,47,0,0,0,149,0,245,0,0,0,189,0,0,0,58,0,206,0,8,0,28,0,247,0,180,0,101,0,208,0,70,0,105,0,0,0,38,0,75,0,189,0,130,0,0,0,90,0,0,0,86,0,129,0,178,0,157,0,193,0,175,0,221,0,33,0,0,0,231,0,113,0,0,0,236,0,223,0,104,0,104,0,0,0,12,0,210,0,172,0,26,0,203,0,11,0,101,0,0,0,104,0,66,0,29,0,0,0,86,0,77,0,42,0,29,0,224,0,195,0,109,0,248,0,195,0,228,0,0,0,221,0,154,0,128,0,11,0,67,0,247,0,71,0,0,0,63,0,168,0,24,0,171,0,157,0,249,0,110,0,181,0,0,0,126,0,0,0,0,0,240,0,89,0,0,0,233,0,51,0,189,0,118,0,55,0,213,0,0,0,37,0,84,0,113,0,130,0,250,0,243,0,77,0,22,0,196,0,92,0,11,0,0,0,41,0,71,0,0,0,0,0,10,0,165,0,78,0,9,0,253,0,0,0,0,0,94,0,116,0,108,0,182,0,0,0,0,0,248,0,0,0,203,0,0,0,44,0,53,0,246,0,81,0,74,0,242,0,198,0,227,0,27,0,243,0,0,0,0,0,117,0,205,0,119,0,40,0,96,0,60,0,212,0,98,0,19,0,58,0,0,0,135,0,0,0,108,0,143,0,242,0,227,0,47,0,158,0,81,0,252,0,84,0,234,0,94,0,158,0,0,0,0,0,45,0,82,0,247,0,207,0,0,0,245,0,89,0,0,0,5,0,0,0,87,0,221,0,255,0,171,0,0,0,131,0,247,0,43,0,0,0,2,0,92,0,23,0,255,0,0,0,23,0,0,0,0,0,0,0,228,0,109,0,232,0,6,0,19,0,26,0,156,0,0,0,228,0,19,0,0,0,95,0,79,0,38,0,189,0,107,0,112,0,0,0,0,0,23,0,102,0,177,0,123,0,186,0,188,0,168,0,235,0,0,0,0,0,0,0,224,0,152,0,67,0,0,0,72,0,0,0,105,0,0,0,14,0,26,0,3,0,102,0,0,0,111,0,39,0,0,0,236,0,18,0,72,0,216,0,32,0,229,0,211,0,21,0,177,0,0,0,80,0,172,0,0,0,50,0,176,0,251,0,159,0,0,0,153,0,186,0,198,0,189,0,240,0,177,0,33,0,0,0,158,0,0,0,34,0,38,0,76,0,29,0,76,0,70,0,141,0,224,0,0,0,170,0,238,0,152,0,127,0,0,0,0,0,246,0,68,0,0,0,154,0,0,0,70,0,11,0,0,0,69,0,185,0,0,0,161,0,39,0,91,0,77,0,129,0,16,0,236,0,17,0,90,0,237,0,79,0,61,0,178,0,0,0,76,0,81,0,0,0,238,0,245,0,135,0,141,0,234,0,138,0,217,0,255,0,157,0,0,0,55,0,247,0,73,0,0,0,115,0,23,0,117,0,75,0,0,0,0,0,93,0,84,0,240,0,0,0,233,0,243,0,60,0,122,0,159,0,203,0,205,0,209,0,92,0,201,0,0,0,91,0,128,0,96,0,214,0,139,0,88,0,255,0,0,0,223,0,0,0,159,0,47,0,47,0,26,0,69,0,0,0,0,0,223,0,110,0,48,0,136,0,92,0,32,0,16,0,247,0,24,0,0,0,99,0,0,0,143,0,0,0,0,0,116,0,109,0,252,0,51,0,78,0,100,0,70,0,136,0,126,0,35,0,22,0,0,0,36,0,207,0,212,0,232,0,0,0,33,0,111,0,99,0,215,0,134,0,56,0,210,0,3,0,165,0,0,0,61,0,0,0,171,0,9,0,10,0,234,0,0,0,63,0,74,0,8,0,198,0,41,0,155,0,178,0,118,0,0,0,141,0,148,0,152,0,40,0,3,0,92,0,53,0,0,0,149,0,2,0,224,0,0,0,109,0,140,0,2,0,0,0,186,0,113,0,79,0,221,0,130,0,117,0,196,0,0,0,141,0,118,0,141,0,134,0,215,0,183,0,246,0,206,0,103,0,24,0,211,0,225,0,120,0,0,0,98,0,0,0,134,0,222,0,59,0,131,0,154,0,33,0,145,0,239,0,22,0,8,0,75,0,212,0,0,0,247,0,47,0,0,0,151,0,0,0,41,0,73,0,156,0,155,0,7,0,0,0,191,0,53,0,139,0,37,0,201,0,255,0,29,0,170,0,0,0,0,0,132,0,0,0,170,0,228,0,122,0,187,0,150,0,0,0,53,0,26,0,180,0,238,0,3,0,4,0,0,0,29,0,155,0,100,0,0,0,141,0,109,0,0,0,161,0,54,0,0,0,102,0,11,0,156,0,54,0,103,0,0,0,112,0,148,0,58,0,82,0,45,0,136,0,93,0,152,0,0,0,102,0,135,0,74,0,111,0,0,0,188,0,144,0,253,0,0,0,253,0,27,0,20,0,0,0,155,0,161,0,10,0,237,0,5,0,0,0,0,0,134,0,133,0,203,0,0,0,209,0,0,0,140,0,59,0,13,0,127,0,0,0,0,0,178,0,0,0,107,0,150,0,88,0,212,0,0,0,118,0,16,0,209,0,53,0,49,0,68,0,202,0,49,0,33,0,223,0,233,0,97,0,0,0,141,0,59,0,192,0,0,0,0,0);
signal scenario_full  : scenario_type := (15,31,13,31,166,31,69,31,125,31,164,31,122,31,215,31,110,31,223,31,223,30,124,31,238,31,37,31,37,30,50,31,23,31,102,31,244,31,94,31,198,31,198,30,105,31,208,31,208,30,223,31,223,30,170,31,126,31,25,31,130,31,4,31,103,31,103,30,234,31,201,31,201,30,21,31,134,31,39,31,1,31,186,31,193,31,179,31,27,31,225,31,54,31,108,31,151,31,151,30,84,31,52,31,81,31,46,31,47,31,47,30,149,31,245,31,245,30,189,31,189,30,58,31,206,31,8,31,28,31,247,31,180,31,101,31,208,31,70,31,105,31,105,30,38,31,75,31,189,31,130,31,130,30,90,31,90,30,86,31,129,31,178,31,157,31,193,31,175,31,221,31,33,31,33,30,231,31,113,31,113,30,236,31,223,31,104,31,104,31,104,30,12,31,210,31,172,31,26,31,203,31,11,31,101,31,101,30,104,31,66,31,29,31,29,30,86,31,77,31,42,31,29,31,224,31,195,31,109,31,248,31,195,31,228,31,228,30,221,31,154,31,128,31,11,31,67,31,247,31,71,31,71,30,63,31,168,31,24,31,171,31,157,31,249,31,110,31,181,31,181,30,126,31,126,30,126,29,240,31,89,31,89,30,233,31,51,31,189,31,118,31,55,31,213,31,213,30,37,31,84,31,113,31,130,31,250,31,243,31,77,31,22,31,196,31,92,31,11,31,11,30,41,31,71,31,71,30,71,29,10,31,165,31,78,31,9,31,253,31,253,30,253,29,94,31,116,31,108,31,182,31,182,30,182,29,248,31,248,30,203,31,203,30,44,31,53,31,246,31,81,31,74,31,242,31,198,31,227,31,27,31,243,31,243,30,243,29,117,31,205,31,119,31,40,31,96,31,60,31,212,31,98,31,19,31,58,31,58,30,135,31,135,30,108,31,143,31,242,31,227,31,47,31,158,31,81,31,252,31,84,31,234,31,94,31,158,31,158,30,158,29,45,31,82,31,247,31,207,31,207,30,245,31,89,31,89,30,5,31,5,30,87,31,221,31,255,31,171,31,171,30,131,31,247,31,43,31,43,30,2,31,92,31,23,31,255,31,255,30,23,31,23,30,23,29,23,28,228,31,109,31,232,31,6,31,19,31,26,31,156,31,156,30,228,31,19,31,19,30,95,31,79,31,38,31,189,31,107,31,112,31,112,30,112,29,23,31,102,31,177,31,123,31,186,31,188,31,168,31,235,31,235,30,235,29,235,28,224,31,152,31,67,31,67,30,72,31,72,30,105,31,105,30,14,31,26,31,3,31,102,31,102,30,111,31,39,31,39,30,236,31,18,31,72,31,216,31,32,31,229,31,211,31,21,31,177,31,177,30,80,31,172,31,172,30,50,31,176,31,251,31,159,31,159,30,153,31,186,31,198,31,189,31,240,31,177,31,33,31,33,30,158,31,158,30,34,31,38,31,76,31,29,31,76,31,70,31,141,31,224,31,224,30,170,31,238,31,152,31,127,31,127,30,127,29,246,31,68,31,68,30,154,31,154,30,70,31,11,31,11,30,69,31,185,31,185,30,161,31,39,31,91,31,77,31,129,31,16,31,236,31,17,31,90,31,237,31,79,31,61,31,178,31,178,30,76,31,81,31,81,30,238,31,245,31,135,31,141,31,234,31,138,31,217,31,255,31,157,31,157,30,55,31,247,31,73,31,73,30,115,31,23,31,117,31,75,31,75,30,75,29,93,31,84,31,240,31,240,30,233,31,243,31,60,31,122,31,159,31,203,31,205,31,209,31,92,31,201,31,201,30,91,31,128,31,96,31,214,31,139,31,88,31,255,31,255,30,223,31,223,30,159,31,47,31,47,31,26,31,69,31,69,30,69,29,223,31,110,31,48,31,136,31,92,31,32,31,16,31,247,31,24,31,24,30,99,31,99,30,143,31,143,30,143,29,116,31,109,31,252,31,51,31,78,31,100,31,70,31,136,31,126,31,35,31,22,31,22,30,36,31,207,31,212,31,232,31,232,30,33,31,111,31,99,31,215,31,134,31,56,31,210,31,3,31,165,31,165,30,61,31,61,30,171,31,9,31,10,31,234,31,234,30,63,31,74,31,8,31,198,31,41,31,155,31,178,31,118,31,118,30,141,31,148,31,152,31,40,31,3,31,92,31,53,31,53,30,149,31,2,31,224,31,224,30,109,31,140,31,2,31,2,30,186,31,113,31,79,31,221,31,130,31,117,31,196,31,196,30,141,31,118,31,141,31,134,31,215,31,183,31,246,31,206,31,103,31,24,31,211,31,225,31,120,31,120,30,98,31,98,30,134,31,222,31,59,31,131,31,154,31,33,31,145,31,239,31,22,31,8,31,75,31,212,31,212,30,247,31,47,31,47,30,151,31,151,30,41,31,73,31,156,31,155,31,7,31,7,30,191,31,53,31,139,31,37,31,201,31,255,31,29,31,170,31,170,30,170,29,132,31,132,30,170,31,228,31,122,31,187,31,150,31,150,30,53,31,26,31,180,31,238,31,3,31,4,31,4,30,29,31,155,31,100,31,100,30,141,31,109,31,109,30,161,31,54,31,54,30,102,31,11,31,156,31,54,31,103,31,103,30,112,31,148,31,58,31,82,31,45,31,136,31,93,31,152,31,152,30,102,31,135,31,74,31,111,31,111,30,188,31,144,31,253,31,253,30,253,31,27,31,20,31,20,30,155,31,161,31,10,31,237,31,5,31,5,30,5,29,134,31,133,31,203,31,203,30,209,31,209,30,140,31,59,31,13,31,127,31,127,30,127,29,178,31,178,30,107,31,150,31,88,31,212,31,212,30,118,31,16,31,209,31,53,31,49,31,68,31,202,31,49,31,33,31,223,31,233,31,97,31,97,30,141,31,59,31,192,31,192,30,192,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
