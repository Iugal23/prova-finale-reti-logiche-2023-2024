-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 736;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,49,0,48,0,247,0,0,0,1,0,127,0,222,0,145,0,10,0,226,0,11,0,0,0,72,0,228,0,89,0,99,0,253,0,0,0,121,0,206,0,43,0,157,0,161,0,196,0,0,0,0,0,158,0,16,0,100,0,127,0,45,0,103,0,0,0,0,0,21,0,141,0,72,0,207,0,44,0,81,0,35,0,167,0,253,0,13,0,6,0,120,0,175,0,0,0,116,0,179,0,216,0,101,0,207,0,194,0,94,0,33,0,246,0,155,0,0,0,37,0,1,0,233,0,51,0,238,0,0,0,0,0,183,0,103,0,0,0,0,0,186,0,245,0,11,0,15,0,7,0,152,0,186,0,91,0,24,0,0,0,214,0,0,0,237,0,219,0,68,0,0,0,20,0,106,0,181,0,56,0,159,0,160,0,0,0,166,0,93,0,182,0,227,0,183,0,58,0,210,0,40,0,27,0,155,0,94,0,191,0,98,0,0,0,98,0,246,0,184,0,35,0,118,0,210,0,10,0,205,0,16,0,11,0,128,0,96,0,0,0,17,0,180,0,216,0,143,0,108,0,0,0,0,0,100,0,241,0,162,0,0,0,0,0,79,0,188,0,224,0,153,0,13,0,105,0,220,0,204,0,23,0,0,0,78,0,45,0,2,0,121,0,249,0,36,0,52,0,173,0,46,0,6,0,76,0,98,0,0,0,0,0,23,0,20,0,121,0,243,0,0,0,66,0,202,0,28,0,110,0,0,0,221,0,154,0,190,0,44,0,0,0,0,0,10,0,0,0,175,0,9,0,0,0,0,0,229,0,0,0,126,0,227,0,224,0,136,0,246,0,62,0,3,0,54,0,160,0,54,0,85,0,84,0,0,0,187,0,146,0,128,0,0,0,133,0,62,0,0,0,5,0,107,0,2,0,80,0,52,0,120,0,0,0,29,0,44,0,0,0,213,0,149,0,67,0,0,0,0,0,187,0,0,0,41,0,215,0,0,0,166,0,164,0,32,0,195,0,28,0,0,0,60,0,24,0,62,0,65,0,147,0,123,0,152,0,182,0,247,0,158,0,140,0,70,0,106,0,244,0,151,0,0,0,168,0,118,0,124,0,0,0,0,0,0,0,140,0,0,0,188,0,168,0,59,0,0,0,37,0,12,0,112,0,115,0,174,0,218,0,173,0,227,0,92,0,4,0,155,0,0,0,126,0,186,0,5,0,143,0,35,0,77,0,0,0,0,0,54,0,0,0,0,0,58,0,38,0,156,0,162,0,143,0,48,0,127,0,0,0,130,0,0,0,153,0,0,0,56,0,4,0,10,0,0,0,120,0,134,0,0,0,248,0,0,0,0,0,0,0,67,0,0,0,33,0,28,0,148,0,0,0,46,0,159,0,76,0,73,0,0,0,232,0,42,0,182,0,0,0,160,0,9,0,55,0,183,0,0,0,232,0,208,0,0,0,153,0,0,0,172,0,0,0,212,0,90,0,240,0,182,0,16,0,173,0,38,0,0,0,66,0,36,0,120,0,136,0,88,0,0,0,0,0,46,0,218,0,66,0,210,0,0,0,0,0,0,0,172,0,94,0,0,0,130,0,22,0,194,0,151,0,26,0,129,0,0,0,33,0,190,0,162,0,137,0,71,0,236,0,0,0,152,0,24,0,48,0,135,0,116,0,28,0,97,0,217,0,0,0,13,0,85,0,231,0,63,0,83,0,234,0,20,0,0,0,29,0,164,0,95,0,251,0,0,0,196,0,151,0,28,0,33,0,153,0,152,0,239,0,129,0,0,0,0,0,211,0,0,0,209,0,76,0,113,0,0,0,248,0,36,0,111,0,204,0,0,0,36,0,155,0,0,0,20,0,58,0,244,0,127,0,172,0,13,0,132,0,0,0,14,0,79,0,183,0,0,0,235,0,207,0,157,0,0,0,0,0,0,0,190,0,144,0,228,0,227,0,128,0,106,0,56,0,35,0,103,0,0,0,69,0,0,0,95,0,0,0,20,0,118,0,52,0,1,0,0,0,2,0,15,0,208,0,239,0,0,0,0,0,50,0,0,0,0,0,1,0,170,0,204,0,49,0,108,0,127,0,0,0,0,0,0,0,0,0,14,0,26,0,36,0,160,0,0,0,88,0,0,0,136,0,159,0,76,0,161,0,0,0,147,0,0,0,190,0,54,0,111,0,0,0,137,0,51,0,185,0,73,0,178,0,0,0,84,0,64,0,158,0,17,0,226,0,80,0,253,0,226,0,11,0,192,0,0,0,57,0,0,0,0,0,110,0,236,0,0,0,70,0,102,0,179,0,130,0,42,0,0,0,50,0,40,0,235,0,50,0,29,0,65,0,148,0,209,0,81,0,9,0,12,0,232,0,228,0,177,0,204,0,0,0,142,0,0,0,71,0,167,0,237,0,19,0,84,0,64,0,220,0,216,0,40,0,219,0,96,0,151,0,217,0,229,0,190,0,131,0,176,0,218,0,45,0,179,0,93,0,133,0,138,0,8,0,37,0,204,0,216,0,0,0,94,0,226,0,37,0,188,0,0,0,49,0,222,0,101,0,162,0,0,0,0,0,32,0,66,0,144,0,123,0,0,0,181,0,194,0,64,0,194,0,0,0,25,0,251,0,72,0,235,0,150,0,0,0,177,0,171,0,0,0,42,0,70,0,0,0,0,0,120,0,0,0,100,0,254,0,134,0,239,0,171,0,70,0,133,0,111,0,0,0,86,0,126,0,86,0,0,0,0,0,249,0,0,0,89,0,0,0,40,0,169,0,38,0,45,0,0,0,196,0,0,0,98,0,0,0,245,0,171,0,0,0,157,0,0,0,0,0,149,0,238,0,155,0,0,0,0,0,147,0,188,0,130,0,141,0,0,0,9,0,7,0,0,0,204,0,132,0,62,0,7,0,12,0,7,0,31,0,167,0,146,0,197,0,43,0,45,0,70,0,7,0,188,0,116,0,0,0,248,0,200,0,95,0,182,0,71,0,129,0,84,0,0,0,28,0,67,0,145,0,251,0,37,0,233,0,0,0,166,0,55,0,38,0,100,0,40,0,158,0,58,0,252,0,0,0,115,0,59,0,192,0,0,0,160,0,0,0,234,0,0,0,177,0,6,0,243,0,15,0,0,0,148,0,239,0,29,0,156,0,0,0,197,0,201,0,51,0,100,0,145,0,229,0,104,0,0,0,108,0,0,0,0,0,162,0,0,0,210,0,0,0,250,0,197,0,164,0,8,0,147,0,130,0,243,0,74,0,199,0,0,0,77,0,0,0,68,0,76,0,149,0,131,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,49,31,48,31,247,31,247,30,1,31,127,31,222,31,145,31,10,31,226,31,11,31,11,30,72,31,228,31,89,31,99,31,253,31,253,30,121,31,206,31,43,31,157,31,161,31,196,31,196,30,196,29,158,31,16,31,100,31,127,31,45,31,103,31,103,30,103,29,21,31,141,31,72,31,207,31,44,31,81,31,35,31,167,31,253,31,13,31,6,31,120,31,175,31,175,30,116,31,179,31,216,31,101,31,207,31,194,31,94,31,33,31,246,31,155,31,155,30,37,31,1,31,233,31,51,31,238,31,238,30,238,29,183,31,103,31,103,30,103,29,186,31,245,31,11,31,15,31,7,31,152,31,186,31,91,31,24,31,24,30,214,31,214,30,237,31,219,31,68,31,68,30,20,31,106,31,181,31,56,31,159,31,160,31,160,30,166,31,93,31,182,31,227,31,183,31,58,31,210,31,40,31,27,31,155,31,94,31,191,31,98,31,98,30,98,31,246,31,184,31,35,31,118,31,210,31,10,31,205,31,16,31,11,31,128,31,96,31,96,30,17,31,180,31,216,31,143,31,108,31,108,30,108,29,100,31,241,31,162,31,162,30,162,29,79,31,188,31,224,31,153,31,13,31,105,31,220,31,204,31,23,31,23,30,78,31,45,31,2,31,121,31,249,31,36,31,52,31,173,31,46,31,6,31,76,31,98,31,98,30,98,29,23,31,20,31,121,31,243,31,243,30,66,31,202,31,28,31,110,31,110,30,221,31,154,31,190,31,44,31,44,30,44,29,10,31,10,30,175,31,9,31,9,30,9,29,229,31,229,30,126,31,227,31,224,31,136,31,246,31,62,31,3,31,54,31,160,31,54,31,85,31,84,31,84,30,187,31,146,31,128,31,128,30,133,31,62,31,62,30,5,31,107,31,2,31,80,31,52,31,120,31,120,30,29,31,44,31,44,30,213,31,149,31,67,31,67,30,67,29,187,31,187,30,41,31,215,31,215,30,166,31,164,31,32,31,195,31,28,31,28,30,60,31,24,31,62,31,65,31,147,31,123,31,152,31,182,31,247,31,158,31,140,31,70,31,106,31,244,31,151,31,151,30,168,31,118,31,124,31,124,30,124,29,124,28,140,31,140,30,188,31,168,31,59,31,59,30,37,31,12,31,112,31,115,31,174,31,218,31,173,31,227,31,92,31,4,31,155,31,155,30,126,31,186,31,5,31,143,31,35,31,77,31,77,30,77,29,54,31,54,30,54,29,58,31,38,31,156,31,162,31,143,31,48,31,127,31,127,30,130,31,130,30,153,31,153,30,56,31,4,31,10,31,10,30,120,31,134,31,134,30,248,31,248,30,248,29,248,28,67,31,67,30,33,31,28,31,148,31,148,30,46,31,159,31,76,31,73,31,73,30,232,31,42,31,182,31,182,30,160,31,9,31,55,31,183,31,183,30,232,31,208,31,208,30,153,31,153,30,172,31,172,30,212,31,90,31,240,31,182,31,16,31,173,31,38,31,38,30,66,31,36,31,120,31,136,31,88,31,88,30,88,29,46,31,218,31,66,31,210,31,210,30,210,29,210,28,172,31,94,31,94,30,130,31,22,31,194,31,151,31,26,31,129,31,129,30,33,31,190,31,162,31,137,31,71,31,236,31,236,30,152,31,24,31,48,31,135,31,116,31,28,31,97,31,217,31,217,30,13,31,85,31,231,31,63,31,83,31,234,31,20,31,20,30,29,31,164,31,95,31,251,31,251,30,196,31,151,31,28,31,33,31,153,31,152,31,239,31,129,31,129,30,129,29,211,31,211,30,209,31,76,31,113,31,113,30,248,31,36,31,111,31,204,31,204,30,36,31,155,31,155,30,20,31,58,31,244,31,127,31,172,31,13,31,132,31,132,30,14,31,79,31,183,31,183,30,235,31,207,31,157,31,157,30,157,29,157,28,190,31,144,31,228,31,227,31,128,31,106,31,56,31,35,31,103,31,103,30,69,31,69,30,95,31,95,30,20,31,118,31,52,31,1,31,1,30,2,31,15,31,208,31,239,31,239,30,239,29,50,31,50,30,50,29,1,31,170,31,204,31,49,31,108,31,127,31,127,30,127,29,127,28,127,27,14,31,26,31,36,31,160,31,160,30,88,31,88,30,136,31,159,31,76,31,161,31,161,30,147,31,147,30,190,31,54,31,111,31,111,30,137,31,51,31,185,31,73,31,178,31,178,30,84,31,64,31,158,31,17,31,226,31,80,31,253,31,226,31,11,31,192,31,192,30,57,31,57,30,57,29,110,31,236,31,236,30,70,31,102,31,179,31,130,31,42,31,42,30,50,31,40,31,235,31,50,31,29,31,65,31,148,31,209,31,81,31,9,31,12,31,232,31,228,31,177,31,204,31,204,30,142,31,142,30,71,31,167,31,237,31,19,31,84,31,64,31,220,31,216,31,40,31,219,31,96,31,151,31,217,31,229,31,190,31,131,31,176,31,218,31,45,31,179,31,93,31,133,31,138,31,8,31,37,31,204,31,216,31,216,30,94,31,226,31,37,31,188,31,188,30,49,31,222,31,101,31,162,31,162,30,162,29,32,31,66,31,144,31,123,31,123,30,181,31,194,31,64,31,194,31,194,30,25,31,251,31,72,31,235,31,150,31,150,30,177,31,171,31,171,30,42,31,70,31,70,30,70,29,120,31,120,30,100,31,254,31,134,31,239,31,171,31,70,31,133,31,111,31,111,30,86,31,126,31,86,31,86,30,86,29,249,31,249,30,89,31,89,30,40,31,169,31,38,31,45,31,45,30,196,31,196,30,98,31,98,30,245,31,171,31,171,30,157,31,157,30,157,29,149,31,238,31,155,31,155,30,155,29,147,31,188,31,130,31,141,31,141,30,9,31,7,31,7,30,204,31,132,31,62,31,7,31,12,31,7,31,31,31,167,31,146,31,197,31,43,31,45,31,70,31,7,31,188,31,116,31,116,30,248,31,200,31,95,31,182,31,71,31,129,31,84,31,84,30,28,31,67,31,145,31,251,31,37,31,233,31,233,30,166,31,55,31,38,31,100,31,40,31,158,31,58,31,252,31,252,30,115,31,59,31,192,31,192,30,160,31,160,30,234,31,234,30,177,31,6,31,243,31,15,31,15,30,148,31,239,31,29,31,156,31,156,30,197,31,201,31,51,31,100,31,145,31,229,31,104,31,104,30,108,31,108,30,108,29,162,31,162,30,210,31,210,30,250,31,197,31,164,31,8,31,147,31,130,31,243,31,74,31,199,31,199,30,77,31,77,30,68,31,76,31,149,31,131,31,131,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
