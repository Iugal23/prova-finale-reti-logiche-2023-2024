-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 634;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,254,0,133,0,170,0,254,0,193,0,20,0,29,0,61,0,40,0,238,0,119,0,111,0,218,0,137,0,0,0,0,0,172,0,246,0,225,0,227,0,202,0,251,0,82,0,25,0,14,0,0,0,104,0,0,0,38,0,248,0,251,0,198,0,210,0,21,0,0,0,238,0,119,0,70,0,175,0,213,0,255,0,191,0,184,0,37,0,0,0,0,0,0,0,221,0,0,0,0,0,3,0,139,0,76,0,200,0,249,0,0,0,204,0,151,0,0,0,149,0,0,0,132,0,30,0,170,0,152,0,205,0,23,0,138,0,0,0,0,0,34,0,157,0,169,0,244,0,175,0,245,0,0,0,129,0,211,0,76,0,192,0,51,0,174,0,147,0,82,0,41,0,167,0,185,0,108,0,208,0,0,0,198,0,157,0,0,0,143,0,33,0,155,0,234,0,102,0,17,0,0,0,206,0,0,0,116,0,130,0,176,0,65,0,0,0,86,0,0,0,167,0,13,0,31,0,253,0,76,0,108,0,85,0,28,0,152,0,205,0,212,0,0,0,184,0,26,0,0,0,76,0,235,0,25,0,203,0,243,0,3,0,59,0,159,0,0,0,0,0,136,0,240,0,34,0,226,0,159,0,143,0,178,0,65,0,229,0,248,0,38,0,225,0,191,0,250,0,113,0,33,0,74,0,41,0,88,0,243,0,126,0,127,0,190,0,73,0,27,0,172,0,124,0,0,0,244,0,197,0,147,0,229,0,157,0,0,0,0,0,107,0,104,0,66,0,32,0,122,0,72,0,183,0,94,0,74,0,0,0,0,0,85,0,119,0,62,0,64,0,0,0,0,0,0,0,203,0,46,0,62,0,150,0,23,0,56,0,131,0,74,0,4,0,0,0,183,0,4,0,0,0,179,0,0,0,147,0,0,0,0,0,176,0,243,0,28,0,0,0,251,0,44,0,105,0,171,0,61,0,12,0,188,0,23,0,71,0,154,0,87,0,166,0,179,0,12,0,34,0,233,0,155,0,11,0,73,0,177,0,81,0,100,0,169,0,191,0,202,0,22,0,0,0,112,0,59,0,148,0,183,0,76,0,72,0,0,0,249,0,217,0,254,0,0,0,25,0,56,0,119,0,41,0,110,0,206,0,153,0,113,0,8,0,51,0,59,0,175,0,0,0,137,0,176,0,219,0,107,0,85,0,182,0,206,0,120,0,49,0,39,0,96,0,68,0,132,0,124,0,195,0,91,0,130,0,0,0,0,0,240,0,149,0,0,0,0,0,72,0,159,0,153,0,0,0,0,0,142,0,165,0,205,0,42,0,110,0,40,0,0,0,203,0,47,0,44,0,74,0,0,0,236,0,12,0,87,0,111,0,35,0,236,0,41,0,93,0,0,0,223,0,66,0,138,0,47,0,164,0,141,0,97,0,0,0,130,0,44,0,48,0,124,0,78,0,174,0,0,0,36,0,117,0,235,0,214,0,0,0,28,0,156,0,217,0,70,0,141,0,0,0,53,0,29,0,105,0,0,0,0,0,57,0,0,0,236,0,12,0,158,0,0,0,172,0,105,0,0,0,0,0,127,0,0,0,124,0,0,0,121,0,0,0,0,0,0,0,13,0,0,0,62,0,62,0,0,0,86,0,53,0,0,0,242,0,219,0,163,0,6,0,167,0,150,0,138,0,152,0,41,0,71,0,172,0,120,0,157,0,146,0,55,0,12,0,0,0,186,0,178,0,54,0,181,0,138,0,233,0,179,0,207,0,0,0,0,0,46,0,94,0,0,0,191,0,0,0,73,0,0,0,181,0,24,0,0,0,70,0,0,0,0,0,64,0,0,0,105,0,154,0,4,0,165,0,133,0,10,0,98,0,0,0,0,0,225,0,139,0,105,0,242,0,0,0,0,0,89,0,148,0,252,0,15,0,50,0,17,0,133,0,242,0,28,0,166,0,12,0,164,0,85,0,42,0,204,0,129,0,35,0,156,0,125,0,250,0,207,0,177,0,26,0,163,0,132,0,140,0,56,0,120,0,247,0,43,0,201,0,162,0,84,0,0,0,218,0,0,0,0,0,10,0,92,0,0,0,154,0,80,0,0,0,226,0,0,0,23,0,0,0,117,0,45,0,7,0,110,0,102,0,0,0,216,0,64,0,88,0,0,0,49,0,49,0,23,0,113,0,0,0,29,0,198,0,189,0,35,0,70,0,205,0,0,0,161,0,0,0,140,0,82,0,236,0,0,0,156,0,112,0,159,0,65,0,7,0,0,0,124,0,84,0,219,0,113,0,53,0,0,0,196,0,21,0,195,0,152,0,68,0,0,0,212,0,32,0,1,0,216,0,132,0,84,0,237,0,44,0,0,0,158,0,89,0,25,0,199,0,246,0,118,0,117,0,9,0,239,0,47,0,8,0,182,0,117,0,31,0,185,0,0,0,203,0,76,0,105,0,0,0,13,0,0,0,53,0,0,0,116,0,181,0,146,0,217,0,77,0,110,0,254,0,37,0,8,0,127,0,200,0,0,0,91,0,9,0,197,0,0,0,132,0,196,0,175,0,0,0,0,0,207,0,0,0,42,0,220,0,168,0,178,0,68,0,149,0,140,0,23,0,0,0,211,0,241,0,156,0,196,0,32,0,0,0,242,0,69,0,0,0,29,0,128,0,189,0,152,0,30,0,0,0,96,0,165,0,0,0,0,0,75,0,95,0,141,0,0,0,0,0,209,0,211,0,198,0,155,0,244,0,249,0,166,0,235,0,163,0,111,0,216,0,250,0,0,0,81,0,202,0,124,0,87,0,253,0,50,0,71,0,55,0,102,0,161,0,0,0,112,0,183,0,180,0);
signal scenario_full  : scenario_type := (68,31,254,31,133,31,170,31,254,31,193,31,20,31,29,31,61,31,40,31,238,31,119,31,111,31,218,31,137,31,137,30,137,29,172,31,246,31,225,31,227,31,202,31,251,31,82,31,25,31,14,31,14,30,104,31,104,30,38,31,248,31,251,31,198,31,210,31,21,31,21,30,238,31,119,31,70,31,175,31,213,31,255,31,191,31,184,31,37,31,37,30,37,29,37,28,221,31,221,30,221,29,3,31,139,31,76,31,200,31,249,31,249,30,204,31,151,31,151,30,149,31,149,30,132,31,30,31,170,31,152,31,205,31,23,31,138,31,138,30,138,29,34,31,157,31,169,31,244,31,175,31,245,31,245,30,129,31,211,31,76,31,192,31,51,31,174,31,147,31,82,31,41,31,167,31,185,31,108,31,208,31,208,30,198,31,157,31,157,30,143,31,33,31,155,31,234,31,102,31,17,31,17,30,206,31,206,30,116,31,130,31,176,31,65,31,65,30,86,31,86,30,167,31,13,31,31,31,253,31,76,31,108,31,85,31,28,31,152,31,205,31,212,31,212,30,184,31,26,31,26,30,76,31,235,31,25,31,203,31,243,31,3,31,59,31,159,31,159,30,159,29,136,31,240,31,34,31,226,31,159,31,143,31,178,31,65,31,229,31,248,31,38,31,225,31,191,31,250,31,113,31,33,31,74,31,41,31,88,31,243,31,126,31,127,31,190,31,73,31,27,31,172,31,124,31,124,30,244,31,197,31,147,31,229,31,157,31,157,30,157,29,107,31,104,31,66,31,32,31,122,31,72,31,183,31,94,31,74,31,74,30,74,29,85,31,119,31,62,31,64,31,64,30,64,29,64,28,203,31,46,31,62,31,150,31,23,31,56,31,131,31,74,31,4,31,4,30,183,31,4,31,4,30,179,31,179,30,147,31,147,30,147,29,176,31,243,31,28,31,28,30,251,31,44,31,105,31,171,31,61,31,12,31,188,31,23,31,71,31,154,31,87,31,166,31,179,31,12,31,34,31,233,31,155,31,11,31,73,31,177,31,81,31,100,31,169,31,191,31,202,31,22,31,22,30,112,31,59,31,148,31,183,31,76,31,72,31,72,30,249,31,217,31,254,31,254,30,25,31,56,31,119,31,41,31,110,31,206,31,153,31,113,31,8,31,51,31,59,31,175,31,175,30,137,31,176,31,219,31,107,31,85,31,182,31,206,31,120,31,49,31,39,31,96,31,68,31,132,31,124,31,195,31,91,31,130,31,130,30,130,29,240,31,149,31,149,30,149,29,72,31,159,31,153,31,153,30,153,29,142,31,165,31,205,31,42,31,110,31,40,31,40,30,203,31,47,31,44,31,74,31,74,30,236,31,12,31,87,31,111,31,35,31,236,31,41,31,93,31,93,30,223,31,66,31,138,31,47,31,164,31,141,31,97,31,97,30,130,31,44,31,48,31,124,31,78,31,174,31,174,30,36,31,117,31,235,31,214,31,214,30,28,31,156,31,217,31,70,31,141,31,141,30,53,31,29,31,105,31,105,30,105,29,57,31,57,30,236,31,12,31,158,31,158,30,172,31,105,31,105,30,105,29,127,31,127,30,124,31,124,30,121,31,121,30,121,29,121,28,13,31,13,30,62,31,62,31,62,30,86,31,53,31,53,30,242,31,219,31,163,31,6,31,167,31,150,31,138,31,152,31,41,31,71,31,172,31,120,31,157,31,146,31,55,31,12,31,12,30,186,31,178,31,54,31,181,31,138,31,233,31,179,31,207,31,207,30,207,29,46,31,94,31,94,30,191,31,191,30,73,31,73,30,181,31,24,31,24,30,70,31,70,30,70,29,64,31,64,30,105,31,154,31,4,31,165,31,133,31,10,31,98,31,98,30,98,29,225,31,139,31,105,31,242,31,242,30,242,29,89,31,148,31,252,31,15,31,50,31,17,31,133,31,242,31,28,31,166,31,12,31,164,31,85,31,42,31,204,31,129,31,35,31,156,31,125,31,250,31,207,31,177,31,26,31,163,31,132,31,140,31,56,31,120,31,247,31,43,31,201,31,162,31,84,31,84,30,218,31,218,30,218,29,10,31,92,31,92,30,154,31,80,31,80,30,226,31,226,30,23,31,23,30,117,31,45,31,7,31,110,31,102,31,102,30,216,31,64,31,88,31,88,30,49,31,49,31,23,31,113,31,113,30,29,31,198,31,189,31,35,31,70,31,205,31,205,30,161,31,161,30,140,31,82,31,236,31,236,30,156,31,112,31,159,31,65,31,7,31,7,30,124,31,84,31,219,31,113,31,53,31,53,30,196,31,21,31,195,31,152,31,68,31,68,30,212,31,32,31,1,31,216,31,132,31,84,31,237,31,44,31,44,30,158,31,89,31,25,31,199,31,246,31,118,31,117,31,9,31,239,31,47,31,8,31,182,31,117,31,31,31,185,31,185,30,203,31,76,31,105,31,105,30,13,31,13,30,53,31,53,30,116,31,181,31,146,31,217,31,77,31,110,31,254,31,37,31,8,31,127,31,200,31,200,30,91,31,9,31,197,31,197,30,132,31,196,31,175,31,175,30,175,29,207,31,207,30,42,31,220,31,168,31,178,31,68,31,149,31,140,31,23,31,23,30,211,31,241,31,156,31,196,31,32,31,32,30,242,31,69,31,69,30,29,31,128,31,189,31,152,31,30,31,30,30,96,31,165,31,165,30,165,29,75,31,95,31,141,31,141,30,141,29,209,31,211,31,198,31,155,31,244,31,249,31,166,31,235,31,163,31,111,31,216,31,250,31,250,30,81,31,202,31,124,31,87,31,253,31,50,31,71,31,55,31,102,31,161,31,161,30,112,31,183,31,180,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
