-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_652 is
end project_tb_652;

architecture project_tb_arch_652 of project_tb_652 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 980;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,0,0,191,0,103,0,12,0,65,0,129,0,100,0,121,0,0,0,33,0,144,0,180,0,15,0,0,0,14,0,2,0,209,0,253,0,100,0,151,0,21,0,249,0,179,0,0,0,24,0,152,0,82,0,228,0,9,0,222,0,102,0,144,0,0,0,67,0,54,0,28,0,203,0,238,0,227,0,0,0,0,0,207,0,45,0,196,0,51,0,122,0,4,0,0,0,122,0,72,0,0,0,111,0,142,0,45,0,112,0,237,0,0,0,0,0,147,0,229,0,39,0,212,0,19,0,0,0,0,0,245,0,87,0,19,0,166,0,63,0,107,0,170,0,0,0,54,0,254,0,22,0,143,0,255,0,134,0,18,0,247,0,0,0,71,0,125,0,9,0,173,0,18,0,74,0,88,0,222,0,48,0,138,0,48,0,186,0,136,0,12,0,0,0,99,0,0,0,173,0,98,0,0,0,187,0,145,0,13,0,119,0,0,0,0,0,62,0,0,0,83,0,254,0,111,0,100,0,211,0,0,0,0,0,119,0,87,0,227,0,94,0,166,0,0,0,56,0,27,0,228,0,0,0,108,0,16,0,0,0,194,0,23,0,106,0,127,0,0,0,0,0,0,0,249,0,0,0,18,0,44,0,93,0,39,0,177,0,225,0,14,0,227,0,141,0,114,0,40,0,0,0,211,0,211,0,0,0,126,0,59,0,6,0,0,0,75,0,0,0,97,0,184,0,36,0,195,0,0,0,22,0,170,0,241,0,174,0,181,0,252,0,95,0,0,0,160,0,0,0,197,0,217,0,208,0,122,0,0,0,0,0,162,0,149,0,82,0,74,0,0,0,7,0,24,0,0,0,236,0,232,0,255,0,105,0,156,0,0,0,18,0,42,0,251,0,251,0,0,0,115,0,0,0,0,0,59,0,232,0,190,0,229,0,83,0,248,0,134,0,96,0,81,0,206,0,147,0,13,0,0,0,136,0,245,0,36,0,246,0,100,0,0,0,196,0,108,0,38,0,227,0,243,0,136,0,11,0,165,0,79,0,244,0,86,0,83,0,237,0,90,0,18,0,149,0,191,0,232,0,140,0,74,0,160,0,243,0,0,0,31,0,225,0,0,0,232,0,42,0,0,0,177,0,49,0,202,0,125,0,17,0,45,0,116,0,255,0,189,0,185,0,0,0,56,0,1,0,246,0,0,0,48,0,0,0,143,0,9,0,69,0,1,0,72,0,0,0,237,0,0,0,0,0,146,0,156,0,67,0,0,0,153,0,122,0,0,0,117,0,155,0,166,0,172,0,132,0,3,0,145,0,167,0,185,0,0,0,0,0,0,0,167,0,71,0,0,0,135,0,0,0,197,0,215,0,221,0,0,0,105,0,0,0,210,0,0,0,6,0,0,0,225,0,119,0,83,0,161,0,233,0,61,0,158,0,236,0,98,0,151,0,107,0,200,0,161,0,132,0,118,0,223,0,255,0,181,0,155,0,62,0,206,0,161,0,234,0,225,0,0,0,100,0,0,0,0,0,156,0,23,0,196,0,213,0,0,0,135,0,0,0,165,0,181,0,150,0,141,0,58,0,130,0,0,0,193,0,146,0,250,0,37,0,4,0,228,0,49,0,171,0,113,0,212,0,226,0,115,0,103,0,164,0,199,0,0,0,84,0,0,0,0,0,0,0,32,0,145,0,82,0,46,0,77,0,154,0,153,0,101,0,0,0,210,0,162,0,0,0,178,0,0,0,175,0,165,0,80,0,74,0,189,0,11,0,110,0,0,0,118,0,81,0,247,0,109,0,144,0,174,0,0,0,94,0,0,0,136,0,255,0,204,0,131,0,149,0,99,0,162,0,153,0,132,0,223,0,0,0,0,0,143,0,58,0,0,0,119,0,0,0,82,0,192,0,245,0,0,0,179,0,46,0,0,0,142,0,46,0,206,0,0,0,172,0,85,0,222,0,0,0,0,0,185,0,176,0,115,0,123,0,117,0,66,0,57,0,188,0,30,0,91,0,39,0,148,0,117,0,169,0,10,0,182,0,12,0,123,0,157,0,89,0,51,0,116,0,3,0,18,0,59,0,223,0,0,0,38,0,176,0,219,0,151,0,227,0,231,0,132,0,20,0,77,0,98,0,247,0,147,0,0,0,218,0,157,0,116,0,78,0,129,0,147,0,108,0,134,0,203,0,156,0,0,0,87,0,0,0,164,0,91,0,35,0,0,0,44,0,0,0,0,0,0,0,0,0,182,0,202,0,0,0,207,0,57,0,10,0,68,0,23,0,242,0,218,0,186,0,170,0,30,0,184,0,149,0,116,0,94,0,225,0,59,0,14,0,0,0,4,0,190,0,162,0,250,0,0,0,131,0,48,0,0,0,144,0,224,0,60,0,88,0,0,0,172,0,0,0,156,0,0,0,37,0,92,0,0,0,72,0,136,0,209,0,120,0,178,0,0,0,0,0,147,0,125,0,81,0,193,0,0,0,221,0,213,0,234,0,211,0,0,0,128,0,25,0,191,0,134,0,0,0,65,0,215,0,0,0,147,0,0,0,0,0,183,0,122,0,0,0,0,0,83,0,0,0,0,0,60,0,222,0,46,0,141,0,114,0,0,0,122,0,0,0,29,0,37,0,232,0,0,0,0,0,162,0,53,0,232,0,0,0,96,0,55,0,110,0,0,0,183,0,183,0,86,0,186,0,41,0,100,0,73,0,230,0,21,0,121,0,127,0,144,0,232,0,239,0,241,0,69,0,190,0,158,0,0,0,178,0,83,0,143,0,0,0,0,0,202,0,0,0,153,0,96,0,124,0,162,0,145,0,156,0,55,0,148,0,184,0,160,0,227,0,234,0,33,0,0,0,119,0,158,0,175,0,243,0,203,0,197,0,0,0,171,0,143,0,46,0,0,0,62,0,2,0,0,0,195,0,0,0,104,0,0,0,205,0,192,0,103,0,36,0,208,0,240,0,0,0,77,0,142,0,151,0,19,0,119,0,75,0,151,0,163,0,142,0,140,0,43,0,3,0,11,0,32,0,251,0,0,0,107,0,152,0,171,0,0,0,0,0,182,0,31,0,133,0,253,0,226,0,98,0,11,0,85,0,183,0,89,0,62,0,88,0,182,0,37,0,136,0,0,0,63,0,232,0,0,0,97,0,68,0,207,0,0,0,47,0,88,0,41,0,137,0,165,0,233,0,144,0,27,0,119,0,237,0,63,0,250,0,193,0,113,0,70,0,184,0,1,0,241,0,37,0,242,0,126,0,253,0,98,0,0,0,0,0,0,0,3,0,109,0,51,0,154,0,187,0,61,0,45,0,232,0,135,0,202,0,0,0,0,0,249,0,40,0,97,0,81,0,181,0,143,0,126,0,216,0,139,0,6,0,1,0,32,0,18,0,113,0,0,0,35,0,111,0,182,0,185,0,94,0,199,0,207,0,7,0,175,0,119,0,151,0,130,0,234,0,152,0,78,0,0,0,231,0,48,0,91,0,144,0,184,0,201,0,101,0,81,0,0,0,13,0,0,0,0,0,108,0,0,0,207,0,105,0,1,0,171,0,149,0,40,0,0,0,212,0,6,0,255,0,184,0,0,0,114,0,30,0,192,0,16,0,192,0,158,0,0,0,60,0,15,0,100,0,0,0,0,0,167,0,210,0,229,0,68,0,182,0,0,0,145,0,48,0,164,0,0,0,245,0,0,0,0,0,120,0,16,0,110,0,98,0,221,0,0,0,0,0,56,0,0,0,28,0,239,0,34,0,57,0,37,0,50,0,236,0,171,0,37,0,0,0,70,0,0,0,0,0,0,0,0,0,165,0,0,0,0,0,34,0,199,0,77,0,74,0,0,0,200,0,0,0,113,0,186,0,0,0,162,0,164,0,109,0,40,0,141,0,0,0,148,0,69,0,0,0,202,0,11,0,213,0,152,0,0,0,17,0,187,0,184,0,0,0,54,0,24,0,85,0,0,0,227,0,83,0,96,0,0,0,26,0,145,0,162,0,0,0,67,0,0,0,2,0,0,0,20,0,83,0,10,0,12,0,90,0,133,0,44,0,14,0,0,0,107,0,110,0,21,0,166,0,48,0,183,0,183,0,156,0,0,0,150,0,210,0,193,0,4,0,203,0,76,0,0,0,122,0,145,0,132,0,0,0,130,0,48,0,0,0,210,0,182,0,124,0,64,0,124,0,0,0,53,0,75,0,226,0,239,0,231,0,63,0,0,0,165,0,52,0,205,0,101,0,34,0,39,0,0,0,246,0,0,0,0,0,157,0,18,0,111,0,135,0,18,0,64,0,0,0,65,0,67,0,169,0,115,0,5,0,95,0,19,0,200,0,26,0,164,0,0,0,42,0,241,0,207,0,239,0,53,0,119,0,214,0,0,0,173,0,155,0);
signal scenario_full  : scenario_type := (149,31,149,30,191,31,103,31,12,31,65,31,129,31,100,31,121,31,121,30,33,31,144,31,180,31,15,31,15,30,14,31,2,31,209,31,253,31,100,31,151,31,21,31,249,31,179,31,179,30,24,31,152,31,82,31,228,31,9,31,222,31,102,31,144,31,144,30,67,31,54,31,28,31,203,31,238,31,227,31,227,30,227,29,207,31,45,31,196,31,51,31,122,31,4,31,4,30,122,31,72,31,72,30,111,31,142,31,45,31,112,31,237,31,237,30,237,29,147,31,229,31,39,31,212,31,19,31,19,30,19,29,245,31,87,31,19,31,166,31,63,31,107,31,170,31,170,30,54,31,254,31,22,31,143,31,255,31,134,31,18,31,247,31,247,30,71,31,125,31,9,31,173,31,18,31,74,31,88,31,222,31,48,31,138,31,48,31,186,31,136,31,12,31,12,30,99,31,99,30,173,31,98,31,98,30,187,31,145,31,13,31,119,31,119,30,119,29,62,31,62,30,83,31,254,31,111,31,100,31,211,31,211,30,211,29,119,31,87,31,227,31,94,31,166,31,166,30,56,31,27,31,228,31,228,30,108,31,16,31,16,30,194,31,23,31,106,31,127,31,127,30,127,29,127,28,249,31,249,30,18,31,44,31,93,31,39,31,177,31,225,31,14,31,227,31,141,31,114,31,40,31,40,30,211,31,211,31,211,30,126,31,59,31,6,31,6,30,75,31,75,30,97,31,184,31,36,31,195,31,195,30,22,31,170,31,241,31,174,31,181,31,252,31,95,31,95,30,160,31,160,30,197,31,217,31,208,31,122,31,122,30,122,29,162,31,149,31,82,31,74,31,74,30,7,31,24,31,24,30,236,31,232,31,255,31,105,31,156,31,156,30,18,31,42,31,251,31,251,31,251,30,115,31,115,30,115,29,59,31,232,31,190,31,229,31,83,31,248,31,134,31,96,31,81,31,206,31,147,31,13,31,13,30,136,31,245,31,36,31,246,31,100,31,100,30,196,31,108,31,38,31,227,31,243,31,136,31,11,31,165,31,79,31,244,31,86,31,83,31,237,31,90,31,18,31,149,31,191,31,232,31,140,31,74,31,160,31,243,31,243,30,31,31,225,31,225,30,232,31,42,31,42,30,177,31,49,31,202,31,125,31,17,31,45,31,116,31,255,31,189,31,185,31,185,30,56,31,1,31,246,31,246,30,48,31,48,30,143,31,9,31,69,31,1,31,72,31,72,30,237,31,237,30,237,29,146,31,156,31,67,31,67,30,153,31,122,31,122,30,117,31,155,31,166,31,172,31,132,31,3,31,145,31,167,31,185,31,185,30,185,29,185,28,167,31,71,31,71,30,135,31,135,30,197,31,215,31,221,31,221,30,105,31,105,30,210,31,210,30,6,31,6,30,225,31,119,31,83,31,161,31,233,31,61,31,158,31,236,31,98,31,151,31,107,31,200,31,161,31,132,31,118,31,223,31,255,31,181,31,155,31,62,31,206,31,161,31,234,31,225,31,225,30,100,31,100,30,100,29,156,31,23,31,196,31,213,31,213,30,135,31,135,30,165,31,181,31,150,31,141,31,58,31,130,31,130,30,193,31,146,31,250,31,37,31,4,31,228,31,49,31,171,31,113,31,212,31,226,31,115,31,103,31,164,31,199,31,199,30,84,31,84,30,84,29,84,28,32,31,145,31,82,31,46,31,77,31,154,31,153,31,101,31,101,30,210,31,162,31,162,30,178,31,178,30,175,31,165,31,80,31,74,31,189,31,11,31,110,31,110,30,118,31,81,31,247,31,109,31,144,31,174,31,174,30,94,31,94,30,136,31,255,31,204,31,131,31,149,31,99,31,162,31,153,31,132,31,223,31,223,30,223,29,143,31,58,31,58,30,119,31,119,30,82,31,192,31,245,31,245,30,179,31,46,31,46,30,142,31,46,31,206,31,206,30,172,31,85,31,222,31,222,30,222,29,185,31,176,31,115,31,123,31,117,31,66,31,57,31,188,31,30,31,91,31,39,31,148,31,117,31,169,31,10,31,182,31,12,31,123,31,157,31,89,31,51,31,116,31,3,31,18,31,59,31,223,31,223,30,38,31,176,31,219,31,151,31,227,31,231,31,132,31,20,31,77,31,98,31,247,31,147,31,147,30,218,31,157,31,116,31,78,31,129,31,147,31,108,31,134,31,203,31,156,31,156,30,87,31,87,30,164,31,91,31,35,31,35,30,44,31,44,30,44,29,44,28,44,27,182,31,202,31,202,30,207,31,57,31,10,31,68,31,23,31,242,31,218,31,186,31,170,31,30,31,184,31,149,31,116,31,94,31,225,31,59,31,14,31,14,30,4,31,190,31,162,31,250,31,250,30,131,31,48,31,48,30,144,31,224,31,60,31,88,31,88,30,172,31,172,30,156,31,156,30,37,31,92,31,92,30,72,31,136,31,209,31,120,31,178,31,178,30,178,29,147,31,125,31,81,31,193,31,193,30,221,31,213,31,234,31,211,31,211,30,128,31,25,31,191,31,134,31,134,30,65,31,215,31,215,30,147,31,147,30,147,29,183,31,122,31,122,30,122,29,83,31,83,30,83,29,60,31,222,31,46,31,141,31,114,31,114,30,122,31,122,30,29,31,37,31,232,31,232,30,232,29,162,31,53,31,232,31,232,30,96,31,55,31,110,31,110,30,183,31,183,31,86,31,186,31,41,31,100,31,73,31,230,31,21,31,121,31,127,31,144,31,232,31,239,31,241,31,69,31,190,31,158,31,158,30,178,31,83,31,143,31,143,30,143,29,202,31,202,30,153,31,96,31,124,31,162,31,145,31,156,31,55,31,148,31,184,31,160,31,227,31,234,31,33,31,33,30,119,31,158,31,175,31,243,31,203,31,197,31,197,30,171,31,143,31,46,31,46,30,62,31,2,31,2,30,195,31,195,30,104,31,104,30,205,31,192,31,103,31,36,31,208,31,240,31,240,30,77,31,142,31,151,31,19,31,119,31,75,31,151,31,163,31,142,31,140,31,43,31,3,31,11,31,32,31,251,31,251,30,107,31,152,31,171,31,171,30,171,29,182,31,31,31,133,31,253,31,226,31,98,31,11,31,85,31,183,31,89,31,62,31,88,31,182,31,37,31,136,31,136,30,63,31,232,31,232,30,97,31,68,31,207,31,207,30,47,31,88,31,41,31,137,31,165,31,233,31,144,31,27,31,119,31,237,31,63,31,250,31,193,31,113,31,70,31,184,31,1,31,241,31,37,31,242,31,126,31,253,31,98,31,98,30,98,29,98,28,3,31,109,31,51,31,154,31,187,31,61,31,45,31,232,31,135,31,202,31,202,30,202,29,249,31,40,31,97,31,81,31,181,31,143,31,126,31,216,31,139,31,6,31,1,31,32,31,18,31,113,31,113,30,35,31,111,31,182,31,185,31,94,31,199,31,207,31,7,31,175,31,119,31,151,31,130,31,234,31,152,31,78,31,78,30,231,31,48,31,91,31,144,31,184,31,201,31,101,31,81,31,81,30,13,31,13,30,13,29,108,31,108,30,207,31,105,31,1,31,171,31,149,31,40,31,40,30,212,31,6,31,255,31,184,31,184,30,114,31,30,31,192,31,16,31,192,31,158,31,158,30,60,31,15,31,100,31,100,30,100,29,167,31,210,31,229,31,68,31,182,31,182,30,145,31,48,31,164,31,164,30,245,31,245,30,245,29,120,31,16,31,110,31,98,31,221,31,221,30,221,29,56,31,56,30,28,31,239,31,34,31,57,31,37,31,50,31,236,31,171,31,37,31,37,30,70,31,70,30,70,29,70,28,70,27,165,31,165,30,165,29,34,31,199,31,77,31,74,31,74,30,200,31,200,30,113,31,186,31,186,30,162,31,164,31,109,31,40,31,141,31,141,30,148,31,69,31,69,30,202,31,11,31,213,31,152,31,152,30,17,31,187,31,184,31,184,30,54,31,24,31,85,31,85,30,227,31,83,31,96,31,96,30,26,31,145,31,162,31,162,30,67,31,67,30,2,31,2,30,20,31,83,31,10,31,12,31,90,31,133,31,44,31,14,31,14,30,107,31,110,31,21,31,166,31,48,31,183,31,183,31,156,31,156,30,150,31,210,31,193,31,4,31,203,31,76,31,76,30,122,31,145,31,132,31,132,30,130,31,48,31,48,30,210,31,182,31,124,31,64,31,124,31,124,30,53,31,75,31,226,31,239,31,231,31,63,31,63,30,165,31,52,31,205,31,101,31,34,31,39,31,39,30,246,31,246,30,246,29,157,31,18,31,111,31,135,31,18,31,64,31,64,30,65,31,67,31,169,31,115,31,5,31,95,31,19,31,200,31,26,31,164,31,164,30,42,31,241,31,207,31,239,31,53,31,119,31,214,31,214,30,173,31,155,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
