-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 930;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (99,0,235,0,0,0,0,0,106,0,74,0,0,0,173,0,167,0,111,0,0,0,129,0,218,0,94,0,243,0,106,0,223,0,0,0,0,0,129,0,198,0,0,0,0,0,106,0,215,0,0,0,94,0,82,0,244,0,0,0,125,0,132,0,11,0,0,0,136,0,43,0,0,0,0,0,219,0,166,0,108,0,111,0,137,0,0,0,164,0,99,0,0,0,87,0,200,0,238,0,0,0,0,0,0,0,99,0,0,0,181,0,125,0,70,0,236,0,46,0,204,0,0,0,181,0,211,0,7,0,251,0,0,0,17,0,173,0,101,0,80,0,121,0,145,0,109,0,230,0,146,0,40,0,183,0,174,0,239,0,163,0,224,0,0,0,159,0,0,0,84,0,0,0,239,0,244,0,0,0,185,0,1,0,3,0,157,0,9,0,93,0,203,0,36,0,40,0,101,0,129,0,176,0,103,0,0,0,238,0,109,0,114,0,0,0,58,0,145,0,18,0,131,0,79,0,40,0,79,0,69,0,0,0,169,0,135,0,106,0,127,0,111,0,151,0,231,0,67,0,0,0,114,0,221,0,173,0,109,0,0,0,192,0,225,0,0,0,104,0,32,0,139,0,59,0,0,0,150,0,5,0,150,0,0,0,34,0,0,0,0,0,0,0,168,0,0,0,6,0,7,0,62,0,132,0,0,0,88,0,13,0,125,0,230,0,0,0,0,0,0,0,0,0,209,0,66,0,0,0,13,0,29,0,123,0,0,0,29,0,194,0,0,0,71,0,183,0,137,0,126,0,177,0,123,0,48,0,179,0,5,0,73,0,239,0,0,0,190,0,143,0,0,0,0,0,192,0,0,0,233,0,188,0,217,0,20,0,219,0,190,0,169,0,87,0,149,0,175,0,205,0,119,0,185,0,61,0,0,0,159,0,254,0,18,0,101,0,133,0,155,0,236,0,222,0,0,0,126,0,253,0,252,0,0,0,23,0,253,0,15,0,253,0,57,0,217,0,43,0,231,0,185,0,242,0,16,0,89,0,36,0,0,0,0,0,111,0,71,0,185,0,192,0,0,0,47,0,221,0,0,0,223,0,181,0,165,0,193,0,101,0,207,0,0,0,22,0,30,0,116,0,90,0,33,0,0,0,31,0,0,0,107,0,16,0,35,0,199,0,252,0,0,0,4,0,195,0,0,0,38,0,136,0,110,0,243,0,0,0,42,0,129,0,189,0,12,0,68,0,2,0,0,0,186,0,249,0,0,0,189,0,166,0,0,0,194,0,0,0,87,0,90,0,214,0,243,0,0,0,0,0,5,0,71,0,203,0,146,0,74,0,235,0,226,0,0,0,141,0,0,0,168,0,123,0,73,0,84,0,0,0,0,0,23,0,255,0,166,0,253,0,233,0,244,0,0,0,142,0,49,0,0,0,5,0,69,0,4,0,248,0,169,0,17,0,0,0,0,0,0,0,0,0,231,0,0,0,0,0,87,0,172,0,39,0,24,0,41,0,6,0,209,0,0,0,244,0,131,0,245,0,155,0,21,0,109,0,69,0,173,0,115,0,0,0,238,0,62,0,198,0,62,0,104,0,0,0,53,0,84,0,201,0,61,0,214,0,179,0,252,0,228,0,167,0,222,0,0,0,133,0,155,0,44,0,43,0,180,0,86,0,0,0,234,0,88,0,188,0,0,0,98,0,233,0,102,0,50,0,0,0,208,0,250,0,0,0,202,0,123,0,0,0,251,0,90,0,0,0,156,0,55,0,123,0,251,0,160,0,41,0,234,0,160,0,173,0,33,0,9,0,60,0,156,0,244,0,248,0,0,0,139,0,161,0,237,0,21,0,222,0,62,0,97,0,81,0,126,0,125,0,249,0,121,0,27,0,69,0,235,0,110,0,228,0,52,0,157,0,0,0,0,0,0,0,99,0,0,0,0,0,193,0,249,0,97,0,0,0,90,0,200,0,94,0,30,0,72,0,129,0,105,0,103,0,164,0,140,0,173,0,22,0,16,0,135,0,0,0,80,0,0,0,0,0,160,0,54,0,0,0,141,0,105,0,249,0,0,0,106,0,0,0,244,0,146,0,155,0,17,0,169,0,0,0,45,0,143,0,0,0,0,0,228,0,145,0,0,0,104,0,177,0,0,0,54,0,125,0,147,0,135,0,74,0,0,0,71,0,205,0,72,0,200,0,0,0,115,0,160,0,122,0,167,0,165,0,184,0,59,0,0,0,31,0,0,0,79,0,137,0,90,0,239,0,39,0,248,0,76,0,91,0,197,0,214,0,233,0,166,0,143,0,82,0,0,0,0,0,137,0,232,0,11,0,46,0,245,0,149,0,83,0,42,0,151,0,89,0,250,0,0,0,0,0,43,0,202,0,14,0,0,0,173,0,205,0,56,0,17,0,50,0,30,0,177,0,193,0,244,0,92,0,122,0,244,0,245,0,134,0,0,0,135,0,172,0,91,0,0,0,0,0,188,0,0,0,166,0,141,0,67,0,166,0,194,0,0,0,235,0,138,0,161,0,14,0,80,0,0,0,217,0,41,0,47,0,197,0,227,0,131,0,86,0,223,0,22,0,241,0,60,0,127,0,152,0,121,0,56,0,206,0,1,0,87,0,67,0,42,0,0,0,0,0,0,0,0,0,27,0,102,0,128,0,4,0,192,0,94,0,248,0,178,0,190,0,142,0,96,0,104,0,0,0,29,0,0,0,165,0,255,0,0,0,52,0,67,0,178,0,103,0,0,0,0,0,0,0,208,0,86,0,196,0,10,0,111,0,1,0,132,0,0,0,0,0,27,0,88,0,189,0,136,0,86,0,10,0,188,0,188,0,226,0,0,0,221,0,215,0,38,0,0,0,182,0,79,0,0,0,239,0,180,0,39,0,30,0,108,0,230,0,0,0,136,0,148,0,242,0,0,0,59,0,243,0,5,0,120,0,156,0,0,0,122,0,16,0,0,0,89,0,58,0,0,0,122,0,0,0,0,0,180,0,0,0,129,0,40,0,255,0,41,0,0,0,55,0,83,0,21,0,0,0,0,0,133,0,83,0,234,0,114,0,43,0,182,0,75,0,0,0,252,0,0,0,61,0,32,0,146,0,227,0,218,0,121,0,124,0,0,0,230,0,179,0,102,0,60,0,96,0,0,0,0,0,127,0,89,0,207,0,0,0,0,0,59,0,168,0,235,0,58,0,45,0,198,0,254,0,0,0,0,0,0,0,15,0,0,0,22,0,148,0,95,0,17,0,51,0,0,0,47,0,226,0,139,0,110,0,191,0,0,0,80,0,0,0,0,0,130,0,110,0,153,0,80,0,0,0,129,0,71,0,43,0,0,0,0,0,251,0,224,0,0,0,187,0,0,0,51,0,201,0,126,0,0,0,6,0,0,0,239,0,76,0,24,0,7,0,158,0,105,0,159,0,126,0,97,0,198,0,16,0,81,0,195,0,57,0,189,0,207,0,17,0,149,0,0,0,69,0,158,0,0,0,194,0,237,0,152,0,0,0,26,0,142,0,226,0,0,0,157,0,118,0,143,0,188,0,0,0,0,0,123,0,0,0,0,0,219,0,255,0,167,0,22,0,80,0,241,0,81,0,92,0,18,0,99,0,120,0,207,0,0,0,0,0,141,0,0,0,0,0,0,0,184,0,114,0,195,0,247,0,0,0,253,0,239,0,225,0,138,0,0,0,56,0,0,0,0,0,47,0,0,0,198,0,0,0,78,0,0,0,194,0,0,0,0,0,10,0,0,0,127,0,15,0,65,0,106,0,0,0,0,0,35,0,199,0,209,0,165,0,0,0,26,0,0,0,18,0,108,0,0,0,0,0,124,0,0,0,164,0,230,0,16,0,153,0,140,0,171,0,60,0,243,0,147,0,0,0,74,0,150,0,100,0,187,0,77,0,104,0,0,0,0,0,0,0,20,0,32,0,30,0,205,0,115,0,217,0,138,0,248,0,253,0,179,0,40,0,214,0,112,0,41,0,82,0,0,0,11,0,174,0,0,0,0,0,74,0,88,0,56,0,56,0,204,0,113,0,241,0,10,0,51,0,21,0,0,0,223,0,192,0,33,0,57,0,158,0,166,0,58,0,104,0,125,0,158,0,116,0,149,0,51,0,132,0,22,0,237,0,128,0,0,0,185,0,147,0,55,0,127,0,0,0);
signal scenario_full  : scenario_type := (99,31,235,31,235,30,235,29,106,31,74,31,74,30,173,31,167,31,111,31,111,30,129,31,218,31,94,31,243,31,106,31,223,31,223,30,223,29,129,31,198,31,198,30,198,29,106,31,215,31,215,30,94,31,82,31,244,31,244,30,125,31,132,31,11,31,11,30,136,31,43,31,43,30,43,29,219,31,166,31,108,31,111,31,137,31,137,30,164,31,99,31,99,30,87,31,200,31,238,31,238,30,238,29,238,28,99,31,99,30,181,31,125,31,70,31,236,31,46,31,204,31,204,30,181,31,211,31,7,31,251,31,251,30,17,31,173,31,101,31,80,31,121,31,145,31,109,31,230,31,146,31,40,31,183,31,174,31,239,31,163,31,224,31,224,30,159,31,159,30,84,31,84,30,239,31,244,31,244,30,185,31,1,31,3,31,157,31,9,31,93,31,203,31,36,31,40,31,101,31,129,31,176,31,103,31,103,30,238,31,109,31,114,31,114,30,58,31,145,31,18,31,131,31,79,31,40,31,79,31,69,31,69,30,169,31,135,31,106,31,127,31,111,31,151,31,231,31,67,31,67,30,114,31,221,31,173,31,109,31,109,30,192,31,225,31,225,30,104,31,32,31,139,31,59,31,59,30,150,31,5,31,150,31,150,30,34,31,34,30,34,29,34,28,168,31,168,30,6,31,7,31,62,31,132,31,132,30,88,31,13,31,125,31,230,31,230,30,230,29,230,28,230,27,209,31,66,31,66,30,13,31,29,31,123,31,123,30,29,31,194,31,194,30,71,31,183,31,137,31,126,31,177,31,123,31,48,31,179,31,5,31,73,31,239,31,239,30,190,31,143,31,143,30,143,29,192,31,192,30,233,31,188,31,217,31,20,31,219,31,190,31,169,31,87,31,149,31,175,31,205,31,119,31,185,31,61,31,61,30,159,31,254,31,18,31,101,31,133,31,155,31,236,31,222,31,222,30,126,31,253,31,252,31,252,30,23,31,253,31,15,31,253,31,57,31,217,31,43,31,231,31,185,31,242,31,16,31,89,31,36,31,36,30,36,29,111,31,71,31,185,31,192,31,192,30,47,31,221,31,221,30,223,31,181,31,165,31,193,31,101,31,207,31,207,30,22,31,30,31,116,31,90,31,33,31,33,30,31,31,31,30,107,31,16,31,35,31,199,31,252,31,252,30,4,31,195,31,195,30,38,31,136,31,110,31,243,31,243,30,42,31,129,31,189,31,12,31,68,31,2,31,2,30,186,31,249,31,249,30,189,31,166,31,166,30,194,31,194,30,87,31,90,31,214,31,243,31,243,30,243,29,5,31,71,31,203,31,146,31,74,31,235,31,226,31,226,30,141,31,141,30,168,31,123,31,73,31,84,31,84,30,84,29,23,31,255,31,166,31,253,31,233,31,244,31,244,30,142,31,49,31,49,30,5,31,69,31,4,31,248,31,169,31,17,31,17,30,17,29,17,28,17,27,231,31,231,30,231,29,87,31,172,31,39,31,24,31,41,31,6,31,209,31,209,30,244,31,131,31,245,31,155,31,21,31,109,31,69,31,173,31,115,31,115,30,238,31,62,31,198,31,62,31,104,31,104,30,53,31,84,31,201,31,61,31,214,31,179,31,252,31,228,31,167,31,222,31,222,30,133,31,155,31,44,31,43,31,180,31,86,31,86,30,234,31,88,31,188,31,188,30,98,31,233,31,102,31,50,31,50,30,208,31,250,31,250,30,202,31,123,31,123,30,251,31,90,31,90,30,156,31,55,31,123,31,251,31,160,31,41,31,234,31,160,31,173,31,33,31,9,31,60,31,156,31,244,31,248,31,248,30,139,31,161,31,237,31,21,31,222,31,62,31,97,31,81,31,126,31,125,31,249,31,121,31,27,31,69,31,235,31,110,31,228,31,52,31,157,31,157,30,157,29,157,28,99,31,99,30,99,29,193,31,249,31,97,31,97,30,90,31,200,31,94,31,30,31,72,31,129,31,105,31,103,31,164,31,140,31,173,31,22,31,16,31,135,31,135,30,80,31,80,30,80,29,160,31,54,31,54,30,141,31,105,31,249,31,249,30,106,31,106,30,244,31,146,31,155,31,17,31,169,31,169,30,45,31,143,31,143,30,143,29,228,31,145,31,145,30,104,31,177,31,177,30,54,31,125,31,147,31,135,31,74,31,74,30,71,31,205,31,72,31,200,31,200,30,115,31,160,31,122,31,167,31,165,31,184,31,59,31,59,30,31,31,31,30,79,31,137,31,90,31,239,31,39,31,248,31,76,31,91,31,197,31,214,31,233,31,166,31,143,31,82,31,82,30,82,29,137,31,232,31,11,31,46,31,245,31,149,31,83,31,42,31,151,31,89,31,250,31,250,30,250,29,43,31,202,31,14,31,14,30,173,31,205,31,56,31,17,31,50,31,30,31,177,31,193,31,244,31,92,31,122,31,244,31,245,31,134,31,134,30,135,31,172,31,91,31,91,30,91,29,188,31,188,30,166,31,141,31,67,31,166,31,194,31,194,30,235,31,138,31,161,31,14,31,80,31,80,30,217,31,41,31,47,31,197,31,227,31,131,31,86,31,223,31,22,31,241,31,60,31,127,31,152,31,121,31,56,31,206,31,1,31,87,31,67,31,42,31,42,30,42,29,42,28,42,27,27,31,102,31,128,31,4,31,192,31,94,31,248,31,178,31,190,31,142,31,96,31,104,31,104,30,29,31,29,30,165,31,255,31,255,30,52,31,67,31,178,31,103,31,103,30,103,29,103,28,208,31,86,31,196,31,10,31,111,31,1,31,132,31,132,30,132,29,27,31,88,31,189,31,136,31,86,31,10,31,188,31,188,31,226,31,226,30,221,31,215,31,38,31,38,30,182,31,79,31,79,30,239,31,180,31,39,31,30,31,108,31,230,31,230,30,136,31,148,31,242,31,242,30,59,31,243,31,5,31,120,31,156,31,156,30,122,31,16,31,16,30,89,31,58,31,58,30,122,31,122,30,122,29,180,31,180,30,129,31,40,31,255,31,41,31,41,30,55,31,83,31,21,31,21,30,21,29,133,31,83,31,234,31,114,31,43,31,182,31,75,31,75,30,252,31,252,30,61,31,32,31,146,31,227,31,218,31,121,31,124,31,124,30,230,31,179,31,102,31,60,31,96,31,96,30,96,29,127,31,89,31,207,31,207,30,207,29,59,31,168,31,235,31,58,31,45,31,198,31,254,31,254,30,254,29,254,28,15,31,15,30,22,31,148,31,95,31,17,31,51,31,51,30,47,31,226,31,139,31,110,31,191,31,191,30,80,31,80,30,80,29,130,31,110,31,153,31,80,31,80,30,129,31,71,31,43,31,43,30,43,29,251,31,224,31,224,30,187,31,187,30,51,31,201,31,126,31,126,30,6,31,6,30,239,31,76,31,24,31,7,31,158,31,105,31,159,31,126,31,97,31,198,31,16,31,81,31,195,31,57,31,189,31,207,31,17,31,149,31,149,30,69,31,158,31,158,30,194,31,237,31,152,31,152,30,26,31,142,31,226,31,226,30,157,31,118,31,143,31,188,31,188,30,188,29,123,31,123,30,123,29,219,31,255,31,167,31,22,31,80,31,241,31,81,31,92,31,18,31,99,31,120,31,207,31,207,30,207,29,141,31,141,30,141,29,141,28,184,31,114,31,195,31,247,31,247,30,253,31,239,31,225,31,138,31,138,30,56,31,56,30,56,29,47,31,47,30,198,31,198,30,78,31,78,30,194,31,194,30,194,29,10,31,10,30,127,31,15,31,65,31,106,31,106,30,106,29,35,31,199,31,209,31,165,31,165,30,26,31,26,30,18,31,108,31,108,30,108,29,124,31,124,30,164,31,230,31,16,31,153,31,140,31,171,31,60,31,243,31,147,31,147,30,74,31,150,31,100,31,187,31,77,31,104,31,104,30,104,29,104,28,20,31,32,31,30,31,205,31,115,31,217,31,138,31,248,31,253,31,179,31,40,31,214,31,112,31,41,31,82,31,82,30,11,31,174,31,174,30,174,29,74,31,88,31,56,31,56,31,204,31,113,31,241,31,10,31,51,31,21,31,21,30,223,31,192,31,33,31,57,31,158,31,166,31,58,31,104,31,125,31,158,31,116,31,149,31,51,31,132,31,22,31,237,31,128,31,128,30,185,31,147,31,55,31,127,31,127,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
