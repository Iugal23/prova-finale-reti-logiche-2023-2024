-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_590 is
end project_tb_590;

architecture project_tb_arch_590 of project_tb_590 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 538;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (18,0,91,0,255,0,0,0,219,0,5,0,61,0,7,0,218,0,176,0,187,0,142,0,237,0,42,0,169,0,0,0,168,0,174,0,0,0,32,0,162,0,88,0,153,0,71,0,0,0,0,0,0,0,182,0,122,0,53,0,82,0,41,0,212,0,156,0,148,0,0,0,0,0,220,0,200,0,52,0,53,0,0,0,136,0,249,0,1,0,0,0,255,0,194,0,49,0,189,0,174,0,233,0,235,0,0,0,228,0,254,0,60,0,195,0,0,0,0,0,38,0,89,0,148,0,193,0,224,0,223,0,0,0,217,0,190,0,244,0,97,0,119,0,152,0,0,0,70,0,0,0,0,0,190,0,149,0,0,0,51,0,12,0,10,0,113,0,136,0,0,0,54,0,38,0,48,0,133,0,94,0,215,0,188,0,86,0,0,0,0,0,14,0,170,0,0,0,0,0,133,0,50,0,0,0,144,0,61,0,255,0,0,0,11,0,0,0,17,0,84,0,0,0,42,0,0,0,106,0,226,0,0,0,0,0,48,0,98,0,79,0,207,0,11,0,162,0,165,0,0,0,173,0,120,0,95,0,195,0,176,0,130,0,252,0,73,0,0,0,115,0,53,0,53,0,166,0,62,0,175,0,250,0,181,0,22,0,103,0,248,0,73,0,155,0,124,0,33,0,105,0,157,0,61,0,176,0,84,0,70,0,0,0,186,0,0,0,87,0,0,0,0,0,0,0,168,0,107,0,0,0,131,0,13,0,191,0,164,0,104,0,44,0,170,0,0,0,3,0,151,0,232,0,6,0,179,0,0,0,80,0,108,0,200,0,12,0,79,0,36,0,0,0,35,0,220,0,0,0,158,0,227,0,122,0,245,0,245,0,163,0,138,0,74,0,37,0,204,0,13,0,156,0,38,0,116,0,72,0,79,0,201,0,26,0,252,0,254,0,32,0,224,0,103,0,0,0,216,0,96,0,0,0,0,0,25,0,0,0,126,0,28,0,215,0,177,0,29,0,46,0,0,0,95,0,230,0,69,0,80,0,96,0,62,0,0,0,202,0,0,0,238,0,0,0,124,0,189,0,164,0,53,0,55,0,233,0,193,0,123,0,92,0,16,0,145,0,128,0,81,0,88,0,112,0,205,0,99,0,145,0,206,0,244,0,143,0,229,0,170,0,247,0,222,0,189,0,173,0,88,0,24,0,167,0,0,0,165,0,29,0,232,0,99,0,146,0,171,0,200,0,0,0,143,0,0,0,128,0,122,0,24,0,62,0,0,0,17,0,198,0,0,0,12,0,135,0,114,0,7,0,101,0,223,0,92,0,114,0,128,0,59,0,56,0,225,0,0,0,171,0,0,0,155,0,0,0,108,0,44,0,98,0,0,0,7,0,114,0,91,0,70,0,0,0,141,0,0,0,0,0,133,0,0,0,115,0,201,0,11,0,172,0,164,0,41,0,236,0,127,0,73,0,108,0,127,0,94,0,31,0,240,0,208,0,135,0,0,0,58,0,0,0,176,0,0,0,58,0,33,0,180,0,0,0,26,0,67,0,0,0,95,0,160,0,249,0,194,0,23,0,0,0,14,0,152,0,199,0,0,0,30,0,200,0,111,0,190,0,70,0,86,0,38,0,0,0,49,0,72,0,0,0,39,0,90,0,247,0,164,0,240,0,218,0,0,0,1,0,200,0,153,0,37,0,0,0,0,0,0,0,188,0,92,0,77,0,158,0,255,0,25,0,0,0,168,0,223,0,0,0,0,0,149,0,220,0,0,0,185,0,8,0,2,0,75,0,0,0,236,0,132,0,138,0,147,0,168,0,0,0,45,0,239,0,221,0,227,0,29,0,189,0,0,0,89,0,29,0,254,0,0,0,184,0,214,0,131,0,6,0,185,0,0,0,50,0,230,0,159,0,123,0,131,0,0,0,8,0,44,0,0,0,43,0,228,0,0,0,124,0,138,0,0,0,73,0,143,0,122,0,236,0,162,0,146,0,86,0,0,0,219,0,0,0,0,0,64,0,207,0,43,0,228,0,213,0,197,0,176,0,81,0,186,0,0,0,233,0,59,0,120,0,124,0,0,0,0,0,79,0,235,0,29,0,93,0,0,0,119,0,0,0,147,0,57,0,0,0,235,0,206,0,57,0,163,0,206,0,0,0,0,0,100,0,162,0,228,0,162,0,42,0,0,0,60,0,203,0,224,0,0,0,117,0,0,0,213,0,56,0,54,0,23,0,58,0,78,0,0,0,34,0,14,0,172,0,133,0,213,0,121,0,0,0,84,0,0,0,146,0,171,0,20,0,205,0,250,0,125,0,230,0,185,0,147,0,183,0,101,0,152,0,0,0,92,0,207,0,19,0,0,0,232,0,230,0,140,0,12,0,0,0,64,0,0,0,0,0,94,0,0,0,251,0);
signal scenario_full  : scenario_type := (18,31,91,31,255,31,255,30,219,31,5,31,61,31,7,31,218,31,176,31,187,31,142,31,237,31,42,31,169,31,169,30,168,31,174,31,174,30,32,31,162,31,88,31,153,31,71,31,71,30,71,29,71,28,182,31,122,31,53,31,82,31,41,31,212,31,156,31,148,31,148,30,148,29,220,31,200,31,52,31,53,31,53,30,136,31,249,31,1,31,1,30,255,31,194,31,49,31,189,31,174,31,233,31,235,31,235,30,228,31,254,31,60,31,195,31,195,30,195,29,38,31,89,31,148,31,193,31,224,31,223,31,223,30,217,31,190,31,244,31,97,31,119,31,152,31,152,30,70,31,70,30,70,29,190,31,149,31,149,30,51,31,12,31,10,31,113,31,136,31,136,30,54,31,38,31,48,31,133,31,94,31,215,31,188,31,86,31,86,30,86,29,14,31,170,31,170,30,170,29,133,31,50,31,50,30,144,31,61,31,255,31,255,30,11,31,11,30,17,31,84,31,84,30,42,31,42,30,106,31,226,31,226,30,226,29,48,31,98,31,79,31,207,31,11,31,162,31,165,31,165,30,173,31,120,31,95,31,195,31,176,31,130,31,252,31,73,31,73,30,115,31,53,31,53,31,166,31,62,31,175,31,250,31,181,31,22,31,103,31,248,31,73,31,155,31,124,31,33,31,105,31,157,31,61,31,176,31,84,31,70,31,70,30,186,31,186,30,87,31,87,30,87,29,87,28,168,31,107,31,107,30,131,31,13,31,191,31,164,31,104,31,44,31,170,31,170,30,3,31,151,31,232,31,6,31,179,31,179,30,80,31,108,31,200,31,12,31,79,31,36,31,36,30,35,31,220,31,220,30,158,31,227,31,122,31,245,31,245,31,163,31,138,31,74,31,37,31,204,31,13,31,156,31,38,31,116,31,72,31,79,31,201,31,26,31,252,31,254,31,32,31,224,31,103,31,103,30,216,31,96,31,96,30,96,29,25,31,25,30,126,31,28,31,215,31,177,31,29,31,46,31,46,30,95,31,230,31,69,31,80,31,96,31,62,31,62,30,202,31,202,30,238,31,238,30,124,31,189,31,164,31,53,31,55,31,233,31,193,31,123,31,92,31,16,31,145,31,128,31,81,31,88,31,112,31,205,31,99,31,145,31,206,31,244,31,143,31,229,31,170,31,247,31,222,31,189,31,173,31,88,31,24,31,167,31,167,30,165,31,29,31,232,31,99,31,146,31,171,31,200,31,200,30,143,31,143,30,128,31,122,31,24,31,62,31,62,30,17,31,198,31,198,30,12,31,135,31,114,31,7,31,101,31,223,31,92,31,114,31,128,31,59,31,56,31,225,31,225,30,171,31,171,30,155,31,155,30,108,31,44,31,98,31,98,30,7,31,114,31,91,31,70,31,70,30,141,31,141,30,141,29,133,31,133,30,115,31,201,31,11,31,172,31,164,31,41,31,236,31,127,31,73,31,108,31,127,31,94,31,31,31,240,31,208,31,135,31,135,30,58,31,58,30,176,31,176,30,58,31,33,31,180,31,180,30,26,31,67,31,67,30,95,31,160,31,249,31,194,31,23,31,23,30,14,31,152,31,199,31,199,30,30,31,200,31,111,31,190,31,70,31,86,31,38,31,38,30,49,31,72,31,72,30,39,31,90,31,247,31,164,31,240,31,218,31,218,30,1,31,200,31,153,31,37,31,37,30,37,29,37,28,188,31,92,31,77,31,158,31,255,31,25,31,25,30,168,31,223,31,223,30,223,29,149,31,220,31,220,30,185,31,8,31,2,31,75,31,75,30,236,31,132,31,138,31,147,31,168,31,168,30,45,31,239,31,221,31,227,31,29,31,189,31,189,30,89,31,29,31,254,31,254,30,184,31,214,31,131,31,6,31,185,31,185,30,50,31,230,31,159,31,123,31,131,31,131,30,8,31,44,31,44,30,43,31,228,31,228,30,124,31,138,31,138,30,73,31,143,31,122,31,236,31,162,31,146,31,86,31,86,30,219,31,219,30,219,29,64,31,207,31,43,31,228,31,213,31,197,31,176,31,81,31,186,31,186,30,233,31,59,31,120,31,124,31,124,30,124,29,79,31,235,31,29,31,93,31,93,30,119,31,119,30,147,31,57,31,57,30,235,31,206,31,57,31,163,31,206,31,206,30,206,29,100,31,162,31,228,31,162,31,42,31,42,30,60,31,203,31,224,31,224,30,117,31,117,30,213,31,56,31,54,31,23,31,58,31,78,31,78,30,34,31,14,31,172,31,133,31,213,31,121,31,121,30,84,31,84,30,146,31,171,31,20,31,205,31,250,31,125,31,230,31,185,31,147,31,183,31,101,31,152,31,152,30,92,31,207,31,19,31,19,30,232,31,230,31,140,31,12,31,12,30,64,31,64,30,64,29,94,31,94,30,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
