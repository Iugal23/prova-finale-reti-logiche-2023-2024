-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 765;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (244,0,158,0,20,0,0,0,96,0,0,0,48,0,91,0,246,0,48,0,85,0,65,0,190,0,0,0,252,0,118,0,0,0,232,0,0,0,108,0,130,0,215,0,2,0,248,0,2,0,0,0,71,0,184,0,188,0,96,0,205,0,41,0,0,0,38,0,0,0,6,0,211,0,238,0,255,0,136,0,0,0,0,0,36,0,215,0,0,0,154,0,0,0,54,0,0,0,69,0,0,0,79,0,150,0,212,0,84,0,24,0,236,0,230,0,0,0,201,0,0,0,0,0,61,0,166,0,232,0,0,0,246,0,4,0,164,0,0,0,154,0,60,0,206,0,225,0,0,0,177,0,21,0,112,0,118,0,123,0,175,0,143,0,0,0,182,0,0,0,0,0,167,0,0,0,43,0,102,0,101,0,112,0,0,0,61,0,158,0,201,0,0,0,148,0,166,0,207,0,0,0,2,0,157,0,173,0,137,0,90,0,189,0,0,0,0,0,73,0,11,0,51,0,30,0,227,0,45,0,112,0,0,0,83,0,52,0,57,0,244,0,165,0,96,0,121,0,126,0,15,0,28,0,0,0,36,0,246,0,0,0,201,0,68,0,106,0,203,0,63,0,55,0,149,0,141,0,123,0,0,0,27,0,32,0,229,0,0,0,249,0,171,0,58,0,196,0,64,0,0,0,117,0,224,0,241,0,0,0,0,0,153,0,205,0,230,0,24,0,46,0,154,0,161,0,237,0,57,0,225,0,10,0,37,0,98,0,204,0,0,0,0,0,0,0,126,0,0,0,59,0,59,0,242,0,212,0,75,0,87,0,60,0,21,0,0,0,221,0,55,0,174,0,46,0,248,0,0,0,164,0,0,0,211,0,147,0,0,0,41,0,0,0,246,0,48,0,0,0,7,0,141,0,19,0,25,0,0,0,215,0,0,0,111,0,251,0,67,0,131,0,110,0,165,0,0,0,0,0,221,0,81,0,49,0,5,0,80,0,0,0,153,0,111,0,0,0,182,0,0,0,169,0,3,0,0,0,73,0,25,0,146,0,47,0,0,0,137,0,0,0,247,0,23,0,215,0,110,0,0,0,127,0,0,0,17,0,218,0,0,0,153,0,160,0,35,0,53,0,77,0,17,0,177,0,0,0,48,0,213,0,182,0,181,0,40,0,0,0,0,0,123,0,0,0,205,0,28,0,126,0,88,0,238,0,94,0,94,0,211,0,214,0,137,0,189,0,191,0,17,0,72,0,38,0,130,0,0,0,0,0,153,0,251,0,90,0,183,0,237,0,105,0,242,0,0,0,0,0,70,0,25,0,120,0,0,0,20,0,85,0,66,0,244,0,19,0,0,0,90,0,0,0,115,0,19,0,108,0,155,0,58,0,0,0,152,0,0,0,39,0,162,0,53,0,0,0,193,0,48,0,0,0,52,0,51,0,92,0,233,0,28,0,15,0,86,0,167,0,126,0,143,0,0,0,121,0,52,0,114,0,55,0,157,0,50,0,123,0,27,0,46,0,182,0,0,0,32,0,216,0,100,0,0,0,25,0,201,0,250,0,145,0,147,0,33,0,167,0,225,0,44,0,131,0,0,0,132,0,126,0,95,0,46,0,81,0,108,0,0,0,93,0,0,0,218,0,255,0,0,0,0,0,193,0,109,0,0,0,254,0,23,0,55,0,254,0,0,0,101,0,35,0,216,0,220,0,0,0,71,0,53,0,0,0,27,0,154,0,177,0,252,0,211,0,245,0,255,0,0,0,128,0,243,0,252,0,158,0,161,0,0,0,97,0,167,0,108,0,0,0,85,0,213,0,202,0,0,0,190,0,253,0,58,0,68,0,54,0,90,0,226,0,37,0,33,0,55,0,0,0,0,0,159,0,0,0,4,0,89,0,144,0,5,0,139,0,22,0,125,0,0,0,216,0,206,0,39,0,228,0,34,0,73,0,226,0,108,0,144,0,130,0,43,0,73,0,199,0,0,0,114,0,123,0,32,0,127,0,245,0,0,0,125,0,35,0,0,0,140,0,241,0,0,0,30,0,0,0,56,0,152,0,0,0,139,0,228,0,234,0,228,0,249,0,0,0,111,0,231,0,84,0,129,0,0,0,120,0,151,0,187,0,0,0,114,0,155,0,101,0,35,0,121,0,211,0,180,0,229,0,252,0,185,0,240,0,188,0,50,0,203,0,168,0,117,0,59,0,58,0,171,0,244,0,0,0,0,0,108,0,0,0,0,0,118,0,163,0,210,0,235,0,0,0,219,0,227,0,119,0,184,0,0,0,59,0,46,0,136,0,214,0,120,0,220,0,76,0,0,0,43,0,226,0,162,0,148,0,105,0,250,0,144,0,193,0,145,0,80,0,0,0,26,0,94,0,252,0,222,0,35,0,27,0,0,0,152,0,177,0,68,0,244,0,0,0,117,0,0,0,177,0,80,0,0,0,0,0,174,0,196,0,0,0,64,0,125,0,0,0,146,0,0,0,0,0,89,0,213,0,162,0,87,0,161,0,99,0,220,0,177,0,0,0,113,0,162,0,25,0,138,0,48,0,225,0,0,0,0,0,126,0,114,0,88,0,90,0,173,0,205,0,103,0,219,0,101,0,0,0,3,0,140,0,0,0,150,0,0,0,0,0,0,0,22,0,0,0,0,0,107,0,148,0,123,0,0,0,64,0,0,0,6,0,157,0,232,0,178,0,54,0,149,0,139,0,116,0,184,0,210,0,57,0,190,0,49,0,84,0,99,0,17,0,76,0,24,0,167,0,89,0,74,0,126,0,42,0,62,0,89,0,107,0,0,0,232,0,4,0,167,0,12,0,177,0,0,0,246,0,0,0,237,0,83,0,219,0,0,0,150,0,102,0,0,0,100,0,90,0,143,0,107,0,218,0,79,0,238,0,144,0,245,0,141,0,46,0,94,0,0,0,254,0,212,0,77,0,1,0,228,0,0,0,10,0,139,0,52,0,22,0,255,0,26,0,207,0,151,0,112,0,153,0,0,0,27,0,0,0,167,0,164,0,0,0,0,0,242,0,190,0,159,0,132,0,0,0,169,0,198,0,252,0,13,0,0,0,113,0,97,0,35,0,130,0,127,0,80,0,82,0,24,0,171,0,36,0,40,0,230,0,0,0,168,0,0,0,197,0,53,0,0,0,193,0,174,0,58,0,232,0,34,0,0,0,30,0,39,0,0,0,51,0,0,0,119,0,199,0,0,0,72,0,155,0,0,0,215,0,128,0,125,0,239,0,227,0,37,0,133,0,16,0,245,0,0,0,0,0,94,0,27,0,141,0,186,0,0,0,180,0,200,0,5,0,148,0,215,0,244,0,100,0,108,0,0,0,233,0,215,0,255,0,0,0,134,0,224,0,242,0,63,0,235,0,121,0,175,0,216,0,24,0,0,0,20,0,206,0,237,0,47,0,118,0,49,0);
signal scenario_full  : scenario_type := (244,31,158,31,20,31,20,30,96,31,96,30,48,31,91,31,246,31,48,31,85,31,65,31,190,31,190,30,252,31,118,31,118,30,232,31,232,30,108,31,130,31,215,31,2,31,248,31,2,31,2,30,71,31,184,31,188,31,96,31,205,31,41,31,41,30,38,31,38,30,6,31,211,31,238,31,255,31,136,31,136,30,136,29,36,31,215,31,215,30,154,31,154,30,54,31,54,30,69,31,69,30,79,31,150,31,212,31,84,31,24,31,236,31,230,31,230,30,201,31,201,30,201,29,61,31,166,31,232,31,232,30,246,31,4,31,164,31,164,30,154,31,60,31,206,31,225,31,225,30,177,31,21,31,112,31,118,31,123,31,175,31,143,31,143,30,182,31,182,30,182,29,167,31,167,30,43,31,102,31,101,31,112,31,112,30,61,31,158,31,201,31,201,30,148,31,166,31,207,31,207,30,2,31,157,31,173,31,137,31,90,31,189,31,189,30,189,29,73,31,11,31,51,31,30,31,227,31,45,31,112,31,112,30,83,31,52,31,57,31,244,31,165,31,96,31,121,31,126,31,15,31,28,31,28,30,36,31,246,31,246,30,201,31,68,31,106,31,203,31,63,31,55,31,149,31,141,31,123,31,123,30,27,31,32,31,229,31,229,30,249,31,171,31,58,31,196,31,64,31,64,30,117,31,224,31,241,31,241,30,241,29,153,31,205,31,230,31,24,31,46,31,154,31,161,31,237,31,57,31,225,31,10,31,37,31,98,31,204,31,204,30,204,29,204,28,126,31,126,30,59,31,59,31,242,31,212,31,75,31,87,31,60,31,21,31,21,30,221,31,55,31,174,31,46,31,248,31,248,30,164,31,164,30,211,31,147,31,147,30,41,31,41,30,246,31,48,31,48,30,7,31,141,31,19,31,25,31,25,30,215,31,215,30,111,31,251,31,67,31,131,31,110,31,165,31,165,30,165,29,221,31,81,31,49,31,5,31,80,31,80,30,153,31,111,31,111,30,182,31,182,30,169,31,3,31,3,30,73,31,25,31,146,31,47,31,47,30,137,31,137,30,247,31,23,31,215,31,110,31,110,30,127,31,127,30,17,31,218,31,218,30,153,31,160,31,35,31,53,31,77,31,17,31,177,31,177,30,48,31,213,31,182,31,181,31,40,31,40,30,40,29,123,31,123,30,205,31,28,31,126,31,88,31,238,31,94,31,94,31,211,31,214,31,137,31,189,31,191,31,17,31,72,31,38,31,130,31,130,30,130,29,153,31,251,31,90,31,183,31,237,31,105,31,242,31,242,30,242,29,70,31,25,31,120,31,120,30,20,31,85,31,66,31,244,31,19,31,19,30,90,31,90,30,115,31,19,31,108,31,155,31,58,31,58,30,152,31,152,30,39,31,162,31,53,31,53,30,193,31,48,31,48,30,52,31,51,31,92,31,233,31,28,31,15,31,86,31,167,31,126,31,143,31,143,30,121,31,52,31,114,31,55,31,157,31,50,31,123,31,27,31,46,31,182,31,182,30,32,31,216,31,100,31,100,30,25,31,201,31,250,31,145,31,147,31,33,31,167,31,225,31,44,31,131,31,131,30,132,31,126,31,95,31,46,31,81,31,108,31,108,30,93,31,93,30,218,31,255,31,255,30,255,29,193,31,109,31,109,30,254,31,23,31,55,31,254,31,254,30,101,31,35,31,216,31,220,31,220,30,71,31,53,31,53,30,27,31,154,31,177,31,252,31,211,31,245,31,255,31,255,30,128,31,243,31,252,31,158,31,161,31,161,30,97,31,167,31,108,31,108,30,85,31,213,31,202,31,202,30,190,31,253,31,58,31,68,31,54,31,90,31,226,31,37,31,33,31,55,31,55,30,55,29,159,31,159,30,4,31,89,31,144,31,5,31,139,31,22,31,125,31,125,30,216,31,206,31,39,31,228,31,34,31,73,31,226,31,108,31,144,31,130,31,43,31,73,31,199,31,199,30,114,31,123,31,32,31,127,31,245,31,245,30,125,31,35,31,35,30,140,31,241,31,241,30,30,31,30,30,56,31,152,31,152,30,139,31,228,31,234,31,228,31,249,31,249,30,111,31,231,31,84,31,129,31,129,30,120,31,151,31,187,31,187,30,114,31,155,31,101,31,35,31,121,31,211,31,180,31,229,31,252,31,185,31,240,31,188,31,50,31,203,31,168,31,117,31,59,31,58,31,171,31,244,31,244,30,244,29,108,31,108,30,108,29,118,31,163,31,210,31,235,31,235,30,219,31,227,31,119,31,184,31,184,30,59,31,46,31,136,31,214,31,120,31,220,31,76,31,76,30,43,31,226,31,162,31,148,31,105,31,250,31,144,31,193,31,145,31,80,31,80,30,26,31,94,31,252,31,222,31,35,31,27,31,27,30,152,31,177,31,68,31,244,31,244,30,117,31,117,30,177,31,80,31,80,30,80,29,174,31,196,31,196,30,64,31,125,31,125,30,146,31,146,30,146,29,89,31,213,31,162,31,87,31,161,31,99,31,220,31,177,31,177,30,113,31,162,31,25,31,138,31,48,31,225,31,225,30,225,29,126,31,114,31,88,31,90,31,173,31,205,31,103,31,219,31,101,31,101,30,3,31,140,31,140,30,150,31,150,30,150,29,150,28,22,31,22,30,22,29,107,31,148,31,123,31,123,30,64,31,64,30,6,31,157,31,232,31,178,31,54,31,149,31,139,31,116,31,184,31,210,31,57,31,190,31,49,31,84,31,99,31,17,31,76,31,24,31,167,31,89,31,74,31,126,31,42,31,62,31,89,31,107,31,107,30,232,31,4,31,167,31,12,31,177,31,177,30,246,31,246,30,237,31,83,31,219,31,219,30,150,31,102,31,102,30,100,31,90,31,143,31,107,31,218,31,79,31,238,31,144,31,245,31,141,31,46,31,94,31,94,30,254,31,212,31,77,31,1,31,228,31,228,30,10,31,139,31,52,31,22,31,255,31,26,31,207,31,151,31,112,31,153,31,153,30,27,31,27,30,167,31,164,31,164,30,164,29,242,31,190,31,159,31,132,31,132,30,169,31,198,31,252,31,13,31,13,30,113,31,97,31,35,31,130,31,127,31,80,31,82,31,24,31,171,31,36,31,40,31,230,31,230,30,168,31,168,30,197,31,53,31,53,30,193,31,174,31,58,31,232,31,34,31,34,30,30,31,39,31,39,30,51,31,51,30,119,31,199,31,199,30,72,31,155,31,155,30,215,31,128,31,125,31,239,31,227,31,37,31,133,31,16,31,245,31,245,30,245,29,94,31,27,31,141,31,186,31,186,30,180,31,200,31,5,31,148,31,215,31,244,31,100,31,108,31,108,30,233,31,215,31,255,31,255,30,134,31,224,31,242,31,63,31,235,31,121,31,175,31,216,31,24,31,24,30,20,31,206,31,237,31,47,31,118,31,49,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
