-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 466;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (32,0,155,0,247,0,148,0,0,0,164,0,121,0,66,0,208,0,130,0,228,0,81,0,138,0,203,0,180,0,89,0,186,0,231,0,47,0,241,0,45,0,57,0,240,0,149,0,107,0,30,0,134,0,222,0,6,0,99,0,0,0,0,0,44,0,167,0,125,0,229,0,11,0,25,0,0,0,13,0,21,0,255,0,239,0,220,0,0,0,58,0,0,0,178,0,0,0,0,0,43,0,84,0,1,0,132,0,210,0,112,0,2,0,0,0,251,0,129,0,25,0,0,0,69,0,207,0,0,0,190,0,201,0,66,0,57,0,69,0,180,0,0,0,24,0,0,0,108,0,91,0,238,0,124,0,0,0,123,0,232,0,200,0,0,0,61,0,30,0,0,0,236,0,113,0,0,0,111,0,76,0,0,0,0,0,240,0,65,0,20,0,159,0,205,0,137,0,74,0,157,0,46,0,0,0,212,0,103,0,0,0,101,0,10,0,0,0,210,0,208,0,117,0,178,0,153,0,196,0,205,0,0,0,202,0,0,0,131,0,185,0,92,0,218,0,241,0,15,0,28,0,193,0,142,0,252,0,19,0,148,0,0,0,0,0,202,0,123,0,0,0,58,0,0,0,190,0,113,0,0,0,0,0,0,0,0,0,112,0,204,0,224,0,19,0,222,0,0,0,174,0,178,0,0,0,182,0,132,0,0,0,135,0,74,0,226,0,206,0,0,0,169,0,33,0,48,0,134,0,204,0,56,0,1,0,165,0,13,0,0,0,172,0,184,0,159,0,208,0,0,0,24,0,0,0,193,0,223,0,111,0,112,0,57,0,0,0,10,0,103,0,0,0,75,0,175,0,0,0,233,0,20,0,0,0,204,0,75,0,0,0,82,0,0,0,199,0,200,0,238,0,143,0,157,0,0,0,176,0,0,0,252,0,0,0,31,0,35,0,119,0,178,0,96,0,0,0,23,0,104,0,160,0,20,0,70,0,40,0,0,0,238,0,124,0,219,0,221,0,146,0,163,0,0,0,138,0,0,0,206,0,119,0,52,0,11,0,166,0,44,0,18,0,200,0,0,0,102,0,55,0,99,0,25,0,47,0,11,0,8,0,146,0,61,0,38,0,174,0,183,0,248,0,161,0,186,0,153,0,0,0,35,0,46,0,179,0,83,0,0,0,169,0,45,0,0,0,85,0,231,0,89,0,0,0,255,0,173,0,46,0,113,0,194,0,51,0,0,0,97,0,90,0,170,0,0,0,15,0,107,0,220,0,0,0,48,0,90,0,185,0,230,0,0,0,12,0,246,0,0,0,162,0,0,0,40,0,164,0,122,0,115,0,91,0,203,0,166,0,155,0,44,0,0,0,233,0,204,0,216,0,0,0,102,0,203,0,214,0,37,0,47,0,238,0,0,0,35,0,0,0,184,0,0,0,186,0,160,0,135,0,199,0,121,0,40,0,158,0,72,0,89,0,90,0,43,0,166,0,69,0,17,0,46,0,0,0,40,0,154,0,138,0,148,0,96,0,209,0,219,0,56,0,236,0,80,0,0,0,178,0,132,0,235,0,123,0,168,0,57,0,143,0,0,0,52,0,148,0,21,0,0,0,47,0,16,0,252,0,152,0,178,0,0,0,0,0,24,0,146,0,0,0,112,0,0,0,251,0,0,0,179,0,146,0,5,0,19,0,122,0,94,0,0,0,38,0,218,0,0,0,84,0,0,0,66,0,212,0,247,0,64,0,166,0,49,0,0,0,96,0,212,0,0,0,190,0,70,0,107,0,231,0,4,0,91,0,33,0,101,0,151,0,31,0,135,0,2,0,0,0,100,0,0,0,156,0,165,0,63,0,183,0,74,0,0,0,162,0,0,0,214,0,117,0,93,0,21,0,238,0,0,0,112,0,143,0,22,0,117,0,39,0,17,0,243,0,0,0,95,0,38,0,182,0,58,0,57,0,180,0,187,0,50,0,42,0,55,0,138,0,221,0,110,0,0,0,232,0,243,0,24,0,100,0,30,0,209,0,183,0,132,0,0,0,122,0,29,0,0,0,0,0,9,0,209,0,172,0,97,0,207,0,43,0,234,0,41,0,105,0);
signal scenario_full  : scenario_type := (32,31,155,31,247,31,148,31,148,30,164,31,121,31,66,31,208,31,130,31,228,31,81,31,138,31,203,31,180,31,89,31,186,31,231,31,47,31,241,31,45,31,57,31,240,31,149,31,107,31,30,31,134,31,222,31,6,31,99,31,99,30,99,29,44,31,167,31,125,31,229,31,11,31,25,31,25,30,13,31,21,31,255,31,239,31,220,31,220,30,58,31,58,30,178,31,178,30,178,29,43,31,84,31,1,31,132,31,210,31,112,31,2,31,2,30,251,31,129,31,25,31,25,30,69,31,207,31,207,30,190,31,201,31,66,31,57,31,69,31,180,31,180,30,24,31,24,30,108,31,91,31,238,31,124,31,124,30,123,31,232,31,200,31,200,30,61,31,30,31,30,30,236,31,113,31,113,30,111,31,76,31,76,30,76,29,240,31,65,31,20,31,159,31,205,31,137,31,74,31,157,31,46,31,46,30,212,31,103,31,103,30,101,31,10,31,10,30,210,31,208,31,117,31,178,31,153,31,196,31,205,31,205,30,202,31,202,30,131,31,185,31,92,31,218,31,241,31,15,31,28,31,193,31,142,31,252,31,19,31,148,31,148,30,148,29,202,31,123,31,123,30,58,31,58,30,190,31,113,31,113,30,113,29,113,28,113,27,112,31,204,31,224,31,19,31,222,31,222,30,174,31,178,31,178,30,182,31,132,31,132,30,135,31,74,31,226,31,206,31,206,30,169,31,33,31,48,31,134,31,204,31,56,31,1,31,165,31,13,31,13,30,172,31,184,31,159,31,208,31,208,30,24,31,24,30,193,31,223,31,111,31,112,31,57,31,57,30,10,31,103,31,103,30,75,31,175,31,175,30,233,31,20,31,20,30,204,31,75,31,75,30,82,31,82,30,199,31,200,31,238,31,143,31,157,31,157,30,176,31,176,30,252,31,252,30,31,31,35,31,119,31,178,31,96,31,96,30,23,31,104,31,160,31,20,31,70,31,40,31,40,30,238,31,124,31,219,31,221,31,146,31,163,31,163,30,138,31,138,30,206,31,119,31,52,31,11,31,166,31,44,31,18,31,200,31,200,30,102,31,55,31,99,31,25,31,47,31,11,31,8,31,146,31,61,31,38,31,174,31,183,31,248,31,161,31,186,31,153,31,153,30,35,31,46,31,179,31,83,31,83,30,169,31,45,31,45,30,85,31,231,31,89,31,89,30,255,31,173,31,46,31,113,31,194,31,51,31,51,30,97,31,90,31,170,31,170,30,15,31,107,31,220,31,220,30,48,31,90,31,185,31,230,31,230,30,12,31,246,31,246,30,162,31,162,30,40,31,164,31,122,31,115,31,91,31,203,31,166,31,155,31,44,31,44,30,233,31,204,31,216,31,216,30,102,31,203,31,214,31,37,31,47,31,238,31,238,30,35,31,35,30,184,31,184,30,186,31,160,31,135,31,199,31,121,31,40,31,158,31,72,31,89,31,90,31,43,31,166,31,69,31,17,31,46,31,46,30,40,31,154,31,138,31,148,31,96,31,209,31,219,31,56,31,236,31,80,31,80,30,178,31,132,31,235,31,123,31,168,31,57,31,143,31,143,30,52,31,148,31,21,31,21,30,47,31,16,31,252,31,152,31,178,31,178,30,178,29,24,31,146,31,146,30,112,31,112,30,251,31,251,30,179,31,146,31,5,31,19,31,122,31,94,31,94,30,38,31,218,31,218,30,84,31,84,30,66,31,212,31,247,31,64,31,166,31,49,31,49,30,96,31,212,31,212,30,190,31,70,31,107,31,231,31,4,31,91,31,33,31,101,31,151,31,31,31,135,31,2,31,2,30,100,31,100,30,156,31,165,31,63,31,183,31,74,31,74,30,162,31,162,30,214,31,117,31,93,31,21,31,238,31,238,30,112,31,143,31,22,31,117,31,39,31,17,31,243,31,243,30,95,31,38,31,182,31,58,31,57,31,180,31,187,31,50,31,42,31,55,31,138,31,221,31,110,31,110,30,232,31,243,31,24,31,100,31,30,31,209,31,183,31,132,31,132,30,122,31,29,31,29,30,29,29,9,31,209,31,172,31,97,31,207,31,43,31,234,31,41,31,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
