-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_22 is
end project_tb_22;

architecture project_tb_arch_22 of project_tb_22 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 834;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,0,0,41,0,79,0,228,0,228,0,108,0,0,0,123,0,87,0,73,0,182,0,229,0,218,0,192,0,142,0,43,0,214,0,63,0,177,0,155,0,200,0,138,0,96,0,201,0,0,0,32,0,0,0,34,0,115,0,181,0,0,0,209,0,5,0,0,0,185,0,233,0,75,0,0,0,0,0,175,0,84,0,231,0,49,0,22,0,0,0,13,0,51,0,2,0,82,0,0,0,241,0,20,0,228,0,238,0,0,0,199,0,117,0,8,0,0,0,198,0,175,0,45,0,246,0,121,0,43,0,0,0,146,0,60,0,159,0,2,0,138,0,8,0,96,0,197,0,0,0,177,0,231,0,154,0,37,0,124,0,216,0,0,0,0,0,0,0,0,0,195,0,104,0,0,0,134,0,195,0,30,0,46,0,126,0,213,0,85,0,224,0,236,0,18,0,125,0,159,0,122,0,0,0,234,0,0,0,93,0,192,0,16,0,255,0,25,0,0,0,247,0,27,0,77,0,198,0,8,0,139,0,0,0,196,0,114,0,0,0,0,0,190,0,130,0,0,0,160,0,14,0,232,0,106,0,67,0,134,0,0,0,83,0,88,0,151,0,201,0,124,0,103,0,227,0,0,0,177,0,210,0,177,0,207,0,233,0,93,0,120,0,0,0,0,0,61,0,59,0,62,0,176,0,82,0,0,0,124,0,0,0,0,0,5,0,48,0,249,0,194,0,0,0,16,0,0,0,32,0,252,0,120,0,188,0,4,0,235,0,83,0,0,0,114,0,229,0,174,0,101,0,0,0,238,0,53,0,0,0,131,0,64,0,255,0,0,0,108,0,98,0,98,0,60,0,0,0,87,0,94,0,239,0,0,0,26,0,216,0,203,0,98,0,94,0,0,0,0,0,133,0,71,0,2,0,52,0,0,0,0,0,158,0,26,0,22,0,216,0,212,0,0,0,150,0,197,0,225,0,126,0,182,0,181,0,126,0,85,0,233,0,178,0,40,0,93,0,124,0,0,0,178,0,0,0,0,0,32,0,104,0,185,0,61,0,68,0,0,0,226,0,51,0,136,0,242,0,20,0,143,0,164,0,62,0,149,0,23,0,245,0,150,0,59,0,21,0,28,0,101,0,58,0,30,0,0,0,123,0,153,0,101,0,24,0,211,0,0,0,87,0,215,0,246,0,183,0,19,0,177,0,24,0,61,0,138,0,183,0,68,0,185,0,233,0,197,0,180,0,76,0,196,0,208,0,31,0,123,0,43,0,79,0,211,0,0,0,73,0,126,0,86,0,72,0,247,0,152,0,84,0,0,0,0,0,0,0,220,0,112,0,0,0,0,0,229,0,27,0,0,0,0,0,0,0,0,0,0,0,212,0,0,0,242,0,98,0,72,0,143,0,0,0,179,0,174,0,191,0,198,0,118,0,147,0,0,0,0,0,165,0,26,0,207,0,85,0,0,0,165,0,4,0,128,0,0,0,0,0,22,0,71,0,109,0,0,0,56,0,183,0,80,0,232,0,66,0,88,0,198,0,68,0,108,0,168,0,41,0,140,0,90,0,151,0,132,0,0,0,154,0,62,0,199,0,203,0,7,0,66,0,0,0,0,0,20,0,0,0,192,0,0,0,0,0,180,0,180,0,131,0,166,0,99,0,69,0,0,0,203,0,12,0,94,0,83,0,0,0,205,0,0,0,139,0,0,0,155,0,84,0,128,0,52,0,199,0,221,0,119,0,46,0,69,0,8,0,0,0,0,0,79,0,149,0,0,0,54,0,231,0,0,0,81,0,0,0,70,0,210,0,0,0,194,0,55,0,10,0,199,0,113,0,220,0,39,0,0,0,166,0,229,0,0,0,110,0,169,0,178,0,92,0,73,0,236,0,17,0,241,0,230,0,56,0,240,0,2,0,239,0,128,0,72,0,42,0,37,0,134,0,241,0,151,0,54,0,139,0,91,0,175,0,63,0,251,0,83,0,106,0,253,0,210,0,0,0,223,0,211,0,194,0,0,0,0,0,233,0,0,0,140,0,115,0,237,0,242,0,138,0,243,0,67,0,179,0,23,0,0,0,14,0,163,0,40,0,225,0,181,0,251,0,0,0,30,0,177,0,0,0,232,0,7,0,232,0,15,0,0,0,208,0,179,0,138,0,174,0,188,0,0,0,0,0,0,0,185,0,165,0,148,0,0,0,167,0,202,0,0,0,52,0,126,0,247,0,11,0,63,0,10,0,0,0,123,0,91,0,117,0,142,0,245,0,46,0,221,0,68,0,236,0,30,0,0,0,148,0,0,0,57,0,0,0,70,0,52,0,0,0,43,0,97,0,45,0,108,0,105,0,12,0,77,0,110,0,100,0,0,0,85,0,54,0,0,0,30,0,0,0,180,0,44,0,146,0,98,0,29,0,0,0,208,0,111,0,254,0,102,0,144,0,134,0,29,0,192,0,92,0,0,0,228,0,240,0,0,0,0,0,217,0,121,0,112,0,197,0,0,0,100,0,0,0,0,0,0,0,121,0,194,0,86,0,0,0,231,0,0,0,184,0,247,0,0,0,129,0,124,0,230,0,215,0,72,0,154,0,78,0,63,0,227,0,0,0,194,0,230,0,102,0,18,0,0,0,86,0,165,0,195,0,218,0,147,0,110,0,253,0,223,0,182,0,128,0,5,0,64,0,80,0,0,0,233,0,10,0,0,0,77,0,120,0,154,0,184,0,62,0,76,0,222,0,242,0,15,0,160,0,101,0,241,0,230,0,107,0,209,0,154,0,153,0,41,0,0,0,56,0,48,0,103,0,139,0,9,0,193,0,88,0,0,0,33,0,0,0,211,0,28,0,29,0,201,0,0,0,141,0,0,0,243,0,112,0,69,0,170,0,188,0,0,0,126,0,145,0,235,0,183,0,8,0,215,0,0,0,165,0,48,0,117,0,0,0,0,0,57,0,175,0,89,0,177,0,0,0,151,0,203,0,68,0,112,0,159,0,136,0,225,0,216,0,250,0,62,0,64,0,4,0,247,0,253,0,0,0,0,0,184,0,77,0,45,0,243,0,109,0,217,0,216,0,78,0,50,0,252,0,0,0,105,0,0,0,90,0,0,0,0,0,84,0,115,0,203,0,42,0,70,0,31,0,194,0,94,0,35,0,0,0,253,0,60,0,0,0,205,0,0,0,28,0,119,0,0,0,158,0,0,0,197,0,116,0,190,0,181,0,201,0,236,0,154,0,107,0,0,0,11,0,0,0,84,0,187,0,228,0,31,0,168,0,140,0,236,0,11,0,166,0,222,0,172,0,208,0,197,0,2,0,21,0,0,0,0,0,175,0,201,0,8,0,50,0,218,0,77,0,69,0,57,0,228,0,181,0,199,0,0,0,232,0,65,0,128,0,207,0,137,0,178,0,191,0,23,0,16,0,28,0,239,0,67,0,96,0,121,0,0,0,127,0,49,0,0,0,217,0,123,0,74,0,20,0,150,0,0,0,0,0,0,0,108,0,130,0,0,0,0,0,254,0,158,0,54,0,0,0,245,0,59,0,0,0,64,0,101,0,0,0,0,0,80,0,222,0,22,0,0,0,255,0,17,0,0,0,15,0,127,0,194,0,254,0,0,0,108,0,0,0,230,0,93,0,0,0,185,0,60,0,172,0,95,0,79,0,139,0,128,0,0,0,151,0,198,0,0,0,149,0,17,0,74,0,170,0,99,0,38,0,0,0,0,0,49,0,75,0,192,0,0,0);
signal scenario_full  : scenario_type := (7,31,7,30,41,31,79,31,228,31,228,31,108,31,108,30,123,31,87,31,73,31,182,31,229,31,218,31,192,31,142,31,43,31,214,31,63,31,177,31,155,31,200,31,138,31,96,31,201,31,201,30,32,31,32,30,34,31,115,31,181,31,181,30,209,31,5,31,5,30,185,31,233,31,75,31,75,30,75,29,175,31,84,31,231,31,49,31,22,31,22,30,13,31,51,31,2,31,82,31,82,30,241,31,20,31,228,31,238,31,238,30,199,31,117,31,8,31,8,30,198,31,175,31,45,31,246,31,121,31,43,31,43,30,146,31,60,31,159,31,2,31,138,31,8,31,96,31,197,31,197,30,177,31,231,31,154,31,37,31,124,31,216,31,216,30,216,29,216,28,216,27,195,31,104,31,104,30,134,31,195,31,30,31,46,31,126,31,213,31,85,31,224,31,236,31,18,31,125,31,159,31,122,31,122,30,234,31,234,30,93,31,192,31,16,31,255,31,25,31,25,30,247,31,27,31,77,31,198,31,8,31,139,31,139,30,196,31,114,31,114,30,114,29,190,31,130,31,130,30,160,31,14,31,232,31,106,31,67,31,134,31,134,30,83,31,88,31,151,31,201,31,124,31,103,31,227,31,227,30,177,31,210,31,177,31,207,31,233,31,93,31,120,31,120,30,120,29,61,31,59,31,62,31,176,31,82,31,82,30,124,31,124,30,124,29,5,31,48,31,249,31,194,31,194,30,16,31,16,30,32,31,252,31,120,31,188,31,4,31,235,31,83,31,83,30,114,31,229,31,174,31,101,31,101,30,238,31,53,31,53,30,131,31,64,31,255,31,255,30,108,31,98,31,98,31,60,31,60,30,87,31,94,31,239,31,239,30,26,31,216,31,203,31,98,31,94,31,94,30,94,29,133,31,71,31,2,31,52,31,52,30,52,29,158,31,26,31,22,31,216,31,212,31,212,30,150,31,197,31,225,31,126,31,182,31,181,31,126,31,85,31,233,31,178,31,40,31,93,31,124,31,124,30,178,31,178,30,178,29,32,31,104,31,185,31,61,31,68,31,68,30,226,31,51,31,136,31,242,31,20,31,143,31,164,31,62,31,149,31,23,31,245,31,150,31,59,31,21,31,28,31,101,31,58,31,30,31,30,30,123,31,153,31,101,31,24,31,211,31,211,30,87,31,215,31,246,31,183,31,19,31,177,31,24,31,61,31,138,31,183,31,68,31,185,31,233,31,197,31,180,31,76,31,196,31,208,31,31,31,123,31,43,31,79,31,211,31,211,30,73,31,126,31,86,31,72,31,247,31,152,31,84,31,84,30,84,29,84,28,220,31,112,31,112,30,112,29,229,31,27,31,27,30,27,29,27,28,27,27,27,26,212,31,212,30,242,31,98,31,72,31,143,31,143,30,179,31,174,31,191,31,198,31,118,31,147,31,147,30,147,29,165,31,26,31,207,31,85,31,85,30,165,31,4,31,128,31,128,30,128,29,22,31,71,31,109,31,109,30,56,31,183,31,80,31,232,31,66,31,88,31,198,31,68,31,108,31,168,31,41,31,140,31,90,31,151,31,132,31,132,30,154,31,62,31,199,31,203,31,7,31,66,31,66,30,66,29,20,31,20,30,192,31,192,30,192,29,180,31,180,31,131,31,166,31,99,31,69,31,69,30,203,31,12,31,94,31,83,31,83,30,205,31,205,30,139,31,139,30,155,31,84,31,128,31,52,31,199,31,221,31,119,31,46,31,69,31,8,31,8,30,8,29,79,31,149,31,149,30,54,31,231,31,231,30,81,31,81,30,70,31,210,31,210,30,194,31,55,31,10,31,199,31,113,31,220,31,39,31,39,30,166,31,229,31,229,30,110,31,169,31,178,31,92,31,73,31,236,31,17,31,241,31,230,31,56,31,240,31,2,31,239,31,128,31,72,31,42,31,37,31,134,31,241,31,151,31,54,31,139,31,91,31,175,31,63,31,251,31,83,31,106,31,253,31,210,31,210,30,223,31,211,31,194,31,194,30,194,29,233,31,233,30,140,31,115,31,237,31,242,31,138,31,243,31,67,31,179,31,23,31,23,30,14,31,163,31,40,31,225,31,181,31,251,31,251,30,30,31,177,31,177,30,232,31,7,31,232,31,15,31,15,30,208,31,179,31,138,31,174,31,188,31,188,30,188,29,188,28,185,31,165,31,148,31,148,30,167,31,202,31,202,30,52,31,126,31,247,31,11,31,63,31,10,31,10,30,123,31,91,31,117,31,142,31,245,31,46,31,221,31,68,31,236,31,30,31,30,30,148,31,148,30,57,31,57,30,70,31,52,31,52,30,43,31,97,31,45,31,108,31,105,31,12,31,77,31,110,31,100,31,100,30,85,31,54,31,54,30,30,31,30,30,180,31,44,31,146,31,98,31,29,31,29,30,208,31,111,31,254,31,102,31,144,31,134,31,29,31,192,31,92,31,92,30,228,31,240,31,240,30,240,29,217,31,121,31,112,31,197,31,197,30,100,31,100,30,100,29,100,28,121,31,194,31,86,31,86,30,231,31,231,30,184,31,247,31,247,30,129,31,124,31,230,31,215,31,72,31,154,31,78,31,63,31,227,31,227,30,194,31,230,31,102,31,18,31,18,30,86,31,165,31,195,31,218,31,147,31,110,31,253,31,223,31,182,31,128,31,5,31,64,31,80,31,80,30,233,31,10,31,10,30,77,31,120,31,154,31,184,31,62,31,76,31,222,31,242,31,15,31,160,31,101,31,241,31,230,31,107,31,209,31,154,31,153,31,41,31,41,30,56,31,48,31,103,31,139,31,9,31,193,31,88,31,88,30,33,31,33,30,211,31,28,31,29,31,201,31,201,30,141,31,141,30,243,31,112,31,69,31,170,31,188,31,188,30,126,31,145,31,235,31,183,31,8,31,215,31,215,30,165,31,48,31,117,31,117,30,117,29,57,31,175,31,89,31,177,31,177,30,151,31,203,31,68,31,112,31,159,31,136,31,225,31,216,31,250,31,62,31,64,31,4,31,247,31,253,31,253,30,253,29,184,31,77,31,45,31,243,31,109,31,217,31,216,31,78,31,50,31,252,31,252,30,105,31,105,30,90,31,90,30,90,29,84,31,115,31,203,31,42,31,70,31,31,31,194,31,94,31,35,31,35,30,253,31,60,31,60,30,205,31,205,30,28,31,119,31,119,30,158,31,158,30,197,31,116,31,190,31,181,31,201,31,236,31,154,31,107,31,107,30,11,31,11,30,84,31,187,31,228,31,31,31,168,31,140,31,236,31,11,31,166,31,222,31,172,31,208,31,197,31,2,31,21,31,21,30,21,29,175,31,201,31,8,31,50,31,218,31,77,31,69,31,57,31,228,31,181,31,199,31,199,30,232,31,65,31,128,31,207,31,137,31,178,31,191,31,23,31,16,31,28,31,239,31,67,31,96,31,121,31,121,30,127,31,49,31,49,30,217,31,123,31,74,31,20,31,150,31,150,30,150,29,150,28,108,31,130,31,130,30,130,29,254,31,158,31,54,31,54,30,245,31,59,31,59,30,64,31,101,31,101,30,101,29,80,31,222,31,22,31,22,30,255,31,17,31,17,30,15,31,127,31,194,31,254,31,254,30,108,31,108,30,230,31,93,31,93,30,185,31,60,31,172,31,95,31,79,31,139,31,128,31,128,30,151,31,198,31,198,30,149,31,17,31,74,31,170,31,99,31,38,31,38,30,38,29,49,31,75,31,192,31,192,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
