-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_597 is
end project_tb_597;

architecture project_tb_arch_597 of project_tb_597 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 543;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,251,0,38,0,237,0,0,0,198,0,216,0,0,0,148,0,60,0,16,0,222,0,0,0,156,0,162,0,197,0,65,0,250,0,251,0,176,0,222,0,7,0,225,0,186,0,202,0,124,0,249,0,247,0,0,0,189,0,117,0,106,0,131,0,244,0,200,0,0,0,0,0,132,0,178,0,168,0,79,0,21,0,131,0,205,0,201,0,182,0,218,0,0,0,187,0,235,0,185,0,164,0,104,0,108,0,116,0,159,0,193,0,221,0,143,0,162,0,195,0,72,0,45,0,252,0,0,0,71,0,13,0,51,0,161,0,0,0,35,0,149,0,88,0,0,0,0,0,171,0,131,0,112,0,205,0,78,0,40,0,144,0,0,0,0,0,165,0,158,0,57,0,110,0,86,0,9,0,207,0,0,0,17,0,15,0,164,0,76,0,64,0,136,0,131,0,220,0,131,0,110,0,149,0,0,0,172,0,23,0,31,0,136,0,35,0,0,0,98,0,166,0,211,0,252,0,0,0,86,0,133,0,80,0,48,0,45,0,0,0,3,0,201,0,0,0,91,0,53,0,148,0,0,0,121,0,18,0,121,0,0,0,230,0,135,0,218,0,17,0,26,0,0,0,6,0,61,0,232,0,173,0,112,0,0,0,141,0,195,0,84,0,191,0,23,0,193,0,0,0,251,0,214,0,29,0,46,0,16,0,9,0,0,0,0,0,235,0,0,0,217,0,127,0,40,0,152,0,89,0,116,0,0,0,241,0,235,0,231,0,220,0,152,0,185,0,97,0,201,0,0,0,0,0,212,0,178,0,131,0,206,0,44,0,200,0,0,0,29,0,155,0,163,0,0,0,161,0,36,0,180,0,190,0,101,0,0,0,0,0,69,0,74,0,0,0,161,0,231,0,105,0,0,0,60,0,49,0,0,0,94,0,69,0,248,0,172,0,17,0,0,0,245,0,132,0,54,0,2,0,235,0,174,0,190,0,246,0,68,0,172,0,201,0,0,0,8,0,21,0,29,0,180,0,0,0,0,0,115,0,197,0,2,0,12,0,0,0,255,0,99,0,222,0,153,0,155,0,0,0,38,0,0,0,96,0,148,0,119,0,51,0,57,0,0,0,184,0,83,0,232,0,29,0,0,0,204,0,68,0,48,0,118,0,232,0,0,0,76,0,104,0,244,0,29,0,152,0,237,0,234,0,236,0,122,0,0,0,165,0,183,0,0,0,227,0,104,0,142,0,131,0,0,0,158,0,11,0,128,0,21,0,238,0,184,0,65,0,115,0,58,0,72,0,171,0,159,0,191,0,176,0,155,0,147,0,38,0,32,0,227,0,46,0,27,0,223,0,0,0,4,0,16,0,147,0,66,0,164,0,0,0,110,0,0,0,189,0,42,0,0,0,110,0,80,0,46,0,172,0,0,0,179,0,100,0,0,0,94,0,40,0,100,0,91,0,148,0,93,0,74,0,99,0,118,0,0,0,207,0,24,0,0,0,216,0,34,0,45,0,47,0,202,0,86,0,0,0,211,0,0,0,100,0,168,0,194,0,86,0,142,0,0,0,0,0,62,0,47,0,103,0,215,0,216,0,154,0,226,0,175,0,0,0,38,0,222,0,252,0,110,0,114,0,131,0,205,0,196,0,131,0,241,0,174,0,9,0,90,0,5,0,0,0,121,0,9,0,11,0,254,0,56,0,1,0,0,0,0,0,73,0,0,0,0,0,200,0,89,0,72,0,46,0,99,0,189,0,35,0,105,0,179,0,66,0,160,0,92,0,122,0,210,0,8,0,0,0,57,0,248,0,77,0,154,0,200,0,117,0,177,0,47,0,0,0,0,0,67,0,29,0,46,0,234,0,166,0,113,0,118,0,134,0,0,0,99,0,175,0,0,0,193,0,82,0,104,0,139,0,228,0,14,0,157,0,160,0,0,0,216,0,130,0,230,0,100,0,0,0,29,0,82,0,3,0,51,0,0,0,120,0,32,0,102,0,0,0,219,0,252,0,28,0,79,0,17,0,137,0,151,0,0,0,72,0,174,0,58,0,0,0,0,0,0,0,13,0,221,0,178,0,194,0,29,0,11,0,87,0,0,0,237,0,0,0,0,0,172,0,186,0,135,0,5,0,45,0,141,0,152,0,49,0,0,0,0,0,11,0,228,0,0,0,9,0,31,0,208,0,58,0,220,0,151,0,0,0,118,0,111,0,31,0,0,0,91,0,0,0,55,0,220,0,35,0,195,0,192,0,191,0,125,0,136,0,6,0,175,0,235,0,224,0,0,0,129,0,165,0,220,0,163,0,142,0,245,0,49,0,0,0,0,0,69,0,108,0,253,0,0,0,196,0,0,0,148,0,161,0,190,0,198,0,0,0,0,0,156,0,212,0,53,0,93,0,146,0,221,0,0,0,82,0,91,0,81,0,219,0,40,0,5,0);
signal scenario_full  : scenario_type := (0,0,251,31,38,31,237,31,237,30,198,31,216,31,216,30,148,31,60,31,16,31,222,31,222,30,156,31,162,31,197,31,65,31,250,31,251,31,176,31,222,31,7,31,225,31,186,31,202,31,124,31,249,31,247,31,247,30,189,31,117,31,106,31,131,31,244,31,200,31,200,30,200,29,132,31,178,31,168,31,79,31,21,31,131,31,205,31,201,31,182,31,218,31,218,30,187,31,235,31,185,31,164,31,104,31,108,31,116,31,159,31,193,31,221,31,143,31,162,31,195,31,72,31,45,31,252,31,252,30,71,31,13,31,51,31,161,31,161,30,35,31,149,31,88,31,88,30,88,29,171,31,131,31,112,31,205,31,78,31,40,31,144,31,144,30,144,29,165,31,158,31,57,31,110,31,86,31,9,31,207,31,207,30,17,31,15,31,164,31,76,31,64,31,136,31,131,31,220,31,131,31,110,31,149,31,149,30,172,31,23,31,31,31,136,31,35,31,35,30,98,31,166,31,211,31,252,31,252,30,86,31,133,31,80,31,48,31,45,31,45,30,3,31,201,31,201,30,91,31,53,31,148,31,148,30,121,31,18,31,121,31,121,30,230,31,135,31,218,31,17,31,26,31,26,30,6,31,61,31,232,31,173,31,112,31,112,30,141,31,195,31,84,31,191,31,23,31,193,31,193,30,251,31,214,31,29,31,46,31,16,31,9,31,9,30,9,29,235,31,235,30,217,31,127,31,40,31,152,31,89,31,116,31,116,30,241,31,235,31,231,31,220,31,152,31,185,31,97,31,201,31,201,30,201,29,212,31,178,31,131,31,206,31,44,31,200,31,200,30,29,31,155,31,163,31,163,30,161,31,36,31,180,31,190,31,101,31,101,30,101,29,69,31,74,31,74,30,161,31,231,31,105,31,105,30,60,31,49,31,49,30,94,31,69,31,248,31,172,31,17,31,17,30,245,31,132,31,54,31,2,31,235,31,174,31,190,31,246,31,68,31,172,31,201,31,201,30,8,31,21,31,29,31,180,31,180,30,180,29,115,31,197,31,2,31,12,31,12,30,255,31,99,31,222,31,153,31,155,31,155,30,38,31,38,30,96,31,148,31,119,31,51,31,57,31,57,30,184,31,83,31,232,31,29,31,29,30,204,31,68,31,48,31,118,31,232,31,232,30,76,31,104,31,244,31,29,31,152,31,237,31,234,31,236,31,122,31,122,30,165,31,183,31,183,30,227,31,104,31,142,31,131,31,131,30,158,31,11,31,128,31,21,31,238,31,184,31,65,31,115,31,58,31,72,31,171,31,159,31,191,31,176,31,155,31,147,31,38,31,32,31,227,31,46,31,27,31,223,31,223,30,4,31,16,31,147,31,66,31,164,31,164,30,110,31,110,30,189,31,42,31,42,30,110,31,80,31,46,31,172,31,172,30,179,31,100,31,100,30,94,31,40,31,100,31,91,31,148,31,93,31,74,31,99,31,118,31,118,30,207,31,24,31,24,30,216,31,34,31,45,31,47,31,202,31,86,31,86,30,211,31,211,30,100,31,168,31,194,31,86,31,142,31,142,30,142,29,62,31,47,31,103,31,215,31,216,31,154,31,226,31,175,31,175,30,38,31,222,31,252,31,110,31,114,31,131,31,205,31,196,31,131,31,241,31,174,31,9,31,90,31,5,31,5,30,121,31,9,31,11,31,254,31,56,31,1,31,1,30,1,29,73,31,73,30,73,29,200,31,89,31,72,31,46,31,99,31,189,31,35,31,105,31,179,31,66,31,160,31,92,31,122,31,210,31,8,31,8,30,57,31,248,31,77,31,154,31,200,31,117,31,177,31,47,31,47,30,47,29,67,31,29,31,46,31,234,31,166,31,113,31,118,31,134,31,134,30,99,31,175,31,175,30,193,31,82,31,104,31,139,31,228,31,14,31,157,31,160,31,160,30,216,31,130,31,230,31,100,31,100,30,29,31,82,31,3,31,51,31,51,30,120,31,32,31,102,31,102,30,219,31,252,31,28,31,79,31,17,31,137,31,151,31,151,30,72,31,174,31,58,31,58,30,58,29,58,28,13,31,221,31,178,31,194,31,29,31,11,31,87,31,87,30,237,31,237,30,237,29,172,31,186,31,135,31,5,31,45,31,141,31,152,31,49,31,49,30,49,29,11,31,228,31,228,30,9,31,31,31,208,31,58,31,220,31,151,31,151,30,118,31,111,31,31,31,31,30,91,31,91,30,55,31,220,31,35,31,195,31,192,31,191,31,125,31,136,31,6,31,175,31,235,31,224,31,224,30,129,31,165,31,220,31,163,31,142,31,245,31,49,31,49,30,49,29,69,31,108,31,253,31,253,30,196,31,196,30,148,31,161,31,190,31,198,31,198,30,198,29,156,31,212,31,53,31,93,31,146,31,221,31,221,30,82,31,91,31,81,31,219,31,40,31,5,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
