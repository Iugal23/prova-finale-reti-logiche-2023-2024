-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 272;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (165,0,8,0,66,0,71,0,123,0,202,0,81,0,72,0,0,0,59,0,0,0,0,0,233,0,39,0,31,0,98,0,79,0,187,0,184,0,165,0,96,0,111,0,218,0,18,0,209,0,0,0,93,0,255,0,80,0,0,0,56,0,81,0,47,0,197,0,0,0,179,0,0,0,49,0,110,0,6,0,137,0,31,0,158,0,0,0,252,0,186,0,0,0,148,0,246,0,34,0,160,0,199,0,49,0,0,0,0,0,123,0,0,0,16,0,105,0,92,0,144,0,0,0,221,0,195,0,211,0,233,0,137,0,145,0,178,0,52,0,148,0,156,0,0,0,0,0,44,0,0,0,122,0,22,0,23,0,172,0,132,0,0,0,131,0,239,0,75,0,78,0,250,0,0,0,0,0,74,0,89,0,0,0,5,0,232,0,41,0,151,0,125,0,218,0,112,0,190,0,138,0,62,0,0,0,178,0,216,0,42,0,183,0,144,0,0,0,153,0,58,0,11,0,177,0,145,0,14,0,50,0,90,0,184,0,140,0,4,0,107,0,175,0,29,0,233,0,184,0,232,0,83,0,56,0,115,0,80,0,144,0,97,0,0,0,242,0,193,0,221,0,0,0,0,0,225,0,50,0,254,0,255,0,0,0,213,0,24,0,0,0,125,0,58,0,160,0,77,0,102,0,111,0,159,0,213,0,117,0,205,0,42,0,0,0,197,0,64,0,218,0,30,0,142,0,70,0,0,0,0,0,38,0,0,0,182,0,94,0,243,0,58,0,90,0,55,0,0,0,139,0,234,0,173,0,250,0,158,0,131,0,0,0,181,0,105,0,240,0,254,0,226,0,90,0,186,0,137,0,141,0,247,0,53,0,85,0,38,0,6,0,152,0,116,0,168,0,209,0,244,0,81,0,111,0,158,0,146,0,139,0,84,0,215,0,233,0,0,0,120,0,0,0,242,0,201,0,101,0,181,0,207,0,215,0,225,0,218,0,0,0,142,0,20,0,0,0,4,0,0,0,36,0,45,0,64,0,68,0,239,0,0,0,0,0,0,0,211,0,218,0,180,0,29,0,0,0,111,0,181,0,40,0,235,0,182,0,125,0,85,0,199,0,13,0,142,0,129,0,192,0,69,0,47,0,179,0,135,0,95,0,123,0,202,0,128,0,195,0,0,0,0,0,38,0,29,0,165,0,113,0,134,0,0,0,117,0,61,0,44,0,144,0);
signal scenario_full  : scenario_type := (165,31,8,31,66,31,71,31,123,31,202,31,81,31,72,31,72,30,59,31,59,30,59,29,233,31,39,31,31,31,98,31,79,31,187,31,184,31,165,31,96,31,111,31,218,31,18,31,209,31,209,30,93,31,255,31,80,31,80,30,56,31,81,31,47,31,197,31,197,30,179,31,179,30,49,31,110,31,6,31,137,31,31,31,158,31,158,30,252,31,186,31,186,30,148,31,246,31,34,31,160,31,199,31,49,31,49,30,49,29,123,31,123,30,16,31,105,31,92,31,144,31,144,30,221,31,195,31,211,31,233,31,137,31,145,31,178,31,52,31,148,31,156,31,156,30,156,29,44,31,44,30,122,31,22,31,23,31,172,31,132,31,132,30,131,31,239,31,75,31,78,31,250,31,250,30,250,29,74,31,89,31,89,30,5,31,232,31,41,31,151,31,125,31,218,31,112,31,190,31,138,31,62,31,62,30,178,31,216,31,42,31,183,31,144,31,144,30,153,31,58,31,11,31,177,31,145,31,14,31,50,31,90,31,184,31,140,31,4,31,107,31,175,31,29,31,233,31,184,31,232,31,83,31,56,31,115,31,80,31,144,31,97,31,97,30,242,31,193,31,221,31,221,30,221,29,225,31,50,31,254,31,255,31,255,30,213,31,24,31,24,30,125,31,58,31,160,31,77,31,102,31,111,31,159,31,213,31,117,31,205,31,42,31,42,30,197,31,64,31,218,31,30,31,142,31,70,31,70,30,70,29,38,31,38,30,182,31,94,31,243,31,58,31,90,31,55,31,55,30,139,31,234,31,173,31,250,31,158,31,131,31,131,30,181,31,105,31,240,31,254,31,226,31,90,31,186,31,137,31,141,31,247,31,53,31,85,31,38,31,6,31,152,31,116,31,168,31,209,31,244,31,81,31,111,31,158,31,146,31,139,31,84,31,215,31,233,31,233,30,120,31,120,30,242,31,201,31,101,31,181,31,207,31,215,31,225,31,218,31,218,30,142,31,20,31,20,30,4,31,4,30,36,31,45,31,64,31,68,31,239,31,239,30,239,29,239,28,211,31,218,31,180,31,29,31,29,30,111,31,181,31,40,31,235,31,182,31,125,31,85,31,199,31,13,31,142,31,129,31,192,31,69,31,47,31,179,31,135,31,95,31,123,31,202,31,128,31,195,31,195,30,195,29,38,31,29,31,165,31,113,31,134,31,134,30,117,31,61,31,44,31,144,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
