-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 469;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,0,0,153,0,0,0,28,0,207,0,220,0,45,0,160,0,229,0,0,0,180,0,201,0,87,0,156,0,191,0,91,0,80,0,0,0,69,0,241,0,159,0,92,0,2,0,136,0,0,0,227,0,158,0,139,0,158,0,36,0,179,0,0,0,249,0,212,0,220,0,13,0,147,0,179,0,85,0,146,0,45,0,5,0,62,0,21,0,55,0,0,0,0,0,0,0,242,0,69,0,222,0,1,0,0,0,223,0,235,0,33,0,0,0,0,0,39,0,206,0,46,0,136,0,7,0,119,0,140,0,164,0,240,0,247,0,0,0,191,0,0,0,0,0,51,0,76,0,224,0,30,0,163,0,40,0,127,0,0,0,155,0,185,0,89,0,139,0,63,0,62,0,228,0,170,0,221,0,170,0,225,0,225,0,176,0,66,0,234,0,129,0,9,0,151,0,73,0,208,0,37,0,97,0,80,0,0,0,0,0,164,0,247,0,27,0,169,0,254,0,6,0,0,0,0,0,157,0,88,0,32,0,234,0,210,0,32,0,242,0,0,0,245,0,62,0,58,0,206,0,149,0,71,0,135,0,0,0,61,0,1,0,0,0,78,0,35,0,130,0,96,0,220,0,119,0,218,0,0,0,247,0,236,0,0,0,0,0,0,0,182,0,156,0,78,0,42,0,72,0,116,0,51,0,243,0,197,0,146,0,0,0,31,0,93,0,56,0,126,0,13,0,14,0,61,0,230,0,0,0,236,0,230,0,138,0,0,0,237,0,0,0,0,0,240,0,159,0,61,0,212,0,69,0,40,0,160,0,63,0,136,0,240,0,168,0,221,0,251,0,0,0,97,0,141,0,228,0,218,0,194,0,64,0,60,0,134,0,45,0,0,0,123,0,0,0,53,0,19,0,188,0,0,0,164,0,133,0,115,0,208,0,190,0,0,0,217,0,0,0,229,0,26,0,154,0,176,0,174,0,183,0,16,0,225,0,14,0,178,0,0,0,0,0,67,0,205,0,31,0,12,0,8,0,234,0,106,0,196,0,167,0,0,0,0,0,0,0,229,0,0,0,239,0,0,0,31,0,161,0,237,0,0,0,0,0,94,0,0,0,0,0,0,0,23,0,103,0,192,0,171,0,80,0,128,0,29,0,64,0,112,0,174,0,84,0,230,0,236,0,98,0,89,0,0,0,79,0,248,0,89,0,245,0,3,0,7,0,211,0,160,0,0,0,203,0,46,0,0,0,251,0,172,0,0,0,218,0,35,0,46,0,205,0,223,0,56,0,12,0,155,0,99,0,181,0,92,0,141,0,0,0,199,0,0,0,227,0,118,0,0,0,154,0,204,0,224,0,88,0,0,0,0,0,0,0,119,0,38,0,76,0,0,0,60,0,0,0,143,0,35,0,110,0,126,0,80,0,214,0,0,0,78,0,224,0,23,0,32,0,214,0,0,0,169,0,123,0,207,0,189,0,168,0,174,0,132,0,188,0,0,0,24,0,108,0,46,0,95,0,11,0,109,0,227,0,49,0,126,0,192,0,121,0,48,0,107,0,0,0,0,0,0,0,200,0,8,0,0,0,0,0,0,0,228,0,29,0,134,0,0,0,0,0,0,0,144,0,0,0,3,0,131,0,0,0,10,0,166,0,99,0,62,0,172,0,0,0,165,0,48,0,56,0,142,0,182,0,253,0,79,0,0,0,0,0,206,0,161,0,0,0,0,0,168,0,32,0,0,0,40,0,157,0,93,0,11,0,0,0,85,0,0,0,167,0,197,0,61,0,0,0,0,0,1,0,242,0,120,0,115,0,6,0,0,0,198,0,0,0,190,0,253,0,0,0,180,0,142,0,165,0,0,0,77,0,225,0,0,0,151,0,74,0,57,0,9,0,194,0,9,0,91,0,7,0,84,0,203,0,172,0,38,0,57,0,244,0,219,0,82,0,0,0,114,0,13,0,207,0,47,0,181,0,160,0,0,0,229,0,171,0,25,0,74,0,0,0,6,0,141,0,171,0,155,0,0,0,0,0,6,0,109,0,147,0,199,0,0,0,0,0,217,0,104,0,63,0,253,0,0,0,145,0,86,0,0,0,0,0,78,0,0,0,62,0);
signal scenario_full  : scenario_type := (128,31,128,30,153,31,153,30,28,31,207,31,220,31,45,31,160,31,229,31,229,30,180,31,201,31,87,31,156,31,191,31,91,31,80,31,80,30,69,31,241,31,159,31,92,31,2,31,136,31,136,30,227,31,158,31,139,31,158,31,36,31,179,31,179,30,249,31,212,31,220,31,13,31,147,31,179,31,85,31,146,31,45,31,5,31,62,31,21,31,55,31,55,30,55,29,55,28,242,31,69,31,222,31,1,31,1,30,223,31,235,31,33,31,33,30,33,29,39,31,206,31,46,31,136,31,7,31,119,31,140,31,164,31,240,31,247,31,247,30,191,31,191,30,191,29,51,31,76,31,224,31,30,31,163,31,40,31,127,31,127,30,155,31,185,31,89,31,139,31,63,31,62,31,228,31,170,31,221,31,170,31,225,31,225,31,176,31,66,31,234,31,129,31,9,31,151,31,73,31,208,31,37,31,97,31,80,31,80,30,80,29,164,31,247,31,27,31,169,31,254,31,6,31,6,30,6,29,157,31,88,31,32,31,234,31,210,31,32,31,242,31,242,30,245,31,62,31,58,31,206,31,149,31,71,31,135,31,135,30,61,31,1,31,1,30,78,31,35,31,130,31,96,31,220,31,119,31,218,31,218,30,247,31,236,31,236,30,236,29,236,28,182,31,156,31,78,31,42,31,72,31,116,31,51,31,243,31,197,31,146,31,146,30,31,31,93,31,56,31,126,31,13,31,14,31,61,31,230,31,230,30,236,31,230,31,138,31,138,30,237,31,237,30,237,29,240,31,159,31,61,31,212,31,69,31,40,31,160,31,63,31,136,31,240,31,168,31,221,31,251,31,251,30,97,31,141,31,228,31,218,31,194,31,64,31,60,31,134,31,45,31,45,30,123,31,123,30,53,31,19,31,188,31,188,30,164,31,133,31,115,31,208,31,190,31,190,30,217,31,217,30,229,31,26,31,154,31,176,31,174,31,183,31,16,31,225,31,14,31,178,31,178,30,178,29,67,31,205,31,31,31,12,31,8,31,234,31,106,31,196,31,167,31,167,30,167,29,167,28,229,31,229,30,239,31,239,30,31,31,161,31,237,31,237,30,237,29,94,31,94,30,94,29,94,28,23,31,103,31,192,31,171,31,80,31,128,31,29,31,64,31,112,31,174,31,84,31,230,31,236,31,98,31,89,31,89,30,79,31,248,31,89,31,245,31,3,31,7,31,211,31,160,31,160,30,203,31,46,31,46,30,251,31,172,31,172,30,218,31,35,31,46,31,205,31,223,31,56,31,12,31,155,31,99,31,181,31,92,31,141,31,141,30,199,31,199,30,227,31,118,31,118,30,154,31,204,31,224,31,88,31,88,30,88,29,88,28,119,31,38,31,76,31,76,30,60,31,60,30,143,31,35,31,110,31,126,31,80,31,214,31,214,30,78,31,224,31,23,31,32,31,214,31,214,30,169,31,123,31,207,31,189,31,168,31,174,31,132,31,188,31,188,30,24,31,108,31,46,31,95,31,11,31,109,31,227,31,49,31,126,31,192,31,121,31,48,31,107,31,107,30,107,29,107,28,200,31,8,31,8,30,8,29,8,28,228,31,29,31,134,31,134,30,134,29,134,28,144,31,144,30,3,31,131,31,131,30,10,31,166,31,99,31,62,31,172,31,172,30,165,31,48,31,56,31,142,31,182,31,253,31,79,31,79,30,79,29,206,31,161,31,161,30,161,29,168,31,32,31,32,30,40,31,157,31,93,31,11,31,11,30,85,31,85,30,167,31,197,31,61,31,61,30,61,29,1,31,242,31,120,31,115,31,6,31,6,30,198,31,198,30,190,31,253,31,253,30,180,31,142,31,165,31,165,30,77,31,225,31,225,30,151,31,74,31,57,31,9,31,194,31,9,31,91,31,7,31,84,31,203,31,172,31,38,31,57,31,244,31,219,31,82,31,82,30,114,31,13,31,207,31,47,31,181,31,160,31,160,30,229,31,171,31,25,31,74,31,74,30,6,31,141,31,171,31,155,31,155,30,155,29,6,31,109,31,147,31,199,31,199,30,199,29,217,31,104,31,63,31,253,31,253,30,145,31,86,31,86,30,86,29,78,31,78,30,62,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
