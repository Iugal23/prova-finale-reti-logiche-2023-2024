-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_198 is
end project_tb_198;

architecture project_tb_arch_198 of project_tb_198 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 491;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,87,0,50,0,150,0,222,0,0,0,246,0,32,0,163,0,81,0,213,0,228,0,45,0,0,0,133,0,0,0,204,0,0,0,228,0,0,0,18,0,0,0,99,0,195,0,121,0,136,0,226,0,143,0,28,0,0,0,242,0,46,0,51,0,138,0,28,0,197,0,83,0,224,0,91,0,45,0,241,0,0,0,174,0,82,0,213,0,198,0,0,0,214,0,43,0,246,0,111,0,0,0,0,0,0,0,98,0,242,0,13,0,0,0,0,0,189,0,202,0,189,0,143,0,174,0,233,0,130,0,0,0,230,0,79,0,173,0,0,0,113,0,46,0,157,0,172,0,0,0,102,0,130,0,3,0,40,0,59,0,116,0,253,0,79,0,180,0,108,0,0,0,206,0,251,0,248,0,0,0,0,0,0,0,166,0,0,0,221,0,131,0,171,0,185,0,143,0,118,0,27,0,234,0,158,0,101,0,219,0,97,0,106,0,0,0,147,0,189,0,73,0,0,0,119,0,17,0,198,0,163,0,0,0,0,0,80,0,0,0,117,0,0,0,189,0,5,0,39,0,0,0,205,0,109,0,24,0,119,0,0,0,238,0,0,0,204,0,147,0,0,0,43,0,0,0,245,0,13,0,29,0,248,0,131,0,69,0,31,0,0,0,0,0,0,0,109,0,224,0,105,0,0,0,0,0,159,0,64,0,0,0,39,0,0,0,226,0,202,0,204,0,160,0,57,0,209,0,213,0,19,0,47,0,131,0,111,0,138,0,87,0,221,0,17,0,125,0,134,0,61,0,169,0,5,0,153,0,164,0,173,0,187,0,215,0,0,0,0,0,0,0,97,0,73,0,20,0,0,0,23,0,0,0,222,0,0,0,0,0,230,0,0,0,0,0,0,0,220,0,131,0,89,0,102,0,23,0,192,0,0,0,134,0,233,0,8,0,212,0,0,0,0,0,0,0,139,0,180,0,0,0,205,0,0,0,35,0,124,0,11,0,120,0,121,0,120,0,173,0,86,0,87,0,181,0,152,0,0,0,137,0,152,0,36,0,196,0,40,0,202,0,30,0,128,0,94,0,81,0,0,0,98,0,64,0,91,0,146,0,18,0,137,0,0,0,0,0,166,0,6,0,165,0,76,0,76,0,0,0,152,0,101,0,36,0,10,0,162,0,186,0,0,0,0,0,237,0,4,0,0,0,239,0,171,0,138,0,209,0,0,0,217,0,185,0,222,0,152,0,88,0,8,0,107,0,0,0,191,0,76,0,22,0,241,0,76,0,239,0,113,0,0,0,0,0,195,0,0,0,227,0,0,0,164,0,51,0,116,0,187,0,114,0,144,0,170,0,0,0,250,0,103,0,95,0,217,0,213,0,139,0,254,0,109,0,0,0,248,0,73,0,192,0,175,0,180,0,175,0,37,0,215,0,0,0,71,0,166,0,158,0,124,0,0,0,169,0,244,0,132,0,0,0,221,0,230,0,178,0,50,0,212,0,210,0,0,0,40,0,2,0,0,0,104,0,68,0,215,0,178,0,137,0,0,0,33,0,22,0,161,0,0,0,150,0,172,0,0,0,51,0,0,0,121,0,0,0,60,0,169,0,80,0,134,0,229,0,186,0,200,0,4,0,0,0,189,0,236,0,0,0,194,0,0,0,130,0,37,0,0,0,0,0,208,0,214,0,0,0,130,0,92,0,0,0,189,0,178,0,127,0,67,0,164,0,12,0,89,0,0,0,226,0,202,0,115,0,233,0,181,0,121,0,0,0,88,0,67,0,50,0,0,0,75,0,89,0,0,0,159,0,0,0,84,0,4,0,13,0,150,0,0,0,185,0,236,0,171,0,18,0,80,0,197,0,66,0,0,0,207,0,159,0,121,0,174,0,42,0,233,0,94,0,196,0,83,0,166,0,72,0,159,0,0,0,150,0,198,0,39,0,182,0,52,0,127,0,0,0,0,0,0,0,225,0,241,0,153,0,20,0,76,0,36,0,162,0,117,0,29,0,32,0,126,0,62,0,122,0,0,0,0,0,91,0,147,0,70,0,247,0,36,0,163,0,84,0,0,0,204,0,0,0,134,0,229,0,154,0,203,0,140,0,232,0,0,0,0,0,197,0,5,0,0,0,51,0,103,0,106,0,36,0,138,0,0,0,184,0,6,0,211,0,0,0,47,0,163,0,0,0,0,0,0,0,134,0,4,0);
signal scenario_full  : scenario_type := (93,31,87,31,50,31,150,31,222,31,222,30,246,31,32,31,163,31,81,31,213,31,228,31,45,31,45,30,133,31,133,30,204,31,204,30,228,31,228,30,18,31,18,30,99,31,195,31,121,31,136,31,226,31,143,31,28,31,28,30,242,31,46,31,51,31,138,31,28,31,197,31,83,31,224,31,91,31,45,31,241,31,241,30,174,31,82,31,213,31,198,31,198,30,214,31,43,31,246,31,111,31,111,30,111,29,111,28,98,31,242,31,13,31,13,30,13,29,189,31,202,31,189,31,143,31,174,31,233,31,130,31,130,30,230,31,79,31,173,31,173,30,113,31,46,31,157,31,172,31,172,30,102,31,130,31,3,31,40,31,59,31,116,31,253,31,79,31,180,31,108,31,108,30,206,31,251,31,248,31,248,30,248,29,248,28,166,31,166,30,221,31,131,31,171,31,185,31,143,31,118,31,27,31,234,31,158,31,101,31,219,31,97,31,106,31,106,30,147,31,189,31,73,31,73,30,119,31,17,31,198,31,163,31,163,30,163,29,80,31,80,30,117,31,117,30,189,31,5,31,39,31,39,30,205,31,109,31,24,31,119,31,119,30,238,31,238,30,204,31,147,31,147,30,43,31,43,30,245,31,13,31,29,31,248,31,131,31,69,31,31,31,31,30,31,29,31,28,109,31,224,31,105,31,105,30,105,29,159,31,64,31,64,30,39,31,39,30,226,31,202,31,204,31,160,31,57,31,209,31,213,31,19,31,47,31,131,31,111,31,138,31,87,31,221,31,17,31,125,31,134,31,61,31,169,31,5,31,153,31,164,31,173,31,187,31,215,31,215,30,215,29,215,28,97,31,73,31,20,31,20,30,23,31,23,30,222,31,222,30,222,29,230,31,230,30,230,29,230,28,220,31,131,31,89,31,102,31,23,31,192,31,192,30,134,31,233,31,8,31,212,31,212,30,212,29,212,28,139,31,180,31,180,30,205,31,205,30,35,31,124,31,11,31,120,31,121,31,120,31,173,31,86,31,87,31,181,31,152,31,152,30,137,31,152,31,36,31,196,31,40,31,202,31,30,31,128,31,94,31,81,31,81,30,98,31,64,31,91,31,146,31,18,31,137,31,137,30,137,29,166,31,6,31,165,31,76,31,76,31,76,30,152,31,101,31,36,31,10,31,162,31,186,31,186,30,186,29,237,31,4,31,4,30,239,31,171,31,138,31,209,31,209,30,217,31,185,31,222,31,152,31,88,31,8,31,107,31,107,30,191,31,76,31,22,31,241,31,76,31,239,31,113,31,113,30,113,29,195,31,195,30,227,31,227,30,164,31,51,31,116,31,187,31,114,31,144,31,170,31,170,30,250,31,103,31,95,31,217,31,213,31,139,31,254,31,109,31,109,30,248,31,73,31,192,31,175,31,180,31,175,31,37,31,215,31,215,30,71,31,166,31,158,31,124,31,124,30,169,31,244,31,132,31,132,30,221,31,230,31,178,31,50,31,212,31,210,31,210,30,40,31,2,31,2,30,104,31,68,31,215,31,178,31,137,31,137,30,33,31,22,31,161,31,161,30,150,31,172,31,172,30,51,31,51,30,121,31,121,30,60,31,169,31,80,31,134,31,229,31,186,31,200,31,4,31,4,30,189,31,236,31,236,30,194,31,194,30,130,31,37,31,37,30,37,29,208,31,214,31,214,30,130,31,92,31,92,30,189,31,178,31,127,31,67,31,164,31,12,31,89,31,89,30,226,31,202,31,115,31,233,31,181,31,121,31,121,30,88,31,67,31,50,31,50,30,75,31,89,31,89,30,159,31,159,30,84,31,4,31,13,31,150,31,150,30,185,31,236,31,171,31,18,31,80,31,197,31,66,31,66,30,207,31,159,31,121,31,174,31,42,31,233,31,94,31,196,31,83,31,166,31,72,31,159,31,159,30,150,31,198,31,39,31,182,31,52,31,127,31,127,30,127,29,127,28,225,31,241,31,153,31,20,31,76,31,36,31,162,31,117,31,29,31,32,31,126,31,62,31,122,31,122,30,122,29,91,31,147,31,70,31,247,31,36,31,163,31,84,31,84,30,204,31,204,30,134,31,229,31,154,31,203,31,140,31,232,31,232,30,232,29,197,31,5,31,5,30,51,31,103,31,106,31,36,31,138,31,138,30,184,31,6,31,211,31,211,30,47,31,163,31,163,30,163,29,163,28,134,31,4,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
