-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_283 is
end project_tb_283;

architecture project_tb_arch_283 of project_tb_283 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 808;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (72,0,225,0,0,0,220,0,143,0,124,0,248,0,154,0,55,0,166,0,30,0,0,0,1,0,247,0,65,0,100,0,0,0,35,0,61,0,162,0,123,0,166,0,213,0,196,0,60,0,216,0,169,0,16,0,136,0,23,0,146,0,86,0,0,0,9,0,153,0,0,0,0,0,195,0,0,0,155,0,167,0,0,0,129,0,48,0,8,0,0,0,0,0,123,0,80,0,0,0,47,0,237,0,101,0,0,0,101,0,121,0,99,0,236,0,242,0,211,0,145,0,37,0,138,0,242,0,222,0,16,0,0,0,54,0,54,0,147,0,108,0,213,0,176,0,0,0,137,0,161,0,0,0,135,0,182,0,149,0,141,0,141,0,0,0,119,0,231,0,0,0,91,0,246,0,155,0,107,0,116,0,63,0,0,0,103,0,150,0,110,0,200,0,42,0,43,0,26,0,79,0,0,0,25,0,126,0,204,0,0,0,114,0,239,0,246,0,59,0,0,0,126,0,0,0,93,0,101,0,103,0,0,0,165,0,89,0,103,0,119,0,229,0,58,0,200,0,182,0,0,0,93,0,70,0,3,0,86,0,158,0,37,0,229,0,240,0,174,0,0,0,210,0,69,0,103,0,0,0,198,0,220,0,0,0,157,0,235,0,0,0,0,0,0,0,234,0,0,0,43,0,20,0,171,0,0,0,251,0,0,0,205,0,223,0,12,0,0,0,65,0,117,0,108,0,85,0,54,0,2,0,190,0,0,0,184,0,46,0,2,0,0,0,95,0,168,0,0,0,13,0,242,0,50,0,2,0,170,0,155,0,0,0,59,0,59,0,60,0,28,0,160,0,65,0,99,0,232,0,0,0,163,0,5,0,77,0,0,0,194,0,0,0,52,0,33,0,0,0,233,0,8,0,91,0,77,0,145,0,6,0,151,0,0,0,42,0,0,0,139,0,135,0,247,0,0,0,0,0,38,0,58,0,0,0,75,0,25,0,216,0,146,0,205,0,63,0,151,0,93,0,4,0,68,0,218,0,58,0,34,0,0,0,7,0,242,0,0,0,208,0,0,0,80,0,131,0,38,0,3,0,250,0,235,0,104,0,242,0,189,0,53,0,109,0,180,0,165,0,37,0,135,0,249,0,0,0,132,0,140,0,226,0,0,0,4,0,0,0,178,0,11,0,141,0,112,0,241,0,111,0,142,0,224,0,117,0,86,0,0,0,0,0,1,0,95,0,127,0,152,0,59,0,62,0,0,0,148,0,147,0,136,0,157,0,108,0,0,0,0,0,136,0,74,0,0,0,0,0,188,0,235,0,0,0,148,0,107,0,172,0,211,0,248,0,0,0,13,0,165,0,41,0,33,0,132,0,95,0,81,0,22,0,236,0,74,0,93,0,155,0,230,0,114,0,117,0,127,0,219,0,237,0,149,0,102,0,88,0,91,0,204,0,121,0,43,0,0,0,0,0,209,0,68,0,251,0,187,0,0,0,139,0,179,0,19,0,52,0,98,0,45,0,127,0,9,0,166,0,134,0,57,0,0,0,53,0,7,0,191,0,150,0,128,0,251,0,170,0,0,0,0,0,0,0,74,0,98,0,215,0,186,0,233,0,43,0,222,0,178,0,141,0,0,0,180,0,167,0,51,0,250,0,254,0,0,0,29,0,24,0,120,0,4,0,207,0,5,0,2,0,157,0,242,0,0,0,122,0,168,0,0,0,161,0,95,0,181,0,104,0,251,0,165,0,248,0,151,0,28,0,40,0,230,0,136,0,112,0,94,0,226,0,210,0,25,0,215,0,14,0,162,0,12,0,70,0,213,0,121,0,83,0,158,0,122,0,164,0,83,0,77,0,44,0,209,0,155,0,0,0,137,0,127,0,12,0,127,0,75,0,240,0,100,0,154,0,69,0,85,0,105,0,11,0,0,0,238,0,194,0,25,0,141,0,19,0,248,0,214,0,106,0,139,0,19,0,153,0,9,0,18,0,48,0,41,0,143,0,249,0,53,0,0,0,116,0,23,0,113,0,160,0,86,0,213,0,17,0,0,0,187,0,110,0,0,0,0,0,94,0,251,0,5,0,177,0,24,0,82,0,175,0,89,0,131,0,0,0,0,0,116,0,123,0,18,0,253,0,189,0,168,0,244,0,130,0,209,0,0,0,91,0,0,0,102,0,79,0,223,0,21,0,212,0,30,0,170,0,0,0,0,0,0,0,0,0,217,0,3,0,67,0,0,0,107,0,174,0,118,0,0,0,180,0,114,0,178,0,151,0,171,0,228,0,0,0,194,0,173,0,250,0,129,0,8,0,188,0,176,0,6,0,205,0,0,0,248,0,100,0,163,0,52,0,44,0,181,0,0,0,110,0,0,0,0,0,95,0,233,0,203,0,122,0,136,0,246,0,177,0,138,0,115,0,169,0,82,0,0,0,110,0,142,0,0,0,0,0,236,0,0,0,20,0,202,0,40,0,15,0,116,0,236,0,0,0,42,0,0,0,110,0,0,0,83,0,56,0,190,0,232,0,44,0,0,0,4,0,0,0,243,0,161,0,171,0,0,0,0,0,244,0,198,0,76,0,49,0,170,0,81,0,206,0,175,0,96,0,88,0,128,0,26,0,20,0,14,0,39,0,0,0,181,0,193,0,164,0,0,0,0,0,249,0,0,0,0,0,92,0,253,0,0,0,0,0,113,0,221,0,93,0,127,0,164,0,92,0,9,0,0,0,242,0,229,0,125,0,180,0,42,0,105,0,135,0,68,0,0,0,109,0,220,0,69,0,156,0,218,0,0,0,237,0,220,0,233,0,69,0,135,0,234,0,0,0,110,0,77,0,0,0,176,0,217,0,198,0,0,0,0,0,206,0,39,0,121,0,28,0,143,0,95,0,70,0,210,0,133,0,45,0,17,0,0,0,193,0,212,0,185,0,198,0,7,0,64,0,163,0,0,0,235,0,0,0,8,0,151,0,22,0,144,0,75,0,76,0,169,0,13,0,240,0,2,0,46,0,136,0,196,0,143,0,102,0,72,0,43,0,8,0,43,0,0,0,96,0,199,0,127,0,0,0,14,0,0,0,28,0,235,0,187,0,0,0,133,0,0,0,0,0,183,0,206,0,50,0,236,0,134,0,15,0,191,0,187,0,67,0,108,0,138,0,104,0,51,0,0,0,57,0,232,0,150,0,0,0,191,0,150,0,0,0,0,0,0,0,247,0,252,0,0,0,31,0,0,0,21,0,39,0,221,0,233,0,89,0,151,0,0,0,0,0,63,0,111,0,47,0,216,0,112,0,186,0,251,0,98,0,61,0,95,0,215,0,108,0,88,0,33,0,36,0,141,0,0,0,0,0,173,0,15,0,207,0,0,0,33,0,84,0,0,0,214,0,0,0,43,0,174,0,44,0,225,0,202,0,0,0,124,0,0,0,0,0,160,0,193,0,56,0,173,0,86,0,0,0,0,0,0,0,59,0,134,0,146,0,235,0,0,0,42,0,187,0,148,0,56,0,75,0,50,0,28,0,23,0,76,0,102,0,241,0,38,0,3,0,210,0,146,0,126,0,0,0,0,0,24,0,85,0,61,0,145,0,246,0,0,0,83,0,2,0,177,0,205,0,95,0,147,0,37,0);
signal scenario_full  : scenario_type := (72,31,225,31,225,30,220,31,143,31,124,31,248,31,154,31,55,31,166,31,30,31,30,30,1,31,247,31,65,31,100,31,100,30,35,31,61,31,162,31,123,31,166,31,213,31,196,31,60,31,216,31,169,31,16,31,136,31,23,31,146,31,86,31,86,30,9,31,153,31,153,30,153,29,195,31,195,30,155,31,167,31,167,30,129,31,48,31,8,31,8,30,8,29,123,31,80,31,80,30,47,31,237,31,101,31,101,30,101,31,121,31,99,31,236,31,242,31,211,31,145,31,37,31,138,31,242,31,222,31,16,31,16,30,54,31,54,31,147,31,108,31,213,31,176,31,176,30,137,31,161,31,161,30,135,31,182,31,149,31,141,31,141,31,141,30,119,31,231,31,231,30,91,31,246,31,155,31,107,31,116,31,63,31,63,30,103,31,150,31,110,31,200,31,42,31,43,31,26,31,79,31,79,30,25,31,126,31,204,31,204,30,114,31,239,31,246,31,59,31,59,30,126,31,126,30,93,31,101,31,103,31,103,30,165,31,89,31,103,31,119,31,229,31,58,31,200,31,182,31,182,30,93,31,70,31,3,31,86,31,158,31,37,31,229,31,240,31,174,31,174,30,210,31,69,31,103,31,103,30,198,31,220,31,220,30,157,31,235,31,235,30,235,29,235,28,234,31,234,30,43,31,20,31,171,31,171,30,251,31,251,30,205,31,223,31,12,31,12,30,65,31,117,31,108,31,85,31,54,31,2,31,190,31,190,30,184,31,46,31,2,31,2,30,95,31,168,31,168,30,13,31,242,31,50,31,2,31,170,31,155,31,155,30,59,31,59,31,60,31,28,31,160,31,65,31,99,31,232,31,232,30,163,31,5,31,77,31,77,30,194,31,194,30,52,31,33,31,33,30,233,31,8,31,91,31,77,31,145,31,6,31,151,31,151,30,42,31,42,30,139,31,135,31,247,31,247,30,247,29,38,31,58,31,58,30,75,31,25,31,216,31,146,31,205,31,63,31,151,31,93,31,4,31,68,31,218,31,58,31,34,31,34,30,7,31,242,31,242,30,208,31,208,30,80,31,131,31,38,31,3,31,250,31,235,31,104,31,242,31,189,31,53,31,109,31,180,31,165,31,37,31,135,31,249,31,249,30,132,31,140,31,226,31,226,30,4,31,4,30,178,31,11,31,141,31,112,31,241,31,111,31,142,31,224,31,117,31,86,31,86,30,86,29,1,31,95,31,127,31,152,31,59,31,62,31,62,30,148,31,147,31,136,31,157,31,108,31,108,30,108,29,136,31,74,31,74,30,74,29,188,31,235,31,235,30,148,31,107,31,172,31,211,31,248,31,248,30,13,31,165,31,41,31,33,31,132,31,95,31,81,31,22,31,236,31,74,31,93,31,155,31,230,31,114,31,117,31,127,31,219,31,237,31,149,31,102,31,88,31,91,31,204,31,121,31,43,31,43,30,43,29,209,31,68,31,251,31,187,31,187,30,139,31,179,31,19,31,52,31,98,31,45,31,127,31,9,31,166,31,134,31,57,31,57,30,53,31,7,31,191,31,150,31,128,31,251,31,170,31,170,30,170,29,170,28,74,31,98,31,215,31,186,31,233,31,43,31,222,31,178,31,141,31,141,30,180,31,167,31,51,31,250,31,254,31,254,30,29,31,24,31,120,31,4,31,207,31,5,31,2,31,157,31,242,31,242,30,122,31,168,31,168,30,161,31,95,31,181,31,104,31,251,31,165,31,248,31,151,31,28,31,40,31,230,31,136,31,112,31,94,31,226,31,210,31,25,31,215,31,14,31,162,31,12,31,70,31,213,31,121,31,83,31,158,31,122,31,164,31,83,31,77,31,44,31,209,31,155,31,155,30,137,31,127,31,12,31,127,31,75,31,240,31,100,31,154,31,69,31,85,31,105,31,11,31,11,30,238,31,194,31,25,31,141,31,19,31,248,31,214,31,106,31,139,31,19,31,153,31,9,31,18,31,48,31,41,31,143,31,249,31,53,31,53,30,116,31,23,31,113,31,160,31,86,31,213,31,17,31,17,30,187,31,110,31,110,30,110,29,94,31,251,31,5,31,177,31,24,31,82,31,175,31,89,31,131,31,131,30,131,29,116,31,123,31,18,31,253,31,189,31,168,31,244,31,130,31,209,31,209,30,91,31,91,30,102,31,79,31,223,31,21,31,212,31,30,31,170,31,170,30,170,29,170,28,170,27,217,31,3,31,67,31,67,30,107,31,174,31,118,31,118,30,180,31,114,31,178,31,151,31,171,31,228,31,228,30,194,31,173,31,250,31,129,31,8,31,188,31,176,31,6,31,205,31,205,30,248,31,100,31,163,31,52,31,44,31,181,31,181,30,110,31,110,30,110,29,95,31,233,31,203,31,122,31,136,31,246,31,177,31,138,31,115,31,169,31,82,31,82,30,110,31,142,31,142,30,142,29,236,31,236,30,20,31,202,31,40,31,15,31,116,31,236,31,236,30,42,31,42,30,110,31,110,30,83,31,56,31,190,31,232,31,44,31,44,30,4,31,4,30,243,31,161,31,171,31,171,30,171,29,244,31,198,31,76,31,49,31,170,31,81,31,206,31,175,31,96,31,88,31,128,31,26,31,20,31,14,31,39,31,39,30,181,31,193,31,164,31,164,30,164,29,249,31,249,30,249,29,92,31,253,31,253,30,253,29,113,31,221,31,93,31,127,31,164,31,92,31,9,31,9,30,242,31,229,31,125,31,180,31,42,31,105,31,135,31,68,31,68,30,109,31,220,31,69,31,156,31,218,31,218,30,237,31,220,31,233,31,69,31,135,31,234,31,234,30,110,31,77,31,77,30,176,31,217,31,198,31,198,30,198,29,206,31,39,31,121,31,28,31,143,31,95,31,70,31,210,31,133,31,45,31,17,31,17,30,193,31,212,31,185,31,198,31,7,31,64,31,163,31,163,30,235,31,235,30,8,31,151,31,22,31,144,31,75,31,76,31,169,31,13,31,240,31,2,31,46,31,136,31,196,31,143,31,102,31,72,31,43,31,8,31,43,31,43,30,96,31,199,31,127,31,127,30,14,31,14,30,28,31,235,31,187,31,187,30,133,31,133,30,133,29,183,31,206,31,50,31,236,31,134,31,15,31,191,31,187,31,67,31,108,31,138,31,104,31,51,31,51,30,57,31,232,31,150,31,150,30,191,31,150,31,150,30,150,29,150,28,247,31,252,31,252,30,31,31,31,30,21,31,39,31,221,31,233,31,89,31,151,31,151,30,151,29,63,31,111,31,47,31,216,31,112,31,186,31,251,31,98,31,61,31,95,31,215,31,108,31,88,31,33,31,36,31,141,31,141,30,141,29,173,31,15,31,207,31,207,30,33,31,84,31,84,30,214,31,214,30,43,31,174,31,44,31,225,31,202,31,202,30,124,31,124,30,124,29,160,31,193,31,56,31,173,31,86,31,86,30,86,29,86,28,59,31,134,31,146,31,235,31,235,30,42,31,187,31,148,31,56,31,75,31,50,31,28,31,23,31,76,31,102,31,241,31,38,31,3,31,210,31,146,31,126,31,126,30,126,29,24,31,85,31,61,31,145,31,246,31,246,30,83,31,2,31,177,31,205,31,95,31,147,31,37,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
