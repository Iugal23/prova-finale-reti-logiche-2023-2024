-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_496 is
end project_tb_496;

architecture project_tb_arch_496 of project_tb_496 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 664;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,237,0,0,0,175,0,244,0,142,0,220,0,52,0,205,0,126,0,22,0,119,0,0,0,201,0,0,0,0,0,107,0,0,0,116,0,166,0,43,0,117,0,194,0,230,0,26,0,112,0,161,0,93,0,5,0,73,0,0,0,189,0,0,0,143,0,239,0,63,0,0,0,114,0,0,0,69,0,48,0,219,0,126,0,110,0,17,0,177,0,53,0,180,0,34,0,0,0,115,0,194,0,170,0,0,0,220,0,114,0,130,0,26,0,0,0,108,0,75,0,198,0,0,0,0,0,2,0,35,0,179,0,23,0,53,0,211,0,161,0,37,0,233,0,255,0,55,0,202,0,154,0,191,0,175,0,114,0,89,0,253,0,71,0,49,0,0,0,0,0,0,0,0,0,154,0,246,0,227,0,210,0,55,0,171,0,0,0,19,0,141,0,248,0,143,0,0,0,161,0,24,0,190,0,66,0,125,0,67,0,94,0,203,0,0,0,146,0,45,0,214,0,156,0,122,0,174,0,199,0,194,0,0,0,52,0,82,0,192,0,56,0,179,0,0,0,111,0,109,0,0,0,149,0,19,0,0,0,54,0,55,0,104,0,199,0,10,0,60,0,104,0,0,0,73,0,0,0,195,0,0,0,0,0,129,0,192,0,0,0,150,0,159,0,0,0,3,0,0,0,0,0,0,0,227,0,203,0,159,0,106,0,244,0,225,0,18,0,225,0,237,0,4,0,162,0,84,0,0,0,0,0,98,0,84,0,249,0,141,0,118,0,121,0,173,0,240,0,167,0,199,0,109,0,117,0,115,0,131,0,175,0,0,0,206,0,6,0,0,0,56,0,0,0,0,0,252,0,144,0,218,0,149,0,25,0,119,0,119,0,183,0,0,0,230,0,6,0,0,0,80,0,204,0,166,0,192,0,29,0,39,0,0,0,30,0,224,0,227,0,106,0,208,0,195,0,76,0,226,0,39,0,0,0,8,0,7,0,34,0,119,0,0,0,251,0,249,0,177,0,164,0,83,0,141,0,216,0,187,0,75,0,0,0,180,0,114,0,157,0,0,0,0,0,28,0,100,0,0,0,211,0,0,0,32,0,0,0,254,0,0,0,27,0,118,0,190,0,186,0,102,0,139,0,72,0,0,0,223,0,186,0,82,0,236,0,247,0,0,0,174,0,113,0,44,0,120,0,21,0,243,0,80,0,0,0,143,0,183,0,120,0,174,0,202,0,119,0,5,0,213,0,0,0,0,0,201,0,154,0,180,0,18,0,145,0,40,0,203,0,7,0,111,0,92,0,169,0,0,0,78,0,10,0,237,0,33,0,240,0,130,0,0,0,252,0,0,0,145,0,55,0,124,0,68,0,0,0,84,0,68,0,219,0,245,0,200,0,6,0,106,0,205,0,217,0,219,0,0,0,3,0,81,0,71,0,0,0,152,0,162,0,0,0,162,0,19,0,192,0,114,0,0,0,95,0,236,0,0,0,217,0,0,0,154,0,233,0,78,0,112,0,198,0,102,0,147,0,99,0,0,0,65,0,0,0,0,0,202,0,30,0,0,0,0,0,0,0,0,0,0,0,147,0,0,0,0,0,33,0,177,0,177,0,100,0,166,0,5,0,0,0,25,0,220,0,98,0,90,0,146,0,95,0,40,0,119,0,0,0,79,0,133,0,22,0,106,0,80,0,243,0,218,0,95,0,0,0,0,0,129,0,114,0,177,0,0,0,0,0,0,0,255,0,214,0,87,0,55,0,255,0,0,0,245,0,85,0,142,0,154,0,15,0,0,0,183,0,0,0,73,0,39,0,0,0,147,0,245,0,183,0,29,0,148,0,114,0,41,0,25,0,0,0,172,0,90,0,85,0,57,0,0,0,163,0,211,0,26,0,91,0,18,0,18,0,59,0,211,0,189,0,0,0,101,0,11,0,218,0,0,0,255,0,119,0,0,0,202,0,130,0,239,0,164,0,77,0,102,0,175,0,32,0,0,0,187,0,15,0,80,0,6,0,135,0,0,0,0,0,156,0,176,0,0,0,108,0,202,0,152,0,205,0,92,0,207,0,251,0,0,0,190,0,103,0,206,0,0,0,6,0,161,0,41,0,105,0,104,0,0,0,253,0,0,0,86,0,174,0,98,0,177,0,75,0,95,0,92,0,78,0,213,0,0,0,0,0,100,0,52,0,40,0,0,0,47,0,179,0,21,0,110,0,0,0,241,0,119,0,207,0,167,0,178,0,220,0,47,0,27,0,107,0,64,0,0,0,96,0,96,0,217,0,190,0,102,0,46,0,162,0,0,0,202,0,0,0,40,0,37,0,222,0,0,0,253,0,177,0,0,0,0,0,0,0,0,0,152,0,218,0,129,0,84,0,253,0,149,0,211,0,79,0,0,0,56,0,173,0,0,0,129,0,84,0,172,0,243,0,248,0,32,0,204,0,39,0,160,0,111,0,0,0,31,0,0,0,0,0,179,0,120,0,176,0,102,0,135,0,47,0,64,0,28,0,230,0,186,0,0,0,106,0,233,0,60,0,222,0,98,0,243,0,44,0,0,0,120,0,200,0,72,0,25,0,64,0,192,0,75,0,84,0,248,0,205,0,218,0,116,0,118,0,107,0,233,0,254,0,239,0,138,0,198,0,0,0,164,0,42,0,44,0,0,0,116,0,40,0,192,0,247,0,175,0,32,0,18,0,0,0,0,0,21,0,221,0,97,0,68,0,235,0,74,0,4,0,180,0,46,0,139,0,193,0,201,0,8,0,119,0,0,0,199,0,224,0,95,0,85,0,97,0,185,0,0,0,207,0,20,0,48,0,0,0,231,0,0,0,96,0,0,0,0,0,94,0,110,0,0,0,0,0,0,0,89,0,185,0,96,0,122,0,221,0,0,0,166,0,31,0,210,0,245,0,6,0,118,0,11,0,31,0,167,0,139,0,121,0,0,0,114,0,220,0,94,0,0,0,176,0,216,0,140,0);
signal scenario_full  : scenario_type := (189,31,237,31,237,30,175,31,244,31,142,31,220,31,52,31,205,31,126,31,22,31,119,31,119,30,201,31,201,30,201,29,107,31,107,30,116,31,166,31,43,31,117,31,194,31,230,31,26,31,112,31,161,31,93,31,5,31,73,31,73,30,189,31,189,30,143,31,239,31,63,31,63,30,114,31,114,30,69,31,48,31,219,31,126,31,110,31,17,31,177,31,53,31,180,31,34,31,34,30,115,31,194,31,170,31,170,30,220,31,114,31,130,31,26,31,26,30,108,31,75,31,198,31,198,30,198,29,2,31,35,31,179,31,23,31,53,31,211,31,161,31,37,31,233,31,255,31,55,31,202,31,154,31,191,31,175,31,114,31,89,31,253,31,71,31,49,31,49,30,49,29,49,28,49,27,154,31,246,31,227,31,210,31,55,31,171,31,171,30,19,31,141,31,248,31,143,31,143,30,161,31,24,31,190,31,66,31,125,31,67,31,94,31,203,31,203,30,146,31,45,31,214,31,156,31,122,31,174,31,199,31,194,31,194,30,52,31,82,31,192,31,56,31,179,31,179,30,111,31,109,31,109,30,149,31,19,31,19,30,54,31,55,31,104,31,199,31,10,31,60,31,104,31,104,30,73,31,73,30,195,31,195,30,195,29,129,31,192,31,192,30,150,31,159,31,159,30,3,31,3,30,3,29,3,28,227,31,203,31,159,31,106,31,244,31,225,31,18,31,225,31,237,31,4,31,162,31,84,31,84,30,84,29,98,31,84,31,249,31,141,31,118,31,121,31,173,31,240,31,167,31,199,31,109,31,117,31,115,31,131,31,175,31,175,30,206,31,6,31,6,30,56,31,56,30,56,29,252,31,144,31,218,31,149,31,25,31,119,31,119,31,183,31,183,30,230,31,6,31,6,30,80,31,204,31,166,31,192,31,29,31,39,31,39,30,30,31,224,31,227,31,106,31,208,31,195,31,76,31,226,31,39,31,39,30,8,31,7,31,34,31,119,31,119,30,251,31,249,31,177,31,164,31,83,31,141,31,216,31,187,31,75,31,75,30,180,31,114,31,157,31,157,30,157,29,28,31,100,31,100,30,211,31,211,30,32,31,32,30,254,31,254,30,27,31,118,31,190,31,186,31,102,31,139,31,72,31,72,30,223,31,186,31,82,31,236,31,247,31,247,30,174,31,113,31,44,31,120,31,21,31,243,31,80,31,80,30,143,31,183,31,120,31,174,31,202,31,119,31,5,31,213,31,213,30,213,29,201,31,154,31,180,31,18,31,145,31,40,31,203,31,7,31,111,31,92,31,169,31,169,30,78,31,10,31,237,31,33,31,240,31,130,31,130,30,252,31,252,30,145,31,55,31,124,31,68,31,68,30,84,31,68,31,219,31,245,31,200,31,6,31,106,31,205,31,217,31,219,31,219,30,3,31,81,31,71,31,71,30,152,31,162,31,162,30,162,31,19,31,192,31,114,31,114,30,95,31,236,31,236,30,217,31,217,30,154,31,233,31,78,31,112,31,198,31,102,31,147,31,99,31,99,30,65,31,65,30,65,29,202,31,30,31,30,30,30,29,30,28,30,27,30,26,147,31,147,30,147,29,33,31,177,31,177,31,100,31,166,31,5,31,5,30,25,31,220,31,98,31,90,31,146,31,95,31,40,31,119,31,119,30,79,31,133,31,22,31,106,31,80,31,243,31,218,31,95,31,95,30,95,29,129,31,114,31,177,31,177,30,177,29,177,28,255,31,214,31,87,31,55,31,255,31,255,30,245,31,85,31,142,31,154,31,15,31,15,30,183,31,183,30,73,31,39,31,39,30,147,31,245,31,183,31,29,31,148,31,114,31,41,31,25,31,25,30,172,31,90,31,85,31,57,31,57,30,163,31,211,31,26,31,91,31,18,31,18,31,59,31,211,31,189,31,189,30,101,31,11,31,218,31,218,30,255,31,119,31,119,30,202,31,130,31,239,31,164,31,77,31,102,31,175,31,32,31,32,30,187,31,15,31,80,31,6,31,135,31,135,30,135,29,156,31,176,31,176,30,108,31,202,31,152,31,205,31,92,31,207,31,251,31,251,30,190,31,103,31,206,31,206,30,6,31,161,31,41,31,105,31,104,31,104,30,253,31,253,30,86,31,174,31,98,31,177,31,75,31,95,31,92,31,78,31,213,31,213,30,213,29,100,31,52,31,40,31,40,30,47,31,179,31,21,31,110,31,110,30,241,31,119,31,207,31,167,31,178,31,220,31,47,31,27,31,107,31,64,31,64,30,96,31,96,31,217,31,190,31,102,31,46,31,162,31,162,30,202,31,202,30,40,31,37,31,222,31,222,30,253,31,177,31,177,30,177,29,177,28,177,27,152,31,218,31,129,31,84,31,253,31,149,31,211,31,79,31,79,30,56,31,173,31,173,30,129,31,84,31,172,31,243,31,248,31,32,31,204,31,39,31,160,31,111,31,111,30,31,31,31,30,31,29,179,31,120,31,176,31,102,31,135,31,47,31,64,31,28,31,230,31,186,31,186,30,106,31,233,31,60,31,222,31,98,31,243,31,44,31,44,30,120,31,200,31,72,31,25,31,64,31,192,31,75,31,84,31,248,31,205,31,218,31,116,31,118,31,107,31,233,31,254,31,239,31,138,31,198,31,198,30,164,31,42,31,44,31,44,30,116,31,40,31,192,31,247,31,175,31,32,31,18,31,18,30,18,29,21,31,221,31,97,31,68,31,235,31,74,31,4,31,180,31,46,31,139,31,193,31,201,31,8,31,119,31,119,30,199,31,224,31,95,31,85,31,97,31,185,31,185,30,207,31,20,31,48,31,48,30,231,31,231,30,96,31,96,30,96,29,94,31,110,31,110,30,110,29,110,28,89,31,185,31,96,31,122,31,221,31,221,30,166,31,31,31,210,31,245,31,6,31,118,31,11,31,31,31,167,31,139,31,121,31,121,30,114,31,220,31,94,31,94,30,176,31,216,31,140,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
