-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 860;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (231,0,39,0,4,0,120,0,0,0,64,0,0,0,0,0,143,0,149,0,120,0,96,0,89,0,234,0,153,0,149,0,178,0,168,0,236,0,184,0,10,0,18,0,220,0,229,0,236,0,160,0,21,0,147,0,167,0,233,0,67,0,241,0,171,0,117,0,135,0,0,0,229,0,97,0,2,0,76,0,10,0,0,0,77,0,217,0,96,0,164,0,0,0,226,0,67,0,30,0,2,0,227,0,240,0,240,0,65,0,31,0,4,0,0,0,115,0,184,0,177,0,0,0,139,0,139,0,122,0,0,0,124,0,252,0,210,0,0,0,247,0,73,0,61,0,3,0,116,0,218,0,112,0,188,0,38,0,163,0,154,0,0,0,131,0,209,0,167,0,74,0,1,0,203,0,23,0,24,0,19,0,12,0,0,0,0,0,25,0,189,0,126,0,108,0,108,0,231,0,129,0,71,0,22,0,222,0,237,0,34,0,122,0,104,0,162,0,0,0,159,0,144,0,28,0,238,0,250,0,125,0,177,0,0,0,0,0,223,0,184,0,200,0,45,0,140,0,146,0,27,0,161,0,162,0,94,0,0,0,15,0,85,0,134,0,77,0,238,0,79,0,155,0,162,0,16,0,221,0,15,0,58,0,71,0,40,0,83,0,220,0,125,0,158,0,247,0,237,0,219,0,155,0,244,0,73,0,82,0,22,0,133,0,104,0,106,0,172,0,175,0,0,0,0,0,214,0,195,0,0,0,0,0,147,0,224,0,0,0,44,0,135,0,115,0,0,0,202,0,106,0,214,0,98,0,0,0,201,0,155,0,191,0,0,0,201,0,138,0,110,0,62,0,138,0,216,0,0,0,138,0,191,0,0,0,144,0,149,0,237,0,15,0,189,0,116,0,104,0,196,0,0,0,171,0,81,0,53,0,81,0,0,0,42,0,13,0,166,0,0,0,223,0,230,0,209,0,70,0,105,0,201,0,235,0,206,0,77,0,216,0,58,0,124,0,109,0,144,0,0,0,174,0,0,0,47,0,127,0,0,0,28,0,0,0,0,0,0,0,23,0,195,0,49,0,213,0,251,0,41,0,0,0,131,0,2,0,39,0,247,0,119,0,158,0,190,0,174,0,220,0,0,0,89,0,131,0,96,0,0,0,0,0,157,0,0,0,192,0,0,0,71,0,0,0,0,0,97,0,53,0,111,0,241,0,0,0,251,0,12,0,142,0,0,0,0,0,0,0,12,0,160,0,251,0,0,0,91,0,192,0,213,0,172,0,228,0,73,0,20,0,232,0,65,0,169,0,94,0,193,0,0,0,245,0,0,0,43,0,0,0,130,0,0,0,219,0,200,0,0,0,91,0,57,0,42,0,106,0,69,0,83,0,49,0,0,0,53,0,217,0,102,0,154,0,193,0,203,0,203,0,27,0,0,0,50,0,107,0,226,0,59,0,131,0,79,0,113,0,153,0,155,0,224,0,96,0,0,0,142,0,51,0,223,0,0,0,233,0,204,0,0,0,128,0,0,0,68,0,107,0,203,0,6,0,87,0,0,0,0,0,92,0,218,0,32,0,239,0,43,0,128,0,61,0,0,0,234,0,177,0,89,0,0,0,163,0,152,0,155,0,16,0,255,0,40,0,143,0,102,0,191,0,175,0,181,0,130,0,207,0,21,0,96,0,154,0,139,0,79,0,138,0,221,0,63,0,0,0,0,0,62,0,0,0,51,0,14,0,55,0,214,0,95,0,30,0,242,0,122,0,242,0,94,0,60,0,211,0,222,0,27,0,251,0,0,0,251,0,250,0,237,0,113,0,177,0,179,0,0,0,46,0,0,0,221,0,194,0,252,0,136,0,82,0,221,0,245,0,178,0,52,0,198,0,201,0,47,0,219,0,249,0,44,0,148,0,78,0,141,0,0,0,1,0,0,0,40,0,0,0,184,0,30,0,0,0,95,0,54,0,62,0,242,0,0,0,88,0,192,0,240,0,234,0,20,0,233,0,139,0,161,0,248,0,155,0,111,0,111,0,0,0,46,0,168,0,0,0,45,0,45,0,36,0,54,0,0,0,6,0,152,0,81,0,131,0,73,0,203,0,83,0,0,0,0,0,0,0,165,0,26,0,233,0,21,0,0,0,74,0,0,0,0,0,14,0,160,0,193,0,228,0,78,0,99,0,126,0,131,0,185,0,0,0,51,0,0,0,143,0,0,0,0,0,179,0,55,0,0,0,124,0,249,0,250,0,0,0,97,0,0,0,26,0,149,0,99,0,224,0,0,0,75,0,100,0,161,0,0,0,79,0,50,0,54,0,74,0,132,0,42,0,60,0,0,0,248,0,193,0,211,0,75,0,22,0,206,0,152,0,0,0,101,0,0,0,41,0,244,0,235,0,27,0,0,0,228,0,0,0,17,0,12,0,21,0,173,0,32,0,19,0,176,0,178,0,92,0,0,0,0,0,195,0,225,0,243,0,87,0,159,0,237,0,111,0,255,0,0,0,0,0,242,0,47,0,229,0,113,0,51,0,0,0,0,0,127,0,208,0,199,0,143,0,254,0,200,0,74,0,225,0,101,0,217,0,0,0,176,0,225,0,0,0,0,0,160,0,177,0,171,0,230,0,93,0,0,0,189,0,200,0,87,0,126,0,22,0,0,0,16,0,95,0,76,0,64,0,219,0,79,0,247,0,14,0,137,0,0,0,9,0,0,0,117,0,117,0,32,0,0,0,0,0,0,0,96,0,0,0,34,0,100,0,228,0,189,0,241,0,0,0,123,0,102,0,97,0,231,0,14,0,218,0,121,0,157,0,152,0,0,0,135,0,6,0,154,0,209,0,33,0,0,0,246,0,17,0,12,0,162,0,115,0,154,0,148,0,16,0,81,0,204,0,132,0,134,0,161,0,153,0,22,0,156,0,0,0,159,0,0,0,217,0,99,0,23,0,220,0,196,0,180,0,30,0,152,0,204,0,0,0,227,0,39,0,224,0,10,0,190,0,120,0,34,0,68,0,206,0,121,0,167,0,237,0,255,0,104,0,114,0,218,0,0,0,48,0,70,0,69,0,148,0,88,0,0,0,0,0,113,0,92,0,200,0,98,0,244,0,90,0,238,0,160,0,0,0,216,0,7,0,0,0,84,0,132,0,0,0,7,0,5,0,0,0,228,0,0,0,0,0,37,0,54,0,170,0,124,0,181,0,160,0,96,0,83,0,169,0,206,0,0,0,129,0,221,0,185,0,179,0,0,0,0,0,208,0,218,0,106,0,86,0,48,0,82,0,205,0,0,0,150,0,0,0,224,0,0,0,0,0,0,0,34,0,0,0,38,0,47,0,192,0,69,0,245,0,83,0,0,0,176,0,0,0,174,0,11,0,0,0,205,0,0,0,0,0,240,0,0,0,0,0,2,0,28,0,96,0,23,0,182,0,0,0,249,0,180,0,3,0,248,0,0,0,221,0,0,0,180,0,83,0,16,0,62,0,187,0,174,0,1,0,105,0,181,0,52,0,0,0,40,0,0,0,182,0,32,0,26,0,0,0,0,0,210,0,179,0,0,0,8,0,113,0,119,0,142,0,176,0,0,0,144,0,0,0,0,0,230,0,36,0,37,0,151,0,206,0,203,0,207,0,0,0,93,0,241,0,0,0,49,0,151,0,0,0,163,0,198,0,121,0,77,0,72,0,221,0,0,0,40,0,42,0,0,0,0,0,24,0,21,0,89,0,87,0,0,0,248,0,0,0,53,0,0,0,163,0,35,0,158,0,33,0,0,0,80,0,138,0,128,0,249,0,160,0,10,0,218,0,0,0,111,0,130,0,60,0,13,0,25,0,233,0,128,0,43,0,186,0,142,0,231,0,0,0);
signal scenario_full  : scenario_type := (231,31,39,31,4,31,120,31,120,30,64,31,64,30,64,29,143,31,149,31,120,31,96,31,89,31,234,31,153,31,149,31,178,31,168,31,236,31,184,31,10,31,18,31,220,31,229,31,236,31,160,31,21,31,147,31,167,31,233,31,67,31,241,31,171,31,117,31,135,31,135,30,229,31,97,31,2,31,76,31,10,31,10,30,77,31,217,31,96,31,164,31,164,30,226,31,67,31,30,31,2,31,227,31,240,31,240,31,65,31,31,31,4,31,4,30,115,31,184,31,177,31,177,30,139,31,139,31,122,31,122,30,124,31,252,31,210,31,210,30,247,31,73,31,61,31,3,31,116,31,218,31,112,31,188,31,38,31,163,31,154,31,154,30,131,31,209,31,167,31,74,31,1,31,203,31,23,31,24,31,19,31,12,31,12,30,12,29,25,31,189,31,126,31,108,31,108,31,231,31,129,31,71,31,22,31,222,31,237,31,34,31,122,31,104,31,162,31,162,30,159,31,144,31,28,31,238,31,250,31,125,31,177,31,177,30,177,29,223,31,184,31,200,31,45,31,140,31,146,31,27,31,161,31,162,31,94,31,94,30,15,31,85,31,134,31,77,31,238,31,79,31,155,31,162,31,16,31,221,31,15,31,58,31,71,31,40,31,83,31,220,31,125,31,158,31,247,31,237,31,219,31,155,31,244,31,73,31,82,31,22,31,133,31,104,31,106,31,172,31,175,31,175,30,175,29,214,31,195,31,195,30,195,29,147,31,224,31,224,30,44,31,135,31,115,31,115,30,202,31,106,31,214,31,98,31,98,30,201,31,155,31,191,31,191,30,201,31,138,31,110,31,62,31,138,31,216,31,216,30,138,31,191,31,191,30,144,31,149,31,237,31,15,31,189,31,116,31,104,31,196,31,196,30,171,31,81,31,53,31,81,31,81,30,42,31,13,31,166,31,166,30,223,31,230,31,209,31,70,31,105,31,201,31,235,31,206,31,77,31,216,31,58,31,124,31,109,31,144,31,144,30,174,31,174,30,47,31,127,31,127,30,28,31,28,30,28,29,28,28,23,31,195,31,49,31,213,31,251,31,41,31,41,30,131,31,2,31,39,31,247,31,119,31,158,31,190,31,174,31,220,31,220,30,89,31,131,31,96,31,96,30,96,29,157,31,157,30,192,31,192,30,71,31,71,30,71,29,97,31,53,31,111,31,241,31,241,30,251,31,12,31,142,31,142,30,142,29,142,28,12,31,160,31,251,31,251,30,91,31,192,31,213,31,172,31,228,31,73,31,20,31,232,31,65,31,169,31,94,31,193,31,193,30,245,31,245,30,43,31,43,30,130,31,130,30,219,31,200,31,200,30,91,31,57,31,42,31,106,31,69,31,83,31,49,31,49,30,53,31,217,31,102,31,154,31,193,31,203,31,203,31,27,31,27,30,50,31,107,31,226,31,59,31,131,31,79,31,113,31,153,31,155,31,224,31,96,31,96,30,142,31,51,31,223,31,223,30,233,31,204,31,204,30,128,31,128,30,68,31,107,31,203,31,6,31,87,31,87,30,87,29,92,31,218,31,32,31,239,31,43,31,128,31,61,31,61,30,234,31,177,31,89,31,89,30,163,31,152,31,155,31,16,31,255,31,40,31,143,31,102,31,191,31,175,31,181,31,130,31,207,31,21,31,96,31,154,31,139,31,79,31,138,31,221,31,63,31,63,30,63,29,62,31,62,30,51,31,14,31,55,31,214,31,95,31,30,31,242,31,122,31,242,31,94,31,60,31,211,31,222,31,27,31,251,31,251,30,251,31,250,31,237,31,113,31,177,31,179,31,179,30,46,31,46,30,221,31,194,31,252,31,136,31,82,31,221,31,245,31,178,31,52,31,198,31,201,31,47,31,219,31,249,31,44,31,148,31,78,31,141,31,141,30,1,31,1,30,40,31,40,30,184,31,30,31,30,30,95,31,54,31,62,31,242,31,242,30,88,31,192,31,240,31,234,31,20,31,233,31,139,31,161,31,248,31,155,31,111,31,111,31,111,30,46,31,168,31,168,30,45,31,45,31,36,31,54,31,54,30,6,31,152,31,81,31,131,31,73,31,203,31,83,31,83,30,83,29,83,28,165,31,26,31,233,31,21,31,21,30,74,31,74,30,74,29,14,31,160,31,193,31,228,31,78,31,99,31,126,31,131,31,185,31,185,30,51,31,51,30,143,31,143,30,143,29,179,31,55,31,55,30,124,31,249,31,250,31,250,30,97,31,97,30,26,31,149,31,99,31,224,31,224,30,75,31,100,31,161,31,161,30,79,31,50,31,54,31,74,31,132,31,42,31,60,31,60,30,248,31,193,31,211,31,75,31,22,31,206,31,152,31,152,30,101,31,101,30,41,31,244,31,235,31,27,31,27,30,228,31,228,30,17,31,12,31,21,31,173,31,32,31,19,31,176,31,178,31,92,31,92,30,92,29,195,31,225,31,243,31,87,31,159,31,237,31,111,31,255,31,255,30,255,29,242,31,47,31,229,31,113,31,51,31,51,30,51,29,127,31,208,31,199,31,143,31,254,31,200,31,74,31,225,31,101,31,217,31,217,30,176,31,225,31,225,30,225,29,160,31,177,31,171,31,230,31,93,31,93,30,189,31,200,31,87,31,126,31,22,31,22,30,16,31,95,31,76,31,64,31,219,31,79,31,247,31,14,31,137,31,137,30,9,31,9,30,117,31,117,31,32,31,32,30,32,29,32,28,96,31,96,30,34,31,100,31,228,31,189,31,241,31,241,30,123,31,102,31,97,31,231,31,14,31,218,31,121,31,157,31,152,31,152,30,135,31,6,31,154,31,209,31,33,31,33,30,246,31,17,31,12,31,162,31,115,31,154,31,148,31,16,31,81,31,204,31,132,31,134,31,161,31,153,31,22,31,156,31,156,30,159,31,159,30,217,31,99,31,23,31,220,31,196,31,180,31,30,31,152,31,204,31,204,30,227,31,39,31,224,31,10,31,190,31,120,31,34,31,68,31,206,31,121,31,167,31,237,31,255,31,104,31,114,31,218,31,218,30,48,31,70,31,69,31,148,31,88,31,88,30,88,29,113,31,92,31,200,31,98,31,244,31,90,31,238,31,160,31,160,30,216,31,7,31,7,30,84,31,132,31,132,30,7,31,5,31,5,30,228,31,228,30,228,29,37,31,54,31,170,31,124,31,181,31,160,31,96,31,83,31,169,31,206,31,206,30,129,31,221,31,185,31,179,31,179,30,179,29,208,31,218,31,106,31,86,31,48,31,82,31,205,31,205,30,150,31,150,30,224,31,224,30,224,29,224,28,34,31,34,30,38,31,47,31,192,31,69,31,245,31,83,31,83,30,176,31,176,30,174,31,11,31,11,30,205,31,205,30,205,29,240,31,240,30,240,29,2,31,28,31,96,31,23,31,182,31,182,30,249,31,180,31,3,31,248,31,248,30,221,31,221,30,180,31,83,31,16,31,62,31,187,31,174,31,1,31,105,31,181,31,52,31,52,30,40,31,40,30,182,31,32,31,26,31,26,30,26,29,210,31,179,31,179,30,8,31,113,31,119,31,142,31,176,31,176,30,144,31,144,30,144,29,230,31,36,31,37,31,151,31,206,31,203,31,207,31,207,30,93,31,241,31,241,30,49,31,151,31,151,30,163,31,198,31,121,31,77,31,72,31,221,31,221,30,40,31,42,31,42,30,42,29,24,31,21,31,89,31,87,31,87,30,248,31,248,30,53,31,53,30,163,31,35,31,158,31,33,31,33,30,80,31,138,31,128,31,249,31,160,31,10,31,218,31,218,30,111,31,130,31,60,31,13,31,25,31,233,31,128,31,43,31,186,31,142,31,231,31,231,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
