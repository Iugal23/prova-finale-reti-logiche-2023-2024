-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_243 is
end project_tb_243;

architecture project_tb_arch_243 of project_tb_243 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 570;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (126,0,23,0,0,0,152,0,24,0,128,0,184,0,64,0,126,0,237,0,139,0,152,0,237,0,154,0,32,0,132,0,253,0,82,0,0,0,135,0,8,0,69,0,252,0,218,0,165,0,143,0,0,0,220,0,0,0,19,0,122,0,0,0,0,0,14,0,0,0,168,0,253,0,29,0,138,0,0,0,177,0,54,0,156,0,127,0,23,0,219,0,65,0,29,0,237,0,176,0,93,0,0,0,58,0,133,0,38,0,0,0,123,0,210,0,70,0,123,0,111,0,231,0,247,0,219,0,123,0,0,0,236,0,48,0,133,0,44,0,200,0,101,0,236,0,136,0,0,0,0,0,0,0,146,0,18,0,230,0,0,0,0,0,12,0,161,0,52,0,147,0,20,0,212,0,4,0,138,0,0,0,52,0,137,0,40,0,245,0,96,0,118,0,251,0,229,0,32,0,106,0,145,0,0,0,170,0,0,0,98,0,0,0,234,0,0,0,108,0,0,0,192,0,64,0,226,0,180,0,0,0,164,0,103,0,87,0,49,0,62,0,30,0,89,0,205,0,9,0,0,0,0,0,28,0,92,0,225,0,141,0,196,0,74,0,0,0,96,0,55,0,0,0,15,0,170,0,155,0,78,0,182,0,2,0,185,0,167,0,0,0,128,0,71,0,165,0,0,0,110,0,127,0,51,0,205,0,134,0,0,0,83,0,0,0,61,0,104,0,110,0,61,0,0,0,30,0,0,0,36,0,0,0,8,0,106,0,108,0,100,0,236,0,22,0,168,0,203,0,6,0,64,0,173,0,189,0,130,0,0,0,138,0,70,0,132,0,0,0,29,0,52,0,134,0,125,0,92,0,93,0,208,0,236,0,158,0,73,0,55,0,229,0,160,0,0,0,170,0,25,0,0,0,141,0,8,0,187,0,160,0,200,0,0,0,134,0,217,0,0,0,14,0,243,0,243,0,0,0,148,0,96,0,58,0,156,0,26,0,0,0,90,0,94,0,128,0,208,0,0,0,219,0,130,0,129,0,0,0,135,0,251,0,227,0,0,0,151,0,156,0,106,0,37,0,0,0,120,0,122,0,0,0,75,0,0,0,5,0,232,0,248,0,244,0,64,0,88,0,215,0,173,0,138,0,0,0,28,0,112,0,0,0,9,0,223,0,42,0,122,0,175,0,0,0,170,0,223,0,3,0,0,0,202,0,78,0,43,0,0,0,0,0,93,0,21,0,30,0,156,0,122,0,92,0,218,0,136,0,0,0,0,0,0,0,61,0,159,0,176,0,117,0,0,0,0,0,80,0,29,0,86,0,168,0,0,0,0,0,68,0,139,0,26,0,0,0,0,0,2,0,140,0,0,0,213,0,83,0,76,0,42,0,84,0,0,0,73,0,210,0,127,0,186,0,206,0,0,0,23,0,130,0,251,0,150,0,36,0,232,0,244,0,90,0,174,0,89,0,220,0,0,0,171,0,159,0,49,0,78,0,179,0,20,0,138,0,2,0,107,0,141,0,144,0,187,0,219,0,226,0,143,0,43,0,0,0,83,0,149,0,147,0,58,0,180,0,254,0,120,0,205,0,150,0,91,0,66,0,74,0,198,0,211,0,201,0,0,0,243,0,0,0,200,0,220,0,252,0,96,0,145,0,214,0,105,0,0,0,187,0,12,0,0,0,13,0,116,0,20,0,158,0,0,0,254,0,18,0,85,0,0,0,210,0,205,0,5,0,0,0,159,0,87,0,0,0,156,0,107,0,17,0,208,0,6,0,170,0,73,0,198,0,0,0,60,0,0,0,8,0,245,0,68,0,252,0,0,0,0,0,85,0,0,0,35,0,179,0,0,0,187,0,52,0,206,0,211,0,106,0,51,0,234,0,36,0,253,0,53,0,119,0,163,0,187,0,132,0,0,0,100,0,76,0,247,0,170,0,0,0,81,0,198,0,214,0,0,0,182,0,235,0,76,0,130,0,140,0,45,0,123,0,23,0,59,0,0,0,36,0,12,0,27,0,31,0,44,0,199,0,121,0,228,0,224,0,173,0,0,0,130,0,161,0,0,0,205,0,105,0,147,0,184,0,113,0,162,0,0,0,135,0,0,0,178,0,255,0,215,0,109,0,225,0,122,0,194,0,0,0,106,0,185,0,57,0,0,0,101,0,0,0,133,0,0,0,160,0,49,0,171,0,72,0,222,0,0,0,118,0,0,0,210,0,3,0,178,0,122,0,0,0,169,0,0,0,0,0,181,0,168,0,93,0,211,0,197,0,59,0,0,0,242,0,13,0,84,0,234,0,144,0,184,0,78,0,0,0,48,0,0,0,242,0,0,0,246,0,132,0,0,0,5,0,199,0,162,0,21,0,169,0,255,0,64,0,68,0,206,0,63,0,226,0,137,0,0,0,0,0,67,0,95,0,0,0,192,0,138,0,144,0,119,0,167,0,121,0,127,0,33,0,0,0,198,0,172,0,9,0,28,0,242,0,0,0,0,0,240,0,123,0,253,0,0,0,53,0,11,0,47,0,110,0,86,0,169,0,186,0,0,0,171,0,106,0,150,0);
signal scenario_full  : scenario_type := (126,31,23,31,23,30,152,31,24,31,128,31,184,31,64,31,126,31,237,31,139,31,152,31,237,31,154,31,32,31,132,31,253,31,82,31,82,30,135,31,8,31,69,31,252,31,218,31,165,31,143,31,143,30,220,31,220,30,19,31,122,31,122,30,122,29,14,31,14,30,168,31,253,31,29,31,138,31,138,30,177,31,54,31,156,31,127,31,23,31,219,31,65,31,29,31,237,31,176,31,93,31,93,30,58,31,133,31,38,31,38,30,123,31,210,31,70,31,123,31,111,31,231,31,247,31,219,31,123,31,123,30,236,31,48,31,133,31,44,31,200,31,101,31,236,31,136,31,136,30,136,29,136,28,146,31,18,31,230,31,230,30,230,29,12,31,161,31,52,31,147,31,20,31,212,31,4,31,138,31,138,30,52,31,137,31,40,31,245,31,96,31,118,31,251,31,229,31,32,31,106,31,145,31,145,30,170,31,170,30,98,31,98,30,234,31,234,30,108,31,108,30,192,31,64,31,226,31,180,31,180,30,164,31,103,31,87,31,49,31,62,31,30,31,89,31,205,31,9,31,9,30,9,29,28,31,92,31,225,31,141,31,196,31,74,31,74,30,96,31,55,31,55,30,15,31,170,31,155,31,78,31,182,31,2,31,185,31,167,31,167,30,128,31,71,31,165,31,165,30,110,31,127,31,51,31,205,31,134,31,134,30,83,31,83,30,61,31,104,31,110,31,61,31,61,30,30,31,30,30,36,31,36,30,8,31,106,31,108,31,100,31,236,31,22,31,168,31,203,31,6,31,64,31,173,31,189,31,130,31,130,30,138,31,70,31,132,31,132,30,29,31,52,31,134,31,125,31,92,31,93,31,208,31,236,31,158,31,73,31,55,31,229,31,160,31,160,30,170,31,25,31,25,30,141,31,8,31,187,31,160,31,200,31,200,30,134,31,217,31,217,30,14,31,243,31,243,31,243,30,148,31,96,31,58,31,156,31,26,31,26,30,90,31,94,31,128,31,208,31,208,30,219,31,130,31,129,31,129,30,135,31,251,31,227,31,227,30,151,31,156,31,106,31,37,31,37,30,120,31,122,31,122,30,75,31,75,30,5,31,232,31,248,31,244,31,64,31,88,31,215,31,173,31,138,31,138,30,28,31,112,31,112,30,9,31,223,31,42,31,122,31,175,31,175,30,170,31,223,31,3,31,3,30,202,31,78,31,43,31,43,30,43,29,93,31,21,31,30,31,156,31,122,31,92,31,218,31,136,31,136,30,136,29,136,28,61,31,159,31,176,31,117,31,117,30,117,29,80,31,29,31,86,31,168,31,168,30,168,29,68,31,139,31,26,31,26,30,26,29,2,31,140,31,140,30,213,31,83,31,76,31,42,31,84,31,84,30,73,31,210,31,127,31,186,31,206,31,206,30,23,31,130,31,251,31,150,31,36,31,232,31,244,31,90,31,174,31,89,31,220,31,220,30,171,31,159,31,49,31,78,31,179,31,20,31,138,31,2,31,107,31,141,31,144,31,187,31,219,31,226,31,143,31,43,31,43,30,83,31,149,31,147,31,58,31,180,31,254,31,120,31,205,31,150,31,91,31,66,31,74,31,198,31,211,31,201,31,201,30,243,31,243,30,200,31,220,31,252,31,96,31,145,31,214,31,105,31,105,30,187,31,12,31,12,30,13,31,116,31,20,31,158,31,158,30,254,31,18,31,85,31,85,30,210,31,205,31,5,31,5,30,159,31,87,31,87,30,156,31,107,31,17,31,208,31,6,31,170,31,73,31,198,31,198,30,60,31,60,30,8,31,245,31,68,31,252,31,252,30,252,29,85,31,85,30,35,31,179,31,179,30,187,31,52,31,206,31,211,31,106,31,51,31,234,31,36,31,253,31,53,31,119,31,163,31,187,31,132,31,132,30,100,31,76,31,247,31,170,31,170,30,81,31,198,31,214,31,214,30,182,31,235,31,76,31,130,31,140,31,45,31,123,31,23,31,59,31,59,30,36,31,12,31,27,31,31,31,44,31,199,31,121,31,228,31,224,31,173,31,173,30,130,31,161,31,161,30,205,31,105,31,147,31,184,31,113,31,162,31,162,30,135,31,135,30,178,31,255,31,215,31,109,31,225,31,122,31,194,31,194,30,106,31,185,31,57,31,57,30,101,31,101,30,133,31,133,30,160,31,49,31,171,31,72,31,222,31,222,30,118,31,118,30,210,31,3,31,178,31,122,31,122,30,169,31,169,30,169,29,181,31,168,31,93,31,211,31,197,31,59,31,59,30,242,31,13,31,84,31,234,31,144,31,184,31,78,31,78,30,48,31,48,30,242,31,242,30,246,31,132,31,132,30,5,31,199,31,162,31,21,31,169,31,255,31,64,31,68,31,206,31,63,31,226,31,137,31,137,30,137,29,67,31,95,31,95,30,192,31,138,31,144,31,119,31,167,31,121,31,127,31,33,31,33,30,198,31,172,31,9,31,28,31,242,31,242,30,242,29,240,31,123,31,253,31,253,30,53,31,11,31,47,31,110,31,86,31,169,31,186,31,186,30,171,31,106,31,150,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
