-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_997 is
end project_tb_997;

architecture project_tb_arch_997 of project_tb_997 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 601;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,251,0,0,0,193,0,0,0,233,0,0,0,184,0,114,0,202,0,54,0,23,0,22,0,186,0,134,0,0,0,89,0,82,0,0,0,130,0,0,0,0,0,193,0,202,0,18,0,224,0,0,0,7,0,2,0,196,0,0,0,5,0,91,0,0,0,0,0,102,0,55,0,37,0,130,0,237,0,100,0,141,0,61,0,0,0,0,0,191,0,141,0,245,0,204,0,0,0,239,0,40,0,209,0,254,0,189,0,0,0,70,0,0,0,55,0,149,0,217,0,188,0,75,0,0,0,176,0,0,0,234,0,0,0,158,0,85,0,0,0,0,0,25,0,161,0,25,0,195,0,0,0,0,0,238,0,0,0,103,0,68,0,0,0,148,0,0,0,110,0,143,0,128,0,223,0,31,0,161,0,0,0,183,0,76,0,110,0,0,0,0,0,183,0,183,0,203,0,21,0,0,0,0,0,189,0,16,0,180,0,214,0,162,0,0,0,181,0,0,0,75,0,87,0,5,0,151,0,140,0,0,0,19,0,25,0,0,0,176,0,0,0,227,0,240,0,0,0,100,0,5,0,72,0,0,0,214,0,10,0,82,0,15,0,80,0,135,0,0,0,245,0,189,0,24,0,106,0,8,0,60,0,172,0,139,0,0,0,0,0,52,0,146,0,83,0,236,0,12,0,50,0,158,0,0,0,130,0,114,0,251,0,205,0,115,0,30,0,85,0,0,0,94,0,9,0,83,0,169,0,88,0,0,0,0,0,0,0,185,0,25,0,70,0,58,0,0,0,66,0,0,0,42,0,49,0,59,0,0,0,0,0,0,0,0,0,118,0,42,0,58,0,166,0,247,0,205,0,154,0,141,0,30,0,111,0,69,0,180,0,40,0,79,0,74,0,171,0,191,0,212,0,151,0,129,0,183,0,81,0,0,0,58,0,162,0,25,0,0,0,205,0,200,0,179,0,231,0,0,0,232,0,63,0,156,0,9,0,0,0,240,0,111,0,200,0,0,0,144,0,0,0,44,0,85,0,253,0,2,0,0,0,11,0,223,0,20,0,0,0,54,0,221,0,0,0,212,0,232,0,93,0,238,0,32,0,21,0,146,0,0,0,0,0,246,0,0,0,107,0,111,0,0,0,187,0,81,0,84,0,31,0,239,0,3,0,163,0,69,0,197,0,237,0,13,0,25,0,32,0,247,0,24,0,178,0,0,0,210,0,90,0,0,0,199,0,38,0,0,0,104,0,0,0,61,0,177,0,69,0,241,0,105,0,108,0,67,0,0,0,154,0,177,0,157,0,110,0,193,0,72,0,0,0,78,0,26,0,155,0,68,0,0,0,161,0,138,0,152,0,97,0,244,0,142,0,35,0,175,0,245,0,0,0,185,0,180,0,0,0,0,0,80,0,54,0,2,0,186,0,0,0,117,0,0,0,90,0,52,0,0,0,29,0,217,0,204,0,76,0,131,0,44,0,68,0,25,0,168,0,0,0,137,0,0,0,246,0,174,0,29,0,192,0,146,0,59,0,46,0,0,0,229,0,112,0,250,0,0,0,72,0,245,0,222,0,153,0,77,0,117,0,11,0,234,0,75,0,84,0,0,0,141,0,4,0,106,0,32,0,97,0,57,0,219,0,122,0,0,0,239,0,0,0,254,0,157,0,0,0,0,0,213,0,0,0,35,0,206,0,82,0,174,0,132,0,43,0,82,0,0,0,192,0,223,0,0,0,32,0,0,0,154,0,168,0,15,0,153,0,179,0,97,0,0,0,0,0,21,0,181,0,63,0,52,0,90,0,0,0,198,0,219,0,0,0,163,0,95,0,8,0,0,0,142,0,196,0,0,0,179,0,143,0,184,0,211,0,165,0,0,0,154,0,146,0,0,0,72,0,184,0,116,0,151,0,95,0,189,0,221,0,0,0,0,0,5,0,172,0,119,0,0,0,119,0,176,0,212,0,193,0,0,0,83,0,102,0,246,0,49,0,0,0,187,0,164,0,159,0,225,0,47,0,170,0,54,0,119,0,237,0,0,0,96,0,0,0,44,0,25,0,164,0,81,0,2,0,0,0,224,0,0,0,125,0,175,0,221,0,245,0,232,0,216,0,209,0,84,0,0,0,0,0,132,0,101,0,152,0,46,0,196,0,99,0,121,0,0,0,161,0,82,0,0,0,30,0,246,0,57,0,79,0,15,0,0,0,70,0,185,0,49,0,189,0,69,0,20,0,63,0,29,0,0,0,40,0,181,0,0,0,184,0,238,0,140,0,51,0,126,0,0,0,0,0,0,0,1,0,0,0,48,0,38,0,172,0,190,0,92,0,204,0,224,0,128,0,51,0,163,0,0,0,0,0,203,0,191,0,0,0,81,0,75,0,0,0,0,0,225,0,154,0,124,0,218,0,4,0,0,0,0,0,193,0,238,0,181,0,93,0,251,0,67,0,52,0,31,0,123,0,0,0,117,0,48,0,254,0,0,0,0,0,70,0,95,0,60,0,0,0,25,0,58,0,23,0,0,0,79,0,163,0,88,0,24,0,198,0,87,0,166,0,0,0,157,0,0,0,149,0,130,0,196,0,100,0,47,0,0,0,63,0,9,0,0,0,0,0,0,0,171,0,72,0,193,0,0,0,0,0,144,0,203,0,122,0,0,0,30,0,178,0,77,0,61,0,0,0,177,0,91,0,107,0,57,0,212,0);
signal scenario_full  : scenario_type := (0,0,251,31,251,30,193,31,193,30,233,31,233,30,184,31,114,31,202,31,54,31,23,31,22,31,186,31,134,31,134,30,89,31,82,31,82,30,130,31,130,30,130,29,193,31,202,31,18,31,224,31,224,30,7,31,2,31,196,31,196,30,5,31,91,31,91,30,91,29,102,31,55,31,37,31,130,31,237,31,100,31,141,31,61,31,61,30,61,29,191,31,141,31,245,31,204,31,204,30,239,31,40,31,209,31,254,31,189,31,189,30,70,31,70,30,55,31,149,31,217,31,188,31,75,31,75,30,176,31,176,30,234,31,234,30,158,31,85,31,85,30,85,29,25,31,161,31,25,31,195,31,195,30,195,29,238,31,238,30,103,31,68,31,68,30,148,31,148,30,110,31,143,31,128,31,223,31,31,31,161,31,161,30,183,31,76,31,110,31,110,30,110,29,183,31,183,31,203,31,21,31,21,30,21,29,189,31,16,31,180,31,214,31,162,31,162,30,181,31,181,30,75,31,87,31,5,31,151,31,140,31,140,30,19,31,25,31,25,30,176,31,176,30,227,31,240,31,240,30,100,31,5,31,72,31,72,30,214,31,10,31,82,31,15,31,80,31,135,31,135,30,245,31,189,31,24,31,106,31,8,31,60,31,172,31,139,31,139,30,139,29,52,31,146,31,83,31,236,31,12,31,50,31,158,31,158,30,130,31,114,31,251,31,205,31,115,31,30,31,85,31,85,30,94,31,9,31,83,31,169,31,88,31,88,30,88,29,88,28,185,31,25,31,70,31,58,31,58,30,66,31,66,30,42,31,49,31,59,31,59,30,59,29,59,28,59,27,118,31,42,31,58,31,166,31,247,31,205,31,154,31,141,31,30,31,111,31,69,31,180,31,40,31,79,31,74,31,171,31,191,31,212,31,151,31,129,31,183,31,81,31,81,30,58,31,162,31,25,31,25,30,205,31,200,31,179,31,231,31,231,30,232,31,63,31,156,31,9,31,9,30,240,31,111,31,200,31,200,30,144,31,144,30,44,31,85,31,253,31,2,31,2,30,11,31,223,31,20,31,20,30,54,31,221,31,221,30,212,31,232,31,93,31,238,31,32,31,21,31,146,31,146,30,146,29,246,31,246,30,107,31,111,31,111,30,187,31,81,31,84,31,31,31,239,31,3,31,163,31,69,31,197,31,237,31,13,31,25,31,32,31,247,31,24,31,178,31,178,30,210,31,90,31,90,30,199,31,38,31,38,30,104,31,104,30,61,31,177,31,69,31,241,31,105,31,108,31,67,31,67,30,154,31,177,31,157,31,110,31,193,31,72,31,72,30,78,31,26,31,155,31,68,31,68,30,161,31,138,31,152,31,97,31,244,31,142,31,35,31,175,31,245,31,245,30,185,31,180,31,180,30,180,29,80,31,54,31,2,31,186,31,186,30,117,31,117,30,90,31,52,31,52,30,29,31,217,31,204,31,76,31,131,31,44,31,68,31,25,31,168,31,168,30,137,31,137,30,246,31,174,31,29,31,192,31,146,31,59,31,46,31,46,30,229,31,112,31,250,31,250,30,72,31,245,31,222,31,153,31,77,31,117,31,11,31,234,31,75,31,84,31,84,30,141,31,4,31,106,31,32,31,97,31,57,31,219,31,122,31,122,30,239,31,239,30,254,31,157,31,157,30,157,29,213,31,213,30,35,31,206,31,82,31,174,31,132,31,43,31,82,31,82,30,192,31,223,31,223,30,32,31,32,30,154,31,168,31,15,31,153,31,179,31,97,31,97,30,97,29,21,31,181,31,63,31,52,31,90,31,90,30,198,31,219,31,219,30,163,31,95,31,8,31,8,30,142,31,196,31,196,30,179,31,143,31,184,31,211,31,165,31,165,30,154,31,146,31,146,30,72,31,184,31,116,31,151,31,95,31,189,31,221,31,221,30,221,29,5,31,172,31,119,31,119,30,119,31,176,31,212,31,193,31,193,30,83,31,102,31,246,31,49,31,49,30,187,31,164,31,159,31,225,31,47,31,170,31,54,31,119,31,237,31,237,30,96,31,96,30,44,31,25,31,164,31,81,31,2,31,2,30,224,31,224,30,125,31,175,31,221,31,245,31,232,31,216,31,209,31,84,31,84,30,84,29,132,31,101,31,152,31,46,31,196,31,99,31,121,31,121,30,161,31,82,31,82,30,30,31,246,31,57,31,79,31,15,31,15,30,70,31,185,31,49,31,189,31,69,31,20,31,63,31,29,31,29,30,40,31,181,31,181,30,184,31,238,31,140,31,51,31,126,31,126,30,126,29,126,28,1,31,1,30,48,31,38,31,172,31,190,31,92,31,204,31,224,31,128,31,51,31,163,31,163,30,163,29,203,31,191,31,191,30,81,31,75,31,75,30,75,29,225,31,154,31,124,31,218,31,4,31,4,30,4,29,193,31,238,31,181,31,93,31,251,31,67,31,52,31,31,31,123,31,123,30,117,31,48,31,254,31,254,30,254,29,70,31,95,31,60,31,60,30,25,31,58,31,23,31,23,30,79,31,163,31,88,31,24,31,198,31,87,31,166,31,166,30,157,31,157,30,149,31,130,31,196,31,100,31,47,31,47,30,63,31,9,31,9,30,9,29,9,28,171,31,72,31,193,31,193,30,193,29,144,31,203,31,122,31,122,30,30,31,178,31,77,31,61,31,61,30,177,31,91,31,107,31,57,31,212,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
