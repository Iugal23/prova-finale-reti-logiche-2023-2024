-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_927 is
end project_tb_927;

architecture project_tb_arch_927 of project_tb_927 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 969;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (63,0,0,0,0,0,129,0,79,0,2,0,163,0,197,0,235,0,0,0,62,0,218,0,79,0,225,0,194,0,166,0,196,0,81,0,66,0,162,0,179,0,0,0,134,0,126,0,224,0,93,0,0,0,213,0,223,0,104,0,145,0,172,0,132,0,229,0,228,0,183,0,184,0,81,0,224,0,226,0,40,0,44,0,2,0,0,0,227,0,162,0,194,0,0,0,171,0,73,0,0,0,134,0,64,0,43,0,103,0,12,0,31,0,91,0,73,0,188,0,231,0,111,0,61,0,37,0,218,0,85,0,129,0,117,0,205,0,30,0,0,0,190,0,245,0,43,0,255,0,205,0,0,0,151,0,0,0,25,0,0,0,89,0,120,0,173,0,233,0,173,0,195,0,8,0,40,0,230,0,227,0,253,0,205,0,0,0,50,0,150,0,0,0,23,0,0,0,112,0,0,0,141,0,216,0,108,0,17,0,147,0,98,0,0,0,77,0,7,0,177,0,72,0,146,0,94,0,131,0,149,0,0,0,114,0,92,0,0,0,174,0,196,0,107,0,0,0,109,0,171,0,192,0,0,0,141,0,52,0,0,0,0,0,176,0,239,0,80,0,231,0,101,0,137,0,164,0,0,0,157,0,0,0,238,0,196,0,86,0,0,0,114,0,34,0,0,0,217,0,149,0,0,0,70,0,0,0,129,0,215,0,225,0,126,0,86,0,213,0,92,0,113,0,199,0,182,0,179,0,137,0,7,0,199,0,206,0,171,0,217,0,181,0,0,0,70,0,47,0,183,0,190,0,181,0,154,0,16,0,215,0,203,0,171,0,0,0,162,0,0,0,122,0,200,0,174,0,0,0,2,0,98,0,136,0,0,0,0,0,189,0,172,0,35,0,143,0,74,0,196,0,126,0,0,0,51,0,0,0,118,0,14,0,0,0,253,0,0,0,43,0,0,0,238,0,226,0,76,0,97,0,160,0,41,0,179,0,10,0,158,0,88,0,194,0,253,0,19,0,0,0,104,0,0,0,52,0,0,0,38,0,170,0,198,0,0,0,57,0,136,0,121,0,100,0,124,0,228,0,226,0,0,0,0,0,20,0,0,0,174,0,205,0,205,0,253,0,100,0,82,0,114,0,79,0,224,0,181,0,0,0,0,0,167,0,244,0,131,0,193,0,196,0,0,0,0,0,249,0,232,0,66,0,154,0,8,0,28,0,82,0,0,0,141,0,56,0,103,0,188,0,236,0,0,0,220,0,0,0,199,0,160,0,121,0,0,0,13,0,136,0,62,0,255,0,153,0,165,0,240,0,19,0,115,0,9,0,182,0,255,0,112,0,60,0,219,0,16,0,83,0,0,0,192,0,36,0,0,0,28,0,66,0,0,0,0,0,49,0,0,0,24,0,91,0,47,0,24,0,142,0,61,0,237,0,248,0,76,0,254,0,248,0,204,0,168,0,102,0,179,0,0,0,171,0,167,0,0,0,0,0,13,0,0,0,72,0,66,0,27,0,16,0,80,0,16,0,209,0,41,0,0,0,0,0,196,0,171,0,112,0,195,0,141,0,40,0,32,0,75,0,43,0,0,0,0,0,167,0,55,0,248,0,103,0,243,0,253,0,56,0,244,0,0,0,0,0,13,0,250,0,0,0,202,0,253,0,198,0,119,0,0,0,43,0,165,0,159,0,145,0,123,0,55,0,21,0,195,0,0,0,179,0,136,0,88,0,84,0,0,0,217,0,0,0,4,0,100,0,0,0,114,0,14,0,165,0,0,0,150,0,0,0,128,0,241,0,0,0,0,0,81,0,80,0,55,0,0,0,0,0,128,0,233,0,11,0,243,0,237,0,27,0,36,0,242,0,192,0,50,0,99,0,0,0,0,0,86,0,43,0,124,0,0,0,0,0,28,0,189,0,153,0,124,0,184,0,0,0,133,0,68,0,229,0,75,0,0,0,0,0,193,0,0,0,0,0,34,0,142,0,30,0,129,0,0,0,171,0,72,0,0,0,0,0,142,0,131,0,35,0,133,0,0,0,148,0,0,0,160,0,139,0,106,0,0,0,0,0,14,0,84,0,69,0,86,0,123,0,0,0,0,0,254,0,165,0,154,0,155,0,203,0,162,0,19,0,103,0,36,0,92,0,225,0,196,0,0,0,83,0,0,0,171,0,243,0,0,0,0,0,28,0,156,0,0,0,97,0,205,0,183,0,93,0,52,0,0,0,26,0,195,0,0,0,0,0,127,0,106,0,168,0,99,0,65,0,194,0,68,0,0,0,28,0,104,0,0,0,201,0,0,0,60,0,17,0,0,0,88,0,253,0,125,0,176,0,24,0,0,0,154,0,0,0,195,0,212,0,102,0,202,0,243,0,244,0,0,0,157,0,7,0,0,0,143,0,29,0,0,0,7,0,0,0,205,0,0,0,0,0,79,0,0,0,123,0,210,0,18,0,160,0,173,0,0,0,84,0,228,0,236,0,109,0,43,0,183,0,0,0,201,0,21,0,15,0,0,0,182,0,84,0,105,0,193,0,91,0,252,0,0,0,15,0,235,0,207,0,202,0,119,0,139,0,115,0,0,0,24,0,31,0,0,0,161,0,0,0,197,0,121,0,65,0,68,0,68,0,221,0,5,0,100,0,247,0,236,0,211,0,166,0,15,0,0,0,146,0,178,0,81,0,122,0,148,0,103,0,166,0,29,0,216,0,0,0,0,0,0,0,207,0,51,0,41,0,74,0,0,0,35,0,155,0,143,0,101,0,242,0,64,0,0,0,252,0,0,0,245,0,0,0,0,0,194,0,45,0,45,0,166,0,122,0,212,0,0,0,183,0,204,0,255,0,253,0,252,0,0,0,136,0,0,0,120,0,133,0,0,0,104,0,158,0,10,0,253,0,84,0,111,0,47,0,215,0,9,0,18,0,111,0,124,0,112,0,0,0,83,0,0,0,0,0,57,0,99,0,158,0,12,0,16,0,197,0,222,0,124,0,77,0,183,0,201,0,24,0,93,0,25,0,49,0,78,0,108,0,245,0,170,0,229,0,34,0,189,0,165,0,28,0,0,0,0,0,52,0,63,0,146,0,213,0,144,0,96,0,226,0,31,0,62,0,0,0,0,0,40,0,88,0,102,0,36,0,0,0,0,0,144,0,101,0,66,0,3,0,0,0,184,0,119,0,163,0,6,0,184,0,247,0,121,0,132,0,70,0,0,0,0,0,161,0,221,0,189,0,104,0,216,0,19,0,80,0,17,0,67,0,60,0,0,0,4,0,66,0,0,0,114,0,176,0,0,0,45,0,73,0,228,0,133,0,0,0,89,0,40,0,207,0,94,0,36,0,194,0,175,0,0,0,153,0,147,0,213,0,95,0,146,0,179,0,11,0,118,0,0,0,47,0,0,0,171,0,67,0,0,0,119,0,83,0,44,0,226,0,0,0,0,0,123,0,0,0,0,0,0,0,185,0,91,0,178,0,206,0,73,0,62,0,218,0,243,0,153,0,57,0,0,0,0,0,217,0,153,0,0,0,93,0,0,0,235,0,183,0,52,0,200,0,0,0,87,0,161,0,0,0,170,0,128,0,214,0,76,0,32,0,65,0,158,0,150,0,89,0,123,0,204,0,79,0,43,0,83,0,203,0,0,0,95,0,254,0,230,0,3,0,216,0,225,0,0,0,76,0,106,0,135,0,159,0,32,0,123,0,46,0,0,0,121,0,0,0,186,0,46,0,0,0,33,0,237,0,144,0,174,0,0,0,245,0,92,0,135,0,91,0,248,0,237,0,252,0,116,0,0,0,231,0,193,0,206,0,225,0,224,0,2,0,0,0,160,0,0,0,81,0,128,0,15,0,0,0,0,0,81,0,173,0,132,0,214,0,0,0,87,0,9,0,150,0,0,0,0,0,62,0,132,0,0,0,156,0,239,0,95,0,0,0,251,0,144,0,0,0,0,0,218,0,142,0,47,0,0,0,240,0,4,0,209,0,151,0,38,0,193,0,104,0,230,0,0,0,12,0,0,0,45,0,198,0,128,0,0,0,137,0,0,0,138,0,238,0,0,0,0,0,59,0,195,0,216,0,44,0,227,0,154,0,41,0,14,0,230,0,81,0,0,0,0,0,49,0,56,0,44,0,9,0,156,0,0,0,0,0,150,0,200,0,0,0,240,0,100,0,215,0,57,0,230,0,102,0,173,0,254,0,86,0,0,0,123,0,122,0,247,0,243,0,170,0,109,0,161,0,224,0,224,0,17,0,2,0,53,0,0,0,146,0,0,0,227,0,0,0,67,0,0,0,145,0,0,0,10,0,0,0,169,0,0,0,83,0,0,0,0,0,0,0,131,0,106,0);
signal scenario_full  : scenario_type := (63,31,63,30,63,29,129,31,79,31,2,31,163,31,197,31,235,31,235,30,62,31,218,31,79,31,225,31,194,31,166,31,196,31,81,31,66,31,162,31,179,31,179,30,134,31,126,31,224,31,93,31,93,30,213,31,223,31,104,31,145,31,172,31,132,31,229,31,228,31,183,31,184,31,81,31,224,31,226,31,40,31,44,31,2,31,2,30,227,31,162,31,194,31,194,30,171,31,73,31,73,30,134,31,64,31,43,31,103,31,12,31,31,31,91,31,73,31,188,31,231,31,111,31,61,31,37,31,218,31,85,31,129,31,117,31,205,31,30,31,30,30,190,31,245,31,43,31,255,31,205,31,205,30,151,31,151,30,25,31,25,30,89,31,120,31,173,31,233,31,173,31,195,31,8,31,40,31,230,31,227,31,253,31,205,31,205,30,50,31,150,31,150,30,23,31,23,30,112,31,112,30,141,31,216,31,108,31,17,31,147,31,98,31,98,30,77,31,7,31,177,31,72,31,146,31,94,31,131,31,149,31,149,30,114,31,92,31,92,30,174,31,196,31,107,31,107,30,109,31,171,31,192,31,192,30,141,31,52,31,52,30,52,29,176,31,239,31,80,31,231,31,101,31,137,31,164,31,164,30,157,31,157,30,238,31,196,31,86,31,86,30,114,31,34,31,34,30,217,31,149,31,149,30,70,31,70,30,129,31,215,31,225,31,126,31,86,31,213,31,92,31,113,31,199,31,182,31,179,31,137,31,7,31,199,31,206,31,171,31,217,31,181,31,181,30,70,31,47,31,183,31,190,31,181,31,154,31,16,31,215,31,203,31,171,31,171,30,162,31,162,30,122,31,200,31,174,31,174,30,2,31,98,31,136,31,136,30,136,29,189,31,172,31,35,31,143,31,74,31,196,31,126,31,126,30,51,31,51,30,118,31,14,31,14,30,253,31,253,30,43,31,43,30,238,31,226,31,76,31,97,31,160,31,41,31,179,31,10,31,158,31,88,31,194,31,253,31,19,31,19,30,104,31,104,30,52,31,52,30,38,31,170,31,198,31,198,30,57,31,136,31,121,31,100,31,124,31,228,31,226,31,226,30,226,29,20,31,20,30,174,31,205,31,205,31,253,31,100,31,82,31,114,31,79,31,224,31,181,31,181,30,181,29,167,31,244,31,131,31,193,31,196,31,196,30,196,29,249,31,232,31,66,31,154,31,8,31,28,31,82,31,82,30,141,31,56,31,103,31,188,31,236,31,236,30,220,31,220,30,199,31,160,31,121,31,121,30,13,31,136,31,62,31,255,31,153,31,165,31,240,31,19,31,115,31,9,31,182,31,255,31,112,31,60,31,219,31,16,31,83,31,83,30,192,31,36,31,36,30,28,31,66,31,66,30,66,29,49,31,49,30,24,31,91,31,47,31,24,31,142,31,61,31,237,31,248,31,76,31,254,31,248,31,204,31,168,31,102,31,179,31,179,30,171,31,167,31,167,30,167,29,13,31,13,30,72,31,66,31,27,31,16,31,80,31,16,31,209,31,41,31,41,30,41,29,196,31,171,31,112,31,195,31,141,31,40,31,32,31,75,31,43,31,43,30,43,29,167,31,55,31,248,31,103,31,243,31,253,31,56,31,244,31,244,30,244,29,13,31,250,31,250,30,202,31,253,31,198,31,119,31,119,30,43,31,165,31,159,31,145,31,123,31,55,31,21,31,195,31,195,30,179,31,136,31,88,31,84,31,84,30,217,31,217,30,4,31,100,31,100,30,114,31,14,31,165,31,165,30,150,31,150,30,128,31,241,31,241,30,241,29,81,31,80,31,55,31,55,30,55,29,128,31,233,31,11,31,243,31,237,31,27,31,36,31,242,31,192,31,50,31,99,31,99,30,99,29,86,31,43,31,124,31,124,30,124,29,28,31,189,31,153,31,124,31,184,31,184,30,133,31,68,31,229,31,75,31,75,30,75,29,193,31,193,30,193,29,34,31,142,31,30,31,129,31,129,30,171,31,72,31,72,30,72,29,142,31,131,31,35,31,133,31,133,30,148,31,148,30,160,31,139,31,106,31,106,30,106,29,14,31,84,31,69,31,86,31,123,31,123,30,123,29,254,31,165,31,154,31,155,31,203,31,162,31,19,31,103,31,36,31,92,31,225,31,196,31,196,30,83,31,83,30,171,31,243,31,243,30,243,29,28,31,156,31,156,30,97,31,205,31,183,31,93,31,52,31,52,30,26,31,195,31,195,30,195,29,127,31,106,31,168,31,99,31,65,31,194,31,68,31,68,30,28,31,104,31,104,30,201,31,201,30,60,31,17,31,17,30,88,31,253,31,125,31,176,31,24,31,24,30,154,31,154,30,195,31,212,31,102,31,202,31,243,31,244,31,244,30,157,31,7,31,7,30,143,31,29,31,29,30,7,31,7,30,205,31,205,30,205,29,79,31,79,30,123,31,210,31,18,31,160,31,173,31,173,30,84,31,228,31,236,31,109,31,43,31,183,31,183,30,201,31,21,31,15,31,15,30,182,31,84,31,105,31,193,31,91,31,252,31,252,30,15,31,235,31,207,31,202,31,119,31,139,31,115,31,115,30,24,31,31,31,31,30,161,31,161,30,197,31,121,31,65,31,68,31,68,31,221,31,5,31,100,31,247,31,236,31,211,31,166,31,15,31,15,30,146,31,178,31,81,31,122,31,148,31,103,31,166,31,29,31,216,31,216,30,216,29,216,28,207,31,51,31,41,31,74,31,74,30,35,31,155,31,143,31,101,31,242,31,64,31,64,30,252,31,252,30,245,31,245,30,245,29,194,31,45,31,45,31,166,31,122,31,212,31,212,30,183,31,204,31,255,31,253,31,252,31,252,30,136,31,136,30,120,31,133,31,133,30,104,31,158,31,10,31,253,31,84,31,111,31,47,31,215,31,9,31,18,31,111,31,124,31,112,31,112,30,83,31,83,30,83,29,57,31,99,31,158,31,12,31,16,31,197,31,222,31,124,31,77,31,183,31,201,31,24,31,93,31,25,31,49,31,78,31,108,31,245,31,170,31,229,31,34,31,189,31,165,31,28,31,28,30,28,29,52,31,63,31,146,31,213,31,144,31,96,31,226,31,31,31,62,31,62,30,62,29,40,31,88,31,102,31,36,31,36,30,36,29,144,31,101,31,66,31,3,31,3,30,184,31,119,31,163,31,6,31,184,31,247,31,121,31,132,31,70,31,70,30,70,29,161,31,221,31,189,31,104,31,216,31,19,31,80,31,17,31,67,31,60,31,60,30,4,31,66,31,66,30,114,31,176,31,176,30,45,31,73,31,228,31,133,31,133,30,89,31,40,31,207,31,94,31,36,31,194,31,175,31,175,30,153,31,147,31,213,31,95,31,146,31,179,31,11,31,118,31,118,30,47,31,47,30,171,31,67,31,67,30,119,31,83,31,44,31,226,31,226,30,226,29,123,31,123,30,123,29,123,28,185,31,91,31,178,31,206,31,73,31,62,31,218,31,243,31,153,31,57,31,57,30,57,29,217,31,153,31,153,30,93,31,93,30,235,31,183,31,52,31,200,31,200,30,87,31,161,31,161,30,170,31,128,31,214,31,76,31,32,31,65,31,158,31,150,31,89,31,123,31,204,31,79,31,43,31,83,31,203,31,203,30,95,31,254,31,230,31,3,31,216,31,225,31,225,30,76,31,106,31,135,31,159,31,32,31,123,31,46,31,46,30,121,31,121,30,186,31,46,31,46,30,33,31,237,31,144,31,174,31,174,30,245,31,92,31,135,31,91,31,248,31,237,31,252,31,116,31,116,30,231,31,193,31,206,31,225,31,224,31,2,31,2,30,160,31,160,30,81,31,128,31,15,31,15,30,15,29,81,31,173,31,132,31,214,31,214,30,87,31,9,31,150,31,150,30,150,29,62,31,132,31,132,30,156,31,239,31,95,31,95,30,251,31,144,31,144,30,144,29,218,31,142,31,47,31,47,30,240,31,4,31,209,31,151,31,38,31,193,31,104,31,230,31,230,30,12,31,12,30,45,31,198,31,128,31,128,30,137,31,137,30,138,31,238,31,238,30,238,29,59,31,195,31,216,31,44,31,227,31,154,31,41,31,14,31,230,31,81,31,81,30,81,29,49,31,56,31,44,31,9,31,156,31,156,30,156,29,150,31,200,31,200,30,240,31,100,31,215,31,57,31,230,31,102,31,173,31,254,31,86,31,86,30,123,31,122,31,247,31,243,31,170,31,109,31,161,31,224,31,224,31,17,31,2,31,53,31,53,30,146,31,146,30,227,31,227,30,67,31,67,30,145,31,145,30,10,31,10,30,169,31,169,30,83,31,83,30,83,29,83,28,131,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
