-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1004;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,120,0,249,0,76,0,0,0,113,0,97,0,0,0,0,0,243,0,0,0,170,0,180,0,179,0,247,0,0,0,8,0,246,0,180,0,70,0,31,0,107,0,10,0,0,0,68,0,157,0,46,0,247,0,223,0,93,0,196,0,135,0,0,0,77,0,191,0,178,0,0,0,0,0,189,0,227,0,167,0,143,0,62,0,145,0,234,0,230,0,40,0,0,0,129,0,12,0,175,0,190,0,0,0,102,0,0,0,0,0,105,0,195,0,207,0,172,0,0,0,237,0,126,0,90,0,0,0,19,0,45,0,244,0,0,0,184,0,0,0,181,0,136,0,137,0,195,0,44,0,166,0,0,0,105,0,0,0,53,0,6,0,0,0,44,0,201,0,89,0,205,0,162,0,0,0,145,0,177,0,27,0,212,0,53,0,0,0,193,0,0,0,95,0,0,0,60,0,221,0,0,0,225,0,107,0,198,0,160,0,163,0,217,0,111,0,246,0,27,0,210,0,114,0,146,0,22,0,61,0,111,0,171,0,243,0,22,0,98,0,0,0,57,0,0,0,75,0,186,0,193,0,159,0,0,0,178,0,81,0,0,0,169,0,194,0,27,0,0,0,106,0,218,0,0,0,129,0,207,0,0,0,150,0,8,0,121,0,142,0,111,0,43,0,237,0,235,0,229,0,253,0,22,0,164,0,168,0,218,0,0,0,219,0,98,0,160,0,92,0,4,0,212,0,0,0,152,0,49,0,0,0,139,0,23,0,243,0,78,0,40,0,0,0,90,0,181,0,193,0,138,0,235,0,144,0,11,0,4,0,58,0,60,0,53,0,87,0,59,0,0,0,200,0,246,0,97,0,75,0,180,0,11,0,49,0,0,0,22,0,0,0,114,0,36,0,0,0,0,0,29,0,84,0,14,0,231,0,29,0,26,0,97,0,139,0,0,0,18,0,179,0,237,0,199,0,200,0,144,0,28,0,107,0,38,0,0,0,0,0,11,0,224,0,231,0,18,0,150,0,60,0,226,0,6,0,0,0,79,0,234,0,182,0,79,0,152,0,231,0,175,0,0,0,6,0,143,0,83,0,163,0,169,0,175,0,223,0,123,0,178,0,104,0,118,0,139,0,174,0,0,0,213,0,0,0,69,0,152,0,55,0,60,0,48,0,0,0,235,0,113,0,132,0,143,0,154,0,249,0,162,0,237,0,88,0,154,0,28,0,171,0,0,0,232,0,0,0,127,0,164,0,0,0,210,0,82,0,60,0,0,0,241,0,0,0,44,0,154,0,238,0,14,0,147,0,124,0,0,0,85,0,105,0,37,0,238,0,77,0,221,0,190,0,136,0,0,0,59,0,104,0,8,0,218,0,168,0,0,0,198,0,152,0,0,0,0,0,84,0,118,0,0,0,61,0,163,0,46,0,247,0,144,0,0,0,224,0,25,0,107,0,0,0,208,0,57,0,0,0,0,0,0,0,32,0,181,0,221,0,65,0,177,0,178,0,0,0,0,0,6,0,218,0,218,0,223,0,127,0,149,0,114,0,58,0,144,0,116,0,208,0,0,0,99,0,155,0,55,0,199,0,0,0,183,0,79,0,102,0,69,0,0,0,213,0,162,0,0,0,172,0,0,0,76,0,0,0,78,0,44,0,0,0,247,0,11,0,223,0,81,0,194,0,145,0,0,0,206,0,196,0,229,0,170,0,81,0,138,0,0,0,6,0,33,0,105,0,0,0,113,0,19,0,0,0,35,0,184,0,146,0,253,0,144,0,216,0,238,0,12,0,231,0,23,0,47,0,138,0,76,0,236,0,0,0,84,0,234,0,185,0,0,0,62,0,14,0,0,0,71,0,0,0,100,0,120,0,107,0,0,0,122,0,0,0,5,0,219,0,221,0,227,0,214,0,24,0,0,0,42,0,0,0,108,0,0,0,55,0,0,0,97,0,10,0,131,0,131,0,0,0,235,0,230,0,183,0,213,0,18,0,159,0,243,0,86,0,232,0,80,0,0,0,0,0,0,0,0,0,0,0,0,0,31,0,221,0,135,0,35,0,64,0,67,0,131,0,0,0,253,0,16,0,57,0,0,0,0,0,85,0,51,0,138,0,61,0,112,0,137,0,89,0,86,0,200,0,70,0,101,0,106,0,178,0,0,0,0,0,138,0,190,0,247,0,133,0,0,0,68,0,133,0,121,0,28,0,6,0,0,0,89,0,0,0,173,0,58,0,62,0,0,0,71,0,154,0,207,0,88,0,76,0,15,0,0,0,52,0,100,0,79,0,192,0,68,0,133,0,128,0,209,0,0,0,160,0,0,0,131,0,213,0,73,0,31,0,166,0,109,0,104,0,232,0,40,0,152,0,80,0,88,0,0,0,252,0,20,0,153,0,60,0,183,0,117,0,108,0,222,0,95,0,123,0,0,0,235,0,122,0,139,0,54,0,49,0,102,0,88,0,54,0,189,0,223,0,0,0,88,0,165,0,193,0,67,0,165,0,172,0,223,0,198,0,244,0,0,0,144,0,0,0,157,0,53,0,37,0,116,0,117,0,172,0,104,0,0,0,159,0,0,0,166,0,245,0,223,0,0,0,122,0,160,0,22,0,198,0,210,0,0,0,0,0,0,0,167,0,14,0,197,0,76,0,129,0,0,0,117,0,0,0,86,0,0,0,0,0,119,0,0,0,147,0,0,0,105,0,33,0,124,0,150,0,220,0,121,0,0,0,170,0,67,0,0,0,0,0,239,0,165,0,0,0,0,0,193,0,28,0,13,0,27,0,0,0,0,0,164,0,98,0,55,0,143,0,140,0,244,0,26,0,0,0,239,0,0,0,107,0,78,0,182,0,147,0,75,0,0,0,241,0,208,0,0,0,173,0,246,0,117,0,81,0,255,0,225,0,214,0,0,0,166,0,0,0,171,0,203,0,129,0,100,0,11,0,0,0,36,0,169,0,197,0,168,0,159,0,0,0,189,0,82,0,36,0,0,0,220,0,127,0,236,0,147,0,112,0,200,0,47,0,0,0,0,0,0,0,0,0,12,0,128,0,172,0,205,0,180,0,0,0,0,0,32,0,231,0,64,0,25,0,245,0,108,0,238,0,27,0,159,0,253,0,141,0,10,0,207,0,202,0,109,0,139,0,0,0,0,0,0,0,188,0,132,0,199,0,0,0,16,0,205,0,0,0,233,0,0,0,0,0,46,0,192,0,0,0,0,0,177,0,45,0,169,0,0,0,0,0,250,0,184,0,144,0,220,0,183,0,154,0,163,0,8,0,0,0,0,0,228,0,42,0,0,0,0,0,244,0,69,0,124,0,0,0,102,0,0,0,78,0,217,0,230,0,204,0,43,0,181,0,160,0,227,0,64,0,249,0,77,0,228,0,0,0,222,0,119,0,201,0,194,0,148,0,205,0,0,0,0,0,0,0,219,0,0,0,120,0,0,0,0,0,205,0,29,0,158,0,1,0,0,0,2,0,0,0,204,0,224,0,49,0,229,0,0,0,255,0,203,0,112,0,153,0,188,0,42,0,171,0,0,0,223,0,148,0,29,0,21,0,35,0,0,0,186,0,140,0,196,0,0,0,12,0,128,0,137,0,212,0,0,0,93,0,141,0,11,0,103,0,0,0,124,0,147,0,98,0,227,0,148,0,121,0,116,0,224,0,160,0,58,0,249,0,59,0,198,0,189,0,223,0,0,0,194,0,0,0,213,0,144,0,229,0,10,0,0,0,109,0,62,0,114,0,0,0,90,0,238,0,123,0,167,0,231,0,82,0,0,0,94,0,201,0,160,0,63,0,83,0,209,0,156,0,52,0,238,0,200,0,0,0,51,0,99,0,18,0,101,0,32,0,33,0,0,0,254,0,142,0,193,0,27,0,187,0,0,0,39,0,150,0,0,0,0,0,240,0,239,0,66,0,41,0,71,0,49,0,0,0,0,0,0,0,0,0,0,0,132,0,254,0,193,0,150,0,34,0,234,0,230,0,223,0,71,0,187,0,64,0,231,0,246,0,10,0,123,0,184,0,215,0,210,0,138,0,37,0,205,0,82,0,0,0,186,0,30,0,134,0,0,0,52,0,67,0,170,0,110,0,53,0,191,0,246,0,81,0,199,0,199,0,97,0,98,0,134,0,23,0,0,0,120,0,101,0,223,0,114,0,145,0,38,0,0,0,198,0,0,0,0,0,42,0,237,0,9,0,107,0,130,0,0,0,0,0,76,0,51,0,25,0,237,0,171,0,107,0,0,0,152,0,246,0,203,0,0,0,68,0,0,0,0,0,63,0,126,0,178,0,213,0,217,0,3,0,124,0,0,0,164,0,148,0,130,0,166,0,140,0,56,0,0,0,33,0,90,0,0,0,249,0,217,0,167,0,204,0,0,0,148,0,76,0,96,0,0,0,173,0,0,0,0,0,150,0,49,0,3,0,109,0,75,0,0,0,14,0,255,0,127,0,68,0,0,0,4,0,105,0,0,0,226,0,81,0,163,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,120,31,249,31,76,31,76,30,113,31,97,31,97,30,97,29,243,31,243,30,170,31,180,31,179,31,247,31,247,30,8,31,246,31,180,31,70,31,31,31,107,31,10,31,10,30,68,31,157,31,46,31,247,31,223,31,93,31,196,31,135,31,135,30,77,31,191,31,178,31,178,30,178,29,189,31,227,31,167,31,143,31,62,31,145,31,234,31,230,31,40,31,40,30,129,31,12,31,175,31,190,31,190,30,102,31,102,30,102,29,105,31,195,31,207,31,172,31,172,30,237,31,126,31,90,31,90,30,19,31,45,31,244,31,244,30,184,31,184,30,181,31,136,31,137,31,195,31,44,31,166,31,166,30,105,31,105,30,53,31,6,31,6,30,44,31,201,31,89,31,205,31,162,31,162,30,145,31,177,31,27,31,212,31,53,31,53,30,193,31,193,30,95,31,95,30,60,31,221,31,221,30,225,31,107,31,198,31,160,31,163,31,217,31,111,31,246,31,27,31,210,31,114,31,146,31,22,31,61,31,111,31,171,31,243,31,22,31,98,31,98,30,57,31,57,30,75,31,186,31,193,31,159,31,159,30,178,31,81,31,81,30,169,31,194,31,27,31,27,30,106,31,218,31,218,30,129,31,207,31,207,30,150,31,8,31,121,31,142,31,111,31,43,31,237,31,235,31,229,31,253,31,22,31,164,31,168,31,218,31,218,30,219,31,98,31,160,31,92,31,4,31,212,31,212,30,152,31,49,31,49,30,139,31,23,31,243,31,78,31,40,31,40,30,90,31,181,31,193,31,138,31,235,31,144,31,11,31,4,31,58,31,60,31,53,31,87,31,59,31,59,30,200,31,246,31,97,31,75,31,180,31,11,31,49,31,49,30,22,31,22,30,114,31,36,31,36,30,36,29,29,31,84,31,14,31,231,31,29,31,26,31,97,31,139,31,139,30,18,31,179,31,237,31,199,31,200,31,144,31,28,31,107,31,38,31,38,30,38,29,11,31,224,31,231,31,18,31,150,31,60,31,226,31,6,31,6,30,79,31,234,31,182,31,79,31,152,31,231,31,175,31,175,30,6,31,143,31,83,31,163,31,169,31,175,31,223,31,123,31,178,31,104,31,118,31,139,31,174,31,174,30,213,31,213,30,69,31,152,31,55,31,60,31,48,31,48,30,235,31,113,31,132,31,143,31,154,31,249,31,162,31,237,31,88,31,154,31,28,31,171,31,171,30,232,31,232,30,127,31,164,31,164,30,210,31,82,31,60,31,60,30,241,31,241,30,44,31,154,31,238,31,14,31,147,31,124,31,124,30,85,31,105,31,37,31,238,31,77,31,221,31,190,31,136,31,136,30,59,31,104,31,8,31,218,31,168,31,168,30,198,31,152,31,152,30,152,29,84,31,118,31,118,30,61,31,163,31,46,31,247,31,144,31,144,30,224,31,25,31,107,31,107,30,208,31,57,31,57,30,57,29,57,28,32,31,181,31,221,31,65,31,177,31,178,31,178,30,178,29,6,31,218,31,218,31,223,31,127,31,149,31,114,31,58,31,144,31,116,31,208,31,208,30,99,31,155,31,55,31,199,31,199,30,183,31,79,31,102,31,69,31,69,30,213,31,162,31,162,30,172,31,172,30,76,31,76,30,78,31,44,31,44,30,247,31,11,31,223,31,81,31,194,31,145,31,145,30,206,31,196,31,229,31,170,31,81,31,138,31,138,30,6,31,33,31,105,31,105,30,113,31,19,31,19,30,35,31,184,31,146,31,253,31,144,31,216,31,238,31,12,31,231,31,23,31,47,31,138,31,76,31,236,31,236,30,84,31,234,31,185,31,185,30,62,31,14,31,14,30,71,31,71,30,100,31,120,31,107,31,107,30,122,31,122,30,5,31,219,31,221,31,227,31,214,31,24,31,24,30,42,31,42,30,108,31,108,30,55,31,55,30,97,31,10,31,131,31,131,31,131,30,235,31,230,31,183,31,213,31,18,31,159,31,243,31,86,31,232,31,80,31,80,30,80,29,80,28,80,27,80,26,80,25,31,31,221,31,135,31,35,31,64,31,67,31,131,31,131,30,253,31,16,31,57,31,57,30,57,29,85,31,51,31,138,31,61,31,112,31,137,31,89,31,86,31,200,31,70,31,101,31,106,31,178,31,178,30,178,29,138,31,190,31,247,31,133,31,133,30,68,31,133,31,121,31,28,31,6,31,6,30,89,31,89,30,173,31,58,31,62,31,62,30,71,31,154,31,207,31,88,31,76,31,15,31,15,30,52,31,100,31,79,31,192,31,68,31,133,31,128,31,209,31,209,30,160,31,160,30,131,31,213,31,73,31,31,31,166,31,109,31,104,31,232,31,40,31,152,31,80,31,88,31,88,30,252,31,20,31,153,31,60,31,183,31,117,31,108,31,222,31,95,31,123,31,123,30,235,31,122,31,139,31,54,31,49,31,102,31,88,31,54,31,189,31,223,31,223,30,88,31,165,31,193,31,67,31,165,31,172,31,223,31,198,31,244,31,244,30,144,31,144,30,157,31,53,31,37,31,116,31,117,31,172,31,104,31,104,30,159,31,159,30,166,31,245,31,223,31,223,30,122,31,160,31,22,31,198,31,210,31,210,30,210,29,210,28,167,31,14,31,197,31,76,31,129,31,129,30,117,31,117,30,86,31,86,30,86,29,119,31,119,30,147,31,147,30,105,31,33,31,124,31,150,31,220,31,121,31,121,30,170,31,67,31,67,30,67,29,239,31,165,31,165,30,165,29,193,31,28,31,13,31,27,31,27,30,27,29,164,31,98,31,55,31,143,31,140,31,244,31,26,31,26,30,239,31,239,30,107,31,78,31,182,31,147,31,75,31,75,30,241,31,208,31,208,30,173,31,246,31,117,31,81,31,255,31,225,31,214,31,214,30,166,31,166,30,171,31,203,31,129,31,100,31,11,31,11,30,36,31,169,31,197,31,168,31,159,31,159,30,189,31,82,31,36,31,36,30,220,31,127,31,236,31,147,31,112,31,200,31,47,31,47,30,47,29,47,28,47,27,12,31,128,31,172,31,205,31,180,31,180,30,180,29,32,31,231,31,64,31,25,31,245,31,108,31,238,31,27,31,159,31,253,31,141,31,10,31,207,31,202,31,109,31,139,31,139,30,139,29,139,28,188,31,132,31,199,31,199,30,16,31,205,31,205,30,233,31,233,30,233,29,46,31,192,31,192,30,192,29,177,31,45,31,169,31,169,30,169,29,250,31,184,31,144,31,220,31,183,31,154,31,163,31,8,31,8,30,8,29,228,31,42,31,42,30,42,29,244,31,69,31,124,31,124,30,102,31,102,30,78,31,217,31,230,31,204,31,43,31,181,31,160,31,227,31,64,31,249,31,77,31,228,31,228,30,222,31,119,31,201,31,194,31,148,31,205,31,205,30,205,29,205,28,219,31,219,30,120,31,120,30,120,29,205,31,29,31,158,31,1,31,1,30,2,31,2,30,204,31,224,31,49,31,229,31,229,30,255,31,203,31,112,31,153,31,188,31,42,31,171,31,171,30,223,31,148,31,29,31,21,31,35,31,35,30,186,31,140,31,196,31,196,30,12,31,128,31,137,31,212,31,212,30,93,31,141,31,11,31,103,31,103,30,124,31,147,31,98,31,227,31,148,31,121,31,116,31,224,31,160,31,58,31,249,31,59,31,198,31,189,31,223,31,223,30,194,31,194,30,213,31,144,31,229,31,10,31,10,30,109,31,62,31,114,31,114,30,90,31,238,31,123,31,167,31,231,31,82,31,82,30,94,31,201,31,160,31,63,31,83,31,209,31,156,31,52,31,238,31,200,31,200,30,51,31,99,31,18,31,101,31,32,31,33,31,33,30,254,31,142,31,193,31,27,31,187,31,187,30,39,31,150,31,150,30,150,29,240,31,239,31,66,31,41,31,71,31,49,31,49,30,49,29,49,28,49,27,49,26,132,31,254,31,193,31,150,31,34,31,234,31,230,31,223,31,71,31,187,31,64,31,231,31,246,31,10,31,123,31,184,31,215,31,210,31,138,31,37,31,205,31,82,31,82,30,186,31,30,31,134,31,134,30,52,31,67,31,170,31,110,31,53,31,191,31,246,31,81,31,199,31,199,31,97,31,98,31,134,31,23,31,23,30,120,31,101,31,223,31,114,31,145,31,38,31,38,30,198,31,198,30,198,29,42,31,237,31,9,31,107,31,130,31,130,30,130,29,76,31,51,31,25,31,237,31,171,31,107,31,107,30,152,31,246,31,203,31,203,30,68,31,68,30,68,29,63,31,126,31,178,31,213,31,217,31,3,31,124,31,124,30,164,31,148,31,130,31,166,31,140,31,56,31,56,30,33,31,90,31,90,30,249,31,217,31,167,31,204,31,204,30,148,31,76,31,96,31,96,30,173,31,173,30,173,29,150,31,49,31,3,31,109,31,75,31,75,30,14,31,255,31,127,31,68,31,68,30,4,31,105,31,105,30,226,31,81,31,163,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
