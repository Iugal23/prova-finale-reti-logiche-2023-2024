-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 874;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (165,0,131,0,148,0,0,0,181,0,3,0,34,0,252,0,35,0,76,0,116,0,7,0,0,0,0,0,245,0,31,0,100,0,52,0,0,0,0,0,99,0,121,0,209,0,0,0,238,0,216,0,138,0,34,0,170,0,82,0,0,0,0,0,248,0,208,0,169,0,198,0,140,0,58,0,5,0,161,0,161,0,27,0,97,0,224,0,238,0,0,0,30,0,0,0,145,0,0,0,22,0,0,0,64,0,83,0,0,0,156,0,147,0,77,0,21,0,184,0,0,0,0,0,16,0,148,0,43,0,0,0,211,0,1,0,10,0,93,0,211,0,91,0,29,0,108,0,132,0,202,0,88,0,0,0,255,0,175,0,61,0,181,0,90,0,104,0,12,0,172,0,0,0,53,0,248,0,0,0,0,0,96,0,171,0,93,0,199,0,0,0,39,0,27,0,53,0,248,0,224,0,187,0,158,0,157,0,58,0,160,0,252,0,63,0,121,0,27,0,159,0,146,0,149,0,254,0,141,0,152,0,17,0,218,0,0,0,92,0,246,0,223,0,23,0,94,0,0,0,1,0,0,0,23,0,237,0,0,0,0,0,0,0,0,0,5,0,43,0,197,0,22,0,231,0,170,0,0,0,0,0,185,0,0,0,14,0,214,0,0,0,0,0,1,0,213,0,0,0,230,0,155,0,237,0,152,0,90,0,145,0,13,0,0,0,43,0,45,0,0,0,62,0,0,0,226,0,1,0,26,0,95,0,225,0,89,0,84,0,37,0,129,0,74,0,215,0,29,0,185,0,244,0,157,0,8,0,50,0,33,0,168,0,51,0,58,0,234,0,156,0,136,0,245,0,97,0,0,0,239,0,0,0,72,0,92,0,147,0,213,0,106,0,119,0,191,0,54,0,199,0,0,0,10,0,0,0,16,0,150,0,170,0,31,0,0,0,51,0,152,0,177,0,243,0,30,0,134,0,153,0,254,0,154,0,0,0,0,0,162,0,233,0,201,0,0,0,44,0,61,0,192,0,119,0,0,0,146,0,0,0,116,0,20,0,0,0,56,0,75,0,20,0,236,0,247,0,241,0,15,0,149,0,0,0,147,0,30,0,0,0,195,0,213,0,97,0,0,0,164,0,79,0,187,0,103,0,241,0,0,0,80,0,21,0,0,0,0,0,78,0,0,0,126,0,0,0,0,0,0,0,224,0,57,0,0,0,5,0,0,0,0,0,66,0,241,0,207,0,93,0,0,0,168,0,26,0,151,0,49,0,2,0,117,0,48,0,218,0,249,0,0,0,45,0,143,0,0,0,212,0,38,0,200,0,219,0,237,0,151,0,188,0,0,0,128,0,2,0,97,0,39,0,80,0,39,0,6,0,0,0,0,0,205,0,4,0,34,0,190,0,219,0,50,0,99,0,0,0,13,0,132,0,111,0,48,0,0,0,36,0,254,0,138,0,77,0,16,0,30,0,183,0,0,0,0,0,0,0,69,0,228,0,23,0,40,0,62,0,90,0,105,0,0,0,0,0,15,0,0,0,156,0,112,0,164,0,161,0,44,0,18,0,184,0,0,0,98,0,221,0,212,0,229,0,41,0,212,0,47,0,92,0,198,0,0,0,159,0,26,0,45,0,193,0,107,0,86,0,0,0,31,0,200,0,131,0,0,0,0,0,57,0,0,0,124,0,0,0,0,0,220,0,169,0,96,0,164,0,120,0,0,0,194,0,41,0,114,0,0,0,80,0,245,0,98,0,69,0,0,0,2,0,36,0,0,0,35,0,79,0,0,0,206,0,192,0,180,0,26,0,62,0,120,0,30,0,13,0,102,0,172,0,4,0,0,0,147,0,0,0,161,0,0,0,245,0,66,0,67,0,8,0,0,0,110,0,17,0,0,0,168,0,68,0,195,0,30,0,92,0,34,0,15,0,113,0,104,0,0,0,231,0,0,0,226,0,0,0,252,0,0,0,0,0,190,0,147,0,109,0,0,0,62,0,120,0,64,0,103,0,17,0,4,0,214,0,198,0,55,0,186,0,229,0,240,0,85,0,116,0,81,0,0,0,148,0,0,0,160,0,124,0,92,0,198,0,172,0,69,0,0,0,248,0,163,0,17,0,128,0,57,0,0,0,0,0,56,0,79,0,184,0,0,0,58,0,0,0,196,0,0,0,0,0,87,0,10,0,178,0,179,0,46,0,58,0,200,0,119,0,0,0,17,0,103,0,49,0,0,0,123,0,55,0,0,0,9,0,187,0,90,0,150,0,93,0,116,0,205,0,126,0,154,0,55,0,229,0,0,0,69,0,0,0,0,0,59,0,227,0,0,0,34,0,239,0,37,0,127,0,113,0,138,0,143,0,0,0,150,0,126,0,92,0,0,0,39,0,27,0,228,0,67,0,206,0,120,0,19,0,8,0,118,0,48,0,174,0,157,0,224,0,36,0,56,0,33,0,242,0,8,0,35,0,34,0,201,0,112,0,0,0,209,0,188,0,233,0,61,0,200,0,0,0,237,0,1,0,2,0,0,0,0,0,0,0,98,0,0,0,73,0,54,0,252,0,175,0,56,0,117,0,117,0,11,0,122,0,136,0,63,0,168,0,0,0,178,0,223,0,240,0,132,0,127,0,0,0,141,0,182,0,0,0,54,0,12,0,0,0,211,0,3,0,132,0,114,0,122,0,250,0,145,0,127,0,124,0,162,0,2,0,224,0,249,0,4,0,59,0,109,0,0,0,74,0,219,0,107,0,8,0,59,0,10,0,216,0,49,0,37,0,249,0,47,0,43,0,4,0,0,0,245,0,84,0,84,0,60,0,0,0,0,0,41,0,237,0,0,0,0,0,197,0,156,0,133,0,196,0,129,0,0,0,0,0,136,0,130,0,54,0,100,0,11,0,129,0,2,0,0,0,24,0,163,0,171,0,133,0,24,0,148,0,55,0,185,0,166,0,5,0,49,0,138,0,136,0,44,0,30,0,65,0,0,0,74,0,19,0,3,0,191,0,163,0,125,0,139,0,0,0,0,0,92,0,76,0,228,0,0,0,2,0,0,0,0,0,58,0,213,0,188,0,26,0,73,0,139,0,0,0,216,0,171,0,59,0,101,0,178,0,116,0,232,0,254,0,134,0,108,0,247,0,228,0,0,0,0,0,25,0,85,0,173,0,88,0,125,0,160,0,112,0,0,0,0,0,83,0,166,0,100,0,0,0,57,0,196,0,0,0,0,0,223,0,0,0,109,0,0,0,201,0,0,0,92,0,107,0,171,0,75,0,167,0,8,0,198,0,0,0,185,0,30,0,127,0,152,0,206,0,84,0,46,0,196,0,0,0,103,0,155,0,81,0,79,0,45,0,219,0,181,0,4,0,142,0,58,0,0,0,226,0,33,0,205,0,39,0,85,0,115,0,148,0,87,0,219,0,153,0,170,0,8,0,154,0,138,0,174,0,76,0,58,0,221,0,134,0,50,0,19,0,0,0,0,0,0,0,218,0,48,0,108,0,158,0,27,0,215,0,252,0,0,0,91,0,43,0,0,0,63,0,22,0,142,0,125,0,68,0,0,0,14,0,243,0,146,0,21,0,0,0,163,0,238,0,235,0,116,0,236,0,231,0,231,0,88,0,162,0,149,0,0,0,219,0,151,0,187,0,0,0,32,0,115,0,0,0,0,0,0,0,0,0,0,0,40,0,41,0,120,0,248,0,201,0,0,0,241,0,200,0,10,0,171,0,254,0,189,0,0,0,231,0,0,0,136,0,119,0,79,0,0,0,0,0,0,0,47,0,165,0,0,0,199,0,55,0,163,0,89,0,103,0,235,0,44,0,118,0,86,0,0,0,95,0,95,0,0,0,0,0,122,0,63,0,8,0,138,0,106,0,102,0,113,0,213,0,0,0,169,0,140,0,202,0,167,0,149,0,0,0,12,0);
signal scenario_full  : scenario_type := (165,31,131,31,148,31,148,30,181,31,3,31,34,31,252,31,35,31,76,31,116,31,7,31,7,30,7,29,245,31,31,31,100,31,52,31,52,30,52,29,99,31,121,31,209,31,209,30,238,31,216,31,138,31,34,31,170,31,82,31,82,30,82,29,248,31,208,31,169,31,198,31,140,31,58,31,5,31,161,31,161,31,27,31,97,31,224,31,238,31,238,30,30,31,30,30,145,31,145,30,22,31,22,30,64,31,83,31,83,30,156,31,147,31,77,31,21,31,184,31,184,30,184,29,16,31,148,31,43,31,43,30,211,31,1,31,10,31,93,31,211,31,91,31,29,31,108,31,132,31,202,31,88,31,88,30,255,31,175,31,61,31,181,31,90,31,104,31,12,31,172,31,172,30,53,31,248,31,248,30,248,29,96,31,171,31,93,31,199,31,199,30,39,31,27,31,53,31,248,31,224,31,187,31,158,31,157,31,58,31,160,31,252,31,63,31,121,31,27,31,159,31,146,31,149,31,254,31,141,31,152,31,17,31,218,31,218,30,92,31,246,31,223,31,23,31,94,31,94,30,1,31,1,30,23,31,237,31,237,30,237,29,237,28,237,27,5,31,43,31,197,31,22,31,231,31,170,31,170,30,170,29,185,31,185,30,14,31,214,31,214,30,214,29,1,31,213,31,213,30,230,31,155,31,237,31,152,31,90,31,145,31,13,31,13,30,43,31,45,31,45,30,62,31,62,30,226,31,1,31,26,31,95,31,225,31,89,31,84,31,37,31,129,31,74,31,215,31,29,31,185,31,244,31,157,31,8,31,50,31,33,31,168,31,51,31,58,31,234,31,156,31,136,31,245,31,97,31,97,30,239,31,239,30,72,31,92,31,147,31,213,31,106,31,119,31,191,31,54,31,199,31,199,30,10,31,10,30,16,31,150,31,170,31,31,31,31,30,51,31,152,31,177,31,243,31,30,31,134,31,153,31,254,31,154,31,154,30,154,29,162,31,233,31,201,31,201,30,44,31,61,31,192,31,119,31,119,30,146,31,146,30,116,31,20,31,20,30,56,31,75,31,20,31,236,31,247,31,241,31,15,31,149,31,149,30,147,31,30,31,30,30,195,31,213,31,97,31,97,30,164,31,79,31,187,31,103,31,241,31,241,30,80,31,21,31,21,30,21,29,78,31,78,30,126,31,126,30,126,29,126,28,224,31,57,31,57,30,5,31,5,30,5,29,66,31,241,31,207,31,93,31,93,30,168,31,26,31,151,31,49,31,2,31,117,31,48,31,218,31,249,31,249,30,45,31,143,31,143,30,212,31,38,31,200,31,219,31,237,31,151,31,188,31,188,30,128,31,2,31,97,31,39,31,80,31,39,31,6,31,6,30,6,29,205,31,4,31,34,31,190,31,219,31,50,31,99,31,99,30,13,31,132,31,111,31,48,31,48,30,36,31,254,31,138,31,77,31,16,31,30,31,183,31,183,30,183,29,183,28,69,31,228,31,23,31,40,31,62,31,90,31,105,31,105,30,105,29,15,31,15,30,156,31,112,31,164,31,161,31,44,31,18,31,184,31,184,30,98,31,221,31,212,31,229,31,41,31,212,31,47,31,92,31,198,31,198,30,159,31,26,31,45,31,193,31,107,31,86,31,86,30,31,31,200,31,131,31,131,30,131,29,57,31,57,30,124,31,124,30,124,29,220,31,169,31,96,31,164,31,120,31,120,30,194,31,41,31,114,31,114,30,80,31,245,31,98,31,69,31,69,30,2,31,36,31,36,30,35,31,79,31,79,30,206,31,192,31,180,31,26,31,62,31,120,31,30,31,13,31,102,31,172,31,4,31,4,30,147,31,147,30,161,31,161,30,245,31,66,31,67,31,8,31,8,30,110,31,17,31,17,30,168,31,68,31,195,31,30,31,92,31,34,31,15,31,113,31,104,31,104,30,231,31,231,30,226,31,226,30,252,31,252,30,252,29,190,31,147,31,109,31,109,30,62,31,120,31,64,31,103,31,17,31,4,31,214,31,198,31,55,31,186,31,229,31,240,31,85,31,116,31,81,31,81,30,148,31,148,30,160,31,124,31,92,31,198,31,172,31,69,31,69,30,248,31,163,31,17,31,128,31,57,31,57,30,57,29,56,31,79,31,184,31,184,30,58,31,58,30,196,31,196,30,196,29,87,31,10,31,178,31,179,31,46,31,58,31,200,31,119,31,119,30,17,31,103,31,49,31,49,30,123,31,55,31,55,30,9,31,187,31,90,31,150,31,93,31,116,31,205,31,126,31,154,31,55,31,229,31,229,30,69,31,69,30,69,29,59,31,227,31,227,30,34,31,239,31,37,31,127,31,113,31,138,31,143,31,143,30,150,31,126,31,92,31,92,30,39,31,27,31,228,31,67,31,206,31,120,31,19,31,8,31,118,31,48,31,174,31,157,31,224,31,36,31,56,31,33,31,242,31,8,31,35,31,34,31,201,31,112,31,112,30,209,31,188,31,233,31,61,31,200,31,200,30,237,31,1,31,2,31,2,30,2,29,2,28,98,31,98,30,73,31,54,31,252,31,175,31,56,31,117,31,117,31,11,31,122,31,136,31,63,31,168,31,168,30,178,31,223,31,240,31,132,31,127,31,127,30,141,31,182,31,182,30,54,31,12,31,12,30,211,31,3,31,132,31,114,31,122,31,250,31,145,31,127,31,124,31,162,31,2,31,224,31,249,31,4,31,59,31,109,31,109,30,74,31,219,31,107,31,8,31,59,31,10,31,216,31,49,31,37,31,249,31,47,31,43,31,4,31,4,30,245,31,84,31,84,31,60,31,60,30,60,29,41,31,237,31,237,30,237,29,197,31,156,31,133,31,196,31,129,31,129,30,129,29,136,31,130,31,54,31,100,31,11,31,129,31,2,31,2,30,24,31,163,31,171,31,133,31,24,31,148,31,55,31,185,31,166,31,5,31,49,31,138,31,136,31,44,31,30,31,65,31,65,30,74,31,19,31,3,31,191,31,163,31,125,31,139,31,139,30,139,29,92,31,76,31,228,31,228,30,2,31,2,30,2,29,58,31,213,31,188,31,26,31,73,31,139,31,139,30,216,31,171,31,59,31,101,31,178,31,116,31,232,31,254,31,134,31,108,31,247,31,228,31,228,30,228,29,25,31,85,31,173,31,88,31,125,31,160,31,112,31,112,30,112,29,83,31,166,31,100,31,100,30,57,31,196,31,196,30,196,29,223,31,223,30,109,31,109,30,201,31,201,30,92,31,107,31,171,31,75,31,167,31,8,31,198,31,198,30,185,31,30,31,127,31,152,31,206,31,84,31,46,31,196,31,196,30,103,31,155,31,81,31,79,31,45,31,219,31,181,31,4,31,142,31,58,31,58,30,226,31,33,31,205,31,39,31,85,31,115,31,148,31,87,31,219,31,153,31,170,31,8,31,154,31,138,31,174,31,76,31,58,31,221,31,134,31,50,31,19,31,19,30,19,29,19,28,218,31,48,31,108,31,158,31,27,31,215,31,252,31,252,30,91,31,43,31,43,30,63,31,22,31,142,31,125,31,68,31,68,30,14,31,243,31,146,31,21,31,21,30,163,31,238,31,235,31,116,31,236,31,231,31,231,31,88,31,162,31,149,31,149,30,219,31,151,31,187,31,187,30,32,31,115,31,115,30,115,29,115,28,115,27,115,26,40,31,41,31,120,31,248,31,201,31,201,30,241,31,200,31,10,31,171,31,254,31,189,31,189,30,231,31,231,30,136,31,119,31,79,31,79,30,79,29,79,28,47,31,165,31,165,30,199,31,55,31,163,31,89,31,103,31,235,31,44,31,118,31,86,31,86,30,95,31,95,31,95,30,95,29,122,31,63,31,8,31,138,31,106,31,102,31,113,31,213,31,213,30,169,31,140,31,202,31,167,31,149,31,149,30,12,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
