-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 242;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,128,0,225,0,25,0,171,0,102,0,166,0,239,0,30,0,161,0,55,0,248,0,0,0,79,0,58,0,225,0,46,0,0,0,138,0,73,0,0,0,0,0,202,0,249,0,62,0,10,0,0,0,0,0,243,0,129,0,0,0,204,0,0,0,0,0,183,0,193,0,0,0,198,0,0,0,0,0,79,0,25,0,141,0,240,0,178,0,0,0,33,0,0,0,5,0,36,0,14,0,42,0,90,0,22,0,11,0,85,0,143,0,0,0,91,0,79,0,27,0,207,0,83,0,219,0,243,0,152,0,170,0,0,0,45,0,226,0,147,0,215,0,171,0,149,0,100,0,4,0,160,0,252,0,125,0,134,0,67,0,43,0,160,0,135,0,92,0,0,0,61,0,0,0,4,0,98,0,233,0,248,0,47,0,208,0,0,0,42,0,241,0,190,0,105,0,128,0,88,0,0,0,109,0,0,0,0,0,171,0,167,0,66,0,171,0,134,0,233,0,199,0,95,0,170,0,103,0,42,0,152,0,186,0,0,0,156,0,26,0,184,0,0,0,13,0,56,0,244,0,115,0,130,0,212,0,46,0,0,0,219,0,138,0,0,0,246,0,81,0,0,0,0,0,0,0,252,0,130,0,0,0,31,0,2,0,0,0,58,0,237,0,82,0,0,0,0,0,132,0,72,0,229,0,218,0,42,0,17,0,230,0,106,0,93,0,62,0,141,0,135,0,0,0,38,0,144,0,210,0,225,0,0,0,110,0,0,0,0,0,2,0,0,0,124,0,0,0,32,0,229,0,131,0,35,0,8,0,29,0,200,0,0,0,24,0,0,0,112,0,0,0,231,0,208,0,0,0,209,0,25,0,10,0,0,0,45,0,96,0,174,0,170,0,0,0,4,0,0,0,134,0,126,0,94,0,209,0,235,0,62,0,218,0,192,0,62,0,225,0,116,0,208,0,250,0,135,0,152,0,0,0,61,0,48,0,0,0,39,0,228,0,243,0,171,0,144,0,175,0,0,0,181,0,0,0,255,0,83,0,0,0,182,0,106,0,235,0,1,0,168,0,0,0,151,0,204,0,189,0,44,0);
signal scenario_full  : scenario_type := (93,31,128,31,225,31,25,31,171,31,102,31,166,31,239,31,30,31,161,31,55,31,248,31,248,30,79,31,58,31,225,31,46,31,46,30,138,31,73,31,73,30,73,29,202,31,249,31,62,31,10,31,10,30,10,29,243,31,129,31,129,30,204,31,204,30,204,29,183,31,193,31,193,30,198,31,198,30,198,29,79,31,25,31,141,31,240,31,178,31,178,30,33,31,33,30,5,31,36,31,14,31,42,31,90,31,22,31,11,31,85,31,143,31,143,30,91,31,79,31,27,31,207,31,83,31,219,31,243,31,152,31,170,31,170,30,45,31,226,31,147,31,215,31,171,31,149,31,100,31,4,31,160,31,252,31,125,31,134,31,67,31,43,31,160,31,135,31,92,31,92,30,61,31,61,30,4,31,98,31,233,31,248,31,47,31,208,31,208,30,42,31,241,31,190,31,105,31,128,31,88,31,88,30,109,31,109,30,109,29,171,31,167,31,66,31,171,31,134,31,233,31,199,31,95,31,170,31,103,31,42,31,152,31,186,31,186,30,156,31,26,31,184,31,184,30,13,31,56,31,244,31,115,31,130,31,212,31,46,31,46,30,219,31,138,31,138,30,246,31,81,31,81,30,81,29,81,28,252,31,130,31,130,30,31,31,2,31,2,30,58,31,237,31,82,31,82,30,82,29,132,31,72,31,229,31,218,31,42,31,17,31,230,31,106,31,93,31,62,31,141,31,135,31,135,30,38,31,144,31,210,31,225,31,225,30,110,31,110,30,110,29,2,31,2,30,124,31,124,30,32,31,229,31,131,31,35,31,8,31,29,31,200,31,200,30,24,31,24,30,112,31,112,30,231,31,208,31,208,30,209,31,25,31,10,31,10,30,45,31,96,31,174,31,170,31,170,30,4,31,4,30,134,31,126,31,94,31,209,31,235,31,62,31,218,31,192,31,62,31,225,31,116,31,208,31,250,31,135,31,152,31,152,30,61,31,48,31,48,30,39,31,228,31,243,31,171,31,144,31,175,31,175,30,181,31,181,30,255,31,83,31,83,30,182,31,106,31,235,31,1,31,168,31,168,30,151,31,204,31,189,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
