-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_786 is
end project_tb_786;

architecture project_tb_arch_786 of project_tb_786 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 851;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (246,0,155,0,103,0,249,0,121,0,51,0,192,0,193,0,221,0,236,0,0,0,107,0,184,0,3,0,0,0,174,0,98,0,175,0,111,0,248,0,32,0,230,0,71,0,227,0,14,0,188,0,234,0,0,0,220,0,255,0,96,0,100,0,238,0,198,0,232,0,172,0,0,0,57,0,10,0,45,0,0,0,97,0,8,0,229,0,252,0,104,0,61,0,0,0,39,0,248,0,158,0,200,0,229,0,252,0,76,0,48,0,11,0,40,0,128,0,0,0,200,0,21,0,91,0,17,0,0,0,79,0,0,0,203,0,0,0,1,0,0,0,246,0,131,0,167,0,0,0,127,0,0,0,14,0,236,0,0,0,0,0,192,0,34,0,54,0,166,0,76,0,206,0,117,0,20,0,31,0,214,0,0,0,57,0,85,0,0,0,86,0,10,0,43,0,119,0,28,0,248,0,0,0,61,0,33,0,0,0,28,0,219,0,24,0,40,0,64,0,206,0,87,0,24,0,0,0,0,0,144,0,197,0,0,0,165,0,130,0,155,0,204,0,155,0,237,0,0,0,0,0,153,0,0,0,13,0,138,0,245,0,214,0,53,0,156,0,145,0,116,0,0,0,0,0,250,0,102,0,177,0,66,0,84,0,42,0,0,0,0,0,0,0,31,0,157,0,118,0,0,0,178,0,0,0,34,0,225,0,39,0,2,0,189,0,199,0,95,0,254,0,0,0,0,0,24,0,147,0,0,0,0,0,222,0,250,0,0,0,224,0,27,0,206,0,181,0,12,0,221,0,91,0,57,0,68,0,106,0,0,0,0,0,242,0,79,0,61,0,246,0,0,0,160,0,199,0,27,0,97,0,191,0,173,0,5,0,233,0,25,0,167,0,0,0,200,0,163,0,68,0,217,0,0,0,197,0,241,0,0,0,0,0,204,0,0,0,158,0,201,0,0,0,219,0,0,0,8,0,243,0,0,0,0,0,185,0,214,0,196,0,147,0,222,0,0,0,142,0,143,0,110,0,226,0,145,0,173,0,189,0,165,0,62,0,175,0,221,0,102,0,115,0,170,0,47,0,55,0,193,0,165,0,120,0,0,0,62,0,47,0,99,0,0,0,114,0,131,0,0,0,63,0,108,0,56,0,3,0,3,0,222,0,32,0,239,0,167,0,106,0,73,0,163,0,118,0,199,0,0,0,44,0,248,0,0,0,186,0,14,0,224,0,118,0,38,0,131,0,128,0,0,0,78,0,0,0,190,0,48,0,89,0,219,0,12,0,0,0,0,0,238,0,159,0,0,0,117,0,252,0,154,0,0,0,0,0,0,0,143,0,170,0,214,0,0,0,154,0,172,0,53,0,146,0,0,0,238,0,56,0,11,0,74,0,0,0,169,0,216,0,87,0,154,0,83,0,144,0,166,0,183,0,242,0,0,0,150,0,250,0,141,0,231,0,212,0,147,0,115,0,102,0,215,0,48,0,166,0,20,0,0,0,0,0,151,0,0,0,249,0,0,0,93,0,177,0,187,0,0,0,67,0,82,0,197,0,83,0,11,0,139,0,232,0,234,0,164,0,0,0,216,0,55,0,0,0,83,0,0,0,34,0,195,0,57,0,187,0,236,0,203,0,72,0,252,0,237,0,25,0,140,0,182,0,254,0,0,0,126,0,58,0,6,0,32,0,58,0,233,0,166,0,178,0,18,0,0,0,0,0,185,0,187,0,209,0,90,0,160,0,250,0,72,0,132,0,199,0,0,0,0,0,161,0,207,0,0,0,21,0,0,0,0,0,60,0,214,0,190,0,0,0,13,0,160,0,72,0,248,0,0,0,0,0,206,0,35,0,196,0,69,0,104,0,119,0,153,0,208,0,110,0,97,0,13,0,144,0,227,0,194,0,233,0,150,0,192,0,38,0,252,0,0,0,20,0,220,0,112,0,240,0,0,0,227,0,1,0,114,0,120,0,229,0,54,0,0,0,215,0,0,0,39,0,221,0,45,0,7,0,77,0,41,0,77,0,220,0,192,0,218,0,90,0,209,0,111,0,51,0,64,0,68,0,0,0,216,0,16,0,0,0,28,0,161,0,118,0,251,0,151,0,240,0,19,0,85,0,26,0,41,0,212,0,0,0,40,0,254,0,249,0,98,0,165,0,157,0,46,0,234,0,87,0,181,0,152,0,238,0,66,0,135,0,176,0,0,0,63,0,205,0,122,0,0,0,92,0,0,0,176,0,194,0,0,0,159,0,67,0,30,0,0,0,179,0,91,0,0,0,104,0,0,0,113,0,212,0,0,0,103,0,205,0,0,0,0,0,244,0,0,0,87,0,19,0,80,0,1,0,13,0,80,0,70,0,0,0,189,0,134,0,0,0,227,0,0,0,31,0,29,0,241,0,77,0,200,0,55,0,128,0,31,0,196,0,251,0,194,0,223,0,200,0,255,0,186,0,45,0,123,0,95,0,54,0,18,0,0,0,88,0,248,0,0,0,0,0,189,0,38,0,0,0,147,0,110,0,182,0,255,0,163,0,240,0,240,0,157,0,0,0,226,0,0,0,60,0,154,0,77,0,99,0,218,0,135,0,90,0,170,0,0,0,0,0,0,0,92,0,0,0,163,0,67,0,0,0,45,0,0,0,82,0,0,0,97,0,0,0,97,0,169,0,36,0,0,0,61,0,0,0,179,0,0,0,251,0,46,0,0,0,125,0,147,0,139,0,228,0,103,0,116,0,0,0,115,0,242,0,175,0,142,0,46,0,94,0,0,0,227,0,78,0,99,0,140,0,16,0,222,0,76,0,175,0,0,0,38,0,14,0,171,0,124,0,64,0,0,0,114,0,25,0,11,0,139,0,207,0,0,0,37,0,11,0,174,0,7,0,164,0,240,0,79,0,0,0,252,0,201,0,0,0,128,0,44,0,183,0,248,0,71,0,192,0,126,0,181,0,227,0,0,0,247,0,197,0,0,0,73,0,0,0,255,0,233,0,250,0,233,0,19,0,0,0,176,0,206,0,150,0,122,0,0,0,0,0,2,0,0,0,178,0,206,0,0,0,93,0,207,0,212,0,211,0,207,0,0,0,138,0,39,0,178,0,92,0,0,0,212,0,0,0,21,0,66,0,255,0,72,0,121,0,158,0,126,0,142,0,0,0,163,0,67,0,139,0,122,0,171,0,0,0,0,0,179,0,74,0,0,0,130,0,18,0,0,0,53,0,0,0,0,0,137,0,30,0,164,0,130,0,0,0,124,0,0,0,135,0,117,0,119,0,110,0,111,0,192,0,60,0,51,0,38,0,45,0,95,0,54,0,172,0,95,0,152,0,163,0,0,0,208,0,0,0,216,0,225,0,0,0,215,0,92,0,190,0,0,0,45,0,0,0,0,0,71,0,197,0,24,0,0,0,218,0,185,0,100,0,64,0,0,0,147,0,20,0,202,0,17,0,186,0,242,0,153,0,250,0,0,0,80,0,17,0,106,0,0,0,19,0,9,0,0,0,0,0,0,0,215,0,152,0,236,0,163,0,79,0,234,0,211,0,247,0,0,0,135,0,114,0,235,0,77,0,0,0,11,0,236,0,0,0,182,0,162,0,1,0,122,0,81,0,135,0,218,0,77,0,231,0,101,0,189,0,132,0,177,0,252,0,251,0,0,0,38,0,7,0,122,0,14,0,6,0,71,0,78,0,230,0,49,0,81,0,0,0,215,0,240,0,0,0,65,0,150,0,0,0,121,0,152,0,0,0,17,0,244,0,73,0,0,0,71,0,154,0,47,0,197,0,43,0,142,0,9,0,217,0,14,0,29,0,254,0,58,0,94,0);
signal scenario_full  : scenario_type := (246,31,155,31,103,31,249,31,121,31,51,31,192,31,193,31,221,31,236,31,236,30,107,31,184,31,3,31,3,30,174,31,98,31,175,31,111,31,248,31,32,31,230,31,71,31,227,31,14,31,188,31,234,31,234,30,220,31,255,31,96,31,100,31,238,31,198,31,232,31,172,31,172,30,57,31,10,31,45,31,45,30,97,31,8,31,229,31,252,31,104,31,61,31,61,30,39,31,248,31,158,31,200,31,229,31,252,31,76,31,48,31,11,31,40,31,128,31,128,30,200,31,21,31,91,31,17,31,17,30,79,31,79,30,203,31,203,30,1,31,1,30,246,31,131,31,167,31,167,30,127,31,127,30,14,31,236,31,236,30,236,29,192,31,34,31,54,31,166,31,76,31,206,31,117,31,20,31,31,31,214,31,214,30,57,31,85,31,85,30,86,31,10,31,43,31,119,31,28,31,248,31,248,30,61,31,33,31,33,30,28,31,219,31,24,31,40,31,64,31,206,31,87,31,24,31,24,30,24,29,144,31,197,31,197,30,165,31,130,31,155,31,204,31,155,31,237,31,237,30,237,29,153,31,153,30,13,31,138,31,245,31,214,31,53,31,156,31,145,31,116,31,116,30,116,29,250,31,102,31,177,31,66,31,84,31,42,31,42,30,42,29,42,28,31,31,157,31,118,31,118,30,178,31,178,30,34,31,225,31,39,31,2,31,189,31,199,31,95,31,254,31,254,30,254,29,24,31,147,31,147,30,147,29,222,31,250,31,250,30,224,31,27,31,206,31,181,31,12,31,221,31,91,31,57,31,68,31,106,31,106,30,106,29,242,31,79,31,61,31,246,31,246,30,160,31,199,31,27,31,97,31,191,31,173,31,5,31,233,31,25,31,167,31,167,30,200,31,163,31,68,31,217,31,217,30,197,31,241,31,241,30,241,29,204,31,204,30,158,31,201,31,201,30,219,31,219,30,8,31,243,31,243,30,243,29,185,31,214,31,196,31,147,31,222,31,222,30,142,31,143,31,110,31,226,31,145,31,173,31,189,31,165,31,62,31,175,31,221,31,102,31,115,31,170,31,47,31,55,31,193,31,165,31,120,31,120,30,62,31,47,31,99,31,99,30,114,31,131,31,131,30,63,31,108,31,56,31,3,31,3,31,222,31,32,31,239,31,167,31,106,31,73,31,163,31,118,31,199,31,199,30,44,31,248,31,248,30,186,31,14,31,224,31,118,31,38,31,131,31,128,31,128,30,78,31,78,30,190,31,48,31,89,31,219,31,12,31,12,30,12,29,238,31,159,31,159,30,117,31,252,31,154,31,154,30,154,29,154,28,143,31,170,31,214,31,214,30,154,31,172,31,53,31,146,31,146,30,238,31,56,31,11,31,74,31,74,30,169,31,216,31,87,31,154,31,83,31,144,31,166,31,183,31,242,31,242,30,150,31,250,31,141,31,231,31,212,31,147,31,115,31,102,31,215,31,48,31,166,31,20,31,20,30,20,29,151,31,151,30,249,31,249,30,93,31,177,31,187,31,187,30,67,31,82,31,197,31,83,31,11,31,139,31,232,31,234,31,164,31,164,30,216,31,55,31,55,30,83,31,83,30,34,31,195,31,57,31,187,31,236,31,203,31,72,31,252,31,237,31,25,31,140,31,182,31,254,31,254,30,126,31,58,31,6,31,32,31,58,31,233,31,166,31,178,31,18,31,18,30,18,29,185,31,187,31,209,31,90,31,160,31,250,31,72,31,132,31,199,31,199,30,199,29,161,31,207,31,207,30,21,31,21,30,21,29,60,31,214,31,190,31,190,30,13,31,160,31,72,31,248,31,248,30,248,29,206,31,35,31,196,31,69,31,104,31,119,31,153,31,208,31,110,31,97,31,13,31,144,31,227,31,194,31,233,31,150,31,192,31,38,31,252,31,252,30,20,31,220,31,112,31,240,31,240,30,227,31,1,31,114,31,120,31,229,31,54,31,54,30,215,31,215,30,39,31,221,31,45,31,7,31,77,31,41,31,77,31,220,31,192,31,218,31,90,31,209,31,111,31,51,31,64,31,68,31,68,30,216,31,16,31,16,30,28,31,161,31,118,31,251,31,151,31,240,31,19,31,85,31,26,31,41,31,212,31,212,30,40,31,254,31,249,31,98,31,165,31,157,31,46,31,234,31,87,31,181,31,152,31,238,31,66,31,135,31,176,31,176,30,63,31,205,31,122,31,122,30,92,31,92,30,176,31,194,31,194,30,159,31,67,31,30,31,30,30,179,31,91,31,91,30,104,31,104,30,113,31,212,31,212,30,103,31,205,31,205,30,205,29,244,31,244,30,87,31,19,31,80,31,1,31,13,31,80,31,70,31,70,30,189,31,134,31,134,30,227,31,227,30,31,31,29,31,241,31,77,31,200,31,55,31,128,31,31,31,196,31,251,31,194,31,223,31,200,31,255,31,186,31,45,31,123,31,95,31,54,31,18,31,18,30,88,31,248,31,248,30,248,29,189,31,38,31,38,30,147,31,110,31,182,31,255,31,163,31,240,31,240,31,157,31,157,30,226,31,226,30,60,31,154,31,77,31,99,31,218,31,135,31,90,31,170,31,170,30,170,29,170,28,92,31,92,30,163,31,67,31,67,30,45,31,45,30,82,31,82,30,97,31,97,30,97,31,169,31,36,31,36,30,61,31,61,30,179,31,179,30,251,31,46,31,46,30,125,31,147,31,139,31,228,31,103,31,116,31,116,30,115,31,242,31,175,31,142,31,46,31,94,31,94,30,227,31,78,31,99,31,140,31,16,31,222,31,76,31,175,31,175,30,38,31,14,31,171,31,124,31,64,31,64,30,114,31,25,31,11,31,139,31,207,31,207,30,37,31,11,31,174,31,7,31,164,31,240,31,79,31,79,30,252,31,201,31,201,30,128,31,44,31,183,31,248,31,71,31,192,31,126,31,181,31,227,31,227,30,247,31,197,31,197,30,73,31,73,30,255,31,233,31,250,31,233,31,19,31,19,30,176,31,206,31,150,31,122,31,122,30,122,29,2,31,2,30,178,31,206,31,206,30,93,31,207,31,212,31,211,31,207,31,207,30,138,31,39,31,178,31,92,31,92,30,212,31,212,30,21,31,66,31,255,31,72,31,121,31,158,31,126,31,142,31,142,30,163,31,67,31,139,31,122,31,171,31,171,30,171,29,179,31,74,31,74,30,130,31,18,31,18,30,53,31,53,30,53,29,137,31,30,31,164,31,130,31,130,30,124,31,124,30,135,31,117,31,119,31,110,31,111,31,192,31,60,31,51,31,38,31,45,31,95,31,54,31,172,31,95,31,152,31,163,31,163,30,208,31,208,30,216,31,225,31,225,30,215,31,92,31,190,31,190,30,45,31,45,30,45,29,71,31,197,31,24,31,24,30,218,31,185,31,100,31,64,31,64,30,147,31,20,31,202,31,17,31,186,31,242,31,153,31,250,31,250,30,80,31,17,31,106,31,106,30,19,31,9,31,9,30,9,29,9,28,215,31,152,31,236,31,163,31,79,31,234,31,211,31,247,31,247,30,135,31,114,31,235,31,77,31,77,30,11,31,236,31,236,30,182,31,162,31,1,31,122,31,81,31,135,31,218,31,77,31,231,31,101,31,189,31,132,31,177,31,252,31,251,31,251,30,38,31,7,31,122,31,14,31,6,31,71,31,78,31,230,31,49,31,81,31,81,30,215,31,240,31,240,30,65,31,150,31,150,30,121,31,152,31,152,30,17,31,244,31,73,31,73,30,71,31,154,31,47,31,197,31,43,31,142,31,9,31,217,31,14,31,29,31,254,31,58,31,94,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
