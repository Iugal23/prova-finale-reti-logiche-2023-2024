-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 350;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (67,0,240,0,145,0,0,0,78,0,169,0,221,0,196,0,0,0,96,0,0,0,56,0,132,0,214,0,55,0,245,0,170,0,93,0,0,0,0,0,0,0,33,0,0,0,149,0,225,0,89,0,108,0,123,0,162,0,150,0,209,0,0,0,87,0,50,0,124,0,0,0,244,0,4,0,246,0,103,0,0,0,0,0,70,0,0,0,105,0,0,0,241,0,0,0,248,0,113,0,129,0,0,0,207,0,127,0,168,0,15,0,0,0,0,0,182,0,0,0,101,0,0,0,110,0,97,0,110,0,157,0,93,0,209,0,228,0,147,0,82,0,250,0,176,0,0,0,220,0,126,0,88,0,0,0,0,0,46,0,144,0,163,0,88,0,0,0,24,0,0,0,0,0,83,0,210,0,182,0,230,0,0,0,84,0,86,0,212,0,59,0,79,0,89,0,204,0,98,0,0,0,248,0,183,0,75,0,10,0,0,0,98,0,38,0,9,0,0,0,27,0,19,0,75,0,161,0,0,0,223,0,25,0,250,0,0,0,218,0,0,0,31,0,0,0,138,0,201,0,179,0,212,0,95,0,189,0,49,0,8,0,0,0,90,0,0,0,187,0,84,0,0,0,0,0,144,0,0,0,69,0,0,0,117,0,155,0,242,0,179,0,206,0,245,0,0,0,214,0,0,0,152,0,73,0,179,0,21,0,203,0,228,0,179,0,162,0,0,0,45,0,173,0,89,0,40,0,90,0,152,0,144,0,97,0,0,0,164,0,22,0,191,0,0,0,99,0,94,0,0,0,0,0,98,0,253,0,0,0,12,0,0,0,192,0,24,0,87,0,195,0,46,0,247,0,252,0,0,0,237,0,53,0,196,0,160,0,128,0,0,0,0,0,173,0,62,0,146,0,83,0,73,0,35,0,69,0,55,0,0,0,248,0,0,0,0,0,180,0,243,0,190,0,0,0,63,0,34,0,47,0,2,0,16,0,127,0,102,0,75,0,178,0,2,0,235,0,103,0,0,0,98,0,0,0,192,0,226,0,252,0,250,0,84,0,239,0,146,0,0,0,25,0,163,0,8,0,81,0,205,0,157,0,0,0,225,0,0,0,0,0,200,0,235,0,34,0,0,0,104,0,232,0,138,0,202,0,190,0,78,0,142,0,48,0,55,0,85,0,205,0,160,0,35,0,0,0,66,0,0,0,60,0,148,0,19,0,111,0,68,0,0,0,76,0,146,0,41,0,244,0,2,0,36,0,0,0,64,0,51,0,14,0,222,0,39,0,151,0,246,0,102,0,196,0,44,0,0,0,15,0,255,0,25,0,90,0,176,0,139,0,31,0,208,0,56,0,164,0,25,0,155,0,0,0,0,0,181,0,153,0,0,0,27,0,210,0,0,0,180,0,116,0,37,0,39,0,102,0,35,0,0,0,126,0,101,0,25,0,48,0,0,0,68,0,31,0,47,0,83,0,0,0,198,0,0,0,38,0,156,0,2,0,92,0,224,0,70,0,228,0,34,0,109,0,170,0,212,0,29,0,207,0,81,0,0,0,94,0,30,0,20,0,0,0,251,0,100,0);
signal scenario_full  : scenario_type := (67,31,240,31,145,31,145,30,78,31,169,31,221,31,196,31,196,30,96,31,96,30,56,31,132,31,214,31,55,31,245,31,170,31,93,31,93,30,93,29,93,28,33,31,33,30,149,31,225,31,89,31,108,31,123,31,162,31,150,31,209,31,209,30,87,31,50,31,124,31,124,30,244,31,4,31,246,31,103,31,103,30,103,29,70,31,70,30,105,31,105,30,241,31,241,30,248,31,113,31,129,31,129,30,207,31,127,31,168,31,15,31,15,30,15,29,182,31,182,30,101,31,101,30,110,31,97,31,110,31,157,31,93,31,209,31,228,31,147,31,82,31,250,31,176,31,176,30,220,31,126,31,88,31,88,30,88,29,46,31,144,31,163,31,88,31,88,30,24,31,24,30,24,29,83,31,210,31,182,31,230,31,230,30,84,31,86,31,212,31,59,31,79,31,89,31,204,31,98,31,98,30,248,31,183,31,75,31,10,31,10,30,98,31,38,31,9,31,9,30,27,31,19,31,75,31,161,31,161,30,223,31,25,31,250,31,250,30,218,31,218,30,31,31,31,30,138,31,201,31,179,31,212,31,95,31,189,31,49,31,8,31,8,30,90,31,90,30,187,31,84,31,84,30,84,29,144,31,144,30,69,31,69,30,117,31,155,31,242,31,179,31,206,31,245,31,245,30,214,31,214,30,152,31,73,31,179,31,21,31,203,31,228,31,179,31,162,31,162,30,45,31,173,31,89,31,40,31,90,31,152,31,144,31,97,31,97,30,164,31,22,31,191,31,191,30,99,31,94,31,94,30,94,29,98,31,253,31,253,30,12,31,12,30,192,31,24,31,87,31,195,31,46,31,247,31,252,31,252,30,237,31,53,31,196,31,160,31,128,31,128,30,128,29,173,31,62,31,146,31,83,31,73,31,35,31,69,31,55,31,55,30,248,31,248,30,248,29,180,31,243,31,190,31,190,30,63,31,34,31,47,31,2,31,16,31,127,31,102,31,75,31,178,31,2,31,235,31,103,31,103,30,98,31,98,30,192,31,226,31,252,31,250,31,84,31,239,31,146,31,146,30,25,31,163,31,8,31,81,31,205,31,157,31,157,30,225,31,225,30,225,29,200,31,235,31,34,31,34,30,104,31,232,31,138,31,202,31,190,31,78,31,142,31,48,31,55,31,85,31,205,31,160,31,35,31,35,30,66,31,66,30,60,31,148,31,19,31,111,31,68,31,68,30,76,31,146,31,41,31,244,31,2,31,36,31,36,30,64,31,51,31,14,31,222,31,39,31,151,31,246,31,102,31,196,31,44,31,44,30,15,31,255,31,25,31,90,31,176,31,139,31,31,31,208,31,56,31,164,31,25,31,155,31,155,30,155,29,181,31,153,31,153,30,27,31,210,31,210,30,180,31,116,31,37,31,39,31,102,31,35,31,35,30,126,31,101,31,25,31,48,31,48,30,68,31,31,31,47,31,83,31,83,30,198,31,198,30,38,31,156,31,2,31,92,31,224,31,70,31,228,31,34,31,109,31,170,31,212,31,29,31,207,31,81,31,81,30,94,31,30,31,20,31,20,30,251,31,100,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
