-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 811;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (73,0,0,0,13,0,214,0,221,0,248,0,116,0,111,0,210,0,253,0,77,0,249,0,136,0,216,0,255,0,143,0,196,0,109,0,245,0,15,0,0,0,62,0,232,0,192,0,0,0,0,0,84,0,173,0,61,0,68,0,26,0,239,0,216,0,93,0,48,0,186,0,90,0,173,0,0,0,16,0,250,0,249,0,231,0,64,0,0,0,63,0,42,0,64,0,136,0,149,0,0,0,152,0,254,0,0,0,161,0,5,0,237,0,112,0,0,0,12,0,244,0,74,0,103,0,248,0,57,0,50,0,30,0,160,0,81,0,166,0,0,0,216,0,0,0,229,0,222,0,101,0,55,0,225,0,0,0,245,0,123,0,219,0,170,0,27,0,150,0,52,0,135,0,86,0,187,0,100,0,191,0,0,0,236,0,181,0,21,0,160,0,0,0,235,0,167,0,125,0,0,0,0,0,7,0,0,0,171,0,136,0,34,0,36,0,223,0,178,0,0,0,117,0,0,0,206,0,43,0,0,0,0,0,46,0,67,0,210,0,0,0,0,0,126,0,68,0,81,0,226,0,155,0,38,0,218,0,252,0,66,0,68,0,182,0,128,0,232,0,229,0,92,0,228,0,152,0,21,0,89,0,69,0,146,0,0,0,73,0,0,0,0,0,109,0,224,0,0,0,100,0,48,0,71,0,242,0,191,0,56,0,211,0,201,0,0,0,14,0,126,0,216,0,252,0,6,0,232,0,33,0,0,0,218,0,81,0,0,0,0,0,186,0,114,0,95,0,246,0,134,0,0,0,136,0,56,0,251,0,94,0,0,0,23,0,0,0,134,0,0,0,222,0,197,0,141,0,165,0,148,0,128,0,178,0,251,0,32,0,80,0,38,0,140,0,0,0,2,0,56,0,191,0,106,0,203,0,0,0,228,0,183,0,36,0,246,0,82,0,0,0,147,0,3,0,88,0,205,0,157,0,0,0,183,0,222,0,27,0,169,0,0,0,182,0,42,0,46,0,0,0,0,0,77,0,24,0,108,0,227,0,193,0,236,0,169,0,140,0,0,0,192,0,44,0,50,0,82,0,114,0,221,0,48,0,38,0,60,0,0,0,0,0,144,0,192,0,64,0,93,0,246,0,86,0,0,0,232,0,95,0,163,0,235,0,246,0,36,0,232,0,48,0,86,0,174,0,0,0,69,0,107,0,229,0,53,0,34,0,76,0,0,0,0,0,216,0,240,0,188,0,168,0,188,0,148,0,239,0,174,0,112,0,0,0,247,0,201,0,91,0,148,0,62,0,80,0,137,0,0,0,0,0,190,0,218,0,201,0,188,0,0,0,129,0,244,0,222,0,176,0,7,0,148,0,99,0,233,0,63,0,189,0,127,0,191,0,179,0,141,0,196,0,0,0,96,0,137,0,30,0,86,0,101,0,99,0,83,0,70,0,99,0,0,0,222,0,0,0,139,0,0,0,50,0,203,0,179,0,67,0,62,0,121,0,116,0,81,0,114,0,154,0,9,0,72,0,156,0,0,0,3,0,172,0,0,0,87,0,161,0,224,0,33,0,151,0,217,0,84,0,203,0,6,0,39,0,222,0,107,0,0,0,75,0,154,0,232,0,21,0,0,0,169,0,52,0,0,0,62,0,232,0,42,0,32,0,68,0,0,0,116,0,52,0,37,0,208,0,111,0,0,0,45,0,182,0,55,0,232,0,58,0,0,0,224,0,228,0,180,0,251,0,0,0,202,0,125,0,225,0,247,0,230,0,94,0,0,0,185,0,221,0,233,0,220,0,102,0,155,0,37,0,107,0,140,0,151,0,0,0,51,0,64,0,105,0,198,0,0,0,43,0,164,0,253,0,182,0,139,0,184,0,55,0,90,0,78,0,214,0,0,0,60,0,0,0,147,0,228,0,224,0,7,0,3,0,148,0,29,0,222,0,91,0,180,0,0,0,146,0,31,0,120,0,212,0,0,0,236,0,7,0,0,0,54,0,0,0,0,0,120,0,16,0,0,0,242,0,254,0,0,0,69,0,218,0,0,0,57,0,234,0,0,0,253,0,7,0,0,0,88,0,147,0,137,0,32,0,176,0,210,0,0,0,213,0,12,0,0,0,0,0,187,0,94,0,0,0,150,0,223,0,246,0,152,0,133,0,154,0,127,0,26,0,66,0,175,0,16,0,0,0,126,0,219,0,235,0,79,0,0,0,0,0,97,0,0,0,173,0,0,0,0,0,87,0,0,0,108,0,80,0,62,0,63,0,224,0,183,0,201,0,174,0,32,0,181,0,25,0,233,0,144,0,90,0,247,0,13,0,130,0,0,0,9,0,0,0,79,0,0,0,47,0,52,0,245,0,95,0,135,0,213,0,210,0,254,0,126,0,221,0,229,0,222,0,66,0,229,0,78,0,121,0,23,0,179,0,84,0,151,0,0,0,68,0,231,0,151,0,213,0,108,0,0,0,0,0,87,0,70,0,220,0,98,0,0,0,217,0,150,0,0,0,80,0,0,0,159,0,238,0,11,0,253,0,0,0,0,0,179,0,151,0,30,0,234,0,48,0,97,0,173,0,128,0,152,0,119,0,4,0,18,0,0,0,176,0,64,0,0,0,253,0,230,0,183,0,62,0,160,0,138,0,222,0,69,0,0,0,58,0,86,0,167,0,252,0,66,0,0,0,229,0,191,0,57,0,33,0,247,0,26,0,127,0,152,0,119,0,254,0,0,0,40,0,205,0,197,0,119,0,70,0,141,0,0,0,143,0,234,0,214,0,123,0,174,0,220,0,141,0,71,0,141,0,139,0,0,0,21,0,0,0,0,0,45,0,48,0,0,0,4,0,245,0,139,0,231,0,250,0,243,0,23,0,147,0,45,0,45,0,126,0,228,0,30,0,0,0,108,0,219,0,213,0,0,0,0,0,0,0,29,0,156,0,112,0,0,0,251,0,130,0,0,0,116,0,0,0,91,0,191,0,2,0,0,0,171,0,0,0,210,0,26,0,0,0,21,0,252,0,37,0,169,0,178,0,235,0,222,0,216,0,110,0,161,0,0,0,246,0,0,0,0,0,158,0,169,0,0,0,41,0,109,0,0,0,107,0,0,0,0,0,0,0,33,0,145,0,6,0,100,0,12,0,241,0,118,0,19,0,0,0,202,0,253,0,176,0,254,0,192,0,118,0,111,0,224,0,224,0,0,0,155,0,20,0,47,0,0,0,66,0,216,0,0,0,67,0,146,0,51,0,0,0,228,0,172,0,0,0,0,0,8,0,254,0,248,0,220,0,221,0,0,0,0,0,229,0,166,0,135,0,67,0,0,0,109,0,0,0,202,0,104,0,33,0,42,0,96,0,229,0,149,0,0,0,102,0,0,0,113,0,0,0,0,0,78,0,255,0,192,0,94,0,40,0,57,0,179,0,181,0,228,0,196,0,124,0,136,0,0,0,7,0,0,0,205,0,248,0,161,0,22,0,28,0,40,0,0,0,108,0,59,0,189,0,0,0,15,0,28,0,189,0,194,0,187,0,124,0,169,0,0,0,205,0,153,0,240,0,143,0,96,0,0,0,241,0,44,0,0,0,249,0,0,0,217,0,158,0,219,0,251,0,76,0,125,0,43,0,99,0,230,0,101,0,58,0);
signal scenario_full  : scenario_type := (73,31,73,30,13,31,214,31,221,31,248,31,116,31,111,31,210,31,253,31,77,31,249,31,136,31,216,31,255,31,143,31,196,31,109,31,245,31,15,31,15,30,62,31,232,31,192,31,192,30,192,29,84,31,173,31,61,31,68,31,26,31,239,31,216,31,93,31,48,31,186,31,90,31,173,31,173,30,16,31,250,31,249,31,231,31,64,31,64,30,63,31,42,31,64,31,136,31,149,31,149,30,152,31,254,31,254,30,161,31,5,31,237,31,112,31,112,30,12,31,244,31,74,31,103,31,248,31,57,31,50,31,30,31,160,31,81,31,166,31,166,30,216,31,216,30,229,31,222,31,101,31,55,31,225,31,225,30,245,31,123,31,219,31,170,31,27,31,150,31,52,31,135,31,86,31,187,31,100,31,191,31,191,30,236,31,181,31,21,31,160,31,160,30,235,31,167,31,125,31,125,30,125,29,7,31,7,30,171,31,136,31,34,31,36,31,223,31,178,31,178,30,117,31,117,30,206,31,43,31,43,30,43,29,46,31,67,31,210,31,210,30,210,29,126,31,68,31,81,31,226,31,155,31,38,31,218,31,252,31,66,31,68,31,182,31,128,31,232,31,229,31,92,31,228,31,152,31,21,31,89,31,69,31,146,31,146,30,73,31,73,30,73,29,109,31,224,31,224,30,100,31,48,31,71,31,242,31,191,31,56,31,211,31,201,31,201,30,14,31,126,31,216,31,252,31,6,31,232,31,33,31,33,30,218,31,81,31,81,30,81,29,186,31,114,31,95,31,246,31,134,31,134,30,136,31,56,31,251,31,94,31,94,30,23,31,23,30,134,31,134,30,222,31,197,31,141,31,165,31,148,31,128,31,178,31,251,31,32,31,80,31,38,31,140,31,140,30,2,31,56,31,191,31,106,31,203,31,203,30,228,31,183,31,36,31,246,31,82,31,82,30,147,31,3,31,88,31,205,31,157,31,157,30,183,31,222,31,27,31,169,31,169,30,182,31,42,31,46,31,46,30,46,29,77,31,24,31,108,31,227,31,193,31,236,31,169,31,140,31,140,30,192,31,44,31,50,31,82,31,114,31,221,31,48,31,38,31,60,31,60,30,60,29,144,31,192,31,64,31,93,31,246,31,86,31,86,30,232,31,95,31,163,31,235,31,246,31,36,31,232,31,48,31,86,31,174,31,174,30,69,31,107,31,229,31,53,31,34,31,76,31,76,30,76,29,216,31,240,31,188,31,168,31,188,31,148,31,239,31,174,31,112,31,112,30,247,31,201,31,91,31,148,31,62,31,80,31,137,31,137,30,137,29,190,31,218,31,201,31,188,31,188,30,129,31,244,31,222,31,176,31,7,31,148,31,99,31,233,31,63,31,189,31,127,31,191,31,179,31,141,31,196,31,196,30,96,31,137,31,30,31,86,31,101,31,99,31,83,31,70,31,99,31,99,30,222,31,222,30,139,31,139,30,50,31,203,31,179,31,67,31,62,31,121,31,116,31,81,31,114,31,154,31,9,31,72,31,156,31,156,30,3,31,172,31,172,30,87,31,161,31,224,31,33,31,151,31,217,31,84,31,203,31,6,31,39,31,222,31,107,31,107,30,75,31,154,31,232,31,21,31,21,30,169,31,52,31,52,30,62,31,232,31,42,31,32,31,68,31,68,30,116,31,52,31,37,31,208,31,111,31,111,30,45,31,182,31,55,31,232,31,58,31,58,30,224,31,228,31,180,31,251,31,251,30,202,31,125,31,225,31,247,31,230,31,94,31,94,30,185,31,221,31,233,31,220,31,102,31,155,31,37,31,107,31,140,31,151,31,151,30,51,31,64,31,105,31,198,31,198,30,43,31,164,31,253,31,182,31,139,31,184,31,55,31,90,31,78,31,214,31,214,30,60,31,60,30,147,31,228,31,224,31,7,31,3,31,148,31,29,31,222,31,91,31,180,31,180,30,146,31,31,31,120,31,212,31,212,30,236,31,7,31,7,30,54,31,54,30,54,29,120,31,16,31,16,30,242,31,254,31,254,30,69,31,218,31,218,30,57,31,234,31,234,30,253,31,7,31,7,30,88,31,147,31,137,31,32,31,176,31,210,31,210,30,213,31,12,31,12,30,12,29,187,31,94,31,94,30,150,31,223,31,246,31,152,31,133,31,154,31,127,31,26,31,66,31,175,31,16,31,16,30,126,31,219,31,235,31,79,31,79,30,79,29,97,31,97,30,173,31,173,30,173,29,87,31,87,30,108,31,80,31,62,31,63,31,224,31,183,31,201,31,174,31,32,31,181,31,25,31,233,31,144,31,90,31,247,31,13,31,130,31,130,30,9,31,9,30,79,31,79,30,47,31,52,31,245,31,95,31,135,31,213,31,210,31,254,31,126,31,221,31,229,31,222,31,66,31,229,31,78,31,121,31,23,31,179,31,84,31,151,31,151,30,68,31,231,31,151,31,213,31,108,31,108,30,108,29,87,31,70,31,220,31,98,31,98,30,217,31,150,31,150,30,80,31,80,30,159,31,238,31,11,31,253,31,253,30,253,29,179,31,151,31,30,31,234,31,48,31,97,31,173,31,128,31,152,31,119,31,4,31,18,31,18,30,176,31,64,31,64,30,253,31,230,31,183,31,62,31,160,31,138,31,222,31,69,31,69,30,58,31,86,31,167,31,252,31,66,31,66,30,229,31,191,31,57,31,33,31,247,31,26,31,127,31,152,31,119,31,254,31,254,30,40,31,205,31,197,31,119,31,70,31,141,31,141,30,143,31,234,31,214,31,123,31,174,31,220,31,141,31,71,31,141,31,139,31,139,30,21,31,21,30,21,29,45,31,48,31,48,30,4,31,245,31,139,31,231,31,250,31,243,31,23,31,147,31,45,31,45,31,126,31,228,31,30,31,30,30,108,31,219,31,213,31,213,30,213,29,213,28,29,31,156,31,112,31,112,30,251,31,130,31,130,30,116,31,116,30,91,31,191,31,2,31,2,30,171,31,171,30,210,31,26,31,26,30,21,31,252,31,37,31,169,31,178,31,235,31,222,31,216,31,110,31,161,31,161,30,246,31,246,30,246,29,158,31,169,31,169,30,41,31,109,31,109,30,107,31,107,30,107,29,107,28,33,31,145,31,6,31,100,31,12,31,241,31,118,31,19,31,19,30,202,31,253,31,176,31,254,31,192,31,118,31,111,31,224,31,224,31,224,30,155,31,20,31,47,31,47,30,66,31,216,31,216,30,67,31,146,31,51,31,51,30,228,31,172,31,172,30,172,29,8,31,254,31,248,31,220,31,221,31,221,30,221,29,229,31,166,31,135,31,67,31,67,30,109,31,109,30,202,31,104,31,33,31,42,31,96,31,229,31,149,31,149,30,102,31,102,30,113,31,113,30,113,29,78,31,255,31,192,31,94,31,40,31,57,31,179,31,181,31,228,31,196,31,124,31,136,31,136,30,7,31,7,30,205,31,248,31,161,31,22,31,28,31,40,31,40,30,108,31,59,31,189,31,189,30,15,31,28,31,189,31,194,31,187,31,124,31,169,31,169,30,205,31,153,31,240,31,143,31,96,31,96,30,241,31,44,31,44,30,249,31,249,30,217,31,158,31,219,31,251,31,76,31,125,31,43,31,99,31,230,31,101,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
