-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 918;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (240,0,251,0,0,0,0,0,11,0,197,0,38,0,70,0,56,0,209,0,71,0,13,0,104,0,162,0,78,0,253,0,124,0,107,0,150,0,129,0,146,0,187,0,248,0,0,0,218,0,94,0,0,0,74,0,188,0,0,0,101,0,154,0,89,0,128,0,0,0,195,0,212,0,174,0,34,0,83,0,15,0,62,0,170,0,0,0,255,0,0,0,25,0,209,0,240,0,53,0,108,0,179,0,121,0,0,0,0,0,241,0,0,0,24,0,238,0,179,0,143,0,244,0,119,0,193,0,245,0,120,0,10,0,79,0,0,0,148,0,0,0,0,0,152,0,89,0,43,0,117,0,50,0,128,0,126,0,174,0,105,0,132,0,0,0,14,0,100,0,0,0,0,0,204,0,0,0,0,0,42,0,183,0,178,0,0,0,191,0,163,0,127,0,76,0,181,0,0,0,17,0,232,0,0,0,129,0,174,0,207,0,125,0,27,0,5,0,210,0,2,0,85,0,221,0,0,0,221,0,225,0,126,0,255,0,0,0,0,0,178,0,0,0,132,0,110,0,230,0,11,0,0,0,0,0,31,0,147,0,44,0,83,0,192,0,61,0,9,0,0,0,17,0,11,0,174,0,178,0,0,0,0,0,156,0,148,0,69,0,0,0,14,0,174,0,178,0,151,0,190,0,109,0,141,0,0,0,76,0,155,0,68,0,166,0,179,0,117,0,113,0,203,0,59,0,147,0,0,0,0,0,30,0,5,0,34,0,90,0,0,0,76,0,59,0,136,0,44,0,60,0,48,0,73,0,82,0,0,0,147,0,201,0,0,0,48,0,107,0,67,0,18,0,112,0,247,0,65,0,97,0,0,0,180,0,246,0,158,0,0,0,92,0,227,0,227,0,203,0,238,0,189,0,0,0,154,0,159,0,121,0,188,0,25,0,122,0,0,0,65,0,0,0,204,0,0,0,0,0,16,0,110,0,13,0,230,0,12,0,29,0,159,0,137,0,30,0,151,0,126,0,56,0,96,0,113,0,0,0,76,0,182,0,0,0,38,0,199,0,108,0,0,0,0,0,0,0,59,0,221,0,222,0,45,0,103,0,192,0,167,0,227,0,226,0,139,0,137,0,0,0,254,0,0,0,182,0,165,0,135,0,147,0,0,0,237,0,69,0,194,0,0,0,0,0,0,0,0,0,156,0,209,0,238,0,10,0,79,0,202,0,180,0,4,0,122,0,227,0,43,0,0,0,0,0,179,0,118,0,204,0,60,0,101,0,92,0,27,0,166,0,121,0,116,0,57,0,108,0,89,0,211,0,137,0,231,0,0,0,0,0,152,0,218,0,133,0,144,0,0,0,167,0,24,0,186,0,218,0,16,0,236,0,17,0,74,0,204,0,222,0,0,0,199,0,106,0,116,0,0,0,0,0,85,0,146,0,217,0,21,0,209,0,148,0,0,0,55,0,0,0,110,0,169,0,0,0,13,0,0,0,0,0,77,0,0,0,207,0,9,0,0,0,113,0,185,0,110,0,0,0,15,0,32,0,144,0,32,0,111,0,39,0,71,0,0,0,126,0,68,0,80,0,0,0,98,0,157,0,0,0,137,0,0,0,227,0,208,0,55,0,128,0,0,0,49,0,70,0,33,0,0,0,194,0,128,0,0,0,0,0,228,0,55,0,222,0,0,0,98,0,62,0,150,0,0,0,35,0,222,0,171,0,225,0,0,0,0,0,195,0,101,0,0,0,247,0,252,0,184,0,22,0,176,0,0,0,0,0,35,0,131,0,0,0,126,0,68,0,205,0,0,0,250,0,58,0,107,0,110,0,221,0,127,0,0,0,54,0,149,0,198,0,0,0,18,0,0,0,0,0,92,0,0,0,8,0,199,0,17,0,224,0,66,0,54,0,114,0,0,0,47,0,41,0,44,0,40,0,40,0,137,0,141,0,87,0,180,0,0,0,56,0,0,0,167,0,2,0,0,0,6,0,232,0,51,0,108,0,229,0,0,0,126,0,19,0,0,0,112,0,0,0,75,0,225,0,203,0,132,0,192,0,115,0,0,0,147,0,0,0,233,0,154,0,0,0,139,0,151,0,246,0,242,0,0,0,80,0,244,0,0,0,104,0,169,0,121,0,242,0,69,0,57,0,138,0,169,0,128,0,208,0,247,0,96,0,56,0,240,0,96,0,147,0,94,0,3,0,151,0,0,0,27,0,103,0,0,0,87,0,30,0,0,0,0,0,106,0,170,0,90,0,63,0,0,0,169,0,0,0,178,0,0,0,9,0,0,0,65,0,129,0,13,0,225,0,255,0,0,0,208,0,0,0,59,0,10,0,0,0,32,0,240,0,138,0,60,0,173,0,20,0,190,0,0,0,0,0,172,0,16,0,129,0,180,0,193,0,167,0,221,0,41,0,77,0,128,0,0,0,232,0,0,0,0,0,142,0,7,0,0,0,167,0,76,0,0,0,83,0,63,0,149,0,224,0,55,0,163,0,118,0,94,0,139,0,216,0,172,0,210,0,72,0,0,0,53,0,49,0,160,0,30,0,23,0,189,0,135,0,0,0,114,0,129,0,159,0,233,0,0,0,163,0,178,0,0,0,218,0,87,0,0,0,0,0,0,0,45,0,0,0,88,0,129,0,0,0,0,0,0,0,143,0,82,0,246,0,203,0,70,0,0,0,138,0,180,0,78,0,0,0,228,0,197,0,155,0,9,0,207,0,72,0,0,0,108,0,121,0,168,0,218,0,0,0,0,0,0,0,197,0,238,0,242,0,216,0,242,0,150,0,0,0,71,0,86,0,106,0,179,0,16,0,99,0,194,0,219,0,63,0,155,0,89,0,216,0,0,0,117,0,20,0,69,0,107,0,209,0,37,0,177,0,38,0,70,0,141,0,246,0,89,0,144,0,240,0,132,0,213,0,0,0,0,0,37,0,138,0,236,0,140,0,89,0,224,0,0,0,192,0,191,0,36,0,125,0,39,0,0,0,0,0,222,0,0,0,96,0,226,0,8,0,165,0,0,0,0,0,200,0,163,0,27,0,0,0,159,0,6,0,0,0,200,0,246,0,202,0,5,0,250,0,227,0,210,0,14,0,129,0,124,0,142,0,61,0,214,0,236,0,104,0,215,0,0,0,53,0,190,0,67,0,5,0,245,0,39,0,0,0,151,0,241,0,139,0,23,0,180,0,0,0,3,0,115,0,23,0,57,0,208,0,39,0,254,0,85,0,36,0,162,0,0,0,0,0,176,0,0,0,10,0,18,0,170,0,18,0,0,0,157,0,11,0,95,0,0,0,0,0,11,0,20,0,23,0,0,0,0,0,63,0,0,0,126,0,189,0,94,0,162,0,125,0,121,0,216,0,166,0,193,0,0,0,178,0,34,0,166,0,87,0,197,0,0,0,160,0,3,0,0,0,151,0,228,0,195,0,76,0,244,0,49,0,135,0,10,0,0,0,78,0,0,0,22,0,201,0,118,0,254,0,214,0,0,0,131,0,126,0,109,0,227,0,247,0,214,0,0,0,0,0,179,0,114,0,74,0,243,0,156,0,0,0,0,0,108,0,0,0,0,0,0,0,0,0,95,0,119,0,161,0,162,0,115,0,192,0,118,0,189,0,226,0,47,0,0,0,0,0,147,0,91,0,147,0,35,0,151,0,0,0,119,0,98,0,141,0,227,0,3,0,100,0,0,0,33,0,11,0,199,0,244,0,239,0,42,0,100,0,110,0,77,0,49,0,0,0,35,0,69,0,0,0,0,0,215,0,35,0,48,0,99,0,208,0,0,0,183,0,0,0,182,0,136,0,232,0,60,0,224,0,13,0,0,0,0,0,139,0,102,0,169,0,130,0,128,0,21,0,97,0,49,0,58,0,0,0,167,0,178,0,152,0,0,0,156,0,0,0,153,0,47,0,61,0,168,0,202,0,132,0,140,0,43,0,0,0,179,0,0,0,247,0,159,0,1,0,147,0,36,0,224,0,0,0,111,0,0,0,210,0,104,0,0,0,81,0,113,0,183,0,0,0,85,0,120,0,144,0,244,0,221,0,107,0,69,0,244,0,198,0,97,0,123,0,182,0,0,0,212,0,213,0,205,0,16,0,77,0,21,0);
signal scenario_full  : scenario_type := (240,31,251,31,251,30,251,29,11,31,197,31,38,31,70,31,56,31,209,31,71,31,13,31,104,31,162,31,78,31,253,31,124,31,107,31,150,31,129,31,146,31,187,31,248,31,248,30,218,31,94,31,94,30,74,31,188,31,188,30,101,31,154,31,89,31,128,31,128,30,195,31,212,31,174,31,34,31,83,31,15,31,62,31,170,31,170,30,255,31,255,30,25,31,209,31,240,31,53,31,108,31,179,31,121,31,121,30,121,29,241,31,241,30,24,31,238,31,179,31,143,31,244,31,119,31,193,31,245,31,120,31,10,31,79,31,79,30,148,31,148,30,148,29,152,31,89,31,43,31,117,31,50,31,128,31,126,31,174,31,105,31,132,31,132,30,14,31,100,31,100,30,100,29,204,31,204,30,204,29,42,31,183,31,178,31,178,30,191,31,163,31,127,31,76,31,181,31,181,30,17,31,232,31,232,30,129,31,174,31,207,31,125,31,27,31,5,31,210,31,2,31,85,31,221,31,221,30,221,31,225,31,126,31,255,31,255,30,255,29,178,31,178,30,132,31,110,31,230,31,11,31,11,30,11,29,31,31,147,31,44,31,83,31,192,31,61,31,9,31,9,30,17,31,11,31,174,31,178,31,178,30,178,29,156,31,148,31,69,31,69,30,14,31,174,31,178,31,151,31,190,31,109,31,141,31,141,30,76,31,155,31,68,31,166,31,179,31,117,31,113,31,203,31,59,31,147,31,147,30,147,29,30,31,5,31,34,31,90,31,90,30,76,31,59,31,136,31,44,31,60,31,48,31,73,31,82,31,82,30,147,31,201,31,201,30,48,31,107,31,67,31,18,31,112,31,247,31,65,31,97,31,97,30,180,31,246,31,158,31,158,30,92,31,227,31,227,31,203,31,238,31,189,31,189,30,154,31,159,31,121,31,188,31,25,31,122,31,122,30,65,31,65,30,204,31,204,30,204,29,16,31,110,31,13,31,230,31,12,31,29,31,159,31,137,31,30,31,151,31,126,31,56,31,96,31,113,31,113,30,76,31,182,31,182,30,38,31,199,31,108,31,108,30,108,29,108,28,59,31,221,31,222,31,45,31,103,31,192,31,167,31,227,31,226,31,139,31,137,31,137,30,254,31,254,30,182,31,165,31,135,31,147,31,147,30,237,31,69,31,194,31,194,30,194,29,194,28,194,27,156,31,209,31,238,31,10,31,79,31,202,31,180,31,4,31,122,31,227,31,43,31,43,30,43,29,179,31,118,31,204,31,60,31,101,31,92,31,27,31,166,31,121,31,116,31,57,31,108,31,89,31,211,31,137,31,231,31,231,30,231,29,152,31,218,31,133,31,144,31,144,30,167,31,24,31,186,31,218,31,16,31,236,31,17,31,74,31,204,31,222,31,222,30,199,31,106,31,116,31,116,30,116,29,85,31,146,31,217,31,21,31,209,31,148,31,148,30,55,31,55,30,110,31,169,31,169,30,13,31,13,30,13,29,77,31,77,30,207,31,9,31,9,30,113,31,185,31,110,31,110,30,15,31,32,31,144,31,32,31,111,31,39,31,71,31,71,30,126,31,68,31,80,31,80,30,98,31,157,31,157,30,137,31,137,30,227,31,208,31,55,31,128,31,128,30,49,31,70,31,33,31,33,30,194,31,128,31,128,30,128,29,228,31,55,31,222,31,222,30,98,31,62,31,150,31,150,30,35,31,222,31,171,31,225,31,225,30,225,29,195,31,101,31,101,30,247,31,252,31,184,31,22,31,176,31,176,30,176,29,35,31,131,31,131,30,126,31,68,31,205,31,205,30,250,31,58,31,107,31,110,31,221,31,127,31,127,30,54,31,149,31,198,31,198,30,18,31,18,30,18,29,92,31,92,30,8,31,199,31,17,31,224,31,66,31,54,31,114,31,114,30,47,31,41,31,44,31,40,31,40,31,137,31,141,31,87,31,180,31,180,30,56,31,56,30,167,31,2,31,2,30,6,31,232,31,51,31,108,31,229,31,229,30,126,31,19,31,19,30,112,31,112,30,75,31,225,31,203,31,132,31,192,31,115,31,115,30,147,31,147,30,233,31,154,31,154,30,139,31,151,31,246,31,242,31,242,30,80,31,244,31,244,30,104,31,169,31,121,31,242,31,69,31,57,31,138,31,169,31,128,31,208,31,247,31,96,31,56,31,240,31,96,31,147,31,94,31,3,31,151,31,151,30,27,31,103,31,103,30,87,31,30,31,30,30,30,29,106,31,170,31,90,31,63,31,63,30,169,31,169,30,178,31,178,30,9,31,9,30,65,31,129,31,13,31,225,31,255,31,255,30,208,31,208,30,59,31,10,31,10,30,32,31,240,31,138,31,60,31,173,31,20,31,190,31,190,30,190,29,172,31,16,31,129,31,180,31,193,31,167,31,221,31,41,31,77,31,128,31,128,30,232,31,232,30,232,29,142,31,7,31,7,30,167,31,76,31,76,30,83,31,63,31,149,31,224,31,55,31,163,31,118,31,94,31,139,31,216,31,172,31,210,31,72,31,72,30,53,31,49,31,160,31,30,31,23,31,189,31,135,31,135,30,114,31,129,31,159,31,233,31,233,30,163,31,178,31,178,30,218,31,87,31,87,30,87,29,87,28,45,31,45,30,88,31,129,31,129,30,129,29,129,28,143,31,82,31,246,31,203,31,70,31,70,30,138,31,180,31,78,31,78,30,228,31,197,31,155,31,9,31,207,31,72,31,72,30,108,31,121,31,168,31,218,31,218,30,218,29,218,28,197,31,238,31,242,31,216,31,242,31,150,31,150,30,71,31,86,31,106,31,179,31,16,31,99,31,194,31,219,31,63,31,155,31,89,31,216,31,216,30,117,31,20,31,69,31,107,31,209,31,37,31,177,31,38,31,70,31,141,31,246,31,89,31,144,31,240,31,132,31,213,31,213,30,213,29,37,31,138,31,236,31,140,31,89,31,224,31,224,30,192,31,191,31,36,31,125,31,39,31,39,30,39,29,222,31,222,30,96,31,226,31,8,31,165,31,165,30,165,29,200,31,163,31,27,31,27,30,159,31,6,31,6,30,200,31,246,31,202,31,5,31,250,31,227,31,210,31,14,31,129,31,124,31,142,31,61,31,214,31,236,31,104,31,215,31,215,30,53,31,190,31,67,31,5,31,245,31,39,31,39,30,151,31,241,31,139,31,23,31,180,31,180,30,3,31,115,31,23,31,57,31,208,31,39,31,254,31,85,31,36,31,162,31,162,30,162,29,176,31,176,30,10,31,18,31,170,31,18,31,18,30,157,31,11,31,95,31,95,30,95,29,11,31,20,31,23,31,23,30,23,29,63,31,63,30,126,31,189,31,94,31,162,31,125,31,121,31,216,31,166,31,193,31,193,30,178,31,34,31,166,31,87,31,197,31,197,30,160,31,3,31,3,30,151,31,228,31,195,31,76,31,244,31,49,31,135,31,10,31,10,30,78,31,78,30,22,31,201,31,118,31,254,31,214,31,214,30,131,31,126,31,109,31,227,31,247,31,214,31,214,30,214,29,179,31,114,31,74,31,243,31,156,31,156,30,156,29,108,31,108,30,108,29,108,28,108,27,95,31,119,31,161,31,162,31,115,31,192,31,118,31,189,31,226,31,47,31,47,30,47,29,147,31,91,31,147,31,35,31,151,31,151,30,119,31,98,31,141,31,227,31,3,31,100,31,100,30,33,31,11,31,199,31,244,31,239,31,42,31,100,31,110,31,77,31,49,31,49,30,35,31,69,31,69,30,69,29,215,31,35,31,48,31,99,31,208,31,208,30,183,31,183,30,182,31,136,31,232,31,60,31,224,31,13,31,13,30,13,29,139,31,102,31,169,31,130,31,128,31,21,31,97,31,49,31,58,31,58,30,167,31,178,31,152,31,152,30,156,31,156,30,153,31,47,31,61,31,168,31,202,31,132,31,140,31,43,31,43,30,179,31,179,30,247,31,159,31,1,31,147,31,36,31,224,31,224,30,111,31,111,30,210,31,104,31,104,30,81,31,113,31,183,31,183,30,85,31,120,31,144,31,244,31,221,31,107,31,69,31,244,31,198,31,97,31,123,31,182,31,182,30,212,31,213,31,205,31,16,31,77,31,21,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
