-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_360 is
end project_tb_360;

architecture project_tb_arch_360 of project_tb_360 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 849;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,178,0,246,0,0,0,25,0,207,0,156,0,56,0,175,0,209,0,87,0,161,0,254,0,54,0,213,0,0,0,0,0,121,0,0,0,0,0,0,0,242,0,188,0,19,0,210,0,142,0,0,0,0,0,211,0,62,0,148,0,64,0,0,0,238,0,0,0,246,0,137,0,0,0,243,0,152,0,130,0,94,0,0,0,0,0,0,0,111,0,199,0,37,0,138,0,249,0,177,0,64,0,170,0,131,0,36,0,57,0,0,0,250,0,121,0,65,0,0,0,152,0,236,0,126,0,0,0,98,0,0,0,0,0,17,0,20,0,0,0,93,0,0,0,78,0,0,0,172,0,0,0,43,0,171,0,238,0,194,0,58,0,148,0,0,0,0,0,0,0,4,0,246,0,0,0,206,0,0,0,23,0,167,0,0,0,121,0,152,0,182,0,36,0,86,0,212,0,0,0,91,0,81,0,185,0,0,0,109,0,58,0,102,0,131,0,0,0,184,0,0,0,160,0,77,0,120,0,47,0,51,0,0,0,0,0,161,0,116,0,165,0,0,0,0,0,236,0,0,0,15,0,213,0,73,0,216,0,212,0,126,0,75,0,57,0,199,0,72,0,0,0,14,0,45,0,33,0,83,0,58,0,182,0,32,0,0,0,0,0,37,0,157,0,17,0,74,0,17,0,48,0,83,0,126,0,0,0,238,0,145,0,2,0,0,0,167,0,192,0,23,0,17,0,232,0,248,0,41,0,129,0,34,0,91,0,63,0,49,0,37,0,29,0,162,0,116,0,77,0,200,0,140,0,136,0,168,0,228,0,24,0,0,0,24,0,0,0,0,0,0,0,48,0,234,0,243,0,192,0,0,0,0,0,154,0,0,0,175,0,234,0,123,0,58,0,0,0,0,0,116,0,0,0,139,0,170,0,47,0,135,0,16,0,107,0,0,0,0,0,97,0,155,0,111,0,38,0,254,0,0,0,149,0,189,0,0,0,218,0,155,0,47,0,0,0,0,0,0,0,25,0,154,0,6,0,146,0,164,0,78,0,91,0,85,0,165,0,0,0,162,0,19,0,31,0,0,0,178,0,1,0,132,0,93,0,141,0,55,0,35,0,35,0,83,0,161,0,69,0,245,0,167,0,244,0,241,0,0,0,0,0,210,0,101,0,74,0,118,0,198,0,0,0,137,0,246,0,13,0,0,0,11,0,155,0,117,0,147,0,136,0,0,0,51,0,0,0,0,0,37,0,138,0,43,0,0,0,55,0,0,0,0,0,0,0,24,0,147,0,174,0,141,0,77,0,241,0,7,0,126,0,202,0,168,0,108,0,216,0,191,0,0,0,41,0,1,0,235,0,127,0,0,0,0,0,0,0,90,0,150,0,61,0,0,0,122,0,212,0,103,0,0,0,34,0,45,0,8,0,148,0,163,0,251,0,148,0,115,0,145,0,0,0,238,0,41,0,0,0,184,0,0,0,83,0,116,0,102,0,0,0,14,0,200,0,191,0,212,0,200,0,31,0,76,0,0,0,187,0,254,0,163,0,0,0,76,0,198,0,0,0,241,0,72,0,0,0,0,0,31,0,184,0,0,0,0,0,235,0,138,0,0,0,0,0,0,0,99,0,192,0,84,0,74,0,92,0,246,0,108,0,122,0,39,0,255,0,230,0,136,0,4,0,226,0,224,0,28,0,0,0,239,0,152,0,11,0,146,0,133,0,113,0,74,0,182,0,5,0,139,0,189,0,0,0,117,0,0,0,157,0,140,0,152,0,37,0,122,0,89,0,0,0,156,0,110,0,149,0,233,0,18,0,112,0,232,0,150,0,0,0,190,0,121,0,69,0,0,0,19,0,100,0,0,0,124,0,8,0,218,0,82,0,2,0,18,0,122,0,146,0,82,0,68,0,175,0,77,0,194,0,46,0,0,0,158,0,180,0,137,0,184,0,150,0,105,0,0,0,0,0,5,0,143,0,90,0,187,0,0,0,35,0,182,0,114,0,222,0,68,0,103,0,56,0,104,0,233,0,102,0,0,0,147,0,174,0,43,0,0,0,131,0,85,0,0,0,0,0,102,0,175,0,237,0,189,0,123,0,167,0,231,0,228,0,20,0,87,0,128,0,192,0,0,0,203,0,179,0,248,0,123,0,195,0,0,0,0,0,0,0,0,0,131,0,57,0,102,0,152,0,118,0,49,0,62,0,167,0,21,0,250,0,12,0,147,0,97,0,146,0,139,0,0,0,0,0,0,0,0,0,86,0,12,0,172,0,0,0,121,0,208,0,0,0,130,0,56,0,135,0,242,0,147,0,188,0,70,0,16,0,22,0,129,0,224,0,245,0,133,0,22,0,0,0,33,0,221,0,238,0,94,0,177,0,167,0,61,0,73,0,0,0,23,0,21,0,154,0,0,0,59,0,159,0,183,0,168,0,242,0,14,0,235,0,66,0,148,0,58,0,3,0,138,0,0,0,0,0,95,0,0,0,0,0,169,0,0,0,46,0,62,0,112,0,11,0,0,0,73,0,212,0,129,0,76,0,255,0,190,0,207,0,50,0,32,0,152,0,66,0,242,0,46,0,174,0,0,0,223,0,0,0,101,0,122,0,43,0,119,0,31,0,33,0,158,0,195,0,65,0,172,0,0,0,80,0,126,0,0,0,247,0,27,0,19,0,81,0,221,0,230,0,156,0,249,0,124,0,91,0,207,0,0,0,247,0,0,0,44,0,8,0,29,0,46,0,131,0,244,0,127,0,19,0,204,0,0,0,227,0,11,0,145,0,212,0,151,0,16,0,0,0,53,0,108,0,120,0,43,0,1,0,66,0,5,0,0,0,117,0,68,0,0,0,98,0,210,0,0,0,70,0,95,0,91,0,85,0,239,0,0,0,221,0,0,0,0,0,81,0,112,0,121,0,103,0,92,0,80,0,83,0,36,0,114,0,0,0,0,0,144,0,84,0,101,0,0,0,54,0,69,0,167,0,0,0,0,0,43,0,175,0,189,0,166,0,0,0,0,0,115,0,144,0,0,0,212,0,84,0,248,0,28,0,0,0,61,0,255,0,99,0,18,0,2,0,21,0,166,0,0,0,30,0,115,0,7,0,0,0,161,0,0,0,20,0,90,0,0,0,54,0,29,0,52,0,157,0,0,0,0,0,132,0,156,0,122,0,180,0,91,0,55,0,51,0,244,0,168,0,72,0,15,0,62,0,121,0,31,0,108,0,164,0,63,0,184,0,209,0,0,0,56,0,0,0,177,0,218,0,0,0,0,0,0,0,171,0,108,0,230,0,0,0,0,0,141,0,40,0,38,0,0,0,35,0,134,0,75,0,41,0,163,0,151,0,121,0,0,0,0,0,115,0,0,0,0,0,240,0,221,0,178,0,110,0,117,0,106,0,173,0,188,0,47,0,62,0,0,0,152,0,109,0,253,0,0,0,232,0,0,0,194,0,72,0,0,0,115,0,0,0,0,0,0,0,158,0,0,0,183,0,177,0,201,0,164,0,75,0,232,0,221,0,0,0,85,0,238,0,0,0,126,0,80,0,186,0,135,0,197,0,92,0,32,0,61,0,162,0,109,0,39,0,0,0,163,0,0,0,63,0,35,0,130,0,61,0,0,0,116,0,0,0,0,0,157,0,133,0,0,0,228,0,148,0,162,0,0,0,130,0,210,0,42,0,146,0,27,0,122,0,0,0,184,0,89,0,146,0,171,0,227,0,251,0,175,0,81,0,8,0,204,0,109,0,15,0,0,0,102,0,146,0,0,0,128,0,20,0,107,0,89,0,90,0,107,0,0,0,4,0,210,0);
signal scenario_full  : scenario_type := (1,31,178,31,246,31,246,30,25,31,207,31,156,31,56,31,175,31,209,31,87,31,161,31,254,31,54,31,213,31,213,30,213,29,121,31,121,30,121,29,121,28,242,31,188,31,19,31,210,31,142,31,142,30,142,29,211,31,62,31,148,31,64,31,64,30,238,31,238,30,246,31,137,31,137,30,243,31,152,31,130,31,94,31,94,30,94,29,94,28,111,31,199,31,37,31,138,31,249,31,177,31,64,31,170,31,131,31,36,31,57,31,57,30,250,31,121,31,65,31,65,30,152,31,236,31,126,31,126,30,98,31,98,30,98,29,17,31,20,31,20,30,93,31,93,30,78,31,78,30,172,31,172,30,43,31,171,31,238,31,194,31,58,31,148,31,148,30,148,29,148,28,4,31,246,31,246,30,206,31,206,30,23,31,167,31,167,30,121,31,152,31,182,31,36,31,86,31,212,31,212,30,91,31,81,31,185,31,185,30,109,31,58,31,102,31,131,31,131,30,184,31,184,30,160,31,77,31,120,31,47,31,51,31,51,30,51,29,161,31,116,31,165,31,165,30,165,29,236,31,236,30,15,31,213,31,73,31,216,31,212,31,126,31,75,31,57,31,199,31,72,31,72,30,14,31,45,31,33,31,83,31,58,31,182,31,32,31,32,30,32,29,37,31,157,31,17,31,74,31,17,31,48,31,83,31,126,31,126,30,238,31,145,31,2,31,2,30,167,31,192,31,23,31,17,31,232,31,248,31,41,31,129,31,34,31,91,31,63,31,49,31,37,31,29,31,162,31,116,31,77,31,200,31,140,31,136,31,168,31,228,31,24,31,24,30,24,31,24,30,24,29,24,28,48,31,234,31,243,31,192,31,192,30,192,29,154,31,154,30,175,31,234,31,123,31,58,31,58,30,58,29,116,31,116,30,139,31,170,31,47,31,135,31,16,31,107,31,107,30,107,29,97,31,155,31,111,31,38,31,254,31,254,30,149,31,189,31,189,30,218,31,155,31,47,31,47,30,47,29,47,28,25,31,154,31,6,31,146,31,164,31,78,31,91,31,85,31,165,31,165,30,162,31,19,31,31,31,31,30,178,31,1,31,132,31,93,31,141,31,55,31,35,31,35,31,83,31,161,31,69,31,245,31,167,31,244,31,241,31,241,30,241,29,210,31,101,31,74,31,118,31,198,31,198,30,137,31,246,31,13,31,13,30,11,31,155,31,117,31,147,31,136,31,136,30,51,31,51,30,51,29,37,31,138,31,43,31,43,30,55,31,55,30,55,29,55,28,24,31,147,31,174,31,141,31,77,31,241,31,7,31,126,31,202,31,168,31,108,31,216,31,191,31,191,30,41,31,1,31,235,31,127,31,127,30,127,29,127,28,90,31,150,31,61,31,61,30,122,31,212,31,103,31,103,30,34,31,45,31,8,31,148,31,163,31,251,31,148,31,115,31,145,31,145,30,238,31,41,31,41,30,184,31,184,30,83,31,116,31,102,31,102,30,14,31,200,31,191,31,212,31,200,31,31,31,76,31,76,30,187,31,254,31,163,31,163,30,76,31,198,31,198,30,241,31,72,31,72,30,72,29,31,31,184,31,184,30,184,29,235,31,138,31,138,30,138,29,138,28,99,31,192,31,84,31,74,31,92,31,246,31,108,31,122,31,39,31,255,31,230,31,136,31,4,31,226,31,224,31,28,31,28,30,239,31,152,31,11,31,146,31,133,31,113,31,74,31,182,31,5,31,139,31,189,31,189,30,117,31,117,30,157,31,140,31,152,31,37,31,122,31,89,31,89,30,156,31,110,31,149,31,233,31,18,31,112,31,232,31,150,31,150,30,190,31,121,31,69,31,69,30,19,31,100,31,100,30,124,31,8,31,218,31,82,31,2,31,18,31,122,31,146,31,82,31,68,31,175,31,77,31,194,31,46,31,46,30,158,31,180,31,137,31,184,31,150,31,105,31,105,30,105,29,5,31,143,31,90,31,187,31,187,30,35,31,182,31,114,31,222,31,68,31,103,31,56,31,104,31,233,31,102,31,102,30,147,31,174,31,43,31,43,30,131,31,85,31,85,30,85,29,102,31,175,31,237,31,189,31,123,31,167,31,231,31,228,31,20,31,87,31,128,31,192,31,192,30,203,31,179,31,248,31,123,31,195,31,195,30,195,29,195,28,195,27,131,31,57,31,102,31,152,31,118,31,49,31,62,31,167,31,21,31,250,31,12,31,147,31,97,31,146,31,139,31,139,30,139,29,139,28,139,27,86,31,12,31,172,31,172,30,121,31,208,31,208,30,130,31,56,31,135,31,242,31,147,31,188,31,70,31,16,31,22,31,129,31,224,31,245,31,133,31,22,31,22,30,33,31,221,31,238,31,94,31,177,31,167,31,61,31,73,31,73,30,23,31,21,31,154,31,154,30,59,31,159,31,183,31,168,31,242,31,14,31,235,31,66,31,148,31,58,31,3,31,138,31,138,30,138,29,95,31,95,30,95,29,169,31,169,30,46,31,62,31,112,31,11,31,11,30,73,31,212,31,129,31,76,31,255,31,190,31,207,31,50,31,32,31,152,31,66,31,242,31,46,31,174,31,174,30,223,31,223,30,101,31,122,31,43,31,119,31,31,31,33,31,158,31,195,31,65,31,172,31,172,30,80,31,126,31,126,30,247,31,27,31,19,31,81,31,221,31,230,31,156,31,249,31,124,31,91,31,207,31,207,30,247,31,247,30,44,31,8,31,29,31,46,31,131,31,244,31,127,31,19,31,204,31,204,30,227,31,11,31,145,31,212,31,151,31,16,31,16,30,53,31,108,31,120,31,43,31,1,31,66,31,5,31,5,30,117,31,68,31,68,30,98,31,210,31,210,30,70,31,95,31,91,31,85,31,239,31,239,30,221,31,221,30,221,29,81,31,112,31,121,31,103,31,92,31,80,31,83,31,36,31,114,31,114,30,114,29,144,31,84,31,101,31,101,30,54,31,69,31,167,31,167,30,167,29,43,31,175,31,189,31,166,31,166,30,166,29,115,31,144,31,144,30,212,31,84,31,248,31,28,31,28,30,61,31,255,31,99,31,18,31,2,31,21,31,166,31,166,30,30,31,115,31,7,31,7,30,161,31,161,30,20,31,90,31,90,30,54,31,29,31,52,31,157,31,157,30,157,29,132,31,156,31,122,31,180,31,91,31,55,31,51,31,244,31,168,31,72,31,15,31,62,31,121,31,31,31,108,31,164,31,63,31,184,31,209,31,209,30,56,31,56,30,177,31,218,31,218,30,218,29,218,28,171,31,108,31,230,31,230,30,230,29,141,31,40,31,38,31,38,30,35,31,134,31,75,31,41,31,163,31,151,31,121,31,121,30,121,29,115,31,115,30,115,29,240,31,221,31,178,31,110,31,117,31,106,31,173,31,188,31,47,31,62,31,62,30,152,31,109,31,253,31,253,30,232,31,232,30,194,31,72,31,72,30,115,31,115,30,115,29,115,28,158,31,158,30,183,31,177,31,201,31,164,31,75,31,232,31,221,31,221,30,85,31,238,31,238,30,126,31,80,31,186,31,135,31,197,31,92,31,32,31,61,31,162,31,109,31,39,31,39,30,163,31,163,30,63,31,35,31,130,31,61,31,61,30,116,31,116,30,116,29,157,31,133,31,133,30,228,31,148,31,162,31,162,30,130,31,210,31,42,31,146,31,27,31,122,31,122,30,184,31,89,31,146,31,171,31,227,31,251,31,175,31,81,31,8,31,204,31,109,31,15,31,15,30,102,31,146,31,146,30,128,31,20,31,107,31,89,31,90,31,107,31,107,30,4,31,210,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
