-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_797 is
end project_tb_797;

architecture project_tb_arch_797 of project_tb_797 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 445;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (67,0,0,0,51,0,62,0,6,0,0,0,0,0,175,0,37,0,183,0,0,0,217,0,0,0,10,0,186,0,57,0,0,0,128,0,159,0,206,0,196,0,253,0,201,0,157,0,108,0,179,0,123,0,254,0,80,0,24,0,50,0,85,0,19,0,223,0,169,0,84,0,100,0,22,0,250,0,175,0,19,0,83,0,205,0,228,0,191,0,221,0,191,0,173,0,41,0,78,0,76,0,0,0,159,0,142,0,15,0,111,0,228,0,0,0,124,0,39,0,74,0,138,0,18,0,53,0,47,0,11,0,244,0,40,0,254,0,165,0,32,0,171,0,154,0,152,0,0,0,156,0,34,0,126,0,241,0,74,0,153,0,54,0,206,0,81,0,197,0,46,0,16,0,181,0,0,0,241,0,206,0,68,0,218,0,0,0,15,0,0,0,25,0,197,0,23,0,208,0,138,0,130,0,0,0,196,0,58,0,215,0,49,0,21,0,239,0,0,0,218,0,187,0,1,0,139,0,147,0,243,0,123,0,76,0,7,0,0,0,174,0,182,0,81,0,240,0,246,0,39,0,5,0,117,0,216,0,126,0,0,0,0,0,46,0,0,0,116,0,200,0,191,0,153,0,51,0,218,0,92,0,210,0,16,0,0,0,195,0,147,0,144,0,119,0,0,0,0,0,96,0,0,0,76,0,222,0,212,0,0,0,96,0,205,0,172,0,0,0,7,0,237,0,109,0,217,0,46,0,143,0,173,0,56,0,9,0,241,0,90,0,64,0,116,0,0,0,130,0,112,0,0,0,0,0,222,0,150,0,0,0,0,0,76,0,182,0,208,0,61,0,19,0,186,0,246,0,191,0,213,0,119,0,0,0,0,0,0,0,0,0,213,0,220,0,44,0,97,0,237,0,120,0,0,0,10,0,55,0,202,0,0,0,0,0,171,0,212,0,85,0,85,0,0,0,161,0,231,0,0,0,234,0,211,0,189,0,85,0,15,0,164,0,136,0,214,0,0,0,3,0,151,0,143,0,0,0,23,0,0,0,29,0,253,0,180,0,146,0,0,0,67,0,132,0,190,0,0,0,5,0,196,0,13,0,193,0,119,0,98,0,243,0,124,0,241,0,79,0,25,0,201,0,101,0,239,0,175,0,70,0,129,0,127,0,78,0,0,0,0,0,174,0,0,0,30,0,0,0,23,0,116,0,0,0,0,0,245,0,110,0,231,0,254,0,197,0,0,0,0,0,0,0,187,0,84,0,214,0,87,0,63,0,184,0,67,0,0,0,37,0,135,0,146,0,33,0,79,0,94,0,0,0,0,0,174,0,0,0,0,0,99,0,0,0,186,0,127,0,138,0,31,0,122,0,252,0,197,0,124,0,208,0,173,0,16,0,0,0,103,0,152,0,242,0,94,0,241,0,147,0,0,0,100,0,50,0,226,0,189,0,0,0,169,0,0,0,27,0,0,0,206,0,212,0,157,0,200,0,39,0,49,0,15,0,0,0,2,0,221,0,122,0,0,0,0,0,0,0,82,0,246,0,38,0,200,0,87,0,0,0,0,0,0,0,247,0,93,0,100,0,91,0,135,0,0,0,214,0,205,0,32,0,178,0,97,0,0,0,0,0,0,0,192,0,239,0,90,0,171,0,214,0,89,0,143,0,143,0,114,0,202,0,133,0,167,0,47,0,148,0,0,0,100,0,157,0,229,0,0,0,207,0,84,0,3,0,130,0,0,0,0,0,0,0,166,0,12,0,143,0,226,0,150,0,30,0,164,0,174,0,152,0,255,0,230,0,111,0,172,0,0,0,254,0,0,0,51,0,162,0,138,0,250,0,0,0,23,0,116,0,239,0,123,0,249,0,109,0,229,0,53,0,126,0,51,0,203,0,59,0,0,0,193,0,182,0,38,0,109,0,75,0,81,0,39,0,149,0,196,0,223,0,48,0,0,0,23,0,242,0,87,0,201,0,60,0,202,0,206,0,135,0,114,0,209,0,0,0);
signal scenario_full  : scenario_type := (67,31,67,30,51,31,62,31,6,31,6,30,6,29,175,31,37,31,183,31,183,30,217,31,217,30,10,31,186,31,57,31,57,30,128,31,159,31,206,31,196,31,253,31,201,31,157,31,108,31,179,31,123,31,254,31,80,31,24,31,50,31,85,31,19,31,223,31,169,31,84,31,100,31,22,31,250,31,175,31,19,31,83,31,205,31,228,31,191,31,221,31,191,31,173,31,41,31,78,31,76,31,76,30,159,31,142,31,15,31,111,31,228,31,228,30,124,31,39,31,74,31,138,31,18,31,53,31,47,31,11,31,244,31,40,31,254,31,165,31,32,31,171,31,154,31,152,31,152,30,156,31,34,31,126,31,241,31,74,31,153,31,54,31,206,31,81,31,197,31,46,31,16,31,181,31,181,30,241,31,206,31,68,31,218,31,218,30,15,31,15,30,25,31,197,31,23,31,208,31,138,31,130,31,130,30,196,31,58,31,215,31,49,31,21,31,239,31,239,30,218,31,187,31,1,31,139,31,147,31,243,31,123,31,76,31,7,31,7,30,174,31,182,31,81,31,240,31,246,31,39,31,5,31,117,31,216,31,126,31,126,30,126,29,46,31,46,30,116,31,200,31,191,31,153,31,51,31,218,31,92,31,210,31,16,31,16,30,195,31,147,31,144,31,119,31,119,30,119,29,96,31,96,30,76,31,222,31,212,31,212,30,96,31,205,31,172,31,172,30,7,31,237,31,109,31,217,31,46,31,143,31,173,31,56,31,9,31,241,31,90,31,64,31,116,31,116,30,130,31,112,31,112,30,112,29,222,31,150,31,150,30,150,29,76,31,182,31,208,31,61,31,19,31,186,31,246,31,191,31,213,31,119,31,119,30,119,29,119,28,119,27,213,31,220,31,44,31,97,31,237,31,120,31,120,30,10,31,55,31,202,31,202,30,202,29,171,31,212,31,85,31,85,31,85,30,161,31,231,31,231,30,234,31,211,31,189,31,85,31,15,31,164,31,136,31,214,31,214,30,3,31,151,31,143,31,143,30,23,31,23,30,29,31,253,31,180,31,146,31,146,30,67,31,132,31,190,31,190,30,5,31,196,31,13,31,193,31,119,31,98,31,243,31,124,31,241,31,79,31,25,31,201,31,101,31,239,31,175,31,70,31,129,31,127,31,78,31,78,30,78,29,174,31,174,30,30,31,30,30,23,31,116,31,116,30,116,29,245,31,110,31,231,31,254,31,197,31,197,30,197,29,197,28,187,31,84,31,214,31,87,31,63,31,184,31,67,31,67,30,37,31,135,31,146,31,33,31,79,31,94,31,94,30,94,29,174,31,174,30,174,29,99,31,99,30,186,31,127,31,138,31,31,31,122,31,252,31,197,31,124,31,208,31,173,31,16,31,16,30,103,31,152,31,242,31,94,31,241,31,147,31,147,30,100,31,50,31,226,31,189,31,189,30,169,31,169,30,27,31,27,30,206,31,212,31,157,31,200,31,39,31,49,31,15,31,15,30,2,31,221,31,122,31,122,30,122,29,122,28,82,31,246,31,38,31,200,31,87,31,87,30,87,29,87,28,247,31,93,31,100,31,91,31,135,31,135,30,214,31,205,31,32,31,178,31,97,31,97,30,97,29,97,28,192,31,239,31,90,31,171,31,214,31,89,31,143,31,143,31,114,31,202,31,133,31,167,31,47,31,148,31,148,30,100,31,157,31,229,31,229,30,207,31,84,31,3,31,130,31,130,30,130,29,130,28,166,31,12,31,143,31,226,31,150,31,30,31,164,31,174,31,152,31,255,31,230,31,111,31,172,31,172,30,254,31,254,30,51,31,162,31,138,31,250,31,250,30,23,31,116,31,239,31,123,31,249,31,109,31,229,31,53,31,126,31,51,31,203,31,59,31,59,30,193,31,182,31,38,31,109,31,75,31,81,31,39,31,149,31,196,31,223,31,48,31,48,30,23,31,242,31,87,31,201,31,60,31,202,31,206,31,135,31,114,31,209,31,209,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
