-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_470 is
end project_tb_470;

architecture project_tb_arch_470 of project_tb_470 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 953;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (26,0,234,0,0,0,139,0,14,0,84,0,203,0,0,0,0,0,66,0,254,0,104,0,0,0,196,0,25,0,173,0,101,0,217,0,124,0,3,0,0,0,75,0,112,0,218,0,125,0,229,0,141,0,60,0,0,0,136,0,164,0,233,0,16,0,92,0,227,0,16,0,93,0,151,0,35,0,167,0,253,0,91,0,70,0,198,0,186,0,0,0,168,0,219,0,71,0,186,0,217,0,230,0,170,0,231,0,164,0,0,0,0,0,69,0,45,0,37,0,174,0,246,0,238,0,0,0,96,0,0,0,215,0,97,0,92,0,212,0,176,0,176,0,156,0,143,0,0,0,67,0,170,0,0,0,109,0,0,0,202,0,0,0,189,0,31,0,172,0,219,0,20,0,249,0,188,0,172,0,79,0,0,0,142,0,106,0,77,0,85,0,43,0,96,0,96,0,135,0,51,0,207,0,253,0,29,0,99,0,47,0,0,0,247,0,120,0,74,0,29,0,164,0,0,0,0,0,187,0,76,0,0,0,168,0,44,0,121,0,240,0,118,0,170,0,140,0,3,0,166,0,142,0,0,0,115,0,0,0,39,0,252,0,156,0,237,0,227,0,237,0,26,0,137,0,87,0,116,0,199,0,221,0,4,0,17,0,179,0,0,0,30,0,0,0,160,0,223,0,212,0,0,0,0,0,239,0,118,0,0,0,97,0,245,0,89,0,0,0,34,0,0,0,197,0,224,0,255,0,77,0,209,0,0,0,136,0,251,0,59,0,79,0,34,0,204,0,0,0,185,0,196,0,32,0,97,0,216,0,211,0,0,0,78,0,104,0,165,0,180,0,116,0,245,0,9,0,0,0,7,0,0,0,219,0,81,0,175,0,99,0,91,0,149,0,0,0,225,0,248,0,234,0,192,0,114,0,0,0,87,0,161,0,0,0,0,0,0,0,156,0,188,0,0,0,153,0,0,0,198,0,24,0,218,0,239,0,180,0,98,0,209,0,0,0,238,0,27,0,253,0,210,0,17,0,68,0,89,0,14,0,128,0,0,0,0,0,132,0,38,0,162,0,0,0,86,0,3,0,149,0,23,0,249,0,69,0,0,0,46,0,232,0,52,0,153,0,106,0,131,0,0,0,49,0,160,0,148,0,218,0,167,0,5,0,28,0,160,0,228,0,0,0,209,0,90,0,247,0,151,0,245,0,209,0,139,0,17,0,195,0,220,0,0,0,226,0,159,0,0,0,120,0,75,0,0,0,76,0,138,0,185,0,0,0,160,0,217,0,254,0,72,0,246,0,134,0,148,0,0,0,16,0,144,0,39,0,0,0,129,0,0,0,200,0,151,0,111,0,54,0,35,0,0,0,22,0,111,0,0,0,180,0,0,0,162,0,98,0,23,0,0,0,224,0,0,0,56,0,76,0,99,0,34,0,21,0,192,0,0,0,168,0,185,0,244,0,95,0,185,0,0,0,131,0,88,0,0,0,131,0,157,0,112,0,0,0,128,0,19,0,103,0,150,0,62,0,178,0,213,0,6,0,207,0,0,0,217,0,243,0,0,0,135,0,217,0,0,0,0,0,0,0,78,0,59,0,187,0,240,0,0,0,114,0,80,0,179,0,56,0,121,0,68,0,0,0,120,0,0,0,17,0,250,0,0,0,185,0,243,0,230,0,169,0,0,0,0,0,123,0,200,0,120,0,35,0,215,0,141,0,202,0,0,0,53,0,0,0,96,0,236,0,237,0,8,0,194,0,187,0,244,0,0,0,119,0,13,0,248,0,95,0,213,0,27,0,255,0,0,0,0,0,224,0,194,0,151,0,110,0,223,0,169,0,157,0,10,0,66,0,0,0,12,0,0,0,213,0,187,0,0,0,203,0,0,0,45,0,0,0,254,0,0,0,193,0,47,0,41,0,0,0,195,0,194,0,171,0,61,0,52,0,247,0,228,0,237,0,35,0,113,0,20,0,254,0,137,0,106,0,230,0,201,0,190,0,170,0,152,0,174,0,144,0,188,0,43,0,125,0,122,0,238,0,76,0,124,0,48,0,43,0,94,0,229,0,139,0,81,0,101,0,0,0,175,0,70,0,186,0,102,0,88,0,211,0,149,0,52,0,0,0,138,0,173,0,25,0,177,0,0,0,202,0,174,0,114,0,10,0,42,0,0,0,0,0,108,0,5,0,0,0,67,0,34,0,98,0,12,0,112,0,50,0,171,0,154,0,126,0,112,0,200,0,200,0,30,0,108,0,234,0,236,0,87,0,0,0,0,0,197,0,114,0,161,0,220,0,105,0,100,0,144,0,2,0,0,0,102,0,13,0,236,0,69,0,124,0,12,0,99,0,98,0,48,0,161,0,82,0,10,0,0,0,116,0,36,0,15,0,251,0,0,0,135,0,153,0,181,0,74,0,0,0,238,0,192,0,0,0,169,0,0,0,140,0,0,0,0,0,239,0,0,0,235,0,210,0,2,0,0,0,0,0,0,0,253,0,226,0,178,0,0,0,0,0,81,0,202,0,215,0,159,0,142,0,0,0,0,0,246,0,0,0,125,0,0,0,228,0,82,0,0,0,193,0,235,0,106,0,0,0,185,0,1,0,0,0,145,0,0,0,204,0,0,0,86,0,91,0,242,0,94,0,135,0,230,0,197,0,73,0,186,0,123,0,0,0,0,0,141,0,153,0,237,0,115,0,81,0,0,0,212,0,95,0,250,0,181,0,58,0,16,0,104,0,193,0,0,0,128,0,97,0,21,0,213,0,219,0,40,0,0,0,0,0,179,0,0,0,241,0,64,0,95,0,12,0,228,0,67,0,44,0,0,0,167,0,0,0,17,0,30,0,141,0,123,0,221,0,81,0,243,0,70,0,6,0,0,0,60,0,48,0,98,0,89,0,0,0,225,0,0,0,223,0,24,0,0,0,169,0,0,0,105,0,0,0,91,0,215,0,0,0,248,0,187,0,79,0,35,0,161,0,234,0,118,0,86,0,50,0,202,0,0,0,0,0,14,0,0,0,0,0,134,0,138,0,48,0,0,0,120,0,80,0,0,0,132,0,246,0,108,0,246,0,76,0,102,0,189,0,47,0,184,0,0,0,97,0,102,0,221,0,165,0,0,0,254,0,151,0,125,0,104,0,108,0,76,0,0,0,0,0,0,0,71,0,157,0,188,0,215,0,220,0,1,0,133,0,0,0,52,0,226,0,193,0,153,0,0,0,237,0,11,0,111,0,141,0,140,0,96,0,127,0,0,0,241,0,238,0,0,0,139,0,0,0,112,0,187,0,242,0,35,0,108,0,138,0,54,0,89,0,58,0,175,0,227,0,47,0,100,0,72,0,44,0,214,0,53,0,224,0,24,0,227,0,60,0,250,0,13,0,170,0,0,0,205,0,204,0,66,0,138,0,172,0,0,0,218,0,3,0,83,0,72,0,53,0,43,0,12,0,205,0,29,0,66,0,205,0,116,0,0,0,0,0,0,0,0,0,0,0,61,0,247,0,12,0,0,0,22,0,0,0,0,0,0,0,113,0,192,0,141,0,5,0,213,0,0,0,48,0,32,0,225,0,0,0,129,0,116,0,136,0,41,0,81,0,0,0,237,0,169,0,53,0,134,0,147,0,83,0,240,0,196,0,61,0,0,0,10,0,66,0,48,0,0,0,25,0,182,0,223,0,0,0,98,0,40,0,178,0,37,0,0,0,255,0,21,0,113,0,61,0,171,0,44,0,218,0,0,0,217,0,214,0,192,0,230,0,237,0,16,0,0,0,147,0,227,0,0,0,0,0,111,0,8,0,75,0,35,0,0,0,0,0,208,0,122,0,143,0,40,0,245,0,0,0,182,0,77,0,177,0,154,0,0,0,107,0,73,0,0,0,27,0,110,0,0,0,150,0,0,0,0,0,216,0,224,0,0,0,65,0,108,0,136,0,211,0,219,0,190,0,197,0,15,0,138,0,87,0,222,0,234,0,0,0,0,0,19,0,4,0,244,0,194,0,0,0,183,0,114,0,0,0,0,0,145,0,121,0,43,0,34,0,108,0,155,0,0,0,123,0,144,0,0,0,81,0,169,0,33,0,68,0,156,0,177,0,228,0,0,0,0,0,0,0,230,0,0,0,230,0,130,0,203,0,222,0,201,0,245,0,140,0,106,0,0,0,242,0,95,0,0,0,253,0,0,0,119,0,199,0,71,0,178,0,21,0,39,0,9,0,236,0,80,0,0,0,111,0,245,0,0,0,211,0,0,0,71,0,114,0,245,0,99,0,191,0,251,0);
signal scenario_full  : scenario_type := (26,31,234,31,234,30,139,31,14,31,84,31,203,31,203,30,203,29,66,31,254,31,104,31,104,30,196,31,25,31,173,31,101,31,217,31,124,31,3,31,3,30,75,31,112,31,218,31,125,31,229,31,141,31,60,31,60,30,136,31,164,31,233,31,16,31,92,31,227,31,16,31,93,31,151,31,35,31,167,31,253,31,91,31,70,31,198,31,186,31,186,30,168,31,219,31,71,31,186,31,217,31,230,31,170,31,231,31,164,31,164,30,164,29,69,31,45,31,37,31,174,31,246,31,238,31,238,30,96,31,96,30,215,31,97,31,92,31,212,31,176,31,176,31,156,31,143,31,143,30,67,31,170,31,170,30,109,31,109,30,202,31,202,30,189,31,31,31,172,31,219,31,20,31,249,31,188,31,172,31,79,31,79,30,142,31,106,31,77,31,85,31,43,31,96,31,96,31,135,31,51,31,207,31,253,31,29,31,99,31,47,31,47,30,247,31,120,31,74,31,29,31,164,31,164,30,164,29,187,31,76,31,76,30,168,31,44,31,121,31,240,31,118,31,170,31,140,31,3,31,166,31,142,31,142,30,115,31,115,30,39,31,252,31,156,31,237,31,227,31,237,31,26,31,137,31,87,31,116,31,199,31,221,31,4,31,17,31,179,31,179,30,30,31,30,30,160,31,223,31,212,31,212,30,212,29,239,31,118,31,118,30,97,31,245,31,89,31,89,30,34,31,34,30,197,31,224,31,255,31,77,31,209,31,209,30,136,31,251,31,59,31,79,31,34,31,204,31,204,30,185,31,196,31,32,31,97,31,216,31,211,31,211,30,78,31,104,31,165,31,180,31,116,31,245,31,9,31,9,30,7,31,7,30,219,31,81,31,175,31,99,31,91,31,149,31,149,30,225,31,248,31,234,31,192,31,114,31,114,30,87,31,161,31,161,30,161,29,161,28,156,31,188,31,188,30,153,31,153,30,198,31,24,31,218,31,239,31,180,31,98,31,209,31,209,30,238,31,27,31,253,31,210,31,17,31,68,31,89,31,14,31,128,31,128,30,128,29,132,31,38,31,162,31,162,30,86,31,3,31,149,31,23,31,249,31,69,31,69,30,46,31,232,31,52,31,153,31,106,31,131,31,131,30,49,31,160,31,148,31,218,31,167,31,5,31,28,31,160,31,228,31,228,30,209,31,90,31,247,31,151,31,245,31,209,31,139,31,17,31,195,31,220,31,220,30,226,31,159,31,159,30,120,31,75,31,75,30,76,31,138,31,185,31,185,30,160,31,217,31,254,31,72,31,246,31,134,31,148,31,148,30,16,31,144,31,39,31,39,30,129,31,129,30,200,31,151,31,111,31,54,31,35,31,35,30,22,31,111,31,111,30,180,31,180,30,162,31,98,31,23,31,23,30,224,31,224,30,56,31,76,31,99,31,34,31,21,31,192,31,192,30,168,31,185,31,244,31,95,31,185,31,185,30,131,31,88,31,88,30,131,31,157,31,112,31,112,30,128,31,19,31,103,31,150,31,62,31,178,31,213,31,6,31,207,31,207,30,217,31,243,31,243,30,135,31,217,31,217,30,217,29,217,28,78,31,59,31,187,31,240,31,240,30,114,31,80,31,179,31,56,31,121,31,68,31,68,30,120,31,120,30,17,31,250,31,250,30,185,31,243,31,230,31,169,31,169,30,169,29,123,31,200,31,120,31,35,31,215,31,141,31,202,31,202,30,53,31,53,30,96,31,236,31,237,31,8,31,194,31,187,31,244,31,244,30,119,31,13,31,248,31,95,31,213,31,27,31,255,31,255,30,255,29,224,31,194,31,151,31,110,31,223,31,169,31,157,31,10,31,66,31,66,30,12,31,12,30,213,31,187,31,187,30,203,31,203,30,45,31,45,30,254,31,254,30,193,31,47,31,41,31,41,30,195,31,194,31,171,31,61,31,52,31,247,31,228,31,237,31,35,31,113,31,20,31,254,31,137,31,106,31,230,31,201,31,190,31,170,31,152,31,174,31,144,31,188,31,43,31,125,31,122,31,238,31,76,31,124,31,48,31,43,31,94,31,229,31,139,31,81,31,101,31,101,30,175,31,70,31,186,31,102,31,88,31,211,31,149,31,52,31,52,30,138,31,173,31,25,31,177,31,177,30,202,31,174,31,114,31,10,31,42,31,42,30,42,29,108,31,5,31,5,30,67,31,34,31,98,31,12,31,112,31,50,31,171,31,154,31,126,31,112,31,200,31,200,31,30,31,108,31,234,31,236,31,87,31,87,30,87,29,197,31,114,31,161,31,220,31,105,31,100,31,144,31,2,31,2,30,102,31,13,31,236,31,69,31,124,31,12,31,99,31,98,31,48,31,161,31,82,31,10,31,10,30,116,31,36,31,15,31,251,31,251,30,135,31,153,31,181,31,74,31,74,30,238,31,192,31,192,30,169,31,169,30,140,31,140,30,140,29,239,31,239,30,235,31,210,31,2,31,2,30,2,29,2,28,253,31,226,31,178,31,178,30,178,29,81,31,202,31,215,31,159,31,142,31,142,30,142,29,246,31,246,30,125,31,125,30,228,31,82,31,82,30,193,31,235,31,106,31,106,30,185,31,1,31,1,30,145,31,145,30,204,31,204,30,86,31,91,31,242,31,94,31,135,31,230,31,197,31,73,31,186,31,123,31,123,30,123,29,141,31,153,31,237,31,115,31,81,31,81,30,212,31,95,31,250,31,181,31,58,31,16,31,104,31,193,31,193,30,128,31,97,31,21,31,213,31,219,31,40,31,40,30,40,29,179,31,179,30,241,31,64,31,95,31,12,31,228,31,67,31,44,31,44,30,167,31,167,30,17,31,30,31,141,31,123,31,221,31,81,31,243,31,70,31,6,31,6,30,60,31,48,31,98,31,89,31,89,30,225,31,225,30,223,31,24,31,24,30,169,31,169,30,105,31,105,30,91,31,215,31,215,30,248,31,187,31,79,31,35,31,161,31,234,31,118,31,86,31,50,31,202,31,202,30,202,29,14,31,14,30,14,29,134,31,138,31,48,31,48,30,120,31,80,31,80,30,132,31,246,31,108,31,246,31,76,31,102,31,189,31,47,31,184,31,184,30,97,31,102,31,221,31,165,31,165,30,254,31,151,31,125,31,104,31,108,31,76,31,76,30,76,29,76,28,71,31,157,31,188,31,215,31,220,31,1,31,133,31,133,30,52,31,226,31,193,31,153,31,153,30,237,31,11,31,111,31,141,31,140,31,96,31,127,31,127,30,241,31,238,31,238,30,139,31,139,30,112,31,187,31,242,31,35,31,108,31,138,31,54,31,89,31,58,31,175,31,227,31,47,31,100,31,72,31,44,31,214,31,53,31,224,31,24,31,227,31,60,31,250,31,13,31,170,31,170,30,205,31,204,31,66,31,138,31,172,31,172,30,218,31,3,31,83,31,72,31,53,31,43,31,12,31,205,31,29,31,66,31,205,31,116,31,116,30,116,29,116,28,116,27,116,26,61,31,247,31,12,31,12,30,22,31,22,30,22,29,22,28,113,31,192,31,141,31,5,31,213,31,213,30,48,31,32,31,225,31,225,30,129,31,116,31,136,31,41,31,81,31,81,30,237,31,169,31,53,31,134,31,147,31,83,31,240,31,196,31,61,31,61,30,10,31,66,31,48,31,48,30,25,31,182,31,223,31,223,30,98,31,40,31,178,31,37,31,37,30,255,31,21,31,113,31,61,31,171,31,44,31,218,31,218,30,217,31,214,31,192,31,230,31,237,31,16,31,16,30,147,31,227,31,227,30,227,29,111,31,8,31,75,31,35,31,35,30,35,29,208,31,122,31,143,31,40,31,245,31,245,30,182,31,77,31,177,31,154,31,154,30,107,31,73,31,73,30,27,31,110,31,110,30,150,31,150,30,150,29,216,31,224,31,224,30,65,31,108,31,136,31,211,31,219,31,190,31,197,31,15,31,138,31,87,31,222,31,234,31,234,30,234,29,19,31,4,31,244,31,194,31,194,30,183,31,114,31,114,30,114,29,145,31,121,31,43,31,34,31,108,31,155,31,155,30,123,31,144,31,144,30,81,31,169,31,33,31,68,31,156,31,177,31,228,31,228,30,228,29,228,28,230,31,230,30,230,31,130,31,203,31,222,31,201,31,245,31,140,31,106,31,106,30,242,31,95,31,95,30,253,31,253,30,119,31,199,31,71,31,178,31,21,31,39,31,9,31,236,31,80,31,80,30,111,31,245,31,245,30,211,31,211,30,71,31,114,31,245,31,99,31,191,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
