-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_195 is
end project_tb_195;

architecture project_tb_arch_195 of project_tb_195 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 251;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,126,0,1,0,0,0,0,0,149,0,27,0,0,0,0,0,0,0,87,0,67,0,91,0,181,0,137,0,17,0,137,0,1,0,140,0,1,0,148,0,77,0,0,0,0,0,150,0,232,0,47,0,0,0,0,0,220,0,57,0,47,0,97,0,5,0,188,0,114,0,89,0,162,0,97,0,249,0,184,0,164,0,209,0,72,0,3,0,166,0,4,0,85,0,6,0,0,0,121,0,88,0,169,0,139,0,185,0,0,0,0,0,233,0,157,0,0,0,176,0,14,0,0,0,0,0,42,0,244,0,251,0,2,0,240,0,95,0,158,0,0,0,36,0,138,0,202,0,3,0,111,0,21,0,194,0,130,0,0,0,49,0,0,0,112,0,244,0,112,0,140,0,139,0,50,0,31,0,253,0,0,0,171,0,58,0,73,0,15,0,0,0,66,0,36,0,235,0,196,0,160,0,63,0,255,0,69,0,231,0,0,0,247,0,8,0,205,0,57,0,1,0,53,0,12,0,116,0,8,0,145,0,0,0,190,0,0,0,2,0,69,0,55,0,98,0,40,0,253,0,169,0,180,0,0,0,117,0,215,0,166,0,99,0,140,0,81,0,128,0,95,0,144,0,176,0,146,0,0,0,0,0,70,0,252,0,222,0,47,0,234,0,244,0,149,0,204,0,0,0,0,0,255,0,235,0,109,0,51,0,136,0,73,0,0,0,0,0,117,0,224,0,50,0,75,0,84,0,57,0,228,0,230,0,0,0,97,0,245,0,0,0,225,0,97,0,3,0,164,0,0,0,192,0,160,0,123,0,64,0,167,0,216,0,19,0,141,0,180,0,0,0,148,0,0,0,45,0,236,0,0,0,98,0,79,0,126,0,0,0,234,0,146,0,58,0,68,0,78,0,151,0,28,0,139,0,0,0,89,0,132,0,154,0,0,0,111,0,91,0,38,0,78,0,0,0,16,0,247,0,0,0,0,0,76,0,0,0,65,0,76,0,0,0,169,0,207,0,235,0,0,0,145,0,9,0,145,0,121,0,0,0,0,0,216,0,237,0,0,0,32,0,29,0,197,0,0,0,0,0,0,0,209,0,82,0,205,0,185,0,0,0,60,0,16,0,133,0,49,0);
signal scenario_full  : scenario_type := (0,0,126,31,1,31,1,30,1,29,149,31,27,31,27,30,27,29,27,28,87,31,67,31,91,31,181,31,137,31,17,31,137,31,1,31,140,31,1,31,148,31,77,31,77,30,77,29,150,31,232,31,47,31,47,30,47,29,220,31,57,31,47,31,97,31,5,31,188,31,114,31,89,31,162,31,97,31,249,31,184,31,164,31,209,31,72,31,3,31,166,31,4,31,85,31,6,31,6,30,121,31,88,31,169,31,139,31,185,31,185,30,185,29,233,31,157,31,157,30,176,31,14,31,14,30,14,29,42,31,244,31,251,31,2,31,240,31,95,31,158,31,158,30,36,31,138,31,202,31,3,31,111,31,21,31,194,31,130,31,130,30,49,31,49,30,112,31,244,31,112,31,140,31,139,31,50,31,31,31,253,31,253,30,171,31,58,31,73,31,15,31,15,30,66,31,36,31,235,31,196,31,160,31,63,31,255,31,69,31,231,31,231,30,247,31,8,31,205,31,57,31,1,31,53,31,12,31,116,31,8,31,145,31,145,30,190,31,190,30,2,31,69,31,55,31,98,31,40,31,253,31,169,31,180,31,180,30,117,31,215,31,166,31,99,31,140,31,81,31,128,31,95,31,144,31,176,31,146,31,146,30,146,29,70,31,252,31,222,31,47,31,234,31,244,31,149,31,204,31,204,30,204,29,255,31,235,31,109,31,51,31,136,31,73,31,73,30,73,29,117,31,224,31,50,31,75,31,84,31,57,31,228,31,230,31,230,30,97,31,245,31,245,30,225,31,97,31,3,31,164,31,164,30,192,31,160,31,123,31,64,31,167,31,216,31,19,31,141,31,180,31,180,30,148,31,148,30,45,31,236,31,236,30,98,31,79,31,126,31,126,30,234,31,146,31,58,31,68,31,78,31,151,31,28,31,139,31,139,30,89,31,132,31,154,31,154,30,111,31,91,31,38,31,78,31,78,30,16,31,247,31,247,30,247,29,76,31,76,30,65,31,76,31,76,30,169,31,207,31,235,31,235,30,145,31,9,31,145,31,121,31,121,30,121,29,216,31,237,31,237,30,32,31,29,31,197,31,197,30,197,29,197,28,209,31,82,31,205,31,185,31,185,30,60,31,16,31,133,31,49,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
