-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 824;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,45,0,226,0,191,0,210,0,149,0,148,0,117,0,0,0,0,0,18,0,0,0,240,0,170,0,215,0,0,0,155,0,0,0,130,0,247,0,62,0,0,0,124,0,81,0,0,0,27,0,178,0,64,0,5,0,106,0,91,0,117,0,83,0,121,0,184,0,233,0,202,0,76,0,0,0,161,0,243,0,94,0,0,0,86,0,33,0,221,0,145,0,188,0,6,0,1,0,180,0,0,0,177,0,65,0,33,0,235,0,93,0,151,0,58,0,0,0,151,0,97,0,84,0,201,0,160,0,39,0,76,0,102,0,216,0,202,0,0,0,76,0,61,0,72,0,0,0,217,0,0,0,67,0,0,0,28,0,20,0,203,0,0,0,187,0,246,0,49,0,0,0,121,0,0,0,0,0,0,0,0,0,83,0,115,0,104,0,224,0,22,0,0,0,146,0,182,0,141,0,217,0,241,0,55,0,148,0,125,0,229,0,132,0,156,0,210,0,0,0,45,0,18,0,0,0,0,0,133,0,30,0,236,0,33,0,10,0,0,0,180,0,145,0,0,0,153,0,171,0,153,0,0,0,20,0,239,0,147,0,50,0,0,0,71,0,0,0,183,0,154,0,33,0,84,0,192,0,112,0,0,0,162,0,222,0,0,0,0,0,142,0,137,0,15,0,131,0,92,0,149,0,36,0,152,0,131,0,208,0,151,0,0,0,75,0,0,0,101,0,33,0,148,0,28,0,196,0,53,0,68,0,121,0,250,0,26,0,0,0,86,0,0,0,18,0,205,0,0,0,139,0,177,0,202,0,184,0,0,0,33,0,133,0,170,0,0,0,22,0,246,0,21,0,53,0,57,0,116,0,0,0,38,0,0,0,0,0,239,0,103,0,65,0,92,0,0,0,0,0,47,0,143,0,200,0,118,0,0,0,4,0,49,0,40,0,193,0,72,0,71,0,107,0,163,0,79,0,148,0,94,0,87,0,243,0,11,0,0,0,53,0,153,0,242,0,63,0,107,0,123,0,73,0,112,0,13,0,0,0,53,0,211,0,166,0,107,0,140,0,229,0,188,0,151,0,123,0,76,0,250,0,0,0,219,0,237,0,58,0,0,0,45,0,121,0,205,0,81,0,221,0,178,0,70,0,94,0,189,0,5,0,0,0,41,0,37,0,32,0,140,0,16,0,0,0,106,0,0,0,0,0,0,0,207,0,59,0,253,0,103,0,197,0,0,0,174,0,115,0,216,0,0,0,0,0,46,0,0,0,47,0,207,0,57,0,0,0,0,0,175,0,232,0,0,0,126,0,175,0,167,0,201,0,0,0,202,0,181,0,104,0,0,0,36,0,219,0,0,0,6,0,2,0,122,0,169,0,167,0,192,0,164,0,130,0,202,0,6,0,44,0,124,0,255,0,220,0,203,0,0,0,111,0,161,0,115,0,130,0,69,0,228,0,113,0,59,0,205,0,66,0,204,0,241,0,232,0,93,0,227,0,0,0,157,0,237,0,0,0,223,0,100,0,21,0,54,0,202,0,85,0,243,0,187,0,160,0,164,0,0,0,190,0,218,0,227,0,146,0,0,0,225,0,245,0,6,0,207,0,110,0,194,0,28,0,49,0,0,0,12,0,80,0,75,0,0,0,0,0,186,0,58,0,0,0,215,0,92,0,129,0,89,0,227,0,67,0,0,0,69,0,7,0,7,0,36,0,67,0,45,0,153,0,165,0,28,0,148,0,253,0,16,0,10,0,71,0,107,0,0,0,184,0,71,0,0,0,5,0,15,0,181,0,49,0,158,0,52,0,143,0,83,0,155,0,5,0,0,0,193,0,0,0,85,0,21,0,155,0,229,0,170,0,193,0,97,0,68,0,243,0,58,0,32,0,37,0,188,0,211,0,186,0,0,0,48,0,114,0,166,0,0,0,0,0,214,0,0,0,160,0,105,0,209,0,45,0,193,0,0,0,38,0,62,0,0,0,205,0,1,0,0,0,56,0,0,0,131,0,0,0,152,0,90,0,234,0,187,0,52,0,62,0,0,0,79,0,134,0,4,0,52,0,121,0,0,0,91,0,176,0,154,0,74,0,108,0,0,0,254,0,0,0,223,0,185,0,171,0,132,0,54,0,241,0,202,0,124,0,162,0,0,0,36,0,187,0,74,0,0,0,230,0,112,0,175,0,56,0,64,0,135,0,0,0,135,0,57,0,221,0,6,0,253,0,156,0,103,0,0,0,0,0,193,0,175,0,166,0,176,0,116,0,8,0,187,0,0,0,103,0,15,0,74,0,220,0,86,0,177,0,18,0,182,0,181,0,58,0,98,0,195,0,237,0,187,0,97,0,201,0,119,0,22,0,174,0,70,0,47,0,225,0,18,0,73,0,188,0,171,0,249,0,120,0,209,0,0,0,0,0,1,0,24,0,155,0,87,0,166,0,6,0,0,0,94,0,163,0,1,0,70,0,155,0,0,0,218,0,0,0,166,0,160,0,233,0,0,0,0,0,95,0,7,0,232,0,0,0,84,0,60,0,155,0,243,0,57,0,250,0,114,0,0,0,202,0,83,0,40,0,231,0,0,0,13,0,163,0,72,0,242,0,241,0,90,0,221,0,86,0,144,0,0,0,128,0,55,0,73,0,0,0,130,0,169,0,217,0,171,0,87,0,252,0,0,0,186,0,19,0,25,0,244,0,0,0,0,0,119,0,81,0,0,0,64,0,132,0,33,0,184,0,0,0,0,0,184,0,184,0,169,0,0,0,94,0,165,0,82,0,47,0,232,0,101,0,0,0,190,0,181,0,78,0,62,0,245,0,0,0,46,0,252,0,46,0,113,0,108,0,214,0,161,0,97,0,198,0,43,0,152,0,0,0,5,0,26,0,228,0,18,0,142,0,0,0,136,0,181,0,186,0,0,0,36,0,100,0,120,0,0,0,134,0,0,0,87,0,47,0,53,0,119,0,19,0,0,0,153,0,111,0,66,0,49,0,71,0,0,0,4,0,249,0,0,0,21,0,117,0,110,0,227,0,215,0,213,0,83,0,203,0,4,0,65,0,225,0,171,0,0,0,83,0,97,0,0,0,16,0,193,0,0,0,194,0,158,0,220,0,119,0,71,0,122,0,151,0,0,0,110,0,0,0,248,0,0,0,183,0,185,0,0,0,151,0,0,0,0,0,37,0,0,0,0,0,97,0,82,0,218,0,0,0,30,0,36,0,0,0,0,0,131,0,0,0,85,0,107,0,125,0,161,0,231,0,134,0,58,0,96,0,68,0,200,0,31,0,57,0,230,0,236,0,0,0,197,0,0,0,219,0,133,0,0,0,0,0,250,0,250,0,120,0,135,0,0,0,163,0,76,0,187,0,0,0,203,0,58,0,196,0,17,0,223,0,40,0,190,0,77,0,15,0,0,0,18,0,0,0,0,0,9,0,0,0,0,0,0,0,209,0,235,0,178,0,100,0,216,0,177,0,143,0,235,0,246,0,168,0,0,0,242,0,202,0,238,0,239,0,127,0,188,0,0,0,182,0,122,0,126,0,118,0,11,0,92,0,182,0,0,0,215,0,178,0,198,0,0,0,0,0,162,0,234,0,12,0,38,0,0,0,20,0,0,0,0,0,80,0,0,0,0,0,217,0,37,0,0,0,0,0,66,0,155,0,0,0,46,0,242,0,4,0,195,0,0,0,147,0,165,0,230,0);
signal scenario_full  : scenario_type := (0,0,45,31,226,31,191,31,210,31,149,31,148,31,117,31,117,30,117,29,18,31,18,30,240,31,170,31,215,31,215,30,155,31,155,30,130,31,247,31,62,31,62,30,124,31,81,31,81,30,27,31,178,31,64,31,5,31,106,31,91,31,117,31,83,31,121,31,184,31,233,31,202,31,76,31,76,30,161,31,243,31,94,31,94,30,86,31,33,31,221,31,145,31,188,31,6,31,1,31,180,31,180,30,177,31,65,31,33,31,235,31,93,31,151,31,58,31,58,30,151,31,97,31,84,31,201,31,160,31,39,31,76,31,102,31,216,31,202,31,202,30,76,31,61,31,72,31,72,30,217,31,217,30,67,31,67,30,28,31,20,31,203,31,203,30,187,31,246,31,49,31,49,30,121,31,121,30,121,29,121,28,121,27,83,31,115,31,104,31,224,31,22,31,22,30,146,31,182,31,141,31,217,31,241,31,55,31,148,31,125,31,229,31,132,31,156,31,210,31,210,30,45,31,18,31,18,30,18,29,133,31,30,31,236,31,33,31,10,31,10,30,180,31,145,31,145,30,153,31,171,31,153,31,153,30,20,31,239,31,147,31,50,31,50,30,71,31,71,30,183,31,154,31,33,31,84,31,192,31,112,31,112,30,162,31,222,31,222,30,222,29,142,31,137,31,15,31,131,31,92,31,149,31,36,31,152,31,131,31,208,31,151,31,151,30,75,31,75,30,101,31,33,31,148,31,28,31,196,31,53,31,68,31,121,31,250,31,26,31,26,30,86,31,86,30,18,31,205,31,205,30,139,31,177,31,202,31,184,31,184,30,33,31,133,31,170,31,170,30,22,31,246,31,21,31,53,31,57,31,116,31,116,30,38,31,38,30,38,29,239,31,103,31,65,31,92,31,92,30,92,29,47,31,143,31,200,31,118,31,118,30,4,31,49,31,40,31,193,31,72,31,71,31,107,31,163,31,79,31,148,31,94,31,87,31,243,31,11,31,11,30,53,31,153,31,242,31,63,31,107,31,123,31,73,31,112,31,13,31,13,30,53,31,211,31,166,31,107,31,140,31,229,31,188,31,151,31,123,31,76,31,250,31,250,30,219,31,237,31,58,31,58,30,45,31,121,31,205,31,81,31,221,31,178,31,70,31,94,31,189,31,5,31,5,30,41,31,37,31,32,31,140,31,16,31,16,30,106,31,106,30,106,29,106,28,207,31,59,31,253,31,103,31,197,31,197,30,174,31,115,31,216,31,216,30,216,29,46,31,46,30,47,31,207,31,57,31,57,30,57,29,175,31,232,31,232,30,126,31,175,31,167,31,201,31,201,30,202,31,181,31,104,31,104,30,36,31,219,31,219,30,6,31,2,31,122,31,169,31,167,31,192,31,164,31,130,31,202,31,6,31,44,31,124,31,255,31,220,31,203,31,203,30,111,31,161,31,115,31,130,31,69,31,228,31,113,31,59,31,205,31,66,31,204,31,241,31,232,31,93,31,227,31,227,30,157,31,237,31,237,30,223,31,100,31,21,31,54,31,202,31,85,31,243,31,187,31,160,31,164,31,164,30,190,31,218,31,227,31,146,31,146,30,225,31,245,31,6,31,207,31,110,31,194,31,28,31,49,31,49,30,12,31,80,31,75,31,75,30,75,29,186,31,58,31,58,30,215,31,92,31,129,31,89,31,227,31,67,31,67,30,69,31,7,31,7,31,36,31,67,31,45,31,153,31,165,31,28,31,148,31,253,31,16,31,10,31,71,31,107,31,107,30,184,31,71,31,71,30,5,31,15,31,181,31,49,31,158,31,52,31,143,31,83,31,155,31,5,31,5,30,193,31,193,30,85,31,21,31,155,31,229,31,170,31,193,31,97,31,68,31,243,31,58,31,32,31,37,31,188,31,211,31,186,31,186,30,48,31,114,31,166,31,166,30,166,29,214,31,214,30,160,31,105,31,209,31,45,31,193,31,193,30,38,31,62,31,62,30,205,31,1,31,1,30,56,31,56,30,131,31,131,30,152,31,90,31,234,31,187,31,52,31,62,31,62,30,79,31,134,31,4,31,52,31,121,31,121,30,91,31,176,31,154,31,74,31,108,31,108,30,254,31,254,30,223,31,185,31,171,31,132,31,54,31,241,31,202,31,124,31,162,31,162,30,36,31,187,31,74,31,74,30,230,31,112,31,175,31,56,31,64,31,135,31,135,30,135,31,57,31,221,31,6,31,253,31,156,31,103,31,103,30,103,29,193,31,175,31,166,31,176,31,116,31,8,31,187,31,187,30,103,31,15,31,74,31,220,31,86,31,177,31,18,31,182,31,181,31,58,31,98,31,195,31,237,31,187,31,97,31,201,31,119,31,22,31,174,31,70,31,47,31,225,31,18,31,73,31,188,31,171,31,249,31,120,31,209,31,209,30,209,29,1,31,24,31,155,31,87,31,166,31,6,31,6,30,94,31,163,31,1,31,70,31,155,31,155,30,218,31,218,30,166,31,160,31,233,31,233,30,233,29,95,31,7,31,232,31,232,30,84,31,60,31,155,31,243,31,57,31,250,31,114,31,114,30,202,31,83,31,40,31,231,31,231,30,13,31,163,31,72,31,242,31,241,31,90,31,221,31,86,31,144,31,144,30,128,31,55,31,73,31,73,30,130,31,169,31,217,31,171,31,87,31,252,31,252,30,186,31,19,31,25,31,244,31,244,30,244,29,119,31,81,31,81,30,64,31,132,31,33,31,184,31,184,30,184,29,184,31,184,31,169,31,169,30,94,31,165,31,82,31,47,31,232,31,101,31,101,30,190,31,181,31,78,31,62,31,245,31,245,30,46,31,252,31,46,31,113,31,108,31,214,31,161,31,97,31,198,31,43,31,152,31,152,30,5,31,26,31,228,31,18,31,142,31,142,30,136,31,181,31,186,31,186,30,36,31,100,31,120,31,120,30,134,31,134,30,87,31,47,31,53,31,119,31,19,31,19,30,153,31,111,31,66,31,49,31,71,31,71,30,4,31,249,31,249,30,21,31,117,31,110,31,227,31,215,31,213,31,83,31,203,31,4,31,65,31,225,31,171,31,171,30,83,31,97,31,97,30,16,31,193,31,193,30,194,31,158,31,220,31,119,31,71,31,122,31,151,31,151,30,110,31,110,30,248,31,248,30,183,31,185,31,185,30,151,31,151,30,151,29,37,31,37,30,37,29,97,31,82,31,218,31,218,30,30,31,36,31,36,30,36,29,131,31,131,30,85,31,107,31,125,31,161,31,231,31,134,31,58,31,96,31,68,31,200,31,31,31,57,31,230,31,236,31,236,30,197,31,197,30,219,31,133,31,133,30,133,29,250,31,250,31,120,31,135,31,135,30,163,31,76,31,187,31,187,30,203,31,58,31,196,31,17,31,223,31,40,31,190,31,77,31,15,31,15,30,18,31,18,30,18,29,9,31,9,30,9,29,9,28,209,31,235,31,178,31,100,31,216,31,177,31,143,31,235,31,246,31,168,31,168,30,242,31,202,31,238,31,239,31,127,31,188,31,188,30,182,31,122,31,126,31,118,31,11,31,92,31,182,31,182,30,215,31,178,31,198,31,198,30,198,29,162,31,234,31,12,31,38,31,38,30,20,31,20,30,20,29,80,31,80,30,80,29,217,31,37,31,37,30,37,29,66,31,155,31,155,30,46,31,242,31,4,31,195,31,195,30,147,31,165,31,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
