-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_863 is
end project_tb_863;

architecture project_tb_arch_863 of project_tb_863 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 340;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (254,0,77,0,0,0,45,0,111,0,157,0,88,0,122,0,85,0,195,0,234,0,212,0,255,0,225,0,190,0,0,0,118,0,155,0,74,0,158,0,225,0,0,0,121,0,5,0,92,0,218,0,159,0,0,0,189,0,169,0,183,0,46,0,107,0,208,0,160,0,75,0,0,0,162,0,135,0,163,0,6,0,51,0,197,0,104,0,157,0,89,0,110,0,199,0,234,0,229,0,183,0,116,0,33,0,20,0,0,0,147,0,121,0,11,0,0,0,15,0,60,0,30,0,32,0,0,0,169,0,181,0,18,0,74,0,158,0,0,0,185,0,0,0,239,0,93,0,121,0,221,0,0,0,252,0,0,0,7,0,196,0,0,0,151,0,88,0,65,0,58,0,0,0,171,0,147,0,0,0,154,0,0,0,33,0,57,0,0,0,230,0,40,0,170,0,94,0,193,0,204,0,0,0,58,0,87,0,180,0,101,0,89,0,15,0,245,0,117,0,14,0,230,0,228,0,41,0,10,0,25,0,190,0,0,0,222,0,0,0,187,0,31,0,253,0,208,0,11,0,0,0,201,0,141,0,244,0,85,0,184,0,201,0,144,0,154,0,244,0,23,0,172,0,25,0,104,0,244,0,17,0,195,0,173,0,200,0,0,0,145,0,196,0,0,0,253,0,203,0,0,0,143,0,0,0,0,0,166,0,107,0,32,0,34,0,153,0,185,0,211,0,204,0,182,0,60,0,0,0,0,0,0,0,56,0,41,0,84,0,124,0,0,0,0,0,185,0,172,0,6,0,0,0,0,0,44,0,191,0,123,0,35,0,0,0,132,0,146,0,107,0,242,0,0,0,0,0,226,0,0,0,0,0,99,0,160,0,251,0,228,0,140,0,159,0,79,0,159,0,21,0,0,0,0,0,0,0,13,0,38,0,250,0,90,0,203,0,165,0,207,0,13,0,0,0,241,0,0,0,59,0,0,0,17,0,222,0,131,0,226,0,0,0,17,0,126,0,191,0,229,0,0,0,59,0,151,0,51,0,132,0,5,0,190,0,152,0,201,0,247,0,116,0,220,0,110,0,98,0,212,0,57,0,237,0,85,0,0,0,156,0,80,0,21,0,243,0,234,0,155,0,215,0,161,0,83,0,0,0,97,0,233,0,31,0,0,0,216,0,81,0,91,0,0,0,0,0,24,0,196,0,181,0,96,0,164,0,0,0,150,0,192,0,124,0,9,0,31,0,127,0,191,0,252,0,189,0,249,0,24,0,52,0,244,0,0,0,0,0,58,0,241,0,105,0,0,0,74,0,144,0,60,0,52,0,13,0,0,0,0,0,29,0,219,0,186,0,46,0,178,0,0,0,92,0,0,0,149,0,17,0,49,0,0,0,140,0,198,0,173,0,129,0,0,0,176,0,156,0,0,0,198,0,24,0,200,0,0,0,239,0,194,0,87,0,0,0,142,0,6,0,68,0,13,0,176,0,0,0,58,0,51,0,147,0,62,0,0,0,185,0,30,0,151,0,196,0,204,0);
signal scenario_full  : scenario_type := (254,31,77,31,77,30,45,31,111,31,157,31,88,31,122,31,85,31,195,31,234,31,212,31,255,31,225,31,190,31,190,30,118,31,155,31,74,31,158,31,225,31,225,30,121,31,5,31,92,31,218,31,159,31,159,30,189,31,169,31,183,31,46,31,107,31,208,31,160,31,75,31,75,30,162,31,135,31,163,31,6,31,51,31,197,31,104,31,157,31,89,31,110,31,199,31,234,31,229,31,183,31,116,31,33,31,20,31,20,30,147,31,121,31,11,31,11,30,15,31,60,31,30,31,32,31,32,30,169,31,181,31,18,31,74,31,158,31,158,30,185,31,185,30,239,31,93,31,121,31,221,31,221,30,252,31,252,30,7,31,196,31,196,30,151,31,88,31,65,31,58,31,58,30,171,31,147,31,147,30,154,31,154,30,33,31,57,31,57,30,230,31,40,31,170,31,94,31,193,31,204,31,204,30,58,31,87,31,180,31,101,31,89,31,15,31,245,31,117,31,14,31,230,31,228,31,41,31,10,31,25,31,190,31,190,30,222,31,222,30,187,31,31,31,253,31,208,31,11,31,11,30,201,31,141,31,244,31,85,31,184,31,201,31,144,31,154,31,244,31,23,31,172,31,25,31,104,31,244,31,17,31,195,31,173,31,200,31,200,30,145,31,196,31,196,30,253,31,203,31,203,30,143,31,143,30,143,29,166,31,107,31,32,31,34,31,153,31,185,31,211,31,204,31,182,31,60,31,60,30,60,29,60,28,56,31,41,31,84,31,124,31,124,30,124,29,185,31,172,31,6,31,6,30,6,29,44,31,191,31,123,31,35,31,35,30,132,31,146,31,107,31,242,31,242,30,242,29,226,31,226,30,226,29,99,31,160,31,251,31,228,31,140,31,159,31,79,31,159,31,21,31,21,30,21,29,21,28,13,31,38,31,250,31,90,31,203,31,165,31,207,31,13,31,13,30,241,31,241,30,59,31,59,30,17,31,222,31,131,31,226,31,226,30,17,31,126,31,191,31,229,31,229,30,59,31,151,31,51,31,132,31,5,31,190,31,152,31,201,31,247,31,116,31,220,31,110,31,98,31,212,31,57,31,237,31,85,31,85,30,156,31,80,31,21,31,243,31,234,31,155,31,215,31,161,31,83,31,83,30,97,31,233,31,31,31,31,30,216,31,81,31,91,31,91,30,91,29,24,31,196,31,181,31,96,31,164,31,164,30,150,31,192,31,124,31,9,31,31,31,127,31,191,31,252,31,189,31,249,31,24,31,52,31,244,31,244,30,244,29,58,31,241,31,105,31,105,30,74,31,144,31,60,31,52,31,13,31,13,30,13,29,29,31,219,31,186,31,46,31,178,31,178,30,92,31,92,30,149,31,17,31,49,31,49,30,140,31,198,31,173,31,129,31,129,30,176,31,156,31,156,30,198,31,24,31,200,31,200,30,239,31,194,31,87,31,87,30,142,31,6,31,68,31,13,31,176,31,176,30,58,31,51,31,147,31,62,31,62,30,185,31,30,31,151,31,196,31,204,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
