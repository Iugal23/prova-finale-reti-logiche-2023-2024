-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_636 is
end project_tb_636;

architecture project_tb_arch_636 of project_tb_636 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 710;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,61,0,198,0,162,0,122,0,23,0,86,0,147,0,64,0,143,0,240,0,0,0,155,0,225,0,238,0,92,0,45,0,162,0,133,0,118,0,246,0,140,0,217,0,172,0,218,0,194,0,81,0,232,0,231,0,93,0,252,0,41,0,30,0,227,0,50,0,210,0,0,0,45,0,242,0,221,0,98,0,175,0,112,0,238,0,41,0,126,0,55,0,249,0,13,0,112,0,41,0,0,0,57,0,0,0,123,0,167,0,0,0,0,0,154,0,0,0,75,0,49,0,152,0,172,0,0,0,186,0,19,0,9,0,36,0,228,0,245,0,50,0,222,0,177,0,52,0,168,0,51,0,125,0,0,0,204,0,24,0,205,0,54,0,133,0,0,0,40,0,0,0,43,0,106,0,96,0,179,0,0,0,166,0,160,0,241,0,199,0,131,0,186,0,2,0,96,0,144,0,6,0,0,0,175,0,231,0,157,0,0,0,176,0,147,0,79,0,148,0,64,0,43,0,135,0,255,0,0,0,0,0,0,0,189,0,126,0,135,0,184,0,47,0,106,0,90,0,163,0,43,0,163,0,170,0,0,0,229,0,5,0,29,0,0,0,172,0,112,0,245,0,139,0,0,0,44,0,36,0,0,0,122,0,0,0,86,0,130,0,83,0,79,0,231,0,157,0,36,0,230,0,2,0,226,0,0,0,2,0,138,0,212,0,161,0,0,0,0,0,94,0,133,0,0,0,163,0,221,0,0,0,18,0,13,0,143,0,140,0,0,0,7,0,169,0,208,0,77,0,0,0,220,0,35,0,3,0,0,0,130,0,123,0,103,0,0,0,0,0,151,0,0,0,16,0,0,0,0,0,130,0,190,0,147,0,198,0,245,0,117,0,79,0,65,0,0,0,252,0,0,0,120,0,144,0,0,0,160,0,42,0,54,0,91,0,0,0,0,0,113,0,38,0,28,0,36,0,0,0,0,0,250,0,98,0,220,0,156,0,21,0,0,0,0,0,157,0,182,0,34,0,93,0,198,0,107,0,254,0,0,0,212,0,0,0,163,0,80,0,123,0,31,0,216,0,63,0,159,0,162,0,0,0,221,0,125,0,104,0,171,0,197,0,65,0,0,0,141,0,21,0,226,0,112,0,230,0,3,0,0,0,27,0,0,0,125,0,204,0,164,0,139,0,108,0,60,0,227,0,30,0,141,0,209,0,56,0,43,0,0,0,0,0,18,0,205,0,96,0,255,0,171,0,187,0,100,0,212,0,0,0,0,0,226,0,50,0,0,0,195,0,79,0,0,0,233,0,80,0,199,0,159,0,0,0,17,0,48,0,9,0,43,0,232,0,29,0,219,0,235,0,130,0,0,0,7,0,222,0,214,0,123,0,85,0,220,0,28,0,4,0,156,0,148,0,126,0,32,0,0,0,20,0,178,0,169,0,0,0,0,0,108,0,11,0,41,0,202,0,227,0,13,0,0,0,113,0,3,0,207,0,88,0,110,0,153,0,0,0,0,0,130,0,53,0,47,0,221,0,70,0,0,0,175,0,251,0,205,0,9,0,60,0,153,0,0,0,149,0,235,0,0,0,188,0,131,0,64,0,152,0,12,0,2,0,136,0,25,0,117,0,244,0,154,0,128,0,208,0,0,0,0,0,133,0,99,0,8,0,0,0,112,0,43,0,117,0,218,0,17,0,13,0,117,0,118,0,229,0,118,0,58,0,223,0,0,0,0,0,55,0,76,0,0,0,37,0,194,0,0,0,81,0,215,0,28,0,0,0,22,0,0,0,0,0,254,0,159,0,108,0,230,0,64,0,121,0,54,0,91,0,228,0,75,0,133,0,0,0,0,0,224,0,0,0,87,0,51,0,121,0,159,0,251,0,0,0,37,0,85,0,183,0,0,0,140,0,0,0,201,0,80,0,225,0,52,0,135,0,94,0,202,0,242,0,0,0,39,0,223,0,4,0,179,0,210,0,32,0,29,0,106,0,19,0,150,0,0,0,141,0,124,0,139,0,0,0,0,0,35,0,18,0,174,0,2,0,182,0,49,0,238,0,136,0,34,0,138,0,154,0,196,0,0,0,123,0,182,0,176,0,0,0,50,0,95,0,98,0,0,0,197,0,148,0,125,0,126,0,37,0,150,0,146,0,214,0,76,0,239,0,141,0,53,0,0,0,41,0,152,0,239,0,0,0,0,0,222,0,67,0,171,0,111,0,186,0,141,0,99,0,31,0,90,0,0,0,206,0,23,0,0,0,0,0,163,0,8,0,0,0,208,0,60,0,137,0,221,0,191,0,0,0,247,0,140,0,82,0,75,0,102,0,38,0,154,0,174,0,142,0,237,0,131,0,172,0,148,0,0,0,171,0,109,0,168,0,213,0,252,0,182,0,91,0,0,0,0,0,74,0,250,0,141,0,50,0,236,0,245,0,59,0,91,0,0,0,103,0,38,0,31,0,0,0,154,0,122,0,51,0,184,0,80,0,177,0,219,0,121,0,59,0,155,0,129,0,0,0,169,0,204,0,250,0,232,0,129,0,37,0,130,0,104,0,102,0,205,0,244,0,148,0,57,0,37,0,249,0,88,0,0,0,0,0,0,0,107,0,231,0,172,0,0,0,45,0,63,0,219,0,240,0,148,0,68,0,0,0,0,0,78,0,38,0,195,0,114,0,28,0,117,0,234,0,142,0,53,0,160,0,13,0,69,0,0,0,0,0,207,0,141,0,202,0,24,0,90,0,228,0,0,0,216,0,10,0,94,0,0,0,17,0,193,0,0,0,3,0,46,0,88,0,0,0,8,0,191,0,47,0,7,0,0,0,0,0,0,0,214,0,199,0,0,0,219,0,79,0,84,0,0,0,128,0,68,0,0,0,0,0,89,0,179,0,243,0,39,0,55,0,151,0,72,0,0,0,73,0,0,0,242,0,237,0,129,0,97,0,0,0,0,0,0,0,255,0,30,0,49,0,196,0,199,0,70,0,203,0,179,0,142,0,30,0,252,0,0,0,64,0,232,0,71,0,199,0,195,0,246,0,123,0,29,0,177,0,200,0,223,0,0,0,233,0,64,0,190,0,253,0,241,0,138,0,98,0,0,0,44,0,35,0,189,0,24,0,32,0,141,0,0,0,39,0,91,0,201,0,0,0,189,0,68,0,3,0,105,0,113,0,67,0,223,0,23,0);
signal scenario_full  : scenario_type := (0,0,61,31,198,31,162,31,122,31,23,31,86,31,147,31,64,31,143,31,240,31,240,30,155,31,225,31,238,31,92,31,45,31,162,31,133,31,118,31,246,31,140,31,217,31,172,31,218,31,194,31,81,31,232,31,231,31,93,31,252,31,41,31,30,31,227,31,50,31,210,31,210,30,45,31,242,31,221,31,98,31,175,31,112,31,238,31,41,31,126,31,55,31,249,31,13,31,112,31,41,31,41,30,57,31,57,30,123,31,167,31,167,30,167,29,154,31,154,30,75,31,49,31,152,31,172,31,172,30,186,31,19,31,9,31,36,31,228,31,245,31,50,31,222,31,177,31,52,31,168,31,51,31,125,31,125,30,204,31,24,31,205,31,54,31,133,31,133,30,40,31,40,30,43,31,106,31,96,31,179,31,179,30,166,31,160,31,241,31,199,31,131,31,186,31,2,31,96,31,144,31,6,31,6,30,175,31,231,31,157,31,157,30,176,31,147,31,79,31,148,31,64,31,43,31,135,31,255,31,255,30,255,29,255,28,189,31,126,31,135,31,184,31,47,31,106,31,90,31,163,31,43,31,163,31,170,31,170,30,229,31,5,31,29,31,29,30,172,31,112,31,245,31,139,31,139,30,44,31,36,31,36,30,122,31,122,30,86,31,130,31,83,31,79,31,231,31,157,31,36,31,230,31,2,31,226,31,226,30,2,31,138,31,212,31,161,31,161,30,161,29,94,31,133,31,133,30,163,31,221,31,221,30,18,31,13,31,143,31,140,31,140,30,7,31,169,31,208,31,77,31,77,30,220,31,35,31,3,31,3,30,130,31,123,31,103,31,103,30,103,29,151,31,151,30,16,31,16,30,16,29,130,31,190,31,147,31,198,31,245,31,117,31,79,31,65,31,65,30,252,31,252,30,120,31,144,31,144,30,160,31,42,31,54,31,91,31,91,30,91,29,113,31,38,31,28,31,36,31,36,30,36,29,250,31,98,31,220,31,156,31,21,31,21,30,21,29,157,31,182,31,34,31,93,31,198,31,107,31,254,31,254,30,212,31,212,30,163,31,80,31,123,31,31,31,216,31,63,31,159,31,162,31,162,30,221,31,125,31,104,31,171,31,197,31,65,31,65,30,141,31,21,31,226,31,112,31,230,31,3,31,3,30,27,31,27,30,125,31,204,31,164,31,139,31,108,31,60,31,227,31,30,31,141,31,209,31,56,31,43,31,43,30,43,29,18,31,205,31,96,31,255,31,171,31,187,31,100,31,212,31,212,30,212,29,226,31,50,31,50,30,195,31,79,31,79,30,233,31,80,31,199,31,159,31,159,30,17,31,48,31,9,31,43,31,232,31,29,31,219,31,235,31,130,31,130,30,7,31,222,31,214,31,123,31,85,31,220,31,28,31,4,31,156,31,148,31,126,31,32,31,32,30,20,31,178,31,169,31,169,30,169,29,108,31,11,31,41,31,202,31,227,31,13,31,13,30,113,31,3,31,207,31,88,31,110,31,153,31,153,30,153,29,130,31,53,31,47,31,221,31,70,31,70,30,175,31,251,31,205,31,9,31,60,31,153,31,153,30,149,31,235,31,235,30,188,31,131,31,64,31,152,31,12,31,2,31,136,31,25,31,117,31,244,31,154,31,128,31,208,31,208,30,208,29,133,31,99,31,8,31,8,30,112,31,43,31,117,31,218,31,17,31,13,31,117,31,118,31,229,31,118,31,58,31,223,31,223,30,223,29,55,31,76,31,76,30,37,31,194,31,194,30,81,31,215,31,28,31,28,30,22,31,22,30,22,29,254,31,159,31,108,31,230,31,64,31,121,31,54,31,91,31,228,31,75,31,133,31,133,30,133,29,224,31,224,30,87,31,51,31,121,31,159,31,251,31,251,30,37,31,85,31,183,31,183,30,140,31,140,30,201,31,80,31,225,31,52,31,135,31,94,31,202,31,242,31,242,30,39,31,223,31,4,31,179,31,210,31,32,31,29,31,106,31,19,31,150,31,150,30,141,31,124,31,139,31,139,30,139,29,35,31,18,31,174,31,2,31,182,31,49,31,238,31,136,31,34,31,138,31,154,31,196,31,196,30,123,31,182,31,176,31,176,30,50,31,95,31,98,31,98,30,197,31,148,31,125,31,126,31,37,31,150,31,146,31,214,31,76,31,239,31,141,31,53,31,53,30,41,31,152,31,239,31,239,30,239,29,222,31,67,31,171,31,111,31,186,31,141,31,99,31,31,31,90,31,90,30,206,31,23,31,23,30,23,29,163,31,8,31,8,30,208,31,60,31,137,31,221,31,191,31,191,30,247,31,140,31,82,31,75,31,102,31,38,31,154,31,174,31,142,31,237,31,131,31,172,31,148,31,148,30,171,31,109,31,168,31,213,31,252,31,182,31,91,31,91,30,91,29,74,31,250,31,141,31,50,31,236,31,245,31,59,31,91,31,91,30,103,31,38,31,31,31,31,30,154,31,122,31,51,31,184,31,80,31,177,31,219,31,121,31,59,31,155,31,129,31,129,30,169,31,204,31,250,31,232,31,129,31,37,31,130,31,104,31,102,31,205,31,244,31,148,31,57,31,37,31,249,31,88,31,88,30,88,29,88,28,107,31,231,31,172,31,172,30,45,31,63,31,219,31,240,31,148,31,68,31,68,30,68,29,78,31,38,31,195,31,114,31,28,31,117,31,234,31,142,31,53,31,160,31,13,31,69,31,69,30,69,29,207,31,141,31,202,31,24,31,90,31,228,31,228,30,216,31,10,31,94,31,94,30,17,31,193,31,193,30,3,31,46,31,88,31,88,30,8,31,191,31,47,31,7,31,7,30,7,29,7,28,214,31,199,31,199,30,219,31,79,31,84,31,84,30,128,31,68,31,68,30,68,29,89,31,179,31,243,31,39,31,55,31,151,31,72,31,72,30,73,31,73,30,242,31,237,31,129,31,97,31,97,30,97,29,97,28,255,31,30,31,49,31,196,31,199,31,70,31,203,31,179,31,142,31,30,31,252,31,252,30,64,31,232,31,71,31,199,31,195,31,246,31,123,31,29,31,177,31,200,31,223,31,223,30,233,31,64,31,190,31,253,31,241,31,138,31,98,31,98,30,44,31,35,31,189,31,24,31,32,31,141,31,141,30,39,31,91,31,201,31,201,30,189,31,68,31,3,31,105,31,113,31,67,31,223,31,23,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
