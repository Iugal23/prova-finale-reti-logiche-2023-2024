-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 653;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (177,0,18,0,171,0,0,0,0,0,26,0,142,0,103,0,139,0,73,0,228,0,87,0,77,0,153,0,5,0,89,0,248,0,48,0,53,0,53,0,144,0,113,0,124,0,180,0,0,0,148,0,0,0,8,0,0,0,108,0,32,0,179,0,12,0,224,0,0,0,70,0,43,0,0,0,119,0,108,0,0,0,157,0,208,0,236,0,12,0,85,0,107,0,114,0,103,0,149,0,41,0,110,0,210,0,0,0,139,0,140,0,0,0,113,0,238,0,0,0,0,0,0,0,0,0,255,0,0,0,248,0,248,0,92,0,63,0,125,0,219,0,0,0,75,0,216,0,244,0,36,0,119,0,106,0,0,0,231,0,84,0,203,0,207,0,60,0,111,0,113,0,37,0,237,0,0,0,0,0,45,0,148,0,5,0,182,0,14,0,210,0,224,0,233,0,0,0,0,0,201,0,38,0,148,0,153,0,43,0,63,0,94,0,223,0,13,0,248,0,198,0,43,0,200,0,109,0,0,0,227,0,190,0,175,0,25,0,0,0,17,0,152,0,64,0,0,0,156,0,241,0,163,0,49,0,173,0,136,0,128,0,0,0,0,0,24,0,222,0,0,0,0,0,212,0,0,0,0,0,36,0,133,0,194,0,197,0,173,0,179,0,3,0,122,0,62,0,0,0,167,0,215,0,95,0,96,0,69,0,0,0,143,0,142,0,173,0,110,0,80,0,96,0,203,0,236,0,116,0,0,0,111,0,105,0,85,0,169,0,228,0,127,0,104,0,0,0,0,0,114,0,181,0,0,0,0,0,49,0,222,0,12,0,0,0,110,0,125,0,0,0,172,0,0,0,2,0,0,0,123,0,0,0,53,0,215,0,9,0,224,0,84,0,153,0,58,0,57,0,0,0,184,0,176,0,134,0,39,0,58,0,0,0,204,0,119,0,223,0,130,0,248,0,4,0,128,0,64,0,71,0,161,0,38,0,113,0,174,0,65,0,0,0,59,0,0,0,145,0,19,0,0,0,0,0,217,0,203,0,174,0,3,0,154,0,127,0,92,0,238,0,70,0,0,0,177,0,203,0,19,0,0,0,0,0,70,0,0,0,0,0,149,0,100,0,0,0,249,0,0,0,237,0,135,0,209,0,1,0,189,0,0,0,186,0,119,0,177,0,46,0,56,0,90,0,254,0,102,0,24,0,4,0,67,0,242,0,202,0,179,0,115,0,126,0,64,0,229,0,0,0,141,0,156,0,79,0,0,0,114,0,153,0,209,0,244,0,2,0,202,0,18,0,0,0,101,0,0,0,92,0,0,0,0,0,215,0,225,0,140,0,0,0,195,0,120,0,204,0,17,0,61,0,0,0,0,0,82,0,0,0,221,0,231,0,108,0,204,0,162,0,163,0,53,0,114,0,202,0,99,0,54,0,253,0,192,0,63,0,0,0,133,0,217,0,35,0,130,0,0,0,237,0,193,0,160,0,0,0,0,0,178,0,191,0,121,0,0,0,190,0,39,0,162,0,157,0,36,0,220,0,0,0,104,0,207,0,61,0,114,0,0,0,40,0,0,0,55,0,36,0,205,0,224,0,200,0,127,0,85,0,237,0,191,0,0,0,21,0,200,0,216,0,245,0,96,0,29,0,133,0,0,0,213,0,46,0,41,0,217,0,0,0,65,0,59,0,232,0,0,0,157,0,63,0,187,0,170,0,34,0,92,0,52,0,171,0,203,0,7,0,194,0,30,0,73,0,186,0,177,0,226,0,91,0,0,0,0,0,0,0,41,0,0,0,7,0,255,0,0,0,223,0,27,0,0,0,237,0,158,0,59,0,88,0,64,0,119,0,184,0,0,0,104,0,0,0,3,0,83,0,13,0,0,0,177,0,9,0,71,0,170,0,0,0,162,0,130,0,9,0,146,0,0,0,220,0,235,0,139,0,189,0,53,0,124,0,101,0,107,0,15,0,69,0,183,0,122,0,14,0,129,0,62,0,195,0,141,0,57,0,167,0,100,0,141,0,38,0,200,0,249,0,86,0,0,0,3,0,240,0,49,0,97,0,155,0,0,0,111,0,214,0,0,0,74,0,244,0,16,0,26,0,186,0,127,0,193,0,157,0,69,0,218,0,85,0,216,0,80,0,161,0,159,0,255,0,253,0,69,0,236,0,0,0,225,0,28,0,7,0,164,0,155,0,0,0,92,0,147,0,0,0,61,0,0,0,247,0,208,0,147,0,237,0,69,0,84,0,0,0,120,0,170,0,218,0,27,0,54,0,135,0,0,0,75,0,0,0,207,0,143,0,77,0,54,0,216,0,39,0,0,0,55,0,43,0,0,0,0,0,192,0,237,0,62,0,232,0,93,0,6,0,181,0,0,0,202,0,0,0,34,0,75,0,0,0,0,0,0,0,243,0,33,0,213,0,0,0,121,0,0,0,0,0,53,0,110,0,186,0,107,0,0,0,249,0,221,0,49,0,75,0,0,0,105,0,0,0,107,0,166,0,191,0,207,0,28,0,0,0,217,0,194,0,0,0,25,0,156,0,74,0,125,0,248,0,36,0,251,0,55,0,229,0,15,0,215,0,15,0,244,0,142,0,0,0,156,0,122,0,119,0,222,0,71,0,8,0,207,0,0,0,121,0,0,0,42,0,49,0,113,0,95,0,224,0,137,0,200,0,0,0,62,0,210,0,97,0,0,0,132,0,41,0,0,0,167,0,0,0,68,0,169,0,2,0,126,0,0,0,0,0,169,0,38,0,0,0,70,0,127,0,72,0,94,0,102,0,185,0,0,0,129,0,0,0,69,0,249,0,247,0,116,0,229,0,228,0,221,0,44,0,0,0,36,0,114,0,34,0,53,0,235,0,24,0,150,0,31,0,119,0,143,0,146,0,239,0,0,0,36,0,101,0,75,0,118,0,48,0,21,0,99,0);
signal scenario_full  : scenario_type := (177,31,18,31,171,31,171,30,171,29,26,31,142,31,103,31,139,31,73,31,228,31,87,31,77,31,153,31,5,31,89,31,248,31,48,31,53,31,53,31,144,31,113,31,124,31,180,31,180,30,148,31,148,30,8,31,8,30,108,31,32,31,179,31,12,31,224,31,224,30,70,31,43,31,43,30,119,31,108,31,108,30,157,31,208,31,236,31,12,31,85,31,107,31,114,31,103,31,149,31,41,31,110,31,210,31,210,30,139,31,140,31,140,30,113,31,238,31,238,30,238,29,238,28,238,27,255,31,255,30,248,31,248,31,92,31,63,31,125,31,219,31,219,30,75,31,216,31,244,31,36,31,119,31,106,31,106,30,231,31,84,31,203,31,207,31,60,31,111,31,113,31,37,31,237,31,237,30,237,29,45,31,148,31,5,31,182,31,14,31,210,31,224,31,233,31,233,30,233,29,201,31,38,31,148,31,153,31,43,31,63,31,94,31,223,31,13,31,248,31,198,31,43,31,200,31,109,31,109,30,227,31,190,31,175,31,25,31,25,30,17,31,152,31,64,31,64,30,156,31,241,31,163,31,49,31,173,31,136,31,128,31,128,30,128,29,24,31,222,31,222,30,222,29,212,31,212,30,212,29,36,31,133,31,194,31,197,31,173,31,179,31,3,31,122,31,62,31,62,30,167,31,215,31,95,31,96,31,69,31,69,30,143,31,142,31,173,31,110,31,80,31,96,31,203,31,236,31,116,31,116,30,111,31,105,31,85,31,169,31,228,31,127,31,104,31,104,30,104,29,114,31,181,31,181,30,181,29,49,31,222,31,12,31,12,30,110,31,125,31,125,30,172,31,172,30,2,31,2,30,123,31,123,30,53,31,215,31,9,31,224,31,84,31,153,31,58,31,57,31,57,30,184,31,176,31,134,31,39,31,58,31,58,30,204,31,119,31,223,31,130,31,248,31,4,31,128,31,64,31,71,31,161,31,38,31,113,31,174,31,65,31,65,30,59,31,59,30,145,31,19,31,19,30,19,29,217,31,203,31,174,31,3,31,154,31,127,31,92,31,238,31,70,31,70,30,177,31,203,31,19,31,19,30,19,29,70,31,70,30,70,29,149,31,100,31,100,30,249,31,249,30,237,31,135,31,209,31,1,31,189,31,189,30,186,31,119,31,177,31,46,31,56,31,90,31,254,31,102,31,24,31,4,31,67,31,242,31,202,31,179,31,115,31,126,31,64,31,229,31,229,30,141,31,156,31,79,31,79,30,114,31,153,31,209,31,244,31,2,31,202,31,18,31,18,30,101,31,101,30,92,31,92,30,92,29,215,31,225,31,140,31,140,30,195,31,120,31,204,31,17,31,61,31,61,30,61,29,82,31,82,30,221,31,231,31,108,31,204,31,162,31,163,31,53,31,114,31,202,31,99,31,54,31,253,31,192,31,63,31,63,30,133,31,217,31,35,31,130,31,130,30,237,31,193,31,160,31,160,30,160,29,178,31,191,31,121,31,121,30,190,31,39,31,162,31,157,31,36,31,220,31,220,30,104,31,207,31,61,31,114,31,114,30,40,31,40,30,55,31,36,31,205,31,224,31,200,31,127,31,85,31,237,31,191,31,191,30,21,31,200,31,216,31,245,31,96,31,29,31,133,31,133,30,213,31,46,31,41,31,217,31,217,30,65,31,59,31,232,31,232,30,157,31,63,31,187,31,170,31,34,31,92,31,52,31,171,31,203,31,7,31,194,31,30,31,73,31,186,31,177,31,226,31,91,31,91,30,91,29,91,28,41,31,41,30,7,31,255,31,255,30,223,31,27,31,27,30,237,31,158,31,59,31,88,31,64,31,119,31,184,31,184,30,104,31,104,30,3,31,83,31,13,31,13,30,177,31,9,31,71,31,170,31,170,30,162,31,130,31,9,31,146,31,146,30,220,31,235,31,139,31,189,31,53,31,124,31,101,31,107,31,15,31,69,31,183,31,122,31,14,31,129,31,62,31,195,31,141,31,57,31,167,31,100,31,141,31,38,31,200,31,249,31,86,31,86,30,3,31,240,31,49,31,97,31,155,31,155,30,111,31,214,31,214,30,74,31,244,31,16,31,26,31,186,31,127,31,193,31,157,31,69,31,218,31,85,31,216,31,80,31,161,31,159,31,255,31,253,31,69,31,236,31,236,30,225,31,28,31,7,31,164,31,155,31,155,30,92,31,147,31,147,30,61,31,61,30,247,31,208,31,147,31,237,31,69,31,84,31,84,30,120,31,170,31,218,31,27,31,54,31,135,31,135,30,75,31,75,30,207,31,143,31,77,31,54,31,216,31,39,31,39,30,55,31,43,31,43,30,43,29,192,31,237,31,62,31,232,31,93,31,6,31,181,31,181,30,202,31,202,30,34,31,75,31,75,30,75,29,75,28,243,31,33,31,213,31,213,30,121,31,121,30,121,29,53,31,110,31,186,31,107,31,107,30,249,31,221,31,49,31,75,31,75,30,105,31,105,30,107,31,166,31,191,31,207,31,28,31,28,30,217,31,194,31,194,30,25,31,156,31,74,31,125,31,248,31,36,31,251,31,55,31,229,31,15,31,215,31,15,31,244,31,142,31,142,30,156,31,122,31,119,31,222,31,71,31,8,31,207,31,207,30,121,31,121,30,42,31,49,31,113,31,95,31,224,31,137,31,200,31,200,30,62,31,210,31,97,31,97,30,132,31,41,31,41,30,167,31,167,30,68,31,169,31,2,31,126,31,126,30,126,29,169,31,38,31,38,30,70,31,127,31,72,31,94,31,102,31,185,31,185,30,129,31,129,30,69,31,249,31,247,31,116,31,229,31,228,31,221,31,44,31,44,30,36,31,114,31,34,31,53,31,235,31,24,31,150,31,31,31,119,31,143,31,146,31,239,31,239,30,36,31,101,31,75,31,118,31,48,31,21,31,99,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
