-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 461;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,104,0,113,0,0,0,252,0,215,0,0,0,103,0,216,0,27,0,228,0,91,0,0,0,210,0,111,0,138,0,110,0,202,0,76,0,0,0,164,0,171,0,137,0,68,0,186,0,113,0,130,0,199,0,0,0,187,0,101,0,195,0,84,0,173,0,47,0,0,0,146,0,150,0,219,0,18,0,1,0,130,0,125,0,2,0,67,0,227,0,0,0,197,0,34,0,101,0,15,0,207,0,142,0,0,0,85,0,225,0,0,0,0,0,34,0,0,0,0,0,14,0,74,0,213,0,123,0,0,0,6,0,56,0,150,0,0,0,49,0,153,0,155,0,0,0,238,0,0,0,0,0,0,0,13,0,159,0,138,0,239,0,150,0,0,0,222,0,204,0,11,0,0,0,0,0,41,0,155,0,201,0,240,0,152,0,152,0,0,0,216,0,227,0,0,0,94,0,49,0,155,0,0,0,0,0,34,0,237,0,146,0,38,0,102,0,240,0,0,0,1,0,147,0,209,0,95,0,79,0,229,0,216,0,137,0,245,0,112,0,225,0,143,0,218,0,4,0,0,0,134,0,0,0,241,0,0,0,157,0,66,0,198,0,53,0,0,0,0,0,204,0,212,0,180,0,219,0,0,0,0,0,26,0,98,0,54,0,131,0,82,0,0,0,4,0,153,0,0,0,95,0,38,0,228,0,159,0,0,0,97,0,4,0,129,0,0,0,30,0,6,0,171,0,41,0,117,0,0,0,10,0,165,0,189,0,25,0,220,0,128,0,186,0,51,0,108,0,0,0,141,0,162,0,208,0,154,0,16,0,164,0,83,0,155,0,126,0,248,0,0,0,142,0,0,0,237,0,241,0,159,0,58,0,177,0,206,0,98,0,127,0,0,0,214,0,13,0,89,0,104,0,0,0,190,0,40,0,217,0,58,0,113,0,0,0,0,0,0,0,0,0,199,0,159,0,61,0,252,0,204,0,177,0,221,0,207,0,167,0,0,0,200,0,170,0,0,0,111,0,99,0,132,0,23,0,6,0,219,0,0,0,15,0,35,0,136,0,156,0,12,0,206,0,245,0,0,0,0,0,212,0,58,0,0,0,165,0,173,0,184,0,52,0,0,0,0,0,82,0,34,0,0,0,60,0,0,0,45,0,6,0,78,0,11,0,111,0,0,0,0,0,0,0,0,0,103,0,158,0,13,0,32,0,69,0,0,0,67,0,90,0,78,0,232,0,135,0,203,0,69,0,0,0,168,0,88,0,116,0,20,0,183,0,239,0,204,0,0,0,163,0,0,0,0,0,147,0,171,0,0,0,0,0,109,0,0,0,124,0,242,0,33,0,203,0,89,0,187,0,97,0,179,0,0,0,235,0,191,0,121,0,241,0,249,0,166,0,0,0,0,0,53,0,0,0,0,0,0,0,254,0,73,0,0,0,68,0,0,0,0,0,197,0,196,0,0,0,219,0,206,0,19,0,184,0,153,0,20,0,0,0,0,0,0,0,9,0,19,0,132,0,0,0,224,0,96,0,118,0,181,0,117,0,199,0,112,0,88,0,117,0,0,0,50,0,0,0,85,0,124,0,23,0,193,0,22,0,24,0,0,0,35,0,33,0,204,0,220,0,42,0,223,0,97,0,107,0,78,0,168,0,21,0,16,0,8,0,112,0,49,0,0,0,37,0,35,0,185,0,227,0,226,0,6,0,163,0,0,0,117,0,107,0,85,0,199,0,87,0,0,0,37,0,64,0,19,0,188,0,85,0,175,0,139,0,168,0,100,0,0,0,202,0,204,0,48,0,149,0,193,0,253,0,0,0,107,0,0,0,149,0,154,0,0,0,0,0,30,0,104,0,96,0,0,0,58,0,0,0,8,0,43,0,0,0,212,0,221,0,0,0,66,0,87,0,187,0,204,0,144,0,200,0,99,0,177,0,0,0,123,0,191,0,15,0,149,0,93,0,55,0,202,0,43,0,122,0,199,0,111,0,235,0,6,0,175,0,255,0,19,0,202,0,229,0,80,0,29,0,181,0,152,0,216,0,46,0,199,0,7,0,254,0,0,0,136,0,0,0);
signal scenario_full  : scenario_type := (0,0,104,31,113,31,113,30,252,31,215,31,215,30,103,31,216,31,27,31,228,31,91,31,91,30,210,31,111,31,138,31,110,31,202,31,76,31,76,30,164,31,171,31,137,31,68,31,186,31,113,31,130,31,199,31,199,30,187,31,101,31,195,31,84,31,173,31,47,31,47,30,146,31,150,31,219,31,18,31,1,31,130,31,125,31,2,31,67,31,227,31,227,30,197,31,34,31,101,31,15,31,207,31,142,31,142,30,85,31,225,31,225,30,225,29,34,31,34,30,34,29,14,31,74,31,213,31,123,31,123,30,6,31,56,31,150,31,150,30,49,31,153,31,155,31,155,30,238,31,238,30,238,29,238,28,13,31,159,31,138,31,239,31,150,31,150,30,222,31,204,31,11,31,11,30,11,29,41,31,155,31,201,31,240,31,152,31,152,31,152,30,216,31,227,31,227,30,94,31,49,31,155,31,155,30,155,29,34,31,237,31,146,31,38,31,102,31,240,31,240,30,1,31,147,31,209,31,95,31,79,31,229,31,216,31,137,31,245,31,112,31,225,31,143,31,218,31,4,31,4,30,134,31,134,30,241,31,241,30,157,31,66,31,198,31,53,31,53,30,53,29,204,31,212,31,180,31,219,31,219,30,219,29,26,31,98,31,54,31,131,31,82,31,82,30,4,31,153,31,153,30,95,31,38,31,228,31,159,31,159,30,97,31,4,31,129,31,129,30,30,31,6,31,171,31,41,31,117,31,117,30,10,31,165,31,189,31,25,31,220,31,128,31,186,31,51,31,108,31,108,30,141,31,162,31,208,31,154,31,16,31,164,31,83,31,155,31,126,31,248,31,248,30,142,31,142,30,237,31,241,31,159,31,58,31,177,31,206,31,98,31,127,31,127,30,214,31,13,31,89,31,104,31,104,30,190,31,40,31,217,31,58,31,113,31,113,30,113,29,113,28,113,27,199,31,159,31,61,31,252,31,204,31,177,31,221,31,207,31,167,31,167,30,200,31,170,31,170,30,111,31,99,31,132,31,23,31,6,31,219,31,219,30,15,31,35,31,136,31,156,31,12,31,206,31,245,31,245,30,245,29,212,31,58,31,58,30,165,31,173,31,184,31,52,31,52,30,52,29,82,31,34,31,34,30,60,31,60,30,45,31,6,31,78,31,11,31,111,31,111,30,111,29,111,28,111,27,103,31,158,31,13,31,32,31,69,31,69,30,67,31,90,31,78,31,232,31,135,31,203,31,69,31,69,30,168,31,88,31,116,31,20,31,183,31,239,31,204,31,204,30,163,31,163,30,163,29,147,31,171,31,171,30,171,29,109,31,109,30,124,31,242,31,33,31,203,31,89,31,187,31,97,31,179,31,179,30,235,31,191,31,121,31,241,31,249,31,166,31,166,30,166,29,53,31,53,30,53,29,53,28,254,31,73,31,73,30,68,31,68,30,68,29,197,31,196,31,196,30,219,31,206,31,19,31,184,31,153,31,20,31,20,30,20,29,20,28,9,31,19,31,132,31,132,30,224,31,96,31,118,31,181,31,117,31,199,31,112,31,88,31,117,31,117,30,50,31,50,30,85,31,124,31,23,31,193,31,22,31,24,31,24,30,35,31,33,31,204,31,220,31,42,31,223,31,97,31,107,31,78,31,168,31,21,31,16,31,8,31,112,31,49,31,49,30,37,31,35,31,185,31,227,31,226,31,6,31,163,31,163,30,117,31,107,31,85,31,199,31,87,31,87,30,37,31,64,31,19,31,188,31,85,31,175,31,139,31,168,31,100,31,100,30,202,31,204,31,48,31,149,31,193,31,253,31,253,30,107,31,107,30,149,31,154,31,154,30,154,29,30,31,104,31,96,31,96,30,58,31,58,30,8,31,43,31,43,30,212,31,221,31,221,30,66,31,87,31,187,31,204,31,144,31,200,31,99,31,177,31,177,30,123,31,191,31,15,31,149,31,93,31,55,31,202,31,43,31,122,31,199,31,111,31,235,31,6,31,175,31,255,31,19,31,202,31,229,31,80,31,29,31,181,31,152,31,216,31,46,31,199,31,7,31,254,31,254,30,136,31,136,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
