-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_602 is
end project_tb_602;

architecture project_tb_arch_602 of project_tb_602 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 300;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (206,0,0,0,0,0,0,0,181,0,144,0,178,0,114,0,42,0,0,0,94,0,0,0,0,0,0,0,240,0,0,0,226,0,144,0,138,0,52,0,0,0,158,0,179,0,163,0,27,0,238,0,68,0,198,0,75,0,0,0,71,0,95,0,161,0,31,0,160,0,142,0,22,0,252,0,63,0,163,0,120,0,0,0,74,0,213,0,0,0,171,0,22,0,229,0,50,0,122,0,33,0,111,0,218,0,31,0,75,0,152,0,50,0,124,0,59,0,141,0,49,0,243,0,204,0,87,0,177,0,215,0,2,0,137,0,52,0,210,0,0,0,104,0,236,0,109,0,248,0,229,0,0,0,210,0,0,0,105,0,101,0,166,0,228,0,0,0,0,0,111,0,0,0,240,0,121,0,156,0,49,0,126,0,43,0,0,0,67,0,211,0,232,0,229,0,86,0,46,0,172,0,42,0,94,0,20,0,0,0,25,0,0,0,247,0,90,0,172,0,0,0,173,0,221,0,56,0,239,0,0,0,43,0,73,0,11,0,160,0,20,0,145,0,132,0,60,0,171,0,28,0,244,0,92,0,54,0,0,0,156,0,12,0,89,0,100,0,87,0,215,0,177,0,225,0,60,0,10,0,67,0,0,0,244,0,217,0,212,0,187,0,0,0,231,0,58,0,0,0,0,0,0,0,0,0,0,0,240,0,213,0,92,0,189,0,50,0,0,0,87,0,40,0,74,0,137,0,0,0,114,0,222,0,54,0,0,0,0,0,194,0,0,0,0,0,158,0,97,0,193,0,1,0,241,0,246,0,161,0,153,0,203,0,0,0,113,0,109,0,216,0,150,0,75,0,0,0,161,0,48,0,72,0,251,0,140,0,88,0,47,0,135,0,215,0,224,0,185,0,0,0,167,0,0,0,210,0,182,0,152,0,156,0,214,0,0,0,120,0,147,0,0,0,0,0,131,0,182,0,102,0,36,0,174,0,1,0,166,0,118,0,88,0,76,0,0,0,165,0,236,0,36,0,0,0,55,0,67,0,0,0,145,0,224,0,0,0,221,0,237,0,179,0,12,0,0,0,144,0,83,0,228,0,0,0,48,0,53,0,0,0,50,0,19,0,0,0,166,0,100,0,93,0,42,0,233,0,122,0,77,0,72,0,147,0,144,0,0,0,185,0,208,0,42,0,76,0,141,0,91,0,0,0,32,0,14,0,36,0,235,0,0,0,250,0,219,0,250,0,198,0,0,0,0,0,116,0,47,0,123,0,4,0,0,0,192,0,28,0,0,0,191,0,0,0,24,0,135,0,136,0,167,0,97,0,185,0,98,0,217,0,158,0,0,0,145,0,212,0);
signal scenario_full  : scenario_type := (206,31,206,30,206,29,206,28,181,31,144,31,178,31,114,31,42,31,42,30,94,31,94,30,94,29,94,28,240,31,240,30,226,31,144,31,138,31,52,31,52,30,158,31,179,31,163,31,27,31,238,31,68,31,198,31,75,31,75,30,71,31,95,31,161,31,31,31,160,31,142,31,22,31,252,31,63,31,163,31,120,31,120,30,74,31,213,31,213,30,171,31,22,31,229,31,50,31,122,31,33,31,111,31,218,31,31,31,75,31,152,31,50,31,124,31,59,31,141,31,49,31,243,31,204,31,87,31,177,31,215,31,2,31,137,31,52,31,210,31,210,30,104,31,236,31,109,31,248,31,229,31,229,30,210,31,210,30,105,31,101,31,166,31,228,31,228,30,228,29,111,31,111,30,240,31,121,31,156,31,49,31,126,31,43,31,43,30,67,31,211,31,232,31,229,31,86,31,46,31,172,31,42,31,94,31,20,31,20,30,25,31,25,30,247,31,90,31,172,31,172,30,173,31,221,31,56,31,239,31,239,30,43,31,73,31,11,31,160,31,20,31,145,31,132,31,60,31,171,31,28,31,244,31,92,31,54,31,54,30,156,31,12,31,89,31,100,31,87,31,215,31,177,31,225,31,60,31,10,31,67,31,67,30,244,31,217,31,212,31,187,31,187,30,231,31,58,31,58,30,58,29,58,28,58,27,58,26,240,31,213,31,92,31,189,31,50,31,50,30,87,31,40,31,74,31,137,31,137,30,114,31,222,31,54,31,54,30,54,29,194,31,194,30,194,29,158,31,97,31,193,31,1,31,241,31,246,31,161,31,153,31,203,31,203,30,113,31,109,31,216,31,150,31,75,31,75,30,161,31,48,31,72,31,251,31,140,31,88,31,47,31,135,31,215,31,224,31,185,31,185,30,167,31,167,30,210,31,182,31,152,31,156,31,214,31,214,30,120,31,147,31,147,30,147,29,131,31,182,31,102,31,36,31,174,31,1,31,166,31,118,31,88,31,76,31,76,30,165,31,236,31,36,31,36,30,55,31,67,31,67,30,145,31,224,31,224,30,221,31,237,31,179,31,12,31,12,30,144,31,83,31,228,31,228,30,48,31,53,31,53,30,50,31,19,31,19,30,166,31,100,31,93,31,42,31,233,31,122,31,77,31,72,31,147,31,144,31,144,30,185,31,208,31,42,31,76,31,141,31,91,31,91,30,32,31,14,31,36,31,235,31,235,30,250,31,219,31,250,31,198,31,198,30,198,29,116,31,47,31,123,31,4,31,4,30,192,31,28,31,28,30,191,31,191,30,24,31,135,31,136,31,167,31,97,31,185,31,98,31,217,31,158,31,158,30,145,31,212,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
