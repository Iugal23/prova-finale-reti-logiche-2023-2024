-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_48 is
end project_tb_48;

architecture project_tb_arch_48 of project_tb_48 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 299;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,180,0,67,0,40,0,164,0,230,0,47,0,171,0,187,0,204,0,79,0,3,0,241,0,58,0,178,0,40,0,165,0,0,0,111,0,248,0,189,0,52,0,14,0,189,0,205,0,235,0,82,0,187,0,0,0,72,0,98,0,0,0,214,0,127,0,102,0,133,0,0,0,0,0,189,0,90,0,43,0,19,0,58,0,157,0,224,0,179,0,163,0,0,0,6,0,0,0,52,0,219,0,0,0,65,0,62,0,212,0,59,0,176,0,20,0,68,0,157,0,70,0,3,0,111,0,103,0,189,0,180,0,0,0,237,0,0,0,0,0,192,0,5,0,0,0,190,0,239,0,42,0,0,0,155,0,92,0,65,0,132,0,39,0,143,0,226,0,66,0,8,0,244,0,24,0,69,0,18,0,0,0,127,0,0,0,77,0,14,0,0,0,187,0,114,0,0,0,50,0,180,0,226,0,48,0,97,0,39,0,0,0,0,0,248,0,0,0,0,0,106,0,21,0,134,0,137,0,230,0,209,0,0,0,247,0,71,0,232,0,212,0,95,0,0,0,0,0,27,0,71,0,0,0,74,0,202,0,0,0,54,0,21,0,141,0,50,0,214,0,220,0,195,0,63,0,77,0,240,0,73,0,0,0,0,0,172,0,211,0,89,0,66,0,232,0,0,0,225,0,24,0,237,0,80,0,0,0,124,0,100,0,35,0,235,0,139,0,0,0,0,0,56,0,135,0,15,0,120,0,0,0,247,0,148,0,219,0,243,0,133,0,63,0,173,0,169,0,191,0,69,0,0,0,0,0,190,0,184,0,158,0,208,0,218,0,210,0,22,0,186,0,45,0,249,0,40,0,0,0,25,0,179,0,224,0,41,0,75,0,0,0,59,0,176,0,76,0,204,0,100,0,26,0,216,0,129,0,0,0,33,0,82,0,0,0,193,0,237,0,0,0,96,0,244,0,164,0,152,0,142,0,174,0,5,0,0,0,182,0,160,0,71,0,123,0,242,0,203,0,255,0,71,0,172,0,0,0,0,0,149,0,91,0,146,0,213,0,125,0,156,0,0,0,63,0,202,0,91,0,113,0,0,0,0,0,166,0,186,0,0,0,142,0,157,0,40,0,252,0,217,0,33,0,219,0,0,0,135,0,192,0,144,0,0,0,205,0,0,0,63,0,0,0,0,0,152,0,129,0,162,0,95,0,203,0,0,0,0,0,91,0,134,0,8,0,0,0,0,0,67,0,229,0,119,0,134,0,209,0,251,0,140,0,88,0,0,0,152,0,160,0,189,0,162,0,133,0,0,0,108,0,141,0,3,0,83,0,153,0,88,0,0,0,203,0);
signal scenario_full  : scenario_type := (35,31,180,31,67,31,40,31,164,31,230,31,47,31,171,31,187,31,204,31,79,31,3,31,241,31,58,31,178,31,40,31,165,31,165,30,111,31,248,31,189,31,52,31,14,31,189,31,205,31,235,31,82,31,187,31,187,30,72,31,98,31,98,30,214,31,127,31,102,31,133,31,133,30,133,29,189,31,90,31,43,31,19,31,58,31,157,31,224,31,179,31,163,31,163,30,6,31,6,30,52,31,219,31,219,30,65,31,62,31,212,31,59,31,176,31,20,31,68,31,157,31,70,31,3,31,111,31,103,31,189,31,180,31,180,30,237,31,237,30,237,29,192,31,5,31,5,30,190,31,239,31,42,31,42,30,155,31,92,31,65,31,132,31,39,31,143,31,226,31,66,31,8,31,244,31,24,31,69,31,18,31,18,30,127,31,127,30,77,31,14,31,14,30,187,31,114,31,114,30,50,31,180,31,226,31,48,31,97,31,39,31,39,30,39,29,248,31,248,30,248,29,106,31,21,31,134,31,137,31,230,31,209,31,209,30,247,31,71,31,232,31,212,31,95,31,95,30,95,29,27,31,71,31,71,30,74,31,202,31,202,30,54,31,21,31,141,31,50,31,214,31,220,31,195,31,63,31,77,31,240,31,73,31,73,30,73,29,172,31,211,31,89,31,66,31,232,31,232,30,225,31,24,31,237,31,80,31,80,30,124,31,100,31,35,31,235,31,139,31,139,30,139,29,56,31,135,31,15,31,120,31,120,30,247,31,148,31,219,31,243,31,133,31,63,31,173,31,169,31,191,31,69,31,69,30,69,29,190,31,184,31,158,31,208,31,218,31,210,31,22,31,186,31,45,31,249,31,40,31,40,30,25,31,179,31,224,31,41,31,75,31,75,30,59,31,176,31,76,31,204,31,100,31,26,31,216,31,129,31,129,30,33,31,82,31,82,30,193,31,237,31,237,30,96,31,244,31,164,31,152,31,142,31,174,31,5,31,5,30,182,31,160,31,71,31,123,31,242,31,203,31,255,31,71,31,172,31,172,30,172,29,149,31,91,31,146,31,213,31,125,31,156,31,156,30,63,31,202,31,91,31,113,31,113,30,113,29,166,31,186,31,186,30,142,31,157,31,40,31,252,31,217,31,33,31,219,31,219,30,135,31,192,31,144,31,144,30,205,31,205,30,63,31,63,30,63,29,152,31,129,31,162,31,95,31,203,31,203,30,203,29,91,31,134,31,8,31,8,30,8,29,67,31,229,31,119,31,134,31,209,31,251,31,140,31,88,31,88,30,152,31,160,31,189,31,162,31,133,31,133,30,108,31,141,31,3,31,83,31,153,31,88,31,88,30,203,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
