-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_149 is
end project_tb_149;

architecture project_tb_arch_149 of project_tb_149 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 685;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (196,0,5,0,22,0,236,0,8,0,101,0,140,0,249,0,133,0,53,0,0,0,101,0,164,0,233,0,128,0,80,0,33,0,213,0,6,0,0,0,179,0,55,0,128,0,228,0,240,0,101,0,67,0,163,0,107,0,0,0,78,0,0,0,222,0,130,0,180,0,182,0,0,0,243,0,0,0,0,0,193,0,166,0,11,0,204,0,19,0,190,0,117,0,5,0,49,0,151,0,73,0,0,0,166,0,232,0,123,0,209,0,0,0,246,0,119,0,207,0,50,0,221,0,46,0,181,0,123,0,0,0,255,0,146,0,143,0,0,0,6,0,151,0,70,0,26,0,223,0,185,0,193,0,163,0,228,0,0,0,141,0,0,0,240,0,241,0,0,0,150,0,0,0,36,0,11,0,0,0,0,0,162,0,211,0,253,0,63,0,0,0,113,0,83,0,0,0,154,0,235,0,0,0,154,0,48,0,56,0,159,0,0,0,237,0,21,0,177,0,187,0,0,0,22,0,138,0,158,0,4,0,73,0,246,0,162,0,18,0,0,0,101,0,73,0,121,0,0,0,0,0,150,0,246,0,209,0,119,0,52,0,221,0,20,0,229,0,0,0,247,0,31,0,113,0,0,0,132,0,212,0,41,0,253,0,120,0,34,0,0,0,196,0,44,0,213,0,55,0,60,0,214,0,115,0,181,0,242,0,233,0,180,0,0,0,0,0,97,0,0,0,170,0,28,0,216,0,143,0,0,0,55,0,68,0,0,0,205,0,0,0,253,0,221,0,44,0,39,0,136,0,153,0,176,0,180,0,105,0,79,0,143,0,0,0,139,0,0,0,176,0,23,0,132,0,172,0,70,0,0,0,236,0,103,0,222,0,2,0,251,0,230,0,185,0,68,0,0,0,0,0,0,0,209,0,0,0,0,0,45,0,0,0,225,0,35,0,81,0,21,0,246,0,161,0,26,0,48,0,18,0,109,0,0,0,69,0,172,0,204,0,228,0,61,0,212,0,41,0,254,0,20,0,0,0,116,0,118,0,61,0,154,0,96,0,119,0,0,0,0,0,131,0,192,0,87,0,101,0,0,0,12,0,0,0,167,0,0,0,149,0,0,0,75,0,192,0,149,0,16,0,90,0,0,0,168,0,50,0,0,0,81,0,0,0,141,0,220,0,0,0,2,0,206,0,223,0,131,0,0,0,250,0,9,0,87,0,229,0,24,0,125,0,145,0,27,0,53,0,226,0,67,0,164,0,205,0,145,0,241,0,244,0,0,0,127,0,172,0,186,0,101,0,132,0,68,0,220,0,183,0,126,0,254,0,235,0,103,0,51,0,252,0,0,0,205,0,211,0,31,0,0,0,73,0,255,0,194,0,163,0,85,0,210,0,0,0,166,0,58,0,23,0,64,0,77,0,135,0,24,0,225,0,208,0,254,0,121,0,0,0,143,0,248,0,0,0,186,0,165,0,131,0,26,0,136,0,0,0,28,0,225,0,199,0,73,0,43,0,0,0,207,0,102,0,171,0,138,0,10,0,105,0,64,0,179,0,98,0,94,0,0,0,0,0,236,0,53,0,0,0,219,0,231,0,0,0,26,0,241,0,61,0,0,0,73,0,55,0,104,0,217,0,100,0,0,0,216,0,32,0,15,0,175,0,165,0,207,0,178,0,153,0,0,0,82,0,13,0,9,0,199,0,165,0,56,0,110,0,237,0,251,0,114,0,67,0,157,0,11,0,184,0,4,0,55,0,255,0,128,0,83,0,96,0,234,0,109,0,31,0,56,0,0,0,136,0,91,0,116,0,0,0,87,0,48,0,132,0,217,0,240,0,145,0,0,0,0,0,86,0,146,0,1,0,0,0,5,0,0,0,73,0,74,0,23,0,0,0,0,0,236,0,135,0,179,0,192,0,223,0,0,0,182,0,0,0,217,0,0,0,13,0,174,0,44,0,106,0,219,0,224,0,0,0,0,0,96,0,0,0,171,0,42,0,170,0,72,0,27,0,31,0,27,0,161,0,225,0,19,0,108,0,206,0,144,0,86,0,0,0,0,0,0,0,132,0,11,0,216,0,0,0,42,0,0,0,113,0,20,0,115,0,0,0,0,0,190,0,137,0,0,0,144,0,0,0,136,0,1,0,81,0,50,0,239,0,249,0,10,0,211,0,96,0,249,0,15,0,0,0,248,0,12,0,0,0,120,0,87,0,59,0,150,0,106,0,134,0,16,0,93,0,190,0,197,0,193,0,0,0,120,0,247,0,0,0,0,0,94,0,78,0,38,0,252,0,115,0,0,0,0,0,0,0,145,0,191,0,227,0,43,0,15,0,134,0,0,0,168,0,0,0,47,0,73,0,31,0,174,0,0,0,159,0,215,0,161,0,135,0,152,0,192,0,243,0,0,0,0,0,142,0,82,0,0,0,70,0,207,0,63,0,104,0,148,0,77,0,55,0,197,0,0,0,0,0,180,0,206,0,69,0,147,0,11,0,132,0,175,0,144,0,14,0,201,0,0,0,245,0,232,0,74,0,38,0,19,0,0,0,21,0,123,0,10,0,0,0,0,0,175,0,52,0,35,0,231,0,135,0,46,0,252,0,165,0,195,0,59,0,0,0,101,0,0,0,40,0,236,0,88,0,181,0,132,0,0,0,0,0,116,0,143,0,0,0,232,0,0,0,0,0,200,0,236,0,212,0,0,0,36,0,172,0,0,0,0,0,41,0,0,0,150,0,19,0,83,0,0,0,185,0,12,0,134,0,20,0,70,0,20,0,28,0,0,0,187,0,72,0,124,0,159,0,0,0,87,0,214,0,66,0,79,0,169,0,221,0,186,0,221,0,203,0,201,0,152,0,104,0,54,0,158,0,147,0,54,0,221,0,65,0,92,0,200,0,102,0,226,0,178,0,0,0,167,0,0,0,255,0,176,0,16,0,122,0,237,0,48,0,42,0,84,0,124,0,92,0,43,0,165,0,155,0,41,0,190,0,245,0,0,0,0,0,204,0,165,0,122,0,79,0,21,0,119,0,205,0,0,0,183,0,129,0,0,0,239,0,12,0,103,0,67,0,0,0,30,0);
signal scenario_full  : scenario_type := (196,31,5,31,22,31,236,31,8,31,101,31,140,31,249,31,133,31,53,31,53,30,101,31,164,31,233,31,128,31,80,31,33,31,213,31,6,31,6,30,179,31,55,31,128,31,228,31,240,31,101,31,67,31,163,31,107,31,107,30,78,31,78,30,222,31,130,31,180,31,182,31,182,30,243,31,243,30,243,29,193,31,166,31,11,31,204,31,19,31,190,31,117,31,5,31,49,31,151,31,73,31,73,30,166,31,232,31,123,31,209,31,209,30,246,31,119,31,207,31,50,31,221,31,46,31,181,31,123,31,123,30,255,31,146,31,143,31,143,30,6,31,151,31,70,31,26,31,223,31,185,31,193,31,163,31,228,31,228,30,141,31,141,30,240,31,241,31,241,30,150,31,150,30,36,31,11,31,11,30,11,29,162,31,211,31,253,31,63,31,63,30,113,31,83,31,83,30,154,31,235,31,235,30,154,31,48,31,56,31,159,31,159,30,237,31,21,31,177,31,187,31,187,30,22,31,138,31,158,31,4,31,73,31,246,31,162,31,18,31,18,30,101,31,73,31,121,31,121,30,121,29,150,31,246,31,209,31,119,31,52,31,221,31,20,31,229,31,229,30,247,31,31,31,113,31,113,30,132,31,212,31,41,31,253,31,120,31,34,31,34,30,196,31,44,31,213,31,55,31,60,31,214,31,115,31,181,31,242,31,233,31,180,31,180,30,180,29,97,31,97,30,170,31,28,31,216,31,143,31,143,30,55,31,68,31,68,30,205,31,205,30,253,31,221,31,44,31,39,31,136,31,153,31,176,31,180,31,105,31,79,31,143,31,143,30,139,31,139,30,176,31,23,31,132,31,172,31,70,31,70,30,236,31,103,31,222,31,2,31,251,31,230,31,185,31,68,31,68,30,68,29,68,28,209,31,209,30,209,29,45,31,45,30,225,31,35,31,81,31,21,31,246,31,161,31,26,31,48,31,18,31,109,31,109,30,69,31,172,31,204,31,228,31,61,31,212,31,41,31,254,31,20,31,20,30,116,31,118,31,61,31,154,31,96,31,119,31,119,30,119,29,131,31,192,31,87,31,101,31,101,30,12,31,12,30,167,31,167,30,149,31,149,30,75,31,192,31,149,31,16,31,90,31,90,30,168,31,50,31,50,30,81,31,81,30,141,31,220,31,220,30,2,31,206,31,223,31,131,31,131,30,250,31,9,31,87,31,229,31,24,31,125,31,145,31,27,31,53,31,226,31,67,31,164,31,205,31,145,31,241,31,244,31,244,30,127,31,172,31,186,31,101,31,132,31,68,31,220,31,183,31,126,31,254,31,235,31,103,31,51,31,252,31,252,30,205,31,211,31,31,31,31,30,73,31,255,31,194,31,163,31,85,31,210,31,210,30,166,31,58,31,23,31,64,31,77,31,135,31,24,31,225,31,208,31,254,31,121,31,121,30,143,31,248,31,248,30,186,31,165,31,131,31,26,31,136,31,136,30,28,31,225,31,199,31,73,31,43,31,43,30,207,31,102,31,171,31,138,31,10,31,105,31,64,31,179,31,98,31,94,31,94,30,94,29,236,31,53,31,53,30,219,31,231,31,231,30,26,31,241,31,61,31,61,30,73,31,55,31,104,31,217,31,100,31,100,30,216,31,32,31,15,31,175,31,165,31,207,31,178,31,153,31,153,30,82,31,13,31,9,31,199,31,165,31,56,31,110,31,237,31,251,31,114,31,67,31,157,31,11,31,184,31,4,31,55,31,255,31,128,31,83,31,96,31,234,31,109,31,31,31,56,31,56,30,136,31,91,31,116,31,116,30,87,31,48,31,132,31,217,31,240,31,145,31,145,30,145,29,86,31,146,31,1,31,1,30,5,31,5,30,73,31,74,31,23,31,23,30,23,29,236,31,135,31,179,31,192,31,223,31,223,30,182,31,182,30,217,31,217,30,13,31,174,31,44,31,106,31,219,31,224,31,224,30,224,29,96,31,96,30,171,31,42,31,170,31,72,31,27,31,31,31,27,31,161,31,225,31,19,31,108,31,206,31,144,31,86,31,86,30,86,29,86,28,132,31,11,31,216,31,216,30,42,31,42,30,113,31,20,31,115,31,115,30,115,29,190,31,137,31,137,30,144,31,144,30,136,31,1,31,81,31,50,31,239,31,249,31,10,31,211,31,96,31,249,31,15,31,15,30,248,31,12,31,12,30,120,31,87,31,59,31,150,31,106,31,134,31,16,31,93,31,190,31,197,31,193,31,193,30,120,31,247,31,247,30,247,29,94,31,78,31,38,31,252,31,115,31,115,30,115,29,115,28,145,31,191,31,227,31,43,31,15,31,134,31,134,30,168,31,168,30,47,31,73,31,31,31,174,31,174,30,159,31,215,31,161,31,135,31,152,31,192,31,243,31,243,30,243,29,142,31,82,31,82,30,70,31,207,31,63,31,104,31,148,31,77,31,55,31,197,31,197,30,197,29,180,31,206,31,69,31,147,31,11,31,132,31,175,31,144,31,14,31,201,31,201,30,245,31,232,31,74,31,38,31,19,31,19,30,21,31,123,31,10,31,10,30,10,29,175,31,52,31,35,31,231,31,135,31,46,31,252,31,165,31,195,31,59,31,59,30,101,31,101,30,40,31,236,31,88,31,181,31,132,31,132,30,132,29,116,31,143,31,143,30,232,31,232,30,232,29,200,31,236,31,212,31,212,30,36,31,172,31,172,30,172,29,41,31,41,30,150,31,19,31,83,31,83,30,185,31,12,31,134,31,20,31,70,31,20,31,28,31,28,30,187,31,72,31,124,31,159,31,159,30,87,31,214,31,66,31,79,31,169,31,221,31,186,31,221,31,203,31,201,31,152,31,104,31,54,31,158,31,147,31,54,31,221,31,65,31,92,31,200,31,102,31,226,31,178,31,178,30,167,31,167,30,255,31,176,31,16,31,122,31,237,31,48,31,42,31,84,31,124,31,92,31,43,31,165,31,155,31,41,31,190,31,245,31,245,30,245,29,204,31,165,31,122,31,79,31,21,31,119,31,205,31,205,30,183,31,129,31,129,30,239,31,12,31,103,31,67,31,67,30,30,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
