-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 410;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (30,0,161,0,173,0,0,0,172,0,207,0,0,0,245,0,247,0,0,0,216,0,0,0,137,0,146,0,247,0,15,0,223,0,249,0,109,0,118,0,16,0,113,0,0,0,77,0,66,0,83,0,0,0,91,0,101,0,0,0,72,0,93,0,1,0,0,0,238,0,75,0,175,0,0,0,41,0,0,0,0,0,56,0,86,0,152,0,181,0,0,0,154,0,205,0,98,0,15,0,118,0,0,0,34,0,0,0,0,0,156,0,24,0,13,0,164,0,165,0,2,0,134,0,115,0,91,0,0,0,159,0,233,0,0,0,0,0,160,0,225,0,210,0,94,0,120,0,122,0,162,0,85,0,31,0,233,0,86,0,0,0,0,0,0,0,165,0,250,0,106,0,171,0,0,0,185,0,175,0,238,0,141,0,16,0,223,0,109,0,14,0,93,0,201,0,36,0,56,0,0,0,53,0,10,0,144,0,198,0,30,0,0,0,184,0,205,0,123,0,181,0,0,0,144,0,224,0,94,0,253,0,123,0,71,0,13,0,179,0,169,0,200,0,5,0,245,0,81,0,142,0,0,0,25,0,59,0,162,0,218,0,188,0,212,0,57,0,188,0,216,0,73,0,179,0,0,0,0,0,131,0,18,0,252,0,93,0,169,0,219,0,0,0,0,0,99,0,0,0,99,0,255,0,48,0,242,0,0,0,155,0,73,0,0,0,2,0,0,0,105,0,0,0,54,0,119,0,222,0,226,0,163,0,203,0,252,0,70,0,165,0,10,0,108,0,0,0,7,0,124,0,6,0,44,0,114,0,0,0,140,0,217,0,236,0,163,0,0,0,143,0,0,0,204,0,137,0,0,0,245,0,145,0,42,0,198,0,0,0,18,0,153,0,19,0,235,0,126,0,176,0,39,0,131,0,28,0,100,0,220,0,36,0,155,0,151,0,0,0,0,0,93,0,235,0,0,0,71,0,0,0,0,0,81,0,0,0,22,0,222,0,53,0,31,0,128,0,92,0,176,0,134,0,216,0,119,0,0,0,21,0,170,0,157,0,2,0,83,0,98,0,42,0,226,0,210,0,241,0,0,0,178,0,0,0,116,0,135,0,0,0,153,0,17,0,17,0,171,0,15,0,175,0,217,0,121,0,0,0,0,0,35,0,255,0,135,0,109,0,0,0,139,0,22,0,70,0,1,0,13,0,129,0,100,0,108,0,23,0,103,0,0,0,0,0,131,0,167,0,229,0,51,0,101,0,100,0,135,0,114,0,156,0,99,0,173,0,0,0,154,0,87,0,98,0,126,0,40,0,233,0,92,0,128,0,24,0,0,0,44,0,5,0,193,0,105,0,35,0,30,0,64,0,73,0,23,0,173,0,208,0,2,0,15,0,107,0,242,0,153,0,0,0,202,0,5,0,156,0,0,0,215,0,165,0,22,0,9,0,123,0,0,0,42,0,204,0,160,0,149,0,0,0,0,0,209,0,221,0,0,0,203,0,168,0,144,0,200,0,138,0,21,0,74,0,83,0,100,0,173,0,109,0,28,0,197,0,95,0,188,0,113,0,137,0,249,0,165,0,233,0,78,0,98,0,216,0,177,0,211,0,119,0,118,0,193,0,225,0,0,0,154,0,197,0,76,0,137,0,37,0,192,0,0,0,0,0,161,0,6,0,77,0,191,0,0,0,142,0,134,0,14,0,68,0,223,0,142,0,53,0,18,0,79,0,64,0,4,0,180,0,154,0,15,0,106,0,183,0,53,0,50,0,219,0,234,0,154,0,200,0,8,0,200,0,7,0,94,0,139,0,231,0,159,0,45,0,169,0,0,0,198,0,0,0,139,0,33,0);
signal scenario_full  : scenario_type := (30,31,161,31,173,31,173,30,172,31,207,31,207,30,245,31,247,31,247,30,216,31,216,30,137,31,146,31,247,31,15,31,223,31,249,31,109,31,118,31,16,31,113,31,113,30,77,31,66,31,83,31,83,30,91,31,101,31,101,30,72,31,93,31,1,31,1,30,238,31,75,31,175,31,175,30,41,31,41,30,41,29,56,31,86,31,152,31,181,31,181,30,154,31,205,31,98,31,15,31,118,31,118,30,34,31,34,30,34,29,156,31,24,31,13,31,164,31,165,31,2,31,134,31,115,31,91,31,91,30,159,31,233,31,233,30,233,29,160,31,225,31,210,31,94,31,120,31,122,31,162,31,85,31,31,31,233,31,86,31,86,30,86,29,86,28,165,31,250,31,106,31,171,31,171,30,185,31,175,31,238,31,141,31,16,31,223,31,109,31,14,31,93,31,201,31,36,31,56,31,56,30,53,31,10,31,144,31,198,31,30,31,30,30,184,31,205,31,123,31,181,31,181,30,144,31,224,31,94,31,253,31,123,31,71,31,13,31,179,31,169,31,200,31,5,31,245,31,81,31,142,31,142,30,25,31,59,31,162,31,218,31,188,31,212,31,57,31,188,31,216,31,73,31,179,31,179,30,179,29,131,31,18,31,252,31,93,31,169,31,219,31,219,30,219,29,99,31,99,30,99,31,255,31,48,31,242,31,242,30,155,31,73,31,73,30,2,31,2,30,105,31,105,30,54,31,119,31,222,31,226,31,163,31,203,31,252,31,70,31,165,31,10,31,108,31,108,30,7,31,124,31,6,31,44,31,114,31,114,30,140,31,217,31,236,31,163,31,163,30,143,31,143,30,204,31,137,31,137,30,245,31,145,31,42,31,198,31,198,30,18,31,153,31,19,31,235,31,126,31,176,31,39,31,131,31,28,31,100,31,220,31,36,31,155,31,151,31,151,30,151,29,93,31,235,31,235,30,71,31,71,30,71,29,81,31,81,30,22,31,222,31,53,31,31,31,128,31,92,31,176,31,134,31,216,31,119,31,119,30,21,31,170,31,157,31,2,31,83,31,98,31,42,31,226,31,210,31,241,31,241,30,178,31,178,30,116,31,135,31,135,30,153,31,17,31,17,31,171,31,15,31,175,31,217,31,121,31,121,30,121,29,35,31,255,31,135,31,109,31,109,30,139,31,22,31,70,31,1,31,13,31,129,31,100,31,108,31,23,31,103,31,103,30,103,29,131,31,167,31,229,31,51,31,101,31,100,31,135,31,114,31,156,31,99,31,173,31,173,30,154,31,87,31,98,31,126,31,40,31,233,31,92,31,128,31,24,31,24,30,44,31,5,31,193,31,105,31,35,31,30,31,64,31,73,31,23,31,173,31,208,31,2,31,15,31,107,31,242,31,153,31,153,30,202,31,5,31,156,31,156,30,215,31,165,31,22,31,9,31,123,31,123,30,42,31,204,31,160,31,149,31,149,30,149,29,209,31,221,31,221,30,203,31,168,31,144,31,200,31,138,31,21,31,74,31,83,31,100,31,173,31,109,31,28,31,197,31,95,31,188,31,113,31,137,31,249,31,165,31,233,31,78,31,98,31,216,31,177,31,211,31,119,31,118,31,193,31,225,31,225,30,154,31,197,31,76,31,137,31,37,31,192,31,192,30,192,29,161,31,6,31,77,31,191,31,191,30,142,31,134,31,14,31,68,31,223,31,142,31,53,31,18,31,79,31,64,31,4,31,180,31,154,31,15,31,106,31,183,31,53,31,50,31,219,31,234,31,154,31,200,31,8,31,200,31,7,31,94,31,139,31,231,31,159,31,45,31,169,31,169,30,198,31,198,30,139,31,33,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
