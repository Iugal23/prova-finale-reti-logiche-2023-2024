-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_624 is
end project_tb_624;

architecture project_tb_arch_624 of project_tb_624 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 499;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (249,0,223,0,210,0,254,0,21,0,97,0,0,0,160,0,81,0,0,0,222,0,118,0,36,0,148,0,151,0,141,0,55,0,215,0,42,0,174,0,192,0,0,0,17,0,237,0,130,0,0,0,35,0,35,0,209,0,237,0,220,0,108,0,74,0,8,0,93,0,249,0,0,0,81,0,190,0,0,0,164,0,0,0,68,0,0,0,228,0,239,0,120,0,245,0,0,0,9,0,0,0,218,0,0,0,140,0,124,0,202,0,99,0,88,0,0,0,0,0,44,0,0,0,203,0,16,0,62,0,0,0,110,0,197,0,157,0,183,0,0,0,65,0,211,0,166,0,219,0,0,0,50,0,198,0,153,0,0,0,70,0,135,0,168,0,0,0,144,0,124,0,0,0,157,0,177,0,77,0,171,0,225,0,144,0,152,0,0,0,240,0,239,0,87,0,145,0,11,0,199,0,218,0,102,0,140,0,88,0,7,0,92,0,0,0,223,0,191,0,0,0,0,0,5,0,94,0,69,0,0,0,19,0,177,0,249,0,208,0,133,0,73,0,117,0,169,0,95,0,0,0,72,0,21,0,143,0,141,0,126,0,0,0,21,0,187,0,85,0,0,0,0,0,122,0,37,0,94,0,0,0,219,0,114,0,0,0,150,0,144,0,199,0,48,0,234,0,0,0,113,0,0,0,61,0,177,0,67,0,0,0,0,0,124,0,56,0,0,0,57,0,0,0,118,0,55,0,237,0,132,0,224,0,57,0,200,0,158,0,17,0,0,0,236,0,99,0,197,0,0,0,122,0,182,0,191,0,58,0,78,0,61,0,134,0,72,0,230,0,56,0,138,0,119,0,14,0,222,0,229,0,229,0,16,0,46,0,0,0,64,0,76,0,53,0,242,0,151,0,246,0,148,0,76,0,234,0,25,0,213,0,181,0,207,0,154,0,101,0,0,0,0,0,0,0,0,0,0,0,170,0,51,0,0,0,43,0,174,0,220,0,51,0,225,0,214,0,159,0,65,0,143,0,0,0,19,0,58,0,232,0,88,0,64,0,107,0,139,0,137,0,130,0,4,0,0,0,39,0,250,0,139,0,20,0,206,0,243,0,117,0,61,0,0,0,86,0,0,0,8,0,99,0,53,0,0,0,92,0,224,0,0,0,0,0,185,0,191,0,251,0,117,0,101,0,184,0,0,0,225,0,249,0,46,0,0,0,0,0,43,0,0,0,98,0,0,0,0,0,206,0,28,0,232,0,211,0,0,0,146,0,0,0,150,0,69,0,50,0,89,0,121,0,0,0,80,0,89,0,56,0,198,0,114,0,58,0,72,0,56,0,208,0,122,0,7,0,254,0,18,0,246,0,185,0,79,0,0,0,71,0,81,0,103,0,98,0,140,0,0,0,65,0,159,0,0,0,129,0,0,0,82,0,231,0,187,0,239,0,83,0,0,0,35,0,0,0,0,0,8,0,216,0,98,0,74,0,255,0,45,0,50,0,0,0,135,0,72,0,169,0,102,0,0,0,3,0,42,0,0,0,39,0,137,0,46,0,0,0,18,0,128,0,72,0,36,0,154,0,34,0,0,0,70,0,96,0,106,0,92,0,65,0,64,0,76,0,0,0,243,0,247,0,117,0,57,0,35,0,78,0,198,0,0,0,2,0,0,0,51,0,0,0,67,0,2,0,245,0,231,0,4,0,130,0,200,0,0,0,0,0,0,0,113,0,74,0,203,0,90,0,91,0,118,0,0,0,67,0,0,0,108,0,50,0,13,0,59,0,131,0,0,0,77,0,2,0,194,0,30,0,0,0,0,0,81,0,168,0,255,0,26,0,113,0,87,0,18,0,0,0,175,0,146,0,215,0,251,0,0,0,39,0,33,0,49,0,219,0,226,0,18,0,235,0,0,0,0,0,124,0,46,0,5,0,254,0,184,0,91,0,150,0,0,0,18,0,35,0,140,0,0,0,87,0,107,0,53,0,182,0,227,0,0,0,215,0,8,0,31,0,60,0,122,0,91,0,240,0,49,0,21,0,0,0,0,0,29,0,233,0,108,0,106,0,135,0,234,0,118,0,156,0,173,0,248,0,125,0,176,0,0,0,105,0,200,0,148,0,168,0,160,0,0,0,177,0,0,0,203,0,157,0,187,0,0,0,0,0,0,0,0,0,139,0,31,0,188,0,181,0,120,0,4,0,141,0,219,0,244,0,210,0,0,0,51,0,122,0,158,0,0,0,121,0,243,0);
signal scenario_full  : scenario_type := (249,31,223,31,210,31,254,31,21,31,97,31,97,30,160,31,81,31,81,30,222,31,118,31,36,31,148,31,151,31,141,31,55,31,215,31,42,31,174,31,192,31,192,30,17,31,237,31,130,31,130,30,35,31,35,31,209,31,237,31,220,31,108,31,74,31,8,31,93,31,249,31,249,30,81,31,190,31,190,30,164,31,164,30,68,31,68,30,228,31,239,31,120,31,245,31,245,30,9,31,9,30,218,31,218,30,140,31,124,31,202,31,99,31,88,31,88,30,88,29,44,31,44,30,203,31,16,31,62,31,62,30,110,31,197,31,157,31,183,31,183,30,65,31,211,31,166,31,219,31,219,30,50,31,198,31,153,31,153,30,70,31,135,31,168,31,168,30,144,31,124,31,124,30,157,31,177,31,77,31,171,31,225,31,144,31,152,31,152,30,240,31,239,31,87,31,145,31,11,31,199,31,218,31,102,31,140,31,88,31,7,31,92,31,92,30,223,31,191,31,191,30,191,29,5,31,94,31,69,31,69,30,19,31,177,31,249,31,208,31,133,31,73,31,117,31,169,31,95,31,95,30,72,31,21,31,143,31,141,31,126,31,126,30,21,31,187,31,85,31,85,30,85,29,122,31,37,31,94,31,94,30,219,31,114,31,114,30,150,31,144,31,199,31,48,31,234,31,234,30,113,31,113,30,61,31,177,31,67,31,67,30,67,29,124,31,56,31,56,30,57,31,57,30,118,31,55,31,237,31,132,31,224,31,57,31,200,31,158,31,17,31,17,30,236,31,99,31,197,31,197,30,122,31,182,31,191,31,58,31,78,31,61,31,134,31,72,31,230,31,56,31,138,31,119,31,14,31,222,31,229,31,229,31,16,31,46,31,46,30,64,31,76,31,53,31,242,31,151,31,246,31,148,31,76,31,234,31,25,31,213,31,181,31,207,31,154,31,101,31,101,30,101,29,101,28,101,27,101,26,170,31,51,31,51,30,43,31,174,31,220,31,51,31,225,31,214,31,159,31,65,31,143,31,143,30,19,31,58,31,232,31,88,31,64,31,107,31,139,31,137,31,130,31,4,31,4,30,39,31,250,31,139,31,20,31,206,31,243,31,117,31,61,31,61,30,86,31,86,30,8,31,99,31,53,31,53,30,92,31,224,31,224,30,224,29,185,31,191,31,251,31,117,31,101,31,184,31,184,30,225,31,249,31,46,31,46,30,46,29,43,31,43,30,98,31,98,30,98,29,206,31,28,31,232,31,211,31,211,30,146,31,146,30,150,31,69,31,50,31,89,31,121,31,121,30,80,31,89,31,56,31,198,31,114,31,58,31,72,31,56,31,208,31,122,31,7,31,254,31,18,31,246,31,185,31,79,31,79,30,71,31,81,31,103,31,98,31,140,31,140,30,65,31,159,31,159,30,129,31,129,30,82,31,231,31,187,31,239,31,83,31,83,30,35,31,35,30,35,29,8,31,216,31,98,31,74,31,255,31,45,31,50,31,50,30,135,31,72,31,169,31,102,31,102,30,3,31,42,31,42,30,39,31,137,31,46,31,46,30,18,31,128,31,72,31,36,31,154,31,34,31,34,30,70,31,96,31,106,31,92,31,65,31,64,31,76,31,76,30,243,31,247,31,117,31,57,31,35,31,78,31,198,31,198,30,2,31,2,30,51,31,51,30,67,31,2,31,245,31,231,31,4,31,130,31,200,31,200,30,200,29,200,28,113,31,74,31,203,31,90,31,91,31,118,31,118,30,67,31,67,30,108,31,50,31,13,31,59,31,131,31,131,30,77,31,2,31,194,31,30,31,30,30,30,29,81,31,168,31,255,31,26,31,113,31,87,31,18,31,18,30,175,31,146,31,215,31,251,31,251,30,39,31,33,31,49,31,219,31,226,31,18,31,235,31,235,30,235,29,124,31,46,31,5,31,254,31,184,31,91,31,150,31,150,30,18,31,35,31,140,31,140,30,87,31,107,31,53,31,182,31,227,31,227,30,215,31,8,31,31,31,60,31,122,31,91,31,240,31,49,31,21,31,21,30,21,29,29,31,233,31,108,31,106,31,135,31,234,31,118,31,156,31,173,31,248,31,125,31,176,31,176,30,105,31,200,31,148,31,168,31,160,31,160,30,177,31,177,30,203,31,157,31,187,31,187,30,187,29,187,28,187,27,139,31,31,31,188,31,181,31,120,31,4,31,141,31,219,31,244,31,210,31,210,30,51,31,122,31,158,31,158,30,121,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
