-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_416 is
end project_tb_416;

architecture project_tb_arch_416 of project_tb_416 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,50,0,0,0,0,0,26,0,83,0,73,0,7,0,135,0,193,0,159,0,49,0,169,0,201,0,73,0,50,0,0,0,26,0,69,0,0,0,158,0,35,0,249,0,217,0,112,0,174,0,126,0,222,0,135,0,35,0,72,0,0,0,3,0,0,0,254,0,102,0,94,0,126,0,191,0,167,0,0,0,27,0,87,0,3,0,0,0,48,0,64,0,0,0,0,0,245,0,53,0,255,0,239,0,119,0,222,0,201,0,11,0,253,0,103,0,187,0,68,0,214,0,0,0,228,0,9,0,45,0,148,0,54,0,158,0,0,0,94,0,132,0,80,0,214,0,1,0,196,0,57,0,52,0,226,0,199,0,251,0,0,0,0,0,30,0,132,0,63,0,211,0,43,0,250,0,0,0,156,0,129,0,0,0,225,0,251,0,81,0,99,0,0,0,0,0,136,0,203,0,213,0,193,0,0,0,0,0,133,0,103,0,195,0,75,0,92,0,41,0,111,0,191,0,59,0,224,0,217,0,12,0,50,0,233,0,250,0,23,0,249,0,38,0,31,0,29,0,231,0,206,0,237,0,165,0,77,0,0,0,161,0,141,0,239,0,80,0,31,0,120,0,119,0,42,0,233,0,12,0,0,0,140,0,62,0,226,0,221,0,0,0,0,0,0,0,69,0,189,0,49,0,107,0,131,0,0,0,0,0,0,0,200,0,121,0,140,0,30,0,247,0,0,0,0,0,0,0,141,0,224,0,38,0,0,0,0,0,83,0,236,0,22,0,89,0,49,0,191,0,125,0,63,0,156,0,247,0,19,0,104,0,19,0,0,0,197,0,181,0,199,0,58,0,187,0,0,0,114,0,115,0,0,0,68,0,247,0,6,0,0,0,0,0,74,0,249,0,0,0,186,0,246,0,0,0,0,0,123,0,54,0,6,0,55,0,111,0,138,0,47,0,44,0,0,0,2,0,74,0,71,0,233,0,136,0,116,0,0,0,141,0,243,0,194,0,0,0,0,0,0,0,64,0,233,0,232,0,138,0,87,0,213,0,17,0,48,0,0,0,47,0,0,0,130,0,0,0,106,0,30,0,80,0,242,0,0,0,0,0,94,0,243,0,122,0,0,0,212,0,0,0,183,0,18,0,60,0,170,0,135,0,50,0,254,0,211,0,131,0,231,0,109,0,253,0,77,0,105,0,14,0,0,0,5,0,86,0,37,0,0,0,79,0,0,0,51,0,143,0,16,0,76,0,39,0,14,0,157,0,0,0,238,0,69,0,220,0,195,0,132,0,243,0,146,0,19,0,246,0,206,0,0,0,0,0,243,0,145,0,181,0,103,0,211,0,156,0,136,0,66,0,91,0,105,0,66,0,46,0,100,0,199,0,125,0,72,0,141,0,143,0,0,0,227,0,137,0,104,0,206,0,4,0,4,0,212,0,20,0,0,0,0,0,141,0,50,0,0,0,6,0,72,0,43,0,0,0,187,0,0,0,200,0,23,0,230,0,45,0,0,0,109,0,13,0,224,0,87,0,173,0,96,0,217,0,239,0,53,0,0,0,51,0,0,0,150,0,0,0,218,0,56,0,244,0,0,0,0,0,0,0,248,0,61,0,21,0,183,0,84,0,196,0,143,0,127,0,0,0,67,0,111,0,161,0,173,0,195,0,0,0,163,0,0,0,81,0,24,0,10,0,169,0,125,0,99,0,0,0,0,0,0,0,174,0,251,0,153,0,27,0,7,0,44,0,0,0,215,0,0,0,95,0,244,0,23,0,77,0,0,0,224,0,215,0,39,0,255,0,139,0,121,0,249,0,238,0,236,0,169,0,88,0,34,0,79,0,218,0,166,0,0,0,5,0,70,0,113,0,24,0,229,0,76,0,114,0,41,0,137,0,198,0,153,0,31,0,188,0,2,0,155,0,27,0,101,0,0,0,98,0,187,0,223,0,76,0,159,0,116,0,155,0,201,0,204,0,12,0,100,0,132,0,71,0,179,0,58,0,93,0,78,0,154,0,137,0,114,0,0,0,0,0,84,0,141,0,112,0,0,0,142,0,128,0,148,0,79,0,114,0,112,0,254,0,0,0,100,0,210,0,76,0,166,0,238,0,37,0,105,0,247,0,122,0,105,0,0,0,204,0,0,0,1,0,226,0,48,0,124,0,248,0,101,0,0,0,27,0,216,0,225,0,0,0,233,0,30,0,191,0,237,0,234,0,33,0,145,0,153,0,116,0,138,0,137,0,0,0,23,0,72,0,238,0,0,0,78,0,0,0,0,0,33,0,208,0,0,0,0,0,220,0,202,0,115,0,105,0,13,0,147,0,153,0,0,0,218,0,65,0,0,0,0,0,154,0,108,0,165,0,15,0,44,0,226,0,250,0,239,0,0,0,0,0,12,0,81,0,171,0,78,0,91,0,207,0,211,0,0,0,134,0,105,0,81,0,72,0,209,0,0,0,16,0,219,0,170,0,0,0,34,0,197,0,0,0,201,0,0,0,52,0,59,0,132,0,124,0,61,0,0,0,64,0,105,0,213,0,62,0,145,0,176,0,86,0,240,0,75,0,198,0,53,0,48,0,222,0,0,0,0,0,0,0,144,0,137,0,245,0,200,0,140,0,209,0,97,0,183,0,44,0,77,0,0,0,0,0,64,0,0,0,0,0,107,0,213,0,234,0,70,0,30,0,69,0,0,0,180,0,240,0,42,0,216,0,197,0,160,0,221,0,0,0,65,0,0,0,190,0,237,0,30,0,144,0,169,0,0,0,140,0,166,0,0,0,0,0,145,0,0,0,76,0,234,0,0,0,187,0,156,0,164,0,167,0,213,0,241,0,89,0,79,0,0,0,0,0,174,0,81,0,93,0,156,0,100,0,250,0,0,0,0,0,133,0,120,0);
signal scenario_full  : scenario_type := (16,31,50,31,50,30,50,29,26,31,83,31,73,31,7,31,135,31,193,31,159,31,49,31,169,31,201,31,73,31,50,31,50,30,26,31,69,31,69,30,158,31,35,31,249,31,217,31,112,31,174,31,126,31,222,31,135,31,35,31,72,31,72,30,3,31,3,30,254,31,102,31,94,31,126,31,191,31,167,31,167,30,27,31,87,31,3,31,3,30,48,31,64,31,64,30,64,29,245,31,53,31,255,31,239,31,119,31,222,31,201,31,11,31,253,31,103,31,187,31,68,31,214,31,214,30,228,31,9,31,45,31,148,31,54,31,158,31,158,30,94,31,132,31,80,31,214,31,1,31,196,31,57,31,52,31,226,31,199,31,251,31,251,30,251,29,30,31,132,31,63,31,211,31,43,31,250,31,250,30,156,31,129,31,129,30,225,31,251,31,81,31,99,31,99,30,99,29,136,31,203,31,213,31,193,31,193,30,193,29,133,31,103,31,195,31,75,31,92,31,41,31,111,31,191,31,59,31,224,31,217,31,12,31,50,31,233,31,250,31,23,31,249,31,38,31,31,31,29,31,231,31,206,31,237,31,165,31,77,31,77,30,161,31,141,31,239,31,80,31,31,31,120,31,119,31,42,31,233,31,12,31,12,30,140,31,62,31,226,31,221,31,221,30,221,29,221,28,69,31,189,31,49,31,107,31,131,31,131,30,131,29,131,28,200,31,121,31,140,31,30,31,247,31,247,30,247,29,247,28,141,31,224,31,38,31,38,30,38,29,83,31,236,31,22,31,89,31,49,31,191,31,125,31,63,31,156,31,247,31,19,31,104,31,19,31,19,30,197,31,181,31,199,31,58,31,187,31,187,30,114,31,115,31,115,30,68,31,247,31,6,31,6,30,6,29,74,31,249,31,249,30,186,31,246,31,246,30,246,29,123,31,54,31,6,31,55,31,111,31,138,31,47,31,44,31,44,30,2,31,74,31,71,31,233,31,136,31,116,31,116,30,141,31,243,31,194,31,194,30,194,29,194,28,64,31,233,31,232,31,138,31,87,31,213,31,17,31,48,31,48,30,47,31,47,30,130,31,130,30,106,31,30,31,80,31,242,31,242,30,242,29,94,31,243,31,122,31,122,30,212,31,212,30,183,31,18,31,60,31,170,31,135,31,50,31,254,31,211,31,131,31,231,31,109,31,253,31,77,31,105,31,14,31,14,30,5,31,86,31,37,31,37,30,79,31,79,30,51,31,143,31,16,31,76,31,39,31,14,31,157,31,157,30,238,31,69,31,220,31,195,31,132,31,243,31,146,31,19,31,246,31,206,31,206,30,206,29,243,31,145,31,181,31,103,31,211,31,156,31,136,31,66,31,91,31,105,31,66,31,46,31,100,31,199,31,125,31,72,31,141,31,143,31,143,30,227,31,137,31,104,31,206,31,4,31,4,31,212,31,20,31,20,30,20,29,141,31,50,31,50,30,6,31,72,31,43,31,43,30,187,31,187,30,200,31,23,31,230,31,45,31,45,30,109,31,13,31,224,31,87,31,173,31,96,31,217,31,239,31,53,31,53,30,51,31,51,30,150,31,150,30,218,31,56,31,244,31,244,30,244,29,244,28,248,31,61,31,21,31,183,31,84,31,196,31,143,31,127,31,127,30,67,31,111,31,161,31,173,31,195,31,195,30,163,31,163,30,81,31,24,31,10,31,169,31,125,31,99,31,99,30,99,29,99,28,174,31,251,31,153,31,27,31,7,31,44,31,44,30,215,31,215,30,95,31,244,31,23,31,77,31,77,30,224,31,215,31,39,31,255,31,139,31,121,31,249,31,238,31,236,31,169,31,88,31,34,31,79,31,218,31,166,31,166,30,5,31,70,31,113,31,24,31,229,31,76,31,114,31,41,31,137,31,198,31,153,31,31,31,188,31,2,31,155,31,27,31,101,31,101,30,98,31,187,31,223,31,76,31,159,31,116,31,155,31,201,31,204,31,12,31,100,31,132,31,71,31,179,31,58,31,93,31,78,31,154,31,137,31,114,31,114,30,114,29,84,31,141,31,112,31,112,30,142,31,128,31,148,31,79,31,114,31,112,31,254,31,254,30,100,31,210,31,76,31,166,31,238,31,37,31,105,31,247,31,122,31,105,31,105,30,204,31,204,30,1,31,226,31,48,31,124,31,248,31,101,31,101,30,27,31,216,31,225,31,225,30,233,31,30,31,191,31,237,31,234,31,33,31,145,31,153,31,116,31,138,31,137,31,137,30,23,31,72,31,238,31,238,30,78,31,78,30,78,29,33,31,208,31,208,30,208,29,220,31,202,31,115,31,105,31,13,31,147,31,153,31,153,30,218,31,65,31,65,30,65,29,154,31,108,31,165,31,15,31,44,31,226,31,250,31,239,31,239,30,239,29,12,31,81,31,171,31,78,31,91,31,207,31,211,31,211,30,134,31,105,31,81,31,72,31,209,31,209,30,16,31,219,31,170,31,170,30,34,31,197,31,197,30,201,31,201,30,52,31,59,31,132,31,124,31,61,31,61,30,64,31,105,31,213,31,62,31,145,31,176,31,86,31,240,31,75,31,198,31,53,31,48,31,222,31,222,30,222,29,222,28,144,31,137,31,245,31,200,31,140,31,209,31,97,31,183,31,44,31,77,31,77,30,77,29,64,31,64,30,64,29,107,31,213,31,234,31,70,31,30,31,69,31,69,30,180,31,240,31,42,31,216,31,197,31,160,31,221,31,221,30,65,31,65,30,190,31,237,31,30,31,144,31,169,31,169,30,140,31,166,31,166,30,166,29,145,31,145,30,76,31,234,31,234,30,187,31,156,31,164,31,167,31,213,31,241,31,89,31,79,31,79,30,79,29,174,31,81,31,93,31,156,31,100,31,250,31,250,30,250,29,133,31,120,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
