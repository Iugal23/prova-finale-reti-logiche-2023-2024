-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_871 is
end project_tb_871;

architecture project_tb_arch_871 of project_tb_871 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 176;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,154,0,0,0,105,0,0,0,42,0,2,0,246,0,204,0,242,0,142,0,124,0,186,0,166,0,133,0,216,0,251,0,93,0,0,0,34,0,33,0,55,0,0,0,0,0,250,0,117,0,186,0,172,0,237,0,244,0,135,0,7,0,171,0,155,0,255,0,2,0,99,0,67,0,34,0,148,0,109,0,114,0,157,0,118,0,144,0,0,0,0,0,39,0,7,0,60,0,31,0,192,0,32,0,202,0,0,0,203,0,159,0,177,0,188,0,0,0,80,0,10,0,200,0,18,0,0,0,177,0,28,0,233,0,136,0,128,0,186,0,43,0,87,0,45,0,103,0,0,0,168,0,0,0,82,0,0,0,14,0,68,0,107,0,0,0,0,0,106,0,119,0,28,0,239,0,121,0,135,0,183,0,82,0,40,0,132,0,218,0,94,0,211,0,128,0,128,0,0,0,119,0,151,0,0,0,122,0,234,0,50,0,32,0,84,0,0,0,72,0,168,0,193,0,0,0,188,0,0,0,97,0,0,0,151,0,0,0,237,0,39,0,109,0,88,0,0,0,43,0,91,0,242,0,160,0,0,0,0,0,211,0,79,0,172,0,0,0,23,0,47,0,136,0,13,0,0,0,0,0,116,0,44,0,0,0,136,0,0,0,111,0,0,0,193,0,163,0,33,0,243,0,198,0,91,0,138,0,174,0,125,0,167,0,10,0,226,0,28,0,0,0,0,0,167,0,198,0,0,0,79,0,165,0,126,0,140,0,201,0,119,0,0,0,145,0,58,0,104,0);
signal scenario_full  : scenario_type := (0,0,154,31,154,30,105,31,105,30,42,31,2,31,246,31,204,31,242,31,142,31,124,31,186,31,166,31,133,31,216,31,251,31,93,31,93,30,34,31,33,31,55,31,55,30,55,29,250,31,117,31,186,31,172,31,237,31,244,31,135,31,7,31,171,31,155,31,255,31,2,31,99,31,67,31,34,31,148,31,109,31,114,31,157,31,118,31,144,31,144,30,144,29,39,31,7,31,60,31,31,31,192,31,32,31,202,31,202,30,203,31,159,31,177,31,188,31,188,30,80,31,10,31,200,31,18,31,18,30,177,31,28,31,233,31,136,31,128,31,186,31,43,31,87,31,45,31,103,31,103,30,168,31,168,30,82,31,82,30,14,31,68,31,107,31,107,30,107,29,106,31,119,31,28,31,239,31,121,31,135,31,183,31,82,31,40,31,132,31,218,31,94,31,211,31,128,31,128,31,128,30,119,31,151,31,151,30,122,31,234,31,50,31,32,31,84,31,84,30,72,31,168,31,193,31,193,30,188,31,188,30,97,31,97,30,151,31,151,30,237,31,39,31,109,31,88,31,88,30,43,31,91,31,242,31,160,31,160,30,160,29,211,31,79,31,172,31,172,30,23,31,47,31,136,31,13,31,13,30,13,29,116,31,44,31,44,30,136,31,136,30,111,31,111,30,193,31,163,31,33,31,243,31,198,31,91,31,138,31,174,31,125,31,167,31,10,31,226,31,28,31,28,30,28,29,167,31,198,31,198,30,79,31,165,31,126,31,140,31,201,31,119,31,119,30,145,31,58,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
