-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_442 is
end project_tb_442;

architecture project_tb_arch_442 of project_tb_442 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 947;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (131,0,75,0,0,0,79,0,0,0,0,0,61,0,49,0,207,0,0,0,0,0,110,0,98,0,0,0,35,0,112,0,59,0,34,0,50,0,147,0,11,0,98,0,63,0,9,0,53,0,156,0,156,0,122,0,24,0,237,0,202,0,168,0,19,0,221,0,128,0,13,0,123,0,144,0,205,0,165,0,108,0,252,0,184,0,9,0,98,0,254,0,238,0,26,0,238,0,85,0,241,0,0,0,26,0,220,0,164,0,246,0,141,0,0,0,87,0,74,0,59,0,163,0,224,0,240,0,0,0,154,0,216,0,177,0,121,0,178,0,0,0,63,0,200,0,147,0,169,0,33,0,73,0,92,0,6,0,139,0,0,0,0,0,154,0,0,0,194,0,132,0,219,0,26,0,219,0,2,0,233,0,164,0,29,0,0,0,254,0,246,0,254,0,0,0,2,0,102,0,0,0,96,0,27,0,0,0,96,0,93,0,0,0,86,0,111,0,237,0,223,0,0,0,150,0,0,0,85,0,61,0,209,0,178,0,218,0,202,0,225,0,40,0,0,0,102,0,220,0,31,0,0,0,107,0,182,0,0,0,237,0,240,0,130,0,173,0,109,0,55,0,16,0,47,0,188,0,129,0,25,0,106,0,76,0,169,0,137,0,247,0,0,0,37,0,20,0,242,0,249,0,248,0,199,0,167,0,5,0,53,0,167,0,226,0,0,0,0,0,249,0,243,0,0,0,226,0,0,0,36,0,11,0,4,0,162,0,118,0,252,0,236,0,0,0,82,0,195,0,0,0,187,0,40,0,187,0,0,0,203,0,238,0,209,0,159,0,183,0,123,0,30,0,0,0,109,0,195,0,241,0,167,0,255,0,192,0,0,0,194,0,150,0,66,0,183,0,91,0,250,0,223,0,0,0,187,0,210,0,4,0,76,0,78,0,236,0,242,0,94,0,37,0,63,0,133,0,106,0,118,0,81,0,214,0,22,0,95,0,241,0,248,0,158,0,191,0,235,0,185,0,229,0,63,0,106,0,205,0,0,0,118,0,123,0,0,0,17,0,34,0,8,0,184,0,0,0,12,0,149,0,102,0,0,0,47,0,211,0,208,0,2,0,222,0,173,0,30,0,0,0,229,0,237,0,124,0,5,0,0,0,90,0,198,0,0,0,149,0,0,0,184,0,138,0,119,0,223,0,243,0,0,0,0,0,0,0,0,0,0,0,133,0,156,0,144,0,0,0,88,0,164,0,150,0,132,0,0,0,9,0,69,0,174,0,70,0,0,0,102,0,0,0,163,0,74,0,240,0,52,0,173,0,73,0,0,0,254,0,201,0,0,0,25,0,228,0,144,0,200,0,5,0,161,0,0,0,0,0,44,0,63,0,0,0,184,0,189,0,30,0,4,0,226,0,97,0,0,0,50,0,162,0,165,0,0,0,66,0,0,0,0,0,41,0,36,0,134,0,0,0,0,0,0,0,0,0,238,0,94,0,115,0,100,0,191,0,138,0,239,0,99,0,0,0,13,0,190,0,153,0,0,0,217,0,34,0,106,0,96,0,0,0,71,0,0,0,158,0,173,0,76,0,12,0,147,0,194,0,0,0,250,0,237,0,5,0,0,0,236,0,65,0,83,0,206,0,130,0,101,0,206,0,241,0,154,0,154,0,118,0,79,0,64,0,0,0,0,0,53,0,192,0,167,0,0,0,0,0,190,0,179,0,61,0,0,0,12,0,108,0,87,0,18,0,207,0,90,0,239,0,27,0,0,0,200,0,0,0,76,0,177,0,18,0,231,0,0,0,124,0,135,0,20,0,117,0,6,0,39,0,252,0,81,0,0,0,170,0,0,0,0,0,76,0,0,0,0,0,145,0,63,0,25,0,15,0,127,0,90,0,0,0,234,0,113,0,90,0,27,0,253,0,184,0,116,0,4,0,138,0,239,0,123,0,160,0,152,0,116,0,238,0,180,0,151,0,42,0,197,0,0,0,97,0,170,0,184,0,237,0,172,0,59,0,160,0,0,0,0,0,47,0,39,0,128,0,63,0,63,0,154,0,11,0,0,0,18,0,26,0,157,0,26,0,0,0,97,0,80,0,191,0,64,0,165,0,21,0,0,0,246,0,232,0,98,0,108,0,254,0,135,0,0,0,138,0,154,0,243,0,45,0,6,0,95,0,136,0,115,0,80,0,115,0,245,0,139,0,183,0,61,0,135,0,92,0,15,0,114,0,18,0,203,0,67,0,251,0,12,0,41,0,27,0,66,0,18,0,0,0,94,0,100,0,124,0,170,0,251,0,122,0,124,0,136,0,235,0,69,0,231,0,108,0,0,0,109,0,0,0,15,0,104,0,0,0,0,0,34,0,20,0,0,0,60,0,188,0,202,0,98,0,52,0,199,0,152,0,33,0,119,0,83,0,86,0,182,0,206,0,152,0,110,0,16,0,52,0,79,0,22,0,90,0,56,0,158,0,0,0,35,0,171,0,235,0,32,0,79,0,30,0,0,0,171,0,155,0,0,0,0,0,125,0,70,0,0,0,90,0,113,0,60,0,192,0,81,0,185,0,0,0,23,0,95,0,216,0,246,0,20,0,98,0,224,0,20,0,0,0,0,0,29,0,28,0,149,0,134,0,0,0,153,0,0,0,6,0,0,0,176,0,0,0,34,0,3,0,225,0,248,0,236,0,35,0,0,0,0,0,139,0,139,0,183,0,67,0,110,0,155,0,23,0,187,0,0,0,0,0,170,0,38,0,215,0,119,0,89,0,107,0,82,0,212,0,149,0,0,0,132,0,0,0,151,0,177,0,85,0,66,0,210,0,0,0,72,0,155,0,120,0,0,0,0,0,0,0,115,0,70,0,152,0,223,0,0,0,0,0,146,0,93,0,187,0,37,0,0,0,115,0,18,0,210,0,88,0,155,0,192,0,198,0,31,0,126,0,174,0,235,0,152,0,16,0,108,0,0,0,0,0,23,0,88,0,75,0,46,0,132,0,248,0,0,0,53,0,0,0,106,0,87,0,0,0,74,0,0,0,37,0,232,0,84,0,229,0,129,0,243,0,224,0,249,0,35,0,0,0,142,0,48,0,54,0,225,0,198,0,192,0,1,0,65,0,25,0,0,0,173,0,175,0,110,0,0,0,0,0,25,0,55,0,242,0,235,0,210,0,68,0,0,0,0,0,136,0,70,0,205,0,220,0,69,0,251,0,243,0,20,0,0,0,148,0,0,0,135,0,14,0,0,0,0,0,88,0,212,0,238,0,127,0,131,0,183,0,22,0,190,0,240,0,0,0,0,0,118,0,134,0,81,0,90,0,6,0,32,0,68,0,0,0,204,0,173,0,211,0,155,0,233,0,249,0,177,0,128,0,63,0,116,0,152,0,120,0,98,0,0,0,217,0,0,0,194,0,196,0,45,0,218,0,80,0,51,0,3,0,239,0,1,0,50,0,0,0,140,0,96,0,32,0,95,0,0,0,254,0,148,0,0,0,171,0,169,0,34,0,184,0,172,0,237,0,57,0,169,0,180,0,241,0,41,0,0,0,223,0,251,0,154,0,237,0,226,0,128,0,89,0,0,0,0,0,134,0,83,0,106,0,146,0,87,0,170,0,253,0,174,0,167,0,179,0,203,0,0,0,195,0,86,0,206,0,38,0,93,0,215,0,100,0,201,0,20,0,110,0,141,0,252,0,121,0,0,0,0,0,57,0,40,0,115,0,0,0,0,0,100,0,68,0,28,0,0,0,237,0,183,0,196,0,0,0,28,0,107,0,14,0,96,0,129,0,0,0,127,0,244,0,0,0,0,0,89,0,33,0,45,0,0,0,24,0,27,0,0,0,161,0,0,0,168,0,238,0,97,0,206,0,0,0,116,0,0,0,28,0,87,0,205,0,0,0,114,0,0,0,0,0,235,0,236,0,118,0,79,0,93,0,121,0,239,0,125,0,46,0,135,0,206,0,179,0,135,0,232,0,55,0,122,0,213,0,118,0,50,0,197,0,32,0,144,0,212,0,239,0,152,0,0,0,106,0,0,0,101,0,177,0,2,0,221,0,141,0,17,0,255,0,139,0,171,0,40,0,48,0,15,0,164,0,0,0,255,0,82,0,115,0,180,0,239,0,124,0,0,0,7,0,142,0,0,0,184,0,120,0,89,0,47,0,0,0,111,0,0,0,56,0,145,0,39,0,0,0,0,0,0,0,0,0,159,0,172,0,0,0,67,0,186,0,36,0,139,0,0,0,100,0);
signal scenario_full  : scenario_type := (131,31,75,31,75,30,79,31,79,30,79,29,61,31,49,31,207,31,207,30,207,29,110,31,98,31,98,30,35,31,112,31,59,31,34,31,50,31,147,31,11,31,98,31,63,31,9,31,53,31,156,31,156,31,122,31,24,31,237,31,202,31,168,31,19,31,221,31,128,31,13,31,123,31,144,31,205,31,165,31,108,31,252,31,184,31,9,31,98,31,254,31,238,31,26,31,238,31,85,31,241,31,241,30,26,31,220,31,164,31,246,31,141,31,141,30,87,31,74,31,59,31,163,31,224,31,240,31,240,30,154,31,216,31,177,31,121,31,178,31,178,30,63,31,200,31,147,31,169,31,33,31,73,31,92,31,6,31,139,31,139,30,139,29,154,31,154,30,194,31,132,31,219,31,26,31,219,31,2,31,233,31,164,31,29,31,29,30,254,31,246,31,254,31,254,30,2,31,102,31,102,30,96,31,27,31,27,30,96,31,93,31,93,30,86,31,111,31,237,31,223,31,223,30,150,31,150,30,85,31,61,31,209,31,178,31,218,31,202,31,225,31,40,31,40,30,102,31,220,31,31,31,31,30,107,31,182,31,182,30,237,31,240,31,130,31,173,31,109,31,55,31,16,31,47,31,188,31,129,31,25,31,106,31,76,31,169,31,137,31,247,31,247,30,37,31,20,31,242,31,249,31,248,31,199,31,167,31,5,31,53,31,167,31,226,31,226,30,226,29,249,31,243,31,243,30,226,31,226,30,36,31,11,31,4,31,162,31,118,31,252,31,236,31,236,30,82,31,195,31,195,30,187,31,40,31,187,31,187,30,203,31,238,31,209,31,159,31,183,31,123,31,30,31,30,30,109,31,195,31,241,31,167,31,255,31,192,31,192,30,194,31,150,31,66,31,183,31,91,31,250,31,223,31,223,30,187,31,210,31,4,31,76,31,78,31,236,31,242,31,94,31,37,31,63,31,133,31,106,31,118,31,81,31,214,31,22,31,95,31,241,31,248,31,158,31,191,31,235,31,185,31,229,31,63,31,106,31,205,31,205,30,118,31,123,31,123,30,17,31,34,31,8,31,184,31,184,30,12,31,149,31,102,31,102,30,47,31,211,31,208,31,2,31,222,31,173,31,30,31,30,30,229,31,237,31,124,31,5,31,5,30,90,31,198,31,198,30,149,31,149,30,184,31,138,31,119,31,223,31,243,31,243,30,243,29,243,28,243,27,243,26,133,31,156,31,144,31,144,30,88,31,164,31,150,31,132,31,132,30,9,31,69,31,174,31,70,31,70,30,102,31,102,30,163,31,74,31,240,31,52,31,173,31,73,31,73,30,254,31,201,31,201,30,25,31,228,31,144,31,200,31,5,31,161,31,161,30,161,29,44,31,63,31,63,30,184,31,189,31,30,31,4,31,226,31,97,31,97,30,50,31,162,31,165,31,165,30,66,31,66,30,66,29,41,31,36,31,134,31,134,30,134,29,134,28,134,27,238,31,94,31,115,31,100,31,191,31,138,31,239,31,99,31,99,30,13,31,190,31,153,31,153,30,217,31,34,31,106,31,96,31,96,30,71,31,71,30,158,31,173,31,76,31,12,31,147,31,194,31,194,30,250,31,237,31,5,31,5,30,236,31,65,31,83,31,206,31,130,31,101,31,206,31,241,31,154,31,154,31,118,31,79,31,64,31,64,30,64,29,53,31,192,31,167,31,167,30,167,29,190,31,179,31,61,31,61,30,12,31,108,31,87,31,18,31,207,31,90,31,239,31,27,31,27,30,200,31,200,30,76,31,177,31,18,31,231,31,231,30,124,31,135,31,20,31,117,31,6,31,39,31,252,31,81,31,81,30,170,31,170,30,170,29,76,31,76,30,76,29,145,31,63,31,25,31,15,31,127,31,90,31,90,30,234,31,113,31,90,31,27,31,253,31,184,31,116,31,4,31,138,31,239,31,123,31,160,31,152,31,116,31,238,31,180,31,151,31,42,31,197,31,197,30,97,31,170,31,184,31,237,31,172,31,59,31,160,31,160,30,160,29,47,31,39,31,128,31,63,31,63,31,154,31,11,31,11,30,18,31,26,31,157,31,26,31,26,30,97,31,80,31,191,31,64,31,165,31,21,31,21,30,246,31,232,31,98,31,108,31,254,31,135,31,135,30,138,31,154,31,243,31,45,31,6,31,95,31,136,31,115,31,80,31,115,31,245,31,139,31,183,31,61,31,135,31,92,31,15,31,114,31,18,31,203,31,67,31,251,31,12,31,41,31,27,31,66,31,18,31,18,30,94,31,100,31,124,31,170,31,251,31,122,31,124,31,136,31,235,31,69,31,231,31,108,31,108,30,109,31,109,30,15,31,104,31,104,30,104,29,34,31,20,31,20,30,60,31,188,31,202,31,98,31,52,31,199,31,152,31,33,31,119,31,83,31,86,31,182,31,206,31,152,31,110,31,16,31,52,31,79,31,22,31,90,31,56,31,158,31,158,30,35,31,171,31,235,31,32,31,79,31,30,31,30,30,171,31,155,31,155,30,155,29,125,31,70,31,70,30,90,31,113,31,60,31,192,31,81,31,185,31,185,30,23,31,95,31,216,31,246,31,20,31,98,31,224,31,20,31,20,30,20,29,29,31,28,31,149,31,134,31,134,30,153,31,153,30,6,31,6,30,176,31,176,30,34,31,3,31,225,31,248,31,236,31,35,31,35,30,35,29,139,31,139,31,183,31,67,31,110,31,155,31,23,31,187,31,187,30,187,29,170,31,38,31,215,31,119,31,89,31,107,31,82,31,212,31,149,31,149,30,132,31,132,30,151,31,177,31,85,31,66,31,210,31,210,30,72,31,155,31,120,31,120,30,120,29,120,28,115,31,70,31,152,31,223,31,223,30,223,29,146,31,93,31,187,31,37,31,37,30,115,31,18,31,210,31,88,31,155,31,192,31,198,31,31,31,126,31,174,31,235,31,152,31,16,31,108,31,108,30,108,29,23,31,88,31,75,31,46,31,132,31,248,31,248,30,53,31,53,30,106,31,87,31,87,30,74,31,74,30,37,31,232,31,84,31,229,31,129,31,243,31,224,31,249,31,35,31,35,30,142,31,48,31,54,31,225,31,198,31,192,31,1,31,65,31,25,31,25,30,173,31,175,31,110,31,110,30,110,29,25,31,55,31,242,31,235,31,210,31,68,31,68,30,68,29,136,31,70,31,205,31,220,31,69,31,251,31,243,31,20,31,20,30,148,31,148,30,135,31,14,31,14,30,14,29,88,31,212,31,238,31,127,31,131,31,183,31,22,31,190,31,240,31,240,30,240,29,118,31,134,31,81,31,90,31,6,31,32,31,68,31,68,30,204,31,173,31,211,31,155,31,233,31,249,31,177,31,128,31,63,31,116,31,152,31,120,31,98,31,98,30,217,31,217,30,194,31,196,31,45,31,218,31,80,31,51,31,3,31,239,31,1,31,50,31,50,30,140,31,96,31,32,31,95,31,95,30,254,31,148,31,148,30,171,31,169,31,34,31,184,31,172,31,237,31,57,31,169,31,180,31,241,31,41,31,41,30,223,31,251,31,154,31,237,31,226,31,128,31,89,31,89,30,89,29,134,31,83,31,106,31,146,31,87,31,170,31,253,31,174,31,167,31,179,31,203,31,203,30,195,31,86,31,206,31,38,31,93,31,215,31,100,31,201,31,20,31,110,31,141,31,252,31,121,31,121,30,121,29,57,31,40,31,115,31,115,30,115,29,100,31,68,31,28,31,28,30,237,31,183,31,196,31,196,30,28,31,107,31,14,31,96,31,129,31,129,30,127,31,244,31,244,30,244,29,89,31,33,31,45,31,45,30,24,31,27,31,27,30,161,31,161,30,168,31,238,31,97,31,206,31,206,30,116,31,116,30,28,31,87,31,205,31,205,30,114,31,114,30,114,29,235,31,236,31,118,31,79,31,93,31,121,31,239,31,125,31,46,31,135,31,206,31,179,31,135,31,232,31,55,31,122,31,213,31,118,31,50,31,197,31,32,31,144,31,212,31,239,31,152,31,152,30,106,31,106,30,101,31,177,31,2,31,221,31,141,31,17,31,255,31,139,31,171,31,40,31,48,31,15,31,164,31,164,30,255,31,82,31,115,31,180,31,239,31,124,31,124,30,7,31,142,31,142,30,184,31,120,31,89,31,47,31,47,30,111,31,111,30,56,31,145,31,39,31,39,30,39,29,39,28,39,27,159,31,172,31,172,30,67,31,186,31,36,31,139,31,139,30,100,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
