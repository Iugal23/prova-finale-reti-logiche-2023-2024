-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 990;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,178,0,25,0,129,0,84,0,29,0,0,0,227,0,0,0,72,0,32,0,164,0,83,0,60,0,150,0,131,0,208,0,194,0,37,0,197,0,23,0,174,0,118,0,3,0,18,0,165,0,84,0,212,0,146,0,230,0,41,0,0,0,38,0,22,0,213,0,213,0,184,0,179,0,47,0,136,0,50,0,246,0,0,0,202,0,115,0,22,0,124,0,120,0,220,0,207,0,61,0,255,0,0,0,0,0,23,0,0,0,0,0,238,0,21,0,170,0,116,0,92,0,228,0,235,0,78,0,73,0,47,0,197,0,4,0,0,0,244,0,0,0,0,0,17,0,0,0,7,0,20,0,88,0,119,0,199,0,0,0,38,0,0,0,0,0,204,0,21,0,0,0,218,0,216,0,0,0,0,0,87,0,181,0,0,0,181,0,160,0,0,0,195,0,134,0,6,0,195,0,39,0,0,0,0,0,161,0,0,0,244,0,243,0,155,0,28,0,56,0,203,0,0,0,0,0,135,0,109,0,0,0,0,0,205,0,0,0,147,0,108,0,226,0,244,0,19,0,129,0,130,0,0,0,34,0,219,0,0,0,118,0,132,0,113,0,0,0,39,0,0,0,126,0,159,0,250,0,114,0,186,0,154,0,52,0,90,0,122,0,0,0,54,0,168,0,190,0,213,0,44,0,102,0,213,0,38,0,94,0,187,0,47,0,131,0,38,0,42,0,79,0,68,0,0,0,69,0,18,0,0,0,0,0,196,0,41,0,55,0,167,0,167,0,202,0,114,0,52,0,0,0,226,0,220,0,0,0,36,0,135,0,47,0,68,0,0,0,0,0,212,0,191,0,0,0,214,0,70,0,204,0,242,0,244,0,0,0,28,0,232,0,163,0,62,0,178,0,170,0,26,0,50,0,108,0,45,0,16,0,79,0,67,0,0,0,16,0,8,0,164,0,78,0,0,0,191,0,91,0,184,0,17,0,0,0,234,0,54,0,114,0,90,0,0,0,192,0,239,0,50,0,251,0,160,0,0,0,0,0,123,0,101,0,0,0,0,0,83,0,250,0,192,0,49,0,195,0,52,0,182,0,247,0,0,0,0,0,6,0,9,0,0,0,6,0,145,0,86,0,98,0,55,0,148,0,75,0,231,0,224,0,142,0,172,0,191,0,0,0,223,0,254,0,0,0,0,0,133,0,245,0,78,0,79,0,0,0,135,0,0,0,131,0,0,0,19,0,213,0,0,0,207,0,18,0,251,0,226,0,28,0,0,0,238,0,66,0,14,0,0,0,0,0,234,0,26,0,83,0,0,0,151,0,200,0,231,0,235,0,0,0,98,0,181,0,162,0,215,0,228,0,76,0,160,0,28,0,87,0,0,0,70,0,0,0,91,0,190,0,16,0,145,0,0,0,116,0,66,0,244,0,30,0,113,0,50,0,0,0,219,0,33,0,0,0,242,0,0,0,33,0,4,0,113,0,0,0,0,0,0,0,1,0,45,0,135,0,0,0,0,0,115,0,195,0,249,0,182,0,71,0,28,0,0,0,1,0,91,0,0,0,0,0,174,0,72,0,132,0,230,0,133,0,0,0,0,0,188,0,21,0,213,0,0,0,211,0,207,0,217,0,124,0,121,0,0,0,0,0,86,0,150,0,0,0,222,0,36,0,0,0,34,0,162,0,0,0,222,0,64,0,33,0,90,0,62,0,202,0,0,0,121,0,38,0,2,0,0,0,151,0,221,0,0,0,129,0,57,0,202,0,252,0,0,0,126,0,30,0,11,0,71,0,111,0,13,0,0,0,50,0,171,0,254,0,211,0,164,0,135,0,0,0,37,0,245,0,234,0,149,0,0,0,0,0,75,0,11,0,17,0,150,0,242,0,168,0,8,0,128,0,130,0,231,0,0,0,163,0,0,0,112,0,0,0,0,0,165,0,0,0,0,0,76,0,42,0,219,0,161,0,222,0,171,0,0,0,163,0,0,0,27,0,245,0,88,0,166,0,192,0,113,0,0,0,173,0,52,0,236,0,202,0,53,0,219,0,32,0,142,0,103,0,132,0,243,0,53,0,244,0,192,0,0,0,219,0,180,0,143,0,105,0,31,0,193,0,130,0,233,0,123,0,224,0,191,0,42,0,0,0,244,0,48,0,61,0,104,0,22,0,89,0,8,0,0,0,86,0,0,0,82,0,238,0,48,0,0,0,235,0,0,0,105,0,0,0,44,0,139,0,16,0,141,0,222,0,45,0,0,0,67,0,211,0,132,0,212,0,125,0,191,0,13,0,167,0,0,0,66,0,243,0,0,0,206,0,112,0,105,0,47,0,125,0,134,0,150,0,178,0,0,0,89,0,0,0,44,0,233,0,31,0,22,0,32,0,162,0,27,0,95,0,185,0,1,0,219,0,44,0,102,0,245,0,0,0,224,0,33,0,0,0,0,0,53,0,0,0,2,0,249,0,0,0,78,0,224,0,77,0,243,0,230,0,127,0,168,0,11,0,91,0,0,0,79,0,0,0,0,0,158,0,0,0,117,0,158,0,162,0,0,0,40,0,235,0,204,0,117,0,155,0,49,0,73,0,48,0,96,0,8,0,64,0,195,0,125,0,57,0,0,0,0,0,44,0,122,0,0,0,210,0,23,0,207,0,0,0,36,0,0,0,60,0,117,0,213,0,173,0,162,0,69,0,193,0,83,0,76,0,0,0,120,0,0,0,0,0,0,0,221,0,187,0,177,0,0,0,123,0,94,0,108,0,36,0,20,0,0,0,0,0,177,0,0,0,12,0,53,0,111,0,0,0,128,0,0,0,97,0,199,0,181,0,136,0,232,0,216,0,0,0,1,0,0,0,229,0,125,0,0,0,186,0,162,0,224,0,89,0,244,0,178,0,62,0,98,0,16,0,69,0,0,0,0,0,141,0,90,0,46,0,90,0,23,0,84,0,112,0,164,0,194,0,92,0,93,0,92,0,131,0,121,0,127,0,161,0,246,0,90,0,167,0,199,0,233,0,115,0,99,0,189,0,104,0,89,0,46,0,0,0,102,0,32,0,74,0,0,0,83,0,102,0,0,0,0,0,36,0,245,0,10,0,142,0,47,0,104,0,243,0,0,0,0,0,123,0,181,0,100,0,169,0,149,0,252,0,211,0,152,0,229,0,118,0,0,0,238,0,142,0,12,0,0,0,125,0,0,0,136,0,243,0,28,0,0,0,213,0,21,0,104,0,112,0,0,0,42,0,0,0,0,0,233,0,10,0,28,0,138,0,158,0,0,0,34,0,41,0,157,0,24,0,0,0,16,0,170,0,0,0,105,0,0,0,37,0,51,0,245,0,0,0,19,0,160,0,97,0,221,0,151,0,238,0,0,0,59,0,211,0,180,0,9,0,160,0,218,0,188,0,54,0,54,0,134,0,180,0,0,0,0,0,96,0,114,0,125,0,230,0,190,0,147,0,0,0,207,0,45,0,13,0,234,0,155,0,253,0,121,0,98,0,144,0,235,0,214,0,254,0,51,0,25,0,17,0,222,0,182,0,220,0,203,0,92,0,99,0,17,0,72,0,229,0,2,0,233,0,140,0,208,0,94,0,0,0,0,0,29,0,115,0,200,0,176,0,83,0,215,0,0,0,47,0,40,0,190,0,165,0,0,0,100,0,131,0,0,0,155,0,0,0,60,0,0,0,7,0,0,0,230,0,251,0,142,0,84,0,34,0,251,0,51,0,188,0,87,0,188,0,181,0,0,0,207,0,163,0,5,0,251,0,0,0,130,0,194,0,108,0,0,0,199,0,0,0,0,0,252,0,0,0,124,0,55,0,25,0,145,0,0,0,141,0,190,0,37,0,121,0,155,0,160,0,249,0,0,0,69,0,171,0,39,0,0,0,250,0,184,0,197,0,0,0,90,0,60,0,118,0,100,0,0,0,62,0,69,0,0,0,5,0,223,0,157,0,27,0,79,0,108,0,0,0,142,0,26,0,37,0,196,0,93,0,196,0,0,0,108,0,167,0,9,0,26,0,160,0,202,0,5,0,61,0,70,0,254,0,85,0,14,0,0,0,157,0,142,0,166,0,56,0,211,0,32,0,0,0,53,0,161,0,0,0,113,0,0,0,0,0,0,0,32,0,0,0,36,0,3,0,144,0,177,0,21,0,72,0,226,0,134,0,91,0,160,0,38,0,128,0,35,0,0,0,215,0,147,0,81,0,16,0,148,0,0,0,233,0,107,0,33,0,233,0,32,0,185,0,184,0,81,0,174,0,0,0,0,0,136,0,57,0,31,0,242,0,174,0,50,0,17,0,16,0,78,0,167,0,0,0,153,0,90,0,0,0,236,0,84,0,0,0,0,0,13,0,64,0,0,0,149,0,120,0,56,0,0,0,237,0,68,0,150,0,0,0,50,0,128,0,87,0,178,0,166,0,101,0,251,0,187,0,238,0);
signal scenario_full  : scenario_type := (0,0,178,31,25,31,129,31,84,31,29,31,29,30,227,31,227,30,72,31,32,31,164,31,83,31,60,31,150,31,131,31,208,31,194,31,37,31,197,31,23,31,174,31,118,31,3,31,18,31,165,31,84,31,212,31,146,31,230,31,41,31,41,30,38,31,22,31,213,31,213,31,184,31,179,31,47,31,136,31,50,31,246,31,246,30,202,31,115,31,22,31,124,31,120,31,220,31,207,31,61,31,255,31,255,30,255,29,23,31,23,30,23,29,238,31,21,31,170,31,116,31,92,31,228,31,235,31,78,31,73,31,47,31,197,31,4,31,4,30,244,31,244,30,244,29,17,31,17,30,7,31,20,31,88,31,119,31,199,31,199,30,38,31,38,30,38,29,204,31,21,31,21,30,218,31,216,31,216,30,216,29,87,31,181,31,181,30,181,31,160,31,160,30,195,31,134,31,6,31,195,31,39,31,39,30,39,29,161,31,161,30,244,31,243,31,155,31,28,31,56,31,203,31,203,30,203,29,135,31,109,31,109,30,109,29,205,31,205,30,147,31,108,31,226,31,244,31,19,31,129,31,130,31,130,30,34,31,219,31,219,30,118,31,132,31,113,31,113,30,39,31,39,30,126,31,159,31,250,31,114,31,186,31,154,31,52,31,90,31,122,31,122,30,54,31,168,31,190,31,213,31,44,31,102,31,213,31,38,31,94,31,187,31,47,31,131,31,38,31,42,31,79,31,68,31,68,30,69,31,18,31,18,30,18,29,196,31,41,31,55,31,167,31,167,31,202,31,114,31,52,31,52,30,226,31,220,31,220,30,36,31,135,31,47,31,68,31,68,30,68,29,212,31,191,31,191,30,214,31,70,31,204,31,242,31,244,31,244,30,28,31,232,31,163,31,62,31,178,31,170,31,26,31,50,31,108,31,45,31,16,31,79,31,67,31,67,30,16,31,8,31,164,31,78,31,78,30,191,31,91,31,184,31,17,31,17,30,234,31,54,31,114,31,90,31,90,30,192,31,239,31,50,31,251,31,160,31,160,30,160,29,123,31,101,31,101,30,101,29,83,31,250,31,192,31,49,31,195,31,52,31,182,31,247,31,247,30,247,29,6,31,9,31,9,30,6,31,145,31,86,31,98,31,55,31,148,31,75,31,231,31,224,31,142,31,172,31,191,31,191,30,223,31,254,31,254,30,254,29,133,31,245,31,78,31,79,31,79,30,135,31,135,30,131,31,131,30,19,31,213,31,213,30,207,31,18,31,251,31,226,31,28,31,28,30,238,31,66,31,14,31,14,30,14,29,234,31,26,31,83,31,83,30,151,31,200,31,231,31,235,31,235,30,98,31,181,31,162,31,215,31,228,31,76,31,160,31,28,31,87,31,87,30,70,31,70,30,91,31,190,31,16,31,145,31,145,30,116,31,66,31,244,31,30,31,113,31,50,31,50,30,219,31,33,31,33,30,242,31,242,30,33,31,4,31,113,31,113,30,113,29,113,28,1,31,45,31,135,31,135,30,135,29,115,31,195,31,249,31,182,31,71,31,28,31,28,30,1,31,91,31,91,30,91,29,174,31,72,31,132,31,230,31,133,31,133,30,133,29,188,31,21,31,213,31,213,30,211,31,207,31,217,31,124,31,121,31,121,30,121,29,86,31,150,31,150,30,222,31,36,31,36,30,34,31,162,31,162,30,222,31,64,31,33,31,90,31,62,31,202,31,202,30,121,31,38,31,2,31,2,30,151,31,221,31,221,30,129,31,57,31,202,31,252,31,252,30,126,31,30,31,11,31,71,31,111,31,13,31,13,30,50,31,171,31,254,31,211,31,164,31,135,31,135,30,37,31,245,31,234,31,149,31,149,30,149,29,75,31,11,31,17,31,150,31,242,31,168,31,8,31,128,31,130,31,231,31,231,30,163,31,163,30,112,31,112,30,112,29,165,31,165,30,165,29,76,31,42,31,219,31,161,31,222,31,171,31,171,30,163,31,163,30,27,31,245,31,88,31,166,31,192,31,113,31,113,30,173,31,52,31,236,31,202,31,53,31,219,31,32,31,142,31,103,31,132,31,243,31,53,31,244,31,192,31,192,30,219,31,180,31,143,31,105,31,31,31,193,31,130,31,233,31,123,31,224,31,191,31,42,31,42,30,244,31,48,31,61,31,104,31,22,31,89,31,8,31,8,30,86,31,86,30,82,31,238,31,48,31,48,30,235,31,235,30,105,31,105,30,44,31,139,31,16,31,141,31,222,31,45,31,45,30,67,31,211,31,132,31,212,31,125,31,191,31,13,31,167,31,167,30,66,31,243,31,243,30,206,31,112,31,105,31,47,31,125,31,134,31,150,31,178,31,178,30,89,31,89,30,44,31,233,31,31,31,22,31,32,31,162,31,27,31,95,31,185,31,1,31,219,31,44,31,102,31,245,31,245,30,224,31,33,31,33,30,33,29,53,31,53,30,2,31,249,31,249,30,78,31,224,31,77,31,243,31,230,31,127,31,168,31,11,31,91,31,91,30,79,31,79,30,79,29,158,31,158,30,117,31,158,31,162,31,162,30,40,31,235,31,204,31,117,31,155,31,49,31,73,31,48,31,96,31,8,31,64,31,195,31,125,31,57,31,57,30,57,29,44,31,122,31,122,30,210,31,23,31,207,31,207,30,36,31,36,30,60,31,117,31,213,31,173,31,162,31,69,31,193,31,83,31,76,31,76,30,120,31,120,30,120,29,120,28,221,31,187,31,177,31,177,30,123,31,94,31,108,31,36,31,20,31,20,30,20,29,177,31,177,30,12,31,53,31,111,31,111,30,128,31,128,30,97,31,199,31,181,31,136,31,232,31,216,31,216,30,1,31,1,30,229,31,125,31,125,30,186,31,162,31,224,31,89,31,244,31,178,31,62,31,98,31,16,31,69,31,69,30,69,29,141,31,90,31,46,31,90,31,23,31,84,31,112,31,164,31,194,31,92,31,93,31,92,31,131,31,121,31,127,31,161,31,246,31,90,31,167,31,199,31,233,31,115,31,99,31,189,31,104,31,89,31,46,31,46,30,102,31,32,31,74,31,74,30,83,31,102,31,102,30,102,29,36,31,245,31,10,31,142,31,47,31,104,31,243,31,243,30,243,29,123,31,181,31,100,31,169,31,149,31,252,31,211,31,152,31,229,31,118,31,118,30,238,31,142,31,12,31,12,30,125,31,125,30,136,31,243,31,28,31,28,30,213,31,21,31,104,31,112,31,112,30,42,31,42,30,42,29,233,31,10,31,28,31,138,31,158,31,158,30,34,31,41,31,157,31,24,31,24,30,16,31,170,31,170,30,105,31,105,30,37,31,51,31,245,31,245,30,19,31,160,31,97,31,221,31,151,31,238,31,238,30,59,31,211,31,180,31,9,31,160,31,218,31,188,31,54,31,54,31,134,31,180,31,180,30,180,29,96,31,114,31,125,31,230,31,190,31,147,31,147,30,207,31,45,31,13,31,234,31,155,31,253,31,121,31,98,31,144,31,235,31,214,31,254,31,51,31,25,31,17,31,222,31,182,31,220,31,203,31,92,31,99,31,17,31,72,31,229,31,2,31,233,31,140,31,208,31,94,31,94,30,94,29,29,31,115,31,200,31,176,31,83,31,215,31,215,30,47,31,40,31,190,31,165,31,165,30,100,31,131,31,131,30,155,31,155,30,60,31,60,30,7,31,7,30,230,31,251,31,142,31,84,31,34,31,251,31,51,31,188,31,87,31,188,31,181,31,181,30,207,31,163,31,5,31,251,31,251,30,130,31,194,31,108,31,108,30,199,31,199,30,199,29,252,31,252,30,124,31,55,31,25,31,145,31,145,30,141,31,190,31,37,31,121,31,155,31,160,31,249,31,249,30,69,31,171,31,39,31,39,30,250,31,184,31,197,31,197,30,90,31,60,31,118,31,100,31,100,30,62,31,69,31,69,30,5,31,223,31,157,31,27,31,79,31,108,31,108,30,142,31,26,31,37,31,196,31,93,31,196,31,196,30,108,31,167,31,9,31,26,31,160,31,202,31,5,31,61,31,70,31,254,31,85,31,14,31,14,30,157,31,142,31,166,31,56,31,211,31,32,31,32,30,53,31,161,31,161,30,113,31,113,30,113,29,113,28,32,31,32,30,36,31,3,31,144,31,177,31,21,31,72,31,226,31,134,31,91,31,160,31,38,31,128,31,35,31,35,30,215,31,147,31,81,31,16,31,148,31,148,30,233,31,107,31,33,31,233,31,32,31,185,31,184,31,81,31,174,31,174,30,174,29,136,31,57,31,31,31,242,31,174,31,50,31,17,31,16,31,78,31,167,31,167,30,153,31,90,31,90,30,236,31,84,31,84,30,84,29,13,31,64,31,64,30,149,31,120,31,56,31,56,30,237,31,68,31,150,31,150,30,50,31,128,31,87,31,178,31,166,31,101,31,251,31,187,31,238,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
