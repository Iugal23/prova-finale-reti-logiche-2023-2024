-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 812;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,0,0,0,0,50,0,194,0,157,0,0,0,117,0,243,0,249,0,0,0,9,0,0,0,55,0,0,0,51,0,164,0,173,0,183,0,116,0,94,0,0,0,70,0,185,0,45,0,168,0,101,0,10,0,146,0,121,0,0,0,27,0,196,0,44,0,88,0,134,0,84,0,63,0,39,0,123,0,224,0,101,0,237,0,0,0,159,0,218,0,0,0,137,0,180,0,198,0,0,0,185,0,139,0,222,0,100,0,0,0,131,0,56,0,0,0,120,0,166,0,6,0,218,0,244,0,154,0,224,0,137,0,184,0,158,0,137,0,16,0,79,0,40,0,253,0,62,0,0,0,0,0,26,0,176,0,251,0,20,0,248,0,158,0,56,0,0,0,0,0,49,0,189,0,0,0,141,0,168,0,131,0,106,0,0,0,177,0,91,0,230,0,131,0,129,0,200,0,31,0,230,0,223,0,80,0,236,0,0,0,0,0,36,0,176,0,216,0,254,0,190,0,0,0,132,0,218,0,0,0,0,0,107,0,115,0,91,0,24,0,15,0,146,0,97,0,180,0,0,0,147,0,0,0,111,0,176,0,169,0,53,0,130,0,1,0,30,0,37,0,233,0,219,0,192,0,68,0,36,0,139,0,87,0,57,0,119,0,229,0,139,0,179,0,245,0,0,0,131,0,185,0,76,0,52,0,137,0,116,0,5,0,56,0,200,0,106,0,139,0,238,0,43,0,216,0,143,0,117,0,0,0,13,0,0,0,121,0,68,0,0,0,172,0,8,0,198,0,184,0,230,0,62,0,14,0,222,0,102,0,46,0,34,0,27,0,0,0,175,0,159,0,236,0,115,0,104,0,239,0,168,0,6,0,203,0,66,0,0,0,0,0,0,0,0,0,0,0,0,0,94,0,92,0,129,0,88,0,0,0,14,0,20,0,178,0,248,0,37,0,0,0,40,0,134,0,68,0,96,0,60,0,85,0,190,0,226,0,0,0,104,0,157,0,50,0,248,0,250,0,166,0,162,0,0,0,221,0,206,0,215,0,121,0,238,0,123,0,4,0,0,0,229,0,28,0,39,0,20,0,0,0,0,0,67,0,69,0,143,0,0,0,48,0,121,0,0,0,0,0,78,0,0,0,44,0,93,0,40,0,127,0,144,0,22,0,218,0,0,0,162,0,249,0,253,0,0,0,161,0,116,0,181,0,38,0,0,0,134,0,88,0,74,0,1,0,0,0,217,0,0,0,43,0,0,0,136,0,181,0,48,0,169,0,90,0,38,0,193,0,154,0,242,0,0,0,49,0,165,0,220,0,0,0,0,0,40,0,8,0,109,0,26,0,189,0,223,0,110,0,196,0,0,0,109,0,236,0,0,0,0,0,71,0,182,0,191,0,201,0,68,0,0,0,130,0,210,0,171,0,0,0,175,0,0,0,120,0,169,0,203,0,4,0,244,0,187,0,72,0,160,0,231,0,147,0,52,0,115,0,113,0,8,0,193,0,189,0,119,0,11,0,102,0,0,0,77,0,224,0,180,0,182,0,0,0,15,0,245,0,113,0,164,0,214,0,133,0,107,0,103,0,0,0,0,0,122,0,0,0,41,0,190,0,34,0,229,0,0,0,173,0,83,0,20,0,97,0,33,0,0,0,62,0,0,0,0,0,0,0,148,0,26,0,149,0,60,0,32,0,1,0,73,0,208,0,72,0,76,0,0,0,0,0,0,0,47,0,205,0,0,0,133,0,214,0,0,0,104,0,9,0,98,0,0,0,220,0,118,0,0,0,7,0,239,0,244,0,0,0,75,0,111,0,185,0,3,0,17,0,73,0,0,0,92,0,79,0,159,0,0,0,215,0,2,0,46,0,95,0,0,0,111,0,151,0,153,0,29,0,90,0,202,0,0,0,15,0,117,0,177,0,39,0,83,0,56,0,41,0,2,0,17,0,173,0,194,0,224,0,13,0,194,0,156,0,232,0,221,0,34,0,0,0,161,0,174,0,0,0,0,0,0,0,183,0,244,0,34,0,93,0,242,0,144,0,0,0,174,0,78,0,168,0,83,0,15,0,242,0,128,0,157,0,0,0,84,0,182,0,232,0,0,0,68,0,142,0,0,0,66,0,8,0,0,0,127,0,116,0,15,0,173,0,174,0,0,0,0,0,16,0,233,0,86,0,165,0,0,0,36,0,0,0,166,0,127,0,71,0,0,0,216,0,25,0,110,0,0,0,0,0,136,0,188,0,148,0,103,0,225,0,27,0,149,0,0,0,186,0,254,0,237,0,252,0,112,0,0,0,205,0,96,0,43,0,0,0,55,0,65,0,183,0,248,0,79,0,236,0,134,0,55,0,153,0,162,0,150,0,0,0,212,0,240,0,234,0,139,0,58,0,218,0,84,0,0,0,0,0,0,0,178,0,19,0,221,0,128,0,148,0,0,0,217,0,227,0,86,0,22,0,194,0,132,0,148,0,106,0,212,0,92,0,98,0,144,0,221,0,176,0,0,0,226,0,124,0,50,0,245,0,52,0,206,0,126,0,0,0,236,0,157,0,0,0,245,0,142,0,124,0,147,0,242,0,41,0,0,0,84,0,98,0,147,0,126,0,82,0,119,0,46,0,161,0,71,0,146,0,0,0,4,0,201,0,0,0,0,0,251,0,157,0,161,0,113,0,134,0,0,0,200,0,31,0,0,0,18,0,14,0,214,0,36,0,125,0,4,0,0,0,0,0,247,0,75,0,199,0,48,0,203,0,102,0,173,0,58,0,68,0,182,0,35,0,40,0,58,0,11,0,220,0,4,0,223,0,34,0,0,0,105,0,149,0,0,0,200,0,158,0,185,0,18,0,141,0,49,0,129,0,221,0,0,0,244,0,25,0,73,0,0,0,94,0,105,0,13,0,30,0,144,0,109,0,115,0,218,0,204,0,69,0,197,0,55,0,185,0,87,0,0,0,41,0,120,0,53,0,134,0,163,0,162,0,201,0,247,0,0,0,239,0,197,0,158,0,95,0,148,0,207,0,206,0,209,0,47,0,184,0,89,0,9,0,248,0,233,0,162,0,49,0,214,0,0,0,0,0,211,0,184,0,235,0,105,0,239,0,85,0,203,0,238,0,7,0,228,0,0,0,87,0,158,0,230,0,173,0,0,0,185,0,5,0,0,0,0,0,193,0,90,0,0,0,158,0,233,0,179,0,94,0,0,0,45,0,46,0,64,0,236,0,253,0,153,0,133,0,56,0,203,0,51,0,70,0,227,0,0,0,207,0,0,0,117,0,105,0,106,0,186,0,168,0,134,0,0,0,68,0,78,0,7,0,181,0,239,0,218,0,228,0,150,0,52,0,246,0,0,0,0,0,86,0,125,0,251,0,151,0,22,0,96,0,151,0,225,0,186,0,112,0,225,0,38,0,111,0,193,0,128,0,80,0,0,0,127,0,54,0,0,0,149,0,4,0,0,0,200,0,85,0,0,0,0,0,103,0,4,0,47,0,60,0,242,0,213,0,181,0,210,0,19,0,54,0,155,0,180,0,246,0,42,0,69,0,69,0,80,0,172,0,35,0,205,0,26,0,157,0,194,0,80,0,217,0,0,0,230,0,38,0,54,0,237,0,246,0,146,0,207,0,145,0,139,0,37,0,64,0);
signal scenario_full  : scenario_type := (147,31,147,30,147,29,50,31,194,31,157,31,157,30,117,31,243,31,249,31,249,30,9,31,9,30,55,31,55,30,51,31,164,31,173,31,183,31,116,31,94,31,94,30,70,31,185,31,45,31,168,31,101,31,10,31,146,31,121,31,121,30,27,31,196,31,44,31,88,31,134,31,84,31,63,31,39,31,123,31,224,31,101,31,237,31,237,30,159,31,218,31,218,30,137,31,180,31,198,31,198,30,185,31,139,31,222,31,100,31,100,30,131,31,56,31,56,30,120,31,166,31,6,31,218,31,244,31,154,31,224,31,137,31,184,31,158,31,137,31,16,31,79,31,40,31,253,31,62,31,62,30,62,29,26,31,176,31,251,31,20,31,248,31,158,31,56,31,56,30,56,29,49,31,189,31,189,30,141,31,168,31,131,31,106,31,106,30,177,31,91,31,230,31,131,31,129,31,200,31,31,31,230,31,223,31,80,31,236,31,236,30,236,29,36,31,176,31,216,31,254,31,190,31,190,30,132,31,218,31,218,30,218,29,107,31,115,31,91,31,24,31,15,31,146,31,97,31,180,31,180,30,147,31,147,30,111,31,176,31,169,31,53,31,130,31,1,31,30,31,37,31,233,31,219,31,192,31,68,31,36,31,139,31,87,31,57,31,119,31,229,31,139,31,179,31,245,31,245,30,131,31,185,31,76,31,52,31,137,31,116,31,5,31,56,31,200,31,106,31,139,31,238,31,43,31,216,31,143,31,117,31,117,30,13,31,13,30,121,31,68,31,68,30,172,31,8,31,198,31,184,31,230,31,62,31,14,31,222,31,102,31,46,31,34,31,27,31,27,30,175,31,159,31,236,31,115,31,104,31,239,31,168,31,6,31,203,31,66,31,66,30,66,29,66,28,66,27,66,26,66,25,94,31,92,31,129,31,88,31,88,30,14,31,20,31,178,31,248,31,37,31,37,30,40,31,134,31,68,31,96,31,60,31,85,31,190,31,226,31,226,30,104,31,157,31,50,31,248,31,250,31,166,31,162,31,162,30,221,31,206,31,215,31,121,31,238,31,123,31,4,31,4,30,229,31,28,31,39,31,20,31,20,30,20,29,67,31,69,31,143,31,143,30,48,31,121,31,121,30,121,29,78,31,78,30,44,31,93,31,40,31,127,31,144,31,22,31,218,31,218,30,162,31,249,31,253,31,253,30,161,31,116,31,181,31,38,31,38,30,134,31,88,31,74,31,1,31,1,30,217,31,217,30,43,31,43,30,136,31,181,31,48,31,169,31,90,31,38,31,193,31,154,31,242,31,242,30,49,31,165,31,220,31,220,30,220,29,40,31,8,31,109,31,26,31,189,31,223,31,110,31,196,31,196,30,109,31,236,31,236,30,236,29,71,31,182,31,191,31,201,31,68,31,68,30,130,31,210,31,171,31,171,30,175,31,175,30,120,31,169,31,203,31,4,31,244,31,187,31,72,31,160,31,231,31,147,31,52,31,115,31,113,31,8,31,193,31,189,31,119,31,11,31,102,31,102,30,77,31,224,31,180,31,182,31,182,30,15,31,245,31,113,31,164,31,214,31,133,31,107,31,103,31,103,30,103,29,122,31,122,30,41,31,190,31,34,31,229,31,229,30,173,31,83,31,20,31,97,31,33,31,33,30,62,31,62,30,62,29,62,28,148,31,26,31,149,31,60,31,32,31,1,31,73,31,208,31,72,31,76,31,76,30,76,29,76,28,47,31,205,31,205,30,133,31,214,31,214,30,104,31,9,31,98,31,98,30,220,31,118,31,118,30,7,31,239,31,244,31,244,30,75,31,111,31,185,31,3,31,17,31,73,31,73,30,92,31,79,31,159,31,159,30,215,31,2,31,46,31,95,31,95,30,111,31,151,31,153,31,29,31,90,31,202,31,202,30,15,31,117,31,177,31,39,31,83,31,56,31,41,31,2,31,17,31,173,31,194,31,224,31,13,31,194,31,156,31,232,31,221,31,34,31,34,30,161,31,174,31,174,30,174,29,174,28,183,31,244,31,34,31,93,31,242,31,144,31,144,30,174,31,78,31,168,31,83,31,15,31,242,31,128,31,157,31,157,30,84,31,182,31,232,31,232,30,68,31,142,31,142,30,66,31,8,31,8,30,127,31,116,31,15,31,173,31,174,31,174,30,174,29,16,31,233,31,86,31,165,31,165,30,36,31,36,30,166,31,127,31,71,31,71,30,216,31,25,31,110,31,110,30,110,29,136,31,188,31,148,31,103,31,225,31,27,31,149,31,149,30,186,31,254,31,237,31,252,31,112,31,112,30,205,31,96,31,43,31,43,30,55,31,65,31,183,31,248,31,79,31,236,31,134,31,55,31,153,31,162,31,150,31,150,30,212,31,240,31,234,31,139,31,58,31,218,31,84,31,84,30,84,29,84,28,178,31,19,31,221,31,128,31,148,31,148,30,217,31,227,31,86,31,22,31,194,31,132,31,148,31,106,31,212,31,92,31,98,31,144,31,221,31,176,31,176,30,226,31,124,31,50,31,245,31,52,31,206,31,126,31,126,30,236,31,157,31,157,30,245,31,142,31,124,31,147,31,242,31,41,31,41,30,84,31,98,31,147,31,126,31,82,31,119,31,46,31,161,31,71,31,146,31,146,30,4,31,201,31,201,30,201,29,251,31,157,31,161,31,113,31,134,31,134,30,200,31,31,31,31,30,18,31,14,31,214,31,36,31,125,31,4,31,4,30,4,29,247,31,75,31,199,31,48,31,203,31,102,31,173,31,58,31,68,31,182,31,35,31,40,31,58,31,11,31,220,31,4,31,223,31,34,31,34,30,105,31,149,31,149,30,200,31,158,31,185,31,18,31,141,31,49,31,129,31,221,31,221,30,244,31,25,31,73,31,73,30,94,31,105,31,13,31,30,31,144,31,109,31,115,31,218,31,204,31,69,31,197,31,55,31,185,31,87,31,87,30,41,31,120,31,53,31,134,31,163,31,162,31,201,31,247,31,247,30,239,31,197,31,158,31,95,31,148,31,207,31,206,31,209,31,47,31,184,31,89,31,9,31,248,31,233,31,162,31,49,31,214,31,214,30,214,29,211,31,184,31,235,31,105,31,239,31,85,31,203,31,238,31,7,31,228,31,228,30,87,31,158,31,230,31,173,31,173,30,185,31,5,31,5,30,5,29,193,31,90,31,90,30,158,31,233,31,179,31,94,31,94,30,45,31,46,31,64,31,236,31,253,31,153,31,133,31,56,31,203,31,51,31,70,31,227,31,227,30,207,31,207,30,117,31,105,31,106,31,186,31,168,31,134,31,134,30,68,31,78,31,7,31,181,31,239,31,218,31,228,31,150,31,52,31,246,31,246,30,246,29,86,31,125,31,251,31,151,31,22,31,96,31,151,31,225,31,186,31,112,31,225,31,38,31,111,31,193,31,128,31,80,31,80,30,127,31,54,31,54,30,149,31,4,31,4,30,200,31,85,31,85,30,85,29,103,31,4,31,47,31,60,31,242,31,213,31,181,31,210,31,19,31,54,31,155,31,180,31,246,31,42,31,69,31,69,31,80,31,172,31,35,31,205,31,26,31,157,31,194,31,80,31,217,31,217,30,230,31,38,31,54,31,237,31,246,31,146,31,207,31,145,31,139,31,37,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
