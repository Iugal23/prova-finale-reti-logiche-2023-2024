-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 968;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,87,0,0,0,172,0,237,0,94,0,51,0,0,0,187,0,0,0,130,0,0,0,59,0,8,0,0,0,48,0,0,0,145,0,191,0,189,0,240,0,71,0,155,0,217,0,55,0,183,0,0,0,0,0,133,0,0,0,173,0,12,0,67,0,52,0,138,0,231,0,92,0,74,0,242,0,158,0,180,0,73,0,77,0,62,0,61,0,109,0,32,0,40,0,175,0,206,0,219,0,0,0,82,0,62,0,232,0,93,0,215,0,76,0,68,0,239,0,5,0,179,0,0,0,201,0,174,0,77,0,124,0,71,0,67,0,165,0,0,0,0,0,0,0,198,0,0,0,40,0,0,0,141,0,0,0,208,0,0,0,37,0,0,0,63,0,52,0,121,0,105,0,208,0,96,0,107,0,23,0,0,0,0,0,234,0,33,0,77,0,223,0,0,0,176,0,255,0,209,0,182,0,57,0,98,0,190,0,81,0,120,0,112,0,203,0,0,0,246,0,241,0,236,0,183,0,212,0,27,0,33,0,95,0,168,0,222,0,0,0,240,0,0,0,0,0,0,0,143,0,0,0,52,0,193,0,35,0,17,0,15,0,219,0,219,0,139,0,125,0,12,0,0,0,35,0,0,0,112,0,78,0,99,0,119,0,241,0,75,0,110,0,129,0,194,0,219,0,85,0,80,0,252,0,0,0,0,0,0,0,46,0,24,0,172,0,184,0,7,0,71,0,0,0,62,0,176,0,206,0,195,0,109,0,236,0,2,0,83,0,59,0,32,0,0,0,131,0,62,0,47,0,181,0,119,0,159,0,0,0,157,0,0,0,0,0,188,0,0,0,127,0,208,0,1,0,72,0,16,0,151,0,247,0,242,0,134,0,189,0,0,0,179,0,143,0,0,0,153,0,8,0,235,0,0,0,0,0,0,0,99,0,137,0,233,0,183,0,2,0,69,0,234,0,0,0,110,0,9,0,19,0,33,0,112,0,122,0,30,0,107,0,247,0,86,0,6,0,129,0,44,0,177,0,0,0,180,0,255,0,58,0,101,0,133,0,18,0,206,0,127,0,0,0,109,0,0,0,187,0,231,0,248,0,246,0,196,0,0,0,0,0,181,0,39,0,167,0,147,0,159,0,0,0,54,0,154,0,2,0,0,0,195,0,0,0,0,0,214,0,82,0,17,0,97,0,21,0,125,0,196,0,104,0,135,0,30,0,0,0,127,0,179,0,0,0,238,0,0,0,0,0,36,0,98,0,0,0,21,0,83,0,185,0,230,0,209,0,196,0,180,0,90,0,138,0,205,0,139,0,46,0,0,0,0,0,48,0,15,0,227,0,16,0,58,0,0,0,123,0,0,0,79,0,123,0,0,0,61,0,222,0,0,0,253,0,0,0,32,0,0,0,77,0,43,0,3,0,166,0,151,0,179,0,0,0,54,0,90,0,93,0,0,0,187,0,0,0,0,0,0,0,0,0,0,0,165,0,246,0,0,0,148,0,198,0,155,0,0,0,253,0,112,0,0,0,23,0,20,0,0,0,196,0,85,0,230,0,131,0,0,0,6,0,59,0,96,0,0,0,248,0,220,0,0,0,123,0,254,0,9,0,225,0,34,0,182,0,160,0,16,0,215,0,104,0,0,0,184,0,203,0,0,0,0,0,0,0,112,0,68,0,0,0,0,0,146,0,102,0,135,0,212,0,253,0,122,0,102,0,58,0,247,0,112,0,217,0,0,0,205,0,74,0,20,0,141,0,219,0,79,0,0,0,77,0,114,0,147,0,0,0,0,0,42,0,135,0,178,0,141,0,244,0,90,0,151,0,21,0,59,0,51,0,118,0,155,0,193,0,193,0,30,0,0,0,118,0,110,0,0,0,0,0,177,0,0,0,0,0,129,0,100,0,236,0,45,0,53,0,181,0,118,0,0,0,59,0,65,0,94,0,243,0,29,0,132,0,138,0,250,0,0,0,176,0,60,0,244,0,67,0,0,0,194,0,246,0,109,0,71,0,164,0,0,0,105,0,0,0,17,0,180,0,50,0,145,0,187,0,179,0,122,0,126,0,233,0,112,0,189,0,0,0,75,0,140,0,0,0,21,0,211,0,31,0,185,0,200,0,128,0,0,0,5,0,245,0,0,0,199,0,163,0,40,0,174,0,106,0,215,0,251,0,19,0,67,0,0,0,57,0,184,0,187,0,64,0,77,0,170,0,247,0,98,0,233,0,0,0,0,0,198,0,198,0,0,0,29,0,238,0,41,0,174,0,54,0,248,0,113,0,46,0,0,0,236,0,81,0,90,0,255,0,63,0,118,0,70,0,0,0,125,0,182,0,153,0,244,0,203,0,44,0,0,0,214,0,0,0,41,0,216,0,151,0,5,0,23,0,228,0,245,0,66,0,0,0,0,0,208,0,218,0,239,0,101,0,0,0,0,0,7,0,179,0,0,0,139,0,18,0,0,0,34,0,252,0,220,0,29,0,0,0,0,0,0,0,125,0,61,0,62,0,31,0,111,0,31,0,224,0,215,0,40,0,0,0,141,0,37,0,132,0,0,0,246,0,213,0,95,0,0,0,155,0,8,0,90,0,69,0,0,0,46,0,0,0,210,0,80,0,131,0,149,0,223,0,82,0,233,0,143,0,232,0,171,0,96,0,216,0,62,0,92,0,121,0,126,0,98,0,35,0,251,0,228,0,23,0,234,0,200,0,179,0,213,0,146,0,0,0,166,0,90,0,238,0,215,0,13,0,0,0,196,0,245,0,0,0,210,0,97,0,121,0,0,0,0,0,218,0,38,0,211,0,190,0,205,0,236,0,123,0,11,0,0,0,53,0,153,0,83,0,28,0,66,0,16,0,104,0,0,0,96,0,3,0,132,0,0,0,67,0,245,0,70,0,200,0,0,0,31,0,151,0,0,0,192,0,216,0,0,0,0,0,52,0,27,0,61,0,0,0,42,0,131,0,0,0,232,0,61,0,0,0,0,0,58,0,0,0,168,0,0,0,54,0,226,0,153,0,193,0,54,0,107,0,0,0,205,0,240,0,231,0,130,0,113,0,98,0,224,0,7,0,219,0,202,0,58,0,0,0,206,0,105,0,232,0,219,0,240,0,22,0,117,0,0,0,85,0,99,0,60,0,248,0,0,0,0,0,201,0,177,0,0,0,217,0,0,0,15,0,53,0,182,0,239,0,29,0,0,0,225,0,91,0,72,0,71,0,187,0,13,0,97,0,65,0,55,0,200,0,76,0,201,0,6,0,0,0,46,0,96,0,51,0,118,0,174,0,136,0,0,0,243,0,201,0,198,0,124,0,0,0,181,0,221,0,52,0,138,0,0,0,0,0,227,0,119,0,0,0,209,0,42,0,0,0,252,0,219,0,0,0,48,0,21,0,71,0,130,0,97,0,0,0,114,0,243,0,0,0,0,0,137,0,153,0,0,0,195,0,0,0,5,0,33,0,38,0,0,0,78,0,0,0,41,0,114,0,0,0,154,0,17,0,37,0,0,0,133,0,208,0,0,0,27,0,219,0,85,0,185,0,83,0,255,0,83,0,229,0,0,0,0,0,221,0,250,0,0,0,169,0,0,0,86,0,0,0,155,0,127,0,156,0,182,0,177,0,181,0,109,0,0,0,108,0,223,0,244,0,71,0,0,0,199,0,0,0,95,0,0,0,96,0,0,0,63,0,111,0,0,0,241,0,251,0,8,0,155,0,58,0,193,0,43,0,229,0,116,0,0,0,46,0,187,0,0,0,135,0,5,0,194,0,129,0,25,0,194,0,157,0,244,0,98,0,102,0,141,0,155,0,194,0,135,0,246,0,14,0,70,0,0,0,201,0,43,0,23,0,125,0,164,0,228,0,231,0,122,0,243,0,251,0,135,0,0,0,0,0,204,0,227,0,149,0,1,0,115,0,39,0,216,0,0,0,23,0,182,0,0,0,68,0,197,0,2,0,0,0,251,0,0,0,0,0,177,0,155,0,1,0,245,0,125,0,33,0,44,0,78,0,190,0,187,0,205,0,146,0,28,0,181,0,165,0,180,0,5,0,48,0,84,0,35,0,194,0,148,0,0,0,204,0,228,0,194,0,190,0,121,0,0,0,59,0,28,0,131,0,240,0,82,0,136,0,0,0,227,0,131,0,96,0,51,0,39,0,100,0,106,0,177,0,85,0,241,0,99,0,220,0,80,0,0,0,152,0,0,0,115,0,0,0,106,0,0,0,251,0,44,0,0,0,153,0,89,0,0,0,37,0,25,0,220,0,0,0,221,0,0,0,18,0,17,0,212,0,198,0,0,0,247,0,214,0,157,0,17,0,0,0,31,0,217,0,80,0,23,0);
signal scenario_full  : scenario_type := (0,0,87,31,87,30,172,31,237,31,94,31,51,31,51,30,187,31,187,30,130,31,130,30,59,31,8,31,8,30,48,31,48,30,145,31,191,31,189,31,240,31,71,31,155,31,217,31,55,31,183,31,183,30,183,29,133,31,133,30,173,31,12,31,67,31,52,31,138,31,231,31,92,31,74,31,242,31,158,31,180,31,73,31,77,31,62,31,61,31,109,31,32,31,40,31,175,31,206,31,219,31,219,30,82,31,62,31,232,31,93,31,215,31,76,31,68,31,239,31,5,31,179,31,179,30,201,31,174,31,77,31,124,31,71,31,67,31,165,31,165,30,165,29,165,28,198,31,198,30,40,31,40,30,141,31,141,30,208,31,208,30,37,31,37,30,63,31,52,31,121,31,105,31,208,31,96,31,107,31,23,31,23,30,23,29,234,31,33,31,77,31,223,31,223,30,176,31,255,31,209,31,182,31,57,31,98,31,190,31,81,31,120,31,112,31,203,31,203,30,246,31,241,31,236,31,183,31,212,31,27,31,33,31,95,31,168,31,222,31,222,30,240,31,240,30,240,29,240,28,143,31,143,30,52,31,193,31,35,31,17,31,15,31,219,31,219,31,139,31,125,31,12,31,12,30,35,31,35,30,112,31,78,31,99,31,119,31,241,31,75,31,110,31,129,31,194,31,219,31,85,31,80,31,252,31,252,30,252,29,252,28,46,31,24,31,172,31,184,31,7,31,71,31,71,30,62,31,176,31,206,31,195,31,109,31,236,31,2,31,83,31,59,31,32,31,32,30,131,31,62,31,47,31,181,31,119,31,159,31,159,30,157,31,157,30,157,29,188,31,188,30,127,31,208,31,1,31,72,31,16,31,151,31,247,31,242,31,134,31,189,31,189,30,179,31,143,31,143,30,153,31,8,31,235,31,235,30,235,29,235,28,99,31,137,31,233,31,183,31,2,31,69,31,234,31,234,30,110,31,9,31,19,31,33,31,112,31,122,31,30,31,107,31,247,31,86,31,6,31,129,31,44,31,177,31,177,30,180,31,255,31,58,31,101,31,133,31,18,31,206,31,127,31,127,30,109,31,109,30,187,31,231,31,248,31,246,31,196,31,196,30,196,29,181,31,39,31,167,31,147,31,159,31,159,30,54,31,154,31,2,31,2,30,195,31,195,30,195,29,214,31,82,31,17,31,97,31,21,31,125,31,196,31,104,31,135,31,30,31,30,30,127,31,179,31,179,30,238,31,238,30,238,29,36,31,98,31,98,30,21,31,83,31,185,31,230,31,209,31,196,31,180,31,90,31,138,31,205,31,139,31,46,31,46,30,46,29,48,31,15,31,227,31,16,31,58,31,58,30,123,31,123,30,79,31,123,31,123,30,61,31,222,31,222,30,253,31,253,30,32,31,32,30,77,31,43,31,3,31,166,31,151,31,179,31,179,30,54,31,90,31,93,31,93,30,187,31,187,30,187,29,187,28,187,27,187,26,165,31,246,31,246,30,148,31,198,31,155,31,155,30,253,31,112,31,112,30,23,31,20,31,20,30,196,31,85,31,230,31,131,31,131,30,6,31,59,31,96,31,96,30,248,31,220,31,220,30,123,31,254,31,9,31,225,31,34,31,182,31,160,31,16,31,215,31,104,31,104,30,184,31,203,31,203,30,203,29,203,28,112,31,68,31,68,30,68,29,146,31,102,31,135,31,212,31,253,31,122,31,102,31,58,31,247,31,112,31,217,31,217,30,205,31,74,31,20,31,141,31,219,31,79,31,79,30,77,31,114,31,147,31,147,30,147,29,42,31,135,31,178,31,141,31,244,31,90,31,151,31,21,31,59,31,51,31,118,31,155,31,193,31,193,31,30,31,30,30,118,31,110,31,110,30,110,29,177,31,177,30,177,29,129,31,100,31,236,31,45,31,53,31,181,31,118,31,118,30,59,31,65,31,94,31,243,31,29,31,132,31,138,31,250,31,250,30,176,31,60,31,244,31,67,31,67,30,194,31,246,31,109,31,71,31,164,31,164,30,105,31,105,30,17,31,180,31,50,31,145,31,187,31,179,31,122,31,126,31,233,31,112,31,189,31,189,30,75,31,140,31,140,30,21,31,211,31,31,31,185,31,200,31,128,31,128,30,5,31,245,31,245,30,199,31,163,31,40,31,174,31,106,31,215,31,251,31,19,31,67,31,67,30,57,31,184,31,187,31,64,31,77,31,170,31,247,31,98,31,233,31,233,30,233,29,198,31,198,31,198,30,29,31,238,31,41,31,174,31,54,31,248,31,113,31,46,31,46,30,236,31,81,31,90,31,255,31,63,31,118,31,70,31,70,30,125,31,182,31,153,31,244,31,203,31,44,31,44,30,214,31,214,30,41,31,216,31,151,31,5,31,23,31,228,31,245,31,66,31,66,30,66,29,208,31,218,31,239,31,101,31,101,30,101,29,7,31,179,31,179,30,139,31,18,31,18,30,34,31,252,31,220,31,29,31,29,30,29,29,29,28,125,31,61,31,62,31,31,31,111,31,31,31,224,31,215,31,40,31,40,30,141,31,37,31,132,31,132,30,246,31,213,31,95,31,95,30,155,31,8,31,90,31,69,31,69,30,46,31,46,30,210,31,80,31,131,31,149,31,223,31,82,31,233,31,143,31,232,31,171,31,96,31,216,31,62,31,92,31,121,31,126,31,98,31,35,31,251,31,228,31,23,31,234,31,200,31,179,31,213,31,146,31,146,30,166,31,90,31,238,31,215,31,13,31,13,30,196,31,245,31,245,30,210,31,97,31,121,31,121,30,121,29,218,31,38,31,211,31,190,31,205,31,236,31,123,31,11,31,11,30,53,31,153,31,83,31,28,31,66,31,16,31,104,31,104,30,96,31,3,31,132,31,132,30,67,31,245,31,70,31,200,31,200,30,31,31,151,31,151,30,192,31,216,31,216,30,216,29,52,31,27,31,61,31,61,30,42,31,131,31,131,30,232,31,61,31,61,30,61,29,58,31,58,30,168,31,168,30,54,31,226,31,153,31,193,31,54,31,107,31,107,30,205,31,240,31,231,31,130,31,113,31,98,31,224,31,7,31,219,31,202,31,58,31,58,30,206,31,105,31,232,31,219,31,240,31,22,31,117,31,117,30,85,31,99,31,60,31,248,31,248,30,248,29,201,31,177,31,177,30,217,31,217,30,15,31,53,31,182,31,239,31,29,31,29,30,225,31,91,31,72,31,71,31,187,31,13,31,97,31,65,31,55,31,200,31,76,31,201,31,6,31,6,30,46,31,96,31,51,31,118,31,174,31,136,31,136,30,243,31,201,31,198,31,124,31,124,30,181,31,221,31,52,31,138,31,138,30,138,29,227,31,119,31,119,30,209,31,42,31,42,30,252,31,219,31,219,30,48,31,21,31,71,31,130,31,97,31,97,30,114,31,243,31,243,30,243,29,137,31,153,31,153,30,195,31,195,30,5,31,33,31,38,31,38,30,78,31,78,30,41,31,114,31,114,30,154,31,17,31,37,31,37,30,133,31,208,31,208,30,27,31,219,31,85,31,185,31,83,31,255,31,83,31,229,31,229,30,229,29,221,31,250,31,250,30,169,31,169,30,86,31,86,30,155,31,127,31,156,31,182,31,177,31,181,31,109,31,109,30,108,31,223,31,244,31,71,31,71,30,199,31,199,30,95,31,95,30,96,31,96,30,63,31,111,31,111,30,241,31,251,31,8,31,155,31,58,31,193,31,43,31,229,31,116,31,116,30,46,31,187,31,187,30,135,31,5,31,194,31,129,31,25,31,194,31,157,31,244,31,98,31,102,31,141,31,155,31,194,31,135,31,246,31,14,31,70,31,70,30,201,31,43,31,23,31,125,31,164,31,228,31,231,31,122,31,243,31,251,31,135,31,135,30,135,29,204,31,227,31,149,31,1,31,115,31,39,31,216,31,216,30,23,31,182,31,182,30,68,31,197,31,2,31,2,30,251,31,251,30,251,29,177,31,155,31,1,31,245,31,125,31,33,31,44,31,78,31,190,31,187,31,205,31,146,31,28,31,181,31,165,31,180,31,5,31,48,31,84,31,35,31,194,31,148,31,148,30,204,31,228,31,194,31,190,31,121,31,121,30,59,31,28,31,131,31,240,31,82,31,136,31,136,30,227,31,131,31,96,31,51,31,39,31,100,31,106,31,177,31,85,31,241,31,99,31,220,31,80,31,80,30,152,31,152,30,115,31,115,30,106,31,106,30,251,31,44,31,44,30,153,31,89,31,89,30,37,31,25,31,220,31,220,30,221,31,221,30,18,31,17,31,212,31,198,31,198,30,247,31,214,31,157,31,17,31,17,30,31,31,217,31,80,31,23,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
