-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 955;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (115,0,199,0,0,0,77,0,0,0,0,0,204,0,14,0,44,0,159,0,48,0,42,0,159,0,233,0,193,0,243,0,164,0,181,0,228,0,170,0,82,0,171,0,207,0,136,0,0,0,120,0,178,0,149,0,203,0,171,0,250,0,66,0,0,0,176,0,163,0,7,0,198,0,5,0,83,0,122,0,24,0,7,0,55,0,18,0,186,0,97,0,24,0,0,0,147,0,27,0,143,0,64,0,0,0,167,0,196,0,119,0,0,0,113,0,134,0,8,0,0,0,0,0,81,0,194,0,49,0,194,0,83,0,145,0,0,0,184,0,19,0,84,0,0,0,0,0,212,0,249,0,0,0,0,0,0,0,94,0,24,0,0,0,132,0,168,0,0,0,0,0,36,0,0,0,0,0,0,0,208,0,0,0,92,0,81,0,204,0,207,0,248,0,11,0,223,0,81,0,84,0,18,0,63,0,133,0,250,0,82,0,82,0,8,0,20,0,232,0,55,0,80,0,101,0,10,0,0,0,221,0,31,0,178,0,147,0,132,0,183,0,92,0,0,0,196,0,86,0,0,0,204,0,92,0,116,0,94,0,246,0,76,0,48,0,90,0,89,0,0,0,0,0,81,0,235,0,98,0,0,0,36,0,65,0,170,0,129,0,218,0,67,0,242,0,203,0,255,0,191,0,159,0,42,0,221,0,30,0,250,0,49,0,199,0,130,0,0,0,101,0,148,0,0,0,24,0,226,0,79,0,86,0,242,0,150,0,247,0,0,0,0,0,84,0,161,0,184,0,209,0,0,0,106,0,0,0,0,0,175,0,235,0,127,0,0,0,199,0,32,0,0,0,64,0,13,0,142,0,71,0,76,0,27,0,206,0,191,0,48,0,0,0,134,0,0,0,53,0,159,0,32,0,151,0,109,0,23,0,0,0,135,0,231,0,0,0,10,0,198,0,0,0,0,0,12,0,217,0,0,0,77,0,69,0,196,0,89,0,129,0,227,0,211,0,33,0,87,0,51,0,0,0,246,0,121,0,72,0,249,0,250,0,198,0,46,0,0,0,62,0,0,0,0,0,233,0,239,0,116,0,13,0,99,0,162,0,0,0,0,0,226,0,64,0,62,0,160,0,0,0,0,0,131,0,248,0,169,0,72,0,49,0,7,0,108,0,25,0,178,0,244,0,36,0,0,0,125,0,58,0,88,0,0,0,210,0,84,0,101,0,105,0,0,0,82,0,41,0,6,0,191,0,95,0,0,0,0,0,0,0,27,0,155,0,0,0,0,0,52,0,180,0,207,0,92,0,195,0,226,0,0,0,215,0,13,0,68,0,244,0,8,0,221,0,0,0,198,0,45,0,218,0,0,0,0,0,61,0,187,0,178,0,230,0,0,0,45,0,35,0,115,0,43,0,48,0,246,0,215,0,13,0,0,0,96,0,0,0,57,0,52,0,30,0,234,0,146,0,0,0,155,0,174,0,80,0,11,0,170,0,93,0,91,0,57,0,0,0,237,0,153,0,235,0,57,0,2,0,91,0,58,0,56,0,208,0,96,0,176,0,169,0,96,0,251,0,169,0,201,0,119,0,252,0,200,0,1,0,6,0,156,0,217,0,63,0,0,0,46,0,125,0,0,0,88,0,81,0,195,0,187,0,183,0,88,0,0,0,0,0,253,0,106,0,9,0,132,0,56,0,220,0,115,0,33,0,153,0,2,0,174,0,87,0,155,0,215,0,110,0,60,0,0,0,30,0,233,0,25,0,47,0,87,0,218,0,251,0,253,0,248,0,204,0,241,0,167,0,0,0,98,0,173,0,0,0,197,0,140,0,0,0,0,0,62,0,36,0,88,0,213,0,17,0,5,0,204,0,119,0,195,0,0,0,102,0,19,0,0,0,149,0,111,0,131,0,167,0,5,0,232,0,153,0,97,0,171,0,169,0,0,0,2,0,220,0,134,0,39,0,140,0,0,0,15,0,19,0,0,0,88,0,125,0,251,0,106,0,220,0,0,0,188,0,180,0,178,0,1,0,0,0,96,0,98,0,0,0,235,0,36,0,204,0,57,0,95,0,33,0,0,0,233,0,0,0,0,0,174,0,0,0,84,0,217,0,138,0,0,0,35,0,0,0,141,0,137,0,143,0,129,0,63,0,150,0,0,0,0,0,0,0,158,0,211,0,92,0,51,0,227,0,0,0,161,0,251,0,207,0,157,0,0,0,0,0,0,0,0,0,36,0,205,0,161,0,149,0,118,0,44,0,0,0,0,0,0,0,165,0,223,0,110,0,242,0,0,0,87,0,10,0,59,0,208,0,0,0,228,0,0,0,118,0,0,0,208,0,45,0,0,0,0,0,82,0,141,0,7,0,199,0,0,0,70,0,134,0,125,0,129,0,0,0,8,0,216,0,64,0,84,0,115,0,238,0,38,0,241,0,105,0,182,0,249,0,128,0,0,0,63,0,7,0,0,0,12,0,189,0,24,0,200,0,84,0,74,0,18,0,0,0,225,0,0,0,21,0,67,0,206,0,93,0,136,0,0,0,242,0,196,0,0,0,60,0,42,0,0,0,179,0,95,0,113,0,188,0,0,0,36,0,206,0,0,0,203,0,0,0,0,0,33,0,235,0,202,0,207,0,226,0,195,0,203,0,154,0,29,0,167,0,0,0,0,0,0,0,0,0,251,0,0,0,4,0,131,0,218,0,73,0,253,0,10,0,239,0,63,0,224,0,15,0,0,0,226,0,103,0,161,0,124,0,19,0,244,0,223,0,60,0,0,0,6,0,148,0,140,0,238,0,0,0,189,0,235,0,10,0,0,0,10,0,17,0,0,0,0,0,199,0,174,0,50,0,49,0,57,0,93,0,92,0,2,0,131,0,0,0,99,0,96,0,25,0,67,0,241,0,114,0,140,0,7,0,226,0,0,0,253,0,204,0,126,0,0,0,181,0,99,0,119,0,157,0,6,0,233,0,39,0,49,0,53,0,157,0,246,0,240,0,239,0,39,0,118,0,146,0,0,0,17,0,95,0,228,0,0,0,112,0,153,0,249,0,115,0,161,0,0,0,69,0,118,0,1,0,215,0,103,0,220,0,160,0,0,0,32,0,0,0,219,0,12,0,16,0,116,0,111,0,0,0,0,0,80,0,0,0,25,0,101,0,144,0,21,0,0,0,88,0,113,0,24,0,172,0,191,0,10,0,0,0,211,0,35,0,0,0,81,0,65,0,170,0,10,0,176,0,2,0,34,0,33,0,220,0,100,0,249,0,124,0,138,0,0,0,0,0,3,0,97,0,0,0,0,0,17,0,159,0,150,0,120,0,0,0,53,0,28,0,0,0,220,0,0,0,10,0,227,0,11,0,177,0,193,0,79,0,91,0,214,0,198,0,0,0,0,0,146,0,0,0,104,0,62,0,104,0,11,0,68,0,27,0,172,0,227,0,120,0,0,0,0,0,201,0,50,0,195,0,47,0,0,0,0,0,200,0,0,0,89,0,23,0,23,0,66,0,135,0,183,0,232,0,21,0,204,0,149,0,47,0,125,0,0,0,165,0,242,0,102,0,126,0,0,0,187,0,0,0,0,0,203,0,0,0,245,0,86,0,167,0,107,0,226,0,243,0,238,0,5,0,136,0,224,0,0,0,0,0,13,0,77,0,251,0,204,0,97,0,126,0,99,0,250,0,0,0,101,0,176,0,101,0,97,0,17,0,0,0,0,0,0,0,99,0,0,0,156,0,56,0,37,0,7,0,25,0,73,0,208,0,205,0,249,0,255,0,232,0,85,0,0,0,76,0,0,0,0,0,246,0,141,0,148,0,191,0,0,0,52,0,63,0,67,0,122,0,24,0,151,0,142,0,33,0,13,0,61,0,239,0,32,0,0,0,11,0,8,0,182,0,5,0,53,0,15,0,20,0,40,0,210,0,172,0,177,0,0,0,133,0,216,0,0,0,89,0,133,0,34,0,78,0,100,0,47,0,142,0,2,0,129,0,0,0,44,0,241,0,36,0,0,0,3,0,81,0,99,0,255,0,16,0,129,0,1,0,51,0,0,0,165,0,253,0,202,0,159,0,154,0,162,0,4,0,110,0,0,0,0,0,182,0,60,0,252,0,0,0,0,0,253,0,198,0,5,0,142,0,0,0,234,0,0,0,0,0,146,0,0,0,246,0,250,0,229,0,0,0,0,0,58,0,5,0,0,0,38,0,0,0,0,0,245,0,168,0,0,0,0,0,0,0,0,0,30,0,157,0,169,0,28,0,241,0,0,0,52,0,20,0,8,0,0,0);
signal scenario_full  : scenario_type := (115,31,199,31,199,30,77,31,77,30,77,29,204,31,14,31,44,31,159,31,48,31,42,31,159,31,233,31,193,31,243,31,164,31,181,31,228,31,170,31,82,31,171,31,207,31,136,31,136,30,120,31,178,31,149,31,203,31,171,31,250,31,66,31,66,30,176,31,163,31,7,31,198,31,5,31,83,31,122,31,24,31,7,31,55,31,18,31,186,31,97,31,24,31,24,30,147,31,27,31,143,31,64,31,64,30,167,31,196,31,119,31,119,30,113,31,134,31,8,31,8,30,8,29,81,31,194,31,49,31,194,31,83,31,145,31,145,30,184,31,19,31,84,31,84,30,84,29,212,31,249,31,249,30,249,29,249,28,94,31,24,31,24,30,132,31,168,31,168,30,168,29,36,31,36,30,36,29,36,28,208,31,208,30,92,31,81,31,204,31,207,31,248,31,11,31,223,31,81,31,84,31,18,31,63,31,133,31,250,31,82,31,82,31,8,31,20,31,232,31,55,31,80,31,101,31,10,31,10,30,221,31,31,31,178,31,147,31,132,31,183,31,92,31,92,30,196,31,86,31,86,30,204,31,92,31,116,31,94,31,246,31,76,31,48,31,90,31,89,31,89,30,89,29,81,31,235,31,98,31,98,30,36,31,65,31,170,31,129,31,218,31,67,31,242,31,203,31,255,31,191,31,159,31,42,31,221,31,30,31,250,31,49,31,199,31,130,31,130,30,101,31,148,31,148,30,24,31,226,31,79,31,86,31,242,31,150,31,247,31,247,30,247,29,84,31,161,31,184,31,209,31,209,30,106,31,106,30,106,29,175,31,235,31,127,31,127,30,199,31,32,31,32,30,64,31,13,31,142,31,71,31,76,31,27,31,206,31,191,31,48,31,48,30,134,31,134,30,53,31,159,31,32,31,151,31,109,31,23,31,23,30,135,31,231,31,231,30,10,31,198,31,198,30,198,29,12,31,217,31,217,30,77,31,69,31,196,31,89,31,129,31,227,31,211,31,33,31,87,31,51,31,51,30,246,31,121,31,72,31,249,31,250,31,198,31,46,31,46,30,62,31,62,30,62,29,233,31,239,31,116,31,13,31,99,31,162,31,162,30,162,29,226,31,64,31,62,31,160,31,160,30,160,29,131,31,248,31,169,31,72,31,49,31,7,31,108,31,25,31,178,31,244,31,36,31,36,30,125,31,58,31,88,31,88,30,210,31,84,31,101,31,105,31,105,30,82,31,41,31,6,31,191,31,95,31,95,30,95,29,95,28,27,31,155,31,155,30,155,29,52,31,180,31,207,31,92,31,195,31,226,31,226,30,215,31,13,31,68,31,244,31,8,31,221,31,221,30,198,31,45,31,218,31,218,30,218,29,61,31,187,31,178,31,230,31,230,30,45,31,35,31,115,31,43,31,48,31,246,31,215,31,13,31,13,30,96,31,96,30,57,31,52,31,30,31,234,31,146,31,146,30,155,31,174,31,80,31,11,31,170,31,93,31,91,31,57,31,57,30,237,31,153,31,235,31,57,31,2,31,91,31,58,31,56,31,208,31,96,31,176,31,169,31,96,31,251,31,169,31,201,31,119,31,252,31,200,31,1,31,6,31,156,31,217,31,63,31,63,30,46,31,125,31,125,30,88,31,81,31,195,31,187,31,183,31,88,31,88,30,88,29,253,31,106,31,9,31,132,31,56,31,220,31,115,31,33,31,153,31,2,31,174,31,87,31,155,31,215,31,110,31,60,31,60,30,30,31,233,31,25,31,47,31,87,31,218,31,251,31,253,31,248,31,204,31,241,31,167,31,167,30,98,31,173,31,173,30,197,31,140,31,140,30,140,29,62,31,36,31,88,31,213,31,17,31,5,31,204,31,119,31,195,31,195,30,102,31,19,31,19,30,149,31,111,31,131,31,167,31,5,31,232,31,153,31,97,31,171,31,169,31,169,30,2,31,220,31,134,31,39,31,140,31,140,30,15,31,19,31,19,30,88,31,125,31,251,31,106,31,220,31,220,30,188,31,180,31,178,31,1,31,1,30,96,31,98,31,98,30,235,31,36,31,204,31,57,31,95,31,33,31,33,30,233,31,233,30,233,29,174,31,174,30,84,31,217,31,138,31,138,30,35,31,35,30,141,31,137,31,143,31,129,31,63,31,150,31,150,30,150,29,150,28,158,31,211,31,92,31,51,31,227,31,227,30,161,31,251,31,207,31,157,31,157,30,157,29,157,28,157,27,36,31,205,31,161,31,149,31,118,31,44,31,44,30,44,29,44,28,165,31,223,31,110,31,242,31,242,30,87,31,10,31,59,31,208,31,208,30,228,31,228,30,118,31,118,30,208,31,45,31,45,30,45,29,82,31,141,31,7,31,199,31,199,30,70,31,134,31,125,31,129,31,129,30,8,31,216,31,64,31,84,31,115,31,238,31,38,31,241,31,105,31,182,31,249,31,128,31,128,30,63,31,7,31,7,30,12,31,189,31,24,31,200,31,84,31,74,31,18,31,18,30,225,31,225,30,21,31,67,31,206,31,93,31,136,31,136,30,242,31,196,31,196,30,60,31,42,31,42,30,179,31,95,31,113,31,188,31,188,30,36,31,206,31,206,30,203,31,203,30,203,29,33,31,235,31,202,31,207,31,226,31,195,31,203,31,154,31,29,31,167,31,167,30,167,29,167,28,167,27,251,31,251,30,4,31,131,31,218,31,73,31,253,31,10,31,239,31,63,31,224,31,15,31,15,30,226,31,103,31,161,31,124,31,19,31,244,31,223,31,60,31,60,30,6,31,148,31,140,31,238,31,238,30,189,31,235,31,10,31,10,30,10,31,17,31,17,30,17,29,199,31,174,31,50,31,49,31,57,31,93,31,92,31,2,31,131,31,131,30,99,31,96,31,25,31,67,31,241,31,114,31,140,31,7,31,226,31,226,30,253,31,204,31,126,31,126,30,181,31,99,31,119,31,157,31,6,31,233,31,39,31,49,31,53,31,157,31,246,31,240,31,239,31,39,31,118,31,146,31,146,30,17,31,95,31,228,31,228,30,112,31,153,31,249,31,115,31,161,31,161,30,69,31,118,31,1,31,215,31,103,31,220,31,160,31,160,30,32,31,32,30,219,31,12,31,16,31,116,31,111,31,111,30,111,29,80,31,80,30,25,31,101,31,144,31,21,31,21,30,88,31,113,31,24,31,172,31,191,31,10,31,10,30,211,31,35,31,35,30,81,31,65,31,170,31,10,31,176,31,2,31,34,31,33,31,220,31,100,31,249,31,124,31,138,31,138,30,138,29,3,31,97,31,97,30,97,29,17,31,159,31,150,31,120,31,120,30,53,31,28,31,28,30,220,31,220,30,10,31,227,31,11,31,177,31,193,31,79,31,91,31,214,31,198,31,198,30,198,29,146,31,146,30,104,31,62,31,104,31,11,31,68,31,27,31,172,31,227,31,120,31,120,30,120,29,201,31,50,31,195,31,47,31,47,30,47,29,200,31,200,30,89,31,23,31,23,31,66,31,135,31,183,31,232,31,21,31,204,31,149,31,47,31,125,31,125,30,165,31,242,31,102,31,126,31,126,30,187,31,187,30,187,29,203,31,203,30,245,31,86,31,167,31,107,31,226,31,243,31,238,31,5,31,136,31,224,31,224,30,224,29,13,31,77,31,251,31,204,31,97,31,126,31,99,31,250,31,250,30,101,31,176,31,101,31,97,31,17,31,17,30,17,29,17,28,99,31,99,30,156,31,56,31,37,31,7,31,25,31,73,31,208,31,205,31,249,31,255,31,232,31,85,31,85,30,76,31,76,30,76,29,246,31,141,31,148,31,191,31,191,30,52,31,63,31,67,31,122,31,24,31,151,31,142,31,33,31,13,31,61,31,239,31,32,31,32,30,11,31,8,31,182,31,5,31,53,31,15,31,20,31,40,31,210,31,172,31,177,31,177,30,133,31,216,31,216,30,89,31,133,31,34,31,78,31,100,31,47,31,142,31,2,31,129,31,129,30,44,31,241,31,36,31,36,30,3,31,81,31,99,31,255,31,16,31,129,31,1,31,51,31,51,30,165,31,253,31,202,31,159,31,154,31,162,31,4,31,110,31,110,30,110,29,182,31,60,31,252,31,252,30,252,29,253,31,198,31,5,31,142,31,142,30,234,31,234,30,234,29,146,31,146,30,246,31,250,31,229,31,229,30,229,29,58,31,5,31,5,30,38,31,38,30,38,29,245,31,168,31,168,30,168,29,168,28,168,27,30,31,157,31,169,31,28,31,241,31,241,30,52,31,20,31,8,31,8,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
