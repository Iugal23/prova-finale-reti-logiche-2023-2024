-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_792 is
end project_tb_792;

architecture project_tb_arch_792 of project_tb_792 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 189;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (144,0,129,0,48,0,96,0,176,0,209,0,0,0,224,0,70,0,18,0,124,0,178,0,141,0,63,0,88,0,0,0,1,0,0,0,102,0,110,0,80,0,171,0,131,0,0,0,0,0,1,0,254,0,0,0,31,0,108,0,0,0,100,0,174,0,66,0,178,0,63,0,19,0,0,0,0,0,69,0,173,0,219,0,124,0,146,0,94,0,149,0,0,0,0,0,173,0,0,0,52,0,141,0,193,0,25,0,199,0,27,0,151,0,122,0,220,0,168,0,125,0,227,0,231,0,185,0,107,0,8,0,128,0,187,0,80,0,52,0,232,0,122,0,0,0,0,0,27,0,33,0,0,0,30,0,8,0,250,0,0,0,182,0,10,0,204,0,188,0,233,0,91,0,91,0,224,0,0,0,83,0,50,0,187,0,206,0,230,0,17,0,252,0,182,0,182,0,202,0,210,0,33,0,145,0,51,0,160,0,10,0,206,0,89,0,145,0,105,0,245,0,165,0,231,0,85,0,222,0,0,0,249,0,78,0,103,0,46,0,73,0,81,0,0,0,20,0,233,0,144,0,162,0,0,0,159,0,87,0,154,0,222,0,0,0,158,0,185,0,29,0,133,0,209,0,33,0,0,0,131,0,44,0,34,0,118,0,122,0,0,0,242,0,120,0,0,0,21,0,0,0,144,0,196,0,187,0,33,0,226,0,78,0,95,0,54,0,93,0,61,0,222,0,77,0,46,0,0,0,218,0,128,0,70,0,0,0,40,0,202,0,167,0,217,0,230,0,71,0,229,0,25,0,25,0,77,0,26,0,242,0,178,0,0,0,0,0,0,0,14,0,203,0,164,0,27,0);
signal scenario_full  : scenario_type := (144,31,129,31,48,31,96,31,176,31,209,31,209,30,224,31,70,31,18,31,124,31,178,31,141,31,63,31,88,31,88,30,1,31,1,30,102,31,110,31,80,31,171,31,131,31,131,30,131,29,1,31,254,31,254,30,31,31,108,31,108,30,100,31,174,31,66,31,178,31,63,31,19,31,19,30,19,29,69,31,173,31,219,31,124,31,146,31,94,31,149,31,149,30,149,29,173,31,173,30,52,31,141,31,193,31,25,31,199,31,27,31,151,31,122,31,220,31,168,31,125,31,227,31,231,31,185,31,107,31,8,31,128,31,187,31,80,31,52,31,232,31,122,31,122,30,122,29,27,31,33,31,33,30,30,31,8,31,250,31,250,30,182,31,10,31,204,31,188,31,233,31,91,31,91,31,224,31,224,30,83,31,50,31,187,31,206,31,230,31,17,31,252,31,182,31,182,31,202,31,210,31,33,31,145,31,51,31,160,31,10,31,206,31,89,31,145,31,105,31,245,31,165,31,231,31,85,31,222,31,222,30,249,31,78,31,103,31,46,31,73,31,81,31,81,30,20,31,233,31,144,31,162,31,162,30,159,31,87,31,154,31,222,31,222,30,158,31,185,31,29,31,133,31,209,31,33,31,33,30,131,31,44,31,34,31,118,31,122,31,122,30,242,31,120,31,120,30,21,31,21,30,144,31,196,31,187,31,33,31,226,31,78,31,95,31,54,31,93,31,61,31,222,31,77,31,46,31,46,30,218,31,128,31,70,31,70,30,40,31,202,31,167,31,217,31,230,31,71,31,229,31,25,31,25,31,77,31,26,31,242,31,178,31,178,30,178,29,178,28,14,31,203,31,164,31,27,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
