-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_868 is
end project_tb_868;

architecture project_tb_arch_868 of project_tb_868 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 861;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (205,0,37,0,69,0,79,0,255,0,102,0,0,0,0,0,140,0,199,0,83,0,176,0,12,0,196,0,194,0,42,0,10,0,137,0,166,0,135,0,128,0,0,0,49,0,58,0,81,0,0,0,40,0,0,0,0,0,0,0,153,0,0,0,0,0,0,0,236,0,203,0,54,0,33,0,163,0,19,0,153,0,24,0,0,0,196,0,119,0,45,0,115,0,0,0,216,0,247,0,72,0,107,0,135,0,47,0,255,0,255,0,0,0,125,0,247,0,77,0,0,0,182,0,41,0,245,0,202,0,0,0,121,0,142,0,0,0,147,0,91,0,220,0,204,0,58,0,218,0,52,0,132,0,193,0,0,0,0,0,136,0,86,0,0,0,102,0,0,0,175,0,56,0,211,0,30,0,141,0,123,0,100,0,0,0,253,0,148,0,70,0,171,0,0,0,0,0,0,0,0,0,56,0,22,0,0,0,131,0,97,0,0,0,77,0,0,0,59,0,112,0,212,0,119,0,82,0,153,0,151,0,137,0,200,0,81,0,200,0,167,0,3,0,142,0,199,0,32,0,177,0,154,0,165,0,0,0,172,0,18,0,216,0,0,0,0,0,41,0,19,0,0,0,96,0,221,0,228,0,224,0,0,0,155,0,0,0,122,0,112,0,142,0,255,0,14,0,231,0,237,0,177,0,207,0,220,0,0,0,39,0,99,0,145,0,166,0,203,0,40,0,194,0,226,0,100,0,255,0,0,0,0,0,0,0,104,0,122,0,156,0,7,0,65,0,175,0,0,0,222,0,186,0,15,0,128,0,247,0,0,0,109,0,6,0,247,0,145,0,105,0,7,0,116,0,37,0,94,0,0,0,72,0,241,0,249,0,15,0,20,0,190,0,145,0,193,0,119,0,23,0,167,0,0,0,0,0,96,0,150,0,0,0,0,0,196,0,0,0,0,0,94,0,194,0,0,0,0,0,0,0,48,0,0,0,57,0,147,0,233,0,202,0,114,0,0,0,144,0,207,0,213,0,113,0,132,0,167,0,229,0,52,0,9,0,0,0,173,0,208,0,232,0,0,0,221,0,0,0,160,0,241,0,117,0,0,0,128,0,0,0,164,0,195,0,72,0,0,0,13,0,117,0,0,0,198,0,7,0,244,0,110,0,245,0,50,0,67,0,0,0,186,0,0,0,107,0,201,0,44,0,239,0,0,0,227,0,0,0,197,0,0,0,0,0,0,0,66,0,123,0,0,0,230,0,211,0,190,0,232,0,56,0,45,0,237,0,237,0,29,0,49,0,239,0,27,0,86,0,57,0,80,0,0,0,86,0,0,0,205,0,97,0,0,0,163,0,187,0,155,0,156,0,40,0,84,0,16,0,233,0,148,0,200,0,196,0,23,0,117,0,61,0,16,0,0,0,133,0,157,0,140,0,15,0,0,0,108,0,3,0,211,0,8,0,98,0,36,0,0,0,0,0,125,0,145,0,0,0,220,0,0,0,43,0,98,0,0,0,10,0,193,0,0,0,134,0,241,0,225,0,135,0,13,0,58,0,0,0,4,0,0,0,1,0,183,0,178,0,117,0,0,0,0,0,96,0,163,0,86,0,34,0,67,0,223,0,133,0,233,0,25,0,187,0,7,0,254,0,14,0,55,0,222,0,181,0,122,0,39,0,205,0,0,0,0,0,73,0,0,0,53,0,119,0,43,0,157,0,233,0,107,0,231,0,59,0,12,0,86,0,171,0,0,0,113,0,248,0,180,0,0,0,14,0,41,0,196,0,2,0,14,0,250,0,167,0,27,0,121,0,168,0,209,0,82,0,19,0,246,0,47,0,117,0,0,0,11,0,0,0,96,0,16,0,190,0,0,0,0,0,0,0,247,0,231,0,123,0,238,0,159,0,17,0,47,0,36,0,197,0,146,0,178,0,16,0,0,0,207,0,46,0,146,0,192,0,0,0,239,0,0,0,160,0,0,0,2,0,214,0,165,0,86,0,16,0,248,0,199,0,96,0,7,0,0,0,187,0,62,0,175,0,16,0,96,0,76,0,69,0,63,0,210,0,0,0,88,0,0,0,0,0,116,0,237,0,4,0,166,0,247,0,0,0,74,0,200,0,0,0,182,0,46,0,64,0,162,0,80,0,170,0,0,0,227,0,86,0,236,0,175,0,0,0,184,0,36,0,58,0,190,0,0,0,0,0,0,0,5,0,77,0,234,0,219,0,186,0,160,0,223,0,95,0,0,0,235,0,0,0,11,0,15,0,0,0,0,0,56,0,232,0,135,0,243,0,92,0,0,0,69,0,139,0,0,0,232,0,240,0,125,0,102,0,89,0,0,0,190,0,27,0,11,0,241,0,104,0,0,0,0,0,55,0,64,0,24,0,80,0,254,0,136,0,132,0,103,0,0,0,36,0,165,0,0,0,92,0,171,0,202,0,39,0,154,0,185,0,250,0,38,0,212,0,93,0,52,0,132,0,205,0,216,0,246,0,46,0,120,0,94,0,82,0,0,0,86,0,47,0,72,0,23,0,0,0,238,0,179,0,84,0,139,0,79,0,13,0,130,0,93,0,0,0,0,0,37,0,75,0,214,0,249,0,0,0,122,0,76,0,168,0,53,0,96,0,174,0,211,0,201,0,246,0,27,0,125,0,127,0,235,0,0,0,0,0,250,0,174,0,175,0,0,0,89,0,98,0,0,0,0,0,45,0,47,0,98,0,0,0,148,0,181,0,13,0,111,0,187,0,123,0,233,0,64,0,142,0,0,0,16,0,117,0,60,0,131,0,99,0,122,0,252,0,0,0,80,0,180,0,241,0,120,0,147,0,99,0,32,0,59,0,106,0,0,0,0,0,0,0,0,0,0,0,93,0,71,0,108,0,72,0,143,0,231,0,57,0,143,0,52,0,48,0,41,0,0,0,219,0,19,0,0,0,0,0,237,0,170,0,11,0,0,0,85,0,190,0,39,0,28,0,68,0,234,0,13,0,249,0,17,0,0,0,0,0,0,0,251,0,0,0,25,0,111,0,0,0,106,0,216,0,180,0,67,0,55,0,192,0,33,0,122,0,68,0,140,0,246,0,247,0,0,0,148,0,93,0,12,0,92,0,226,0,74,0,218,0,72,0,106,0,143,0,16,0,0,0,0,0,0,0,101,0,0,0,253,0,163,0,93,0,207,0,172,0,0,0,220,0,0,0,93,0,203,0,76,0,139,0,136,0,137,0,0,0,48,0,71,0,211,0,252,0,78,0,35,0,0,0,0,0,109,0,74,0,116,0,43,0,112,0,20,0,75,0,130,0,0,0,0,0,32,0,36,0,21,0,6,0,13,0,92,0,0,0,165,0,0,0,0,0,81,0,100,0,0,0,0,0,45,0,26,0,0,0,226,0,107,0,97,0,198,0,215,0,197,0,156,0,195,0,35,0,24,0,103,0,212,0,67,0,62,0,140,0,231,0,154,0,0,0,94,0,56,0,226,0,17,0,232,0,62,0,0,0,89,0,38,0,39,0,126,0,124,0,56,0,96,0,206,0,169,0,115,0,103,0,100,0,0,0,148,0,193,0,173,0,0,0,248,0,204,0,154,0,0,0,168,0,86,0,168,0,0,0,2,0,80,0,5,0,0,0,215,0,127,0,15,0,50,0,0,0,170,0,184,0,17,0,86,0,27,0,97,0,121,0,158,0,94,0,119,0,181,0,0,0,95,0,0,0,159,0,0,0,86,0,26,0,56,0,24,0,138,0,201,0,244,0,51,0,225,0,253,0,207,0,211,0,207,0,250,0,31,0,112,0,195,0,0,0,36,0,0,0,235,0,119,0,233,0,0,0,197,0,48,0,244,0,197,0,175,0,0,0,166,0,125,0);
signal scenario_full  : scenario_type := (205,31,37,31,69,31,79,31,255,31,102,31,102,30,102,29,140,31,199,31,83,31,176,31,12,31,196,31,194,31,42,31,10,31,137,31,166,31,135,31,128,31,128,30,49,31,58,31,81,31,81,30,40,31,40,30,40,29,40,28,153,31,153,30,153,29,153,28,236,31,203,31,54,31,33,31,163,31,19,31,153,31,24,31,24,30,196,31,119,31,45,31,115,31,115,30,216,31,247,31,72,31,107,31,135,31,47,31,255,31,255,31,255,30,125,31,247,31,77,31,77,30,182,31,41,31,245,31,202,31,202,30,121,31,142,31,142,30,147,31,91,31,220,31,204,31,58,31,218,31,52,31,132,31,193,31,193,30,193,29,136,31,86,31,86,30,102,31,102,30,175,31,56,31,211,31,30,31,141,31,123,31,100,31,100,30,253,31,148,31,70,31,171,31,171,30,171,29,171,28,171,27,56,31,22,31,22,30,131,31,97,31,97,30,77,31,77,30,59,31,112,31,212,31,119,31,82,31,153,31,151,31,137,31,200,31,81,31,200,31,167,31,3,31,142,31,199,31,32,31,177,31,154,31,165,31,165,30,172,31,18,31,216,31,216,30,216,29,41,31,19,31,19,30,96,31,221,31,228,31,224,31,224,30,155,31,155,30,122,31,112,31,142,31,255,31,14,31,231,31,237,31,177,31,207,31,220,31,220,30,39,31,99,31,145,31,166,31,203,31,40,31,194,31,226,31,100,31,255,31,255,30,255,29,255,28,104,31,122,31,156,31,7,31,65,31,175,31,175,30,222,31,186,31,15,31,128,31,247,31,247,30,109,31,6,31,247,31,145,31,105,31,7,31,116,31,37,31,94,31,94,30,72,31,241,31,249,31,15,31,20,31,190,31,145,31,193,31,119,31,23,31,167,31,167,30,167,29,96,31,150,31,150,30,150,29,196,31,196,30,196,29,94,31,194,31,194,30,194,29,194,28,48,31,48,30,57,31,147,31,233,31,202,31,114,31,114,30,144,31,207,31,213,31,113,31,132,31,167,31,229,31,52,31,9,31,9,30,173,31,208,31,232,31,232,30,221,31,221,30,160,31,241,31,117,31,117,30,128,31,128,30,164,31,195,31,72,31,72,30,13,31,117,31,117,30,198,31,7,31,244,31,110,31,245,31,50,31,67,31,67,30,186,31,186,30,107,31,201,31,44,31,239,31,239,30,227,31,227,30,197,31,197,30,197,29,197,28,66,31,123,31,123,30,230,31,211,31,190,31,232,31,56,31,45,31,237,31,237,31,29,31,49,31,239,31,27,31,86,31,57,31,80,31,80,30,86,31,86,30,205,31,97,31,97,30,163,31,187,31,155,31,156,31,40,31,84,31,16,31,233,31,148,31,200,31,196,31,23,31,117,31,61,31,16,31,16,30,133,31,157,31,140,31,15,31,15,30,108,31,3,31,211,31,8,31,98,31,36,31,36,30,36,29,125,31,145,31,145,30,220,31,220,30,43,31,98,31,98,30,10,31,193,31,193,30,134,31,241,31,225,31,135,31,13,31,58,31,58,30,4,31,4,30,1,31,183,31,178,31,117,31,117,30,117,29,96,31,163,31,86,31,34,31,67,31,223,31,133,31,233,31,25,31,187,31,7,31,254,31,14,31,55,31,222,31,181,31,122,31,39,31,205,31,205,30,205,29,73,31,73,30,53,31,119,31,43,31,157,31,233,31,107,31,231,31,59,31,12,31,86,31,171,31,171,30,113,31,248,31,180,31,180,30,14,31,41,31,196,31,2,31,14,31,250,31,167,31,27,31,121,31,168,31,209,31,82,31,19,31,246,31,47,31,117,31,117,30,11,31,11,30,96,31,16,31,190,31,190,30,190,29,190,28,247,31,231,31,123,31,238,31,159,31,17,31,47,31,36,31,197,31,146,31,178,31,16,31,16,30,207,31,46,31,146,31,192,31,192,30,239,31,239,30,160,31,160,30,2,31,214,31,165,31,86,31,16,31,248,31,199,31,96,31,7,31,7,30,187,31,62,31,175,31,16,31,96,31,76,31,69,31,63,31,210,31,210,30,88,31,88,30,88,29,116,31,237,31,4,31,166,31,247,31,247,30,74,31,200,31,200,30,182,31,46,31,64,31,162,31,80,31,170,31,170,30,227,31,86,31,236,31,175,31,175,30,184,31,36,31,58,31,190,31,190,30,190,29,190,28,5,31,77,31,234,31,219,31,186,31,160,31,223,31,95,31,95,30,235,31,235,30,11,31,15,31,15,30,15,29,56,31,232,31,135,31,243,31,92,31,92,30,69,31,139,31,139,30,232,31,240,31,125,31,102,31,89,31,89,30,190,31,27,31,11,31,241,31,104,31,104,30,104,29,55,31,64,31,24,31,80,31,254,31,136,31,132,31,103,31,103,30,36,31,165,31,165,30,92,31,171,31,202,31,39,31,154,31,185,31,250,31,38,31,212,31,93,31,52,31,132,31,205,31,216,31,246,31,46,31,120,31,94,31,82,31,82,30,86,31,47,31,72,31,23,31,23,30,238,31,179,31,84,31,139,31,79,31,13,31,130,31,93,31,93,30,93,29,37,31,75,31,214,31,249,31,249,30,122,31,76,31,168,31,53,31,96,31,174,31,211,31,201,31,246,31,27,31,125,31,127,31,235,31,235,30,235,29,250,31,174,31,175,31,175,30,89,31,98,31,98,30,98,29,45,31,47,31,98,31,98,30,148,31,181,31,13,31,111,31,187,31,123,31,233,31,64,31,142,31,142,30,16,31,117,31,60,31,131,31,99,31,122,31,252,31,252,30,80,31,180,31,241,31,120,31,147,31,99,31,32,31,59,31,106,31,106,30,106,29,106,28,106,27,106,26,93,31,71,31,108,31,72,31,143,31,231,31,57,31,143,31,52,31,48,31,41,31,41,30,219,31,19,31,19,30,19,29,237,31,170,31,11,31,11,30,85,31,190,31,39,31,28,31,68,31,234,31,13,31,249,31,17,31,17,30,17,29,17,28,251,31,251,30,25,31,111,31,111,30,106,31,216,31,180,31,67,31,55,31,192,31,33,31,122,31,68,31,140,31,246,31,247,31,247,30,148,31,93,31,12,31,92,31,226,31,74,31,218,31,72,31,106,31,143,31,16,31,16,30,16,29,16,28,101,31,101,30,253,31,163,31,93,31,207,31,172,31,172,30,220,31,220,30,93,31,203,31,76,31,139,31,136,31,137,31,137,30,48,31,71,31,211,31,252,31,78,31,35,31,35,30,35,29,109,31,74,31,116,31,43,31,112,31,20,31,75,31,130,31,130,30,130,29,32,31,36,31,21,31,6,31,13,31,92,31,92,30,165,31,165,30,165,29,81,31,100,31,100,30,100,29,45,31,26,31,26,30,226,31,107,31,97,31,198,31,215,31,197,31,156,31,195,31,35,31,24,31,103,31,212,31,67,31,62,31,140,31,231,31,154,31,154,30,94,31,56,31,226,31,17,31,232,31,62,31,62,30,89,31,38,31,39,31,126,31,124,31,56,31,96,31,206,31,169,31,115,31,103,31,100,31,100,30,148,31,193,31,173,31,173,30,248,31,204,31,154,31,154,30,168,31,86,31,168,31,168,30,2,31,80,31,5,31,5,30,215,31,127,31,15,31,50,31,50,30,170,31,184,31,17,31,86,31,27,31,97,31,121,31,158,31,94,31,119,31,181,31,181,30,95,31,95,30,159,31,159,30,86,31,26,31,56,31,24,31,138,31,201,31,244,31,51,31,225,31,253,31,207,31,211,31,207,31,250,31,31,31,112,31,195,31,195,30,36,31,36,30,235,31,119,31,233,31,233,30,197,31,48,31,244,31,197,31,175,31,175,30,166,31,125,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
