-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 458;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (190,0,195,0,119,0,198,0,45,0,57,0,0,0,211,0,185,0,77,0,212,0,249,0,164,0,211,0,0,0,0,0,29,0,149,0,88,0,145,0,5,0,0,0,108,0,134,0,161,0,231,0,0,0,118,0,22,0,106,0,69,0,196,0,62,0,55,0,255,0,158,0,31,0,138,0,227,0,24,0,251,0,44,0,117,0,253,0,185,0,118,0,253,0,9,0,34,0,197,0,86,0,211,0,159,0,121,0,0,0,0,0,0,0,77,0,57,0,0,0,115,0,158,0,224,0,176,0,122,0,207,0,83,0,203,0,148,0,253,0,245,0,225,0,0,0,28,0,0,0,151,0,219,0,220,0,49,0,181,0,140,0,121,0,90,0,78,0,227,0,97,0,70,0,253,0,47,0,222,0,243,0,96,0,178,0,3,0,97,0,243,0,71,0,0,0,137,0,19,0,0,0,0,0,0,0,84,0,0,0,0,0,0,0,18,0,210,0,0,0,47,0,160,0,106,0,0,0,148,0,139,0,39,0,137,0,225,0,60,0,61,0,232,0,58,0,251,0,10,0,0,0,0,0,189,0,120,0,0,0,0,0,184,0,120,0,0,0,0,0,254,0,37,0,0,0,88,0,3,0,3,0,4,0,215,0,238,0,32,0,45,0,0,0,126,0,182,0,0,0,77,0,45,0,75,0,241,0,231,0,200,0,207,0,149,0,213,0,214,0,45,0,56,0,54,0,187,0,142,0,7,0,194,0,0,0,224,0,237,0,211,0,180,0,203,0,0,0,40,0,17,0,0,0,0,0,97,0,43,0,0,0,10,0,112,0,203,0,144,0,0,0,101,0,234,0,112,0,84,0,254,0,0,0,0,0,0,0,207,0,184,0,116,0,204,0,56,0,0,0,168,0,0,0,0,0,245,0,236,0,185,0,13,0,0,0,241,0,0,0,110,0,112,0,45,0,254,0,94,0,247,0,230,0,216,0,80,0,39,0,32,0,136,0,67,0,124,0,34,0,129,0,179,0,36,0,86,0,0,0,17,0,131,0,62,0,200,0,56,0,0,0,0,0,197,0,86,0,133,0,205,0,92,0,100,0,0,0,173,0,167,0,89,0,0,0,103,0,168,0,223,0,108,0,194,0,143,0,0,0,100,0,207,0,167,0,0,0,200,0,143,0,67,0,61,0,0,0,0,0,97,0,23,0,210,0,134,0,0,0,68,0,223,0,47,0,203,0,36,0,105,0,0,0,189,0,116,0,172,0,178,0,239,0,211,0,238,0,0,0,93,0,198,0,77,0,119,0,38,0,173,0,248,0,0,0,203,0,184,0,246,0,121,0,182,0,149,0,235,0,11,0,216,0,247,0,0,0,27,0,0,0,84,0,0,0,171,0,246,0,0,0,182,0,52,0,0,0,96,0,59,0,244,0,252,0,26,0,157,0,27,0,121,0,10,0,0,0,133,0,206,0,232,0,177,0,204,0,0,0,171,0,72,0,117,0,0,0,59,0,0,0,0,0,229,0,0,0,12,0,250,0,0,0,0,0,0,0,117,0,0,0,38,0,224,0,65,0,99,0,122,0,38,0,204,0,0,0,240,0,176,0,0,0,242,0,83,0,223,0,102,0,131,0,172,0,88,0,66,0,174,0,29,0,0,0,161,0,25,0,145,0,11,0,178,0,104,0,84,0,4,0,0,0,1,0,110,0,0,0,70,0,0,0,51,0,78,0,36,0,0,0,0,0,133,0,95,0,0,0,0,0,251,0,166,0,0,0,68,0,195,0,189,0,64,0,0,0,0,0,138,0,211,0,92,0,119,0,0,0,252,0,136,0,45,0,110,0,23,0,113,0,0,0,0,0,245,0,3,0,75,0,209,0,130,0,106,0,32,0,125,0,147,0,0,0,205,0,0,0,217,0,0,0,0,0,155,0,5,0,215,0,164,0,0,0,160,0,26,0,8,0,171,0,0,0,0,0,53,0,80,0,0,0,33,0,105,0,203,0,109,0,156,0,0,0,39,0,252,0,251,0,0,0,92,0,41,0,248,0,173,0,113,0,44,0);
signal scenario_full  : scenario_type := (190,31,195,31,119,31,198,31,45,31,57,31,57,30,211,31,185,31,77,31,212,31,249,31,164,31,211,31,211,30,211,29,29,31,149,31,88,31,145,31,5,31,5,30,108,31,134,31,161,31,231,31,231,30,118,31,22,31,106,31,69,31,196,31,62,31,55,31,255,31,158,31,31,31,138,31,227,31,24,31,251,31,44,31,117,31,253,31,185,31,118,31,253,31,9,31,34,31,197,31,86,31,211,31,159,31,121,31,121,30,121,29,121,28,77,31,57,31,57,30,115,31,158,31,224,31,176,31,122,31,207,31,83,31,203,31,148,31,253,31,245,31,225,31,225,30,28,31,28,30,151,31,219,31,220,31,49,31,181,31,140,31,121,31,90,31,78,31,227,31,97,31,70,31,253,31,47,31,222,31,243,31,96,31,178,31,3,31,97,31,243,31,71,31,71,30,137,31,19,31,19,30,19,29,19,28,84,31,84,30,84,29,84,28,18,31,210,31,210,30,47,31,160,31,106,31,106,30,148,31,139,31,39,31,137,31,225,31,60,31,61,31,232,31,58,31,251,31,10,31,10,30,10,29,189,31,120,31,120,30,120,29,184,31,120,31,120,30,120,29,254,31,37,31,37,30,88,31,3,31,3,31,4,31,215,31,238,31,32,31,45,31,45,30,126,31,182,31,182,30,77,31,45,31,75,31,241,31,231,31,200,31,207,31,149,31,213,31,214,31,45,31,56,31,54,31,187,31,142,31,7,31,194,31,194,30,224,31,237,31,211,31,180,31,203,31,203,30,40,31,17,31,17,30,17,29,97,31,43,31,43,30,10,31,112,31,203,31,144,31,144,30,101,31,234,31,112,31,84,31,254,31,254,30,254,29,254,28,207,31,184,31,116,31,204,31,56,31,56,30,168,31,168,30,168,29,245,31,236,31,185,31,13,31,13,30,241,31,241,30,110,31,112,31,45,31,254,31,94,31,247,31,230,31,216,31,80,31,39,31,32,31,136,31,67,31,124,31,34,31,129,31,179,31,36,31,86,31,86,30,17,31,131,31,62,31,200,31,56,31,56,30,56,29,197,31,86,31,133,31,205,31,92,31,100,31,100,30,173,31,167,31,89,31,89,30,103,31,168,31,223,31,108,31,194,31,143,31,143,30,100,31,207,31,167,31,167,30,200,31,143,31,67,31,61,31,61,30,61,29,97,31,23,31,210,31,134,31,134,30,68,31,223,31,47,31,203,31,36,31,105,31,105,30,189,31,116,31,172,31,178,31,239,31,211,31,238,31,238,30,93,31,198,31,77,31,119,31,38,31,173,31,248,31,248,30,203,31,184,31,246,31,121,31,182,31,149,31,235,31,11,31,216,31,247,31,247,30,27,31,27,30,84,31,84,30,171,31,246,31,246,30,182,31,52,31,52,30,96,31,59,31,244,31,252,31,26,31,157,31,27,31,121,31,10,31,10,30,133,31,206,31,232,31,177,31,204,31,204,30,171,31,72,31,117,31,117,30,59,31,59,30,59,29,229,31,229,30,12,31,250,31,250,30,250,29,250,28,117,31,117,30,38,31,224,31,65,31,99,31,122,31,38,31,204,31,204,30,240,31,176,31,176,30,242,31,83,31,223,31,102,31,131,31,172,31,88,31,66,31,174,31,29,31,29,30,161,31,25,31,145,31,11,31,178,31,104,31,84,31,4,31,4,30,1,31,110,31,110,30,70,31,70,30,51,31,78,31,36,31,36,30,36,29,133,31,95,31,95,30,95,29,251,31,166,31,166,30,68,31,195,31,189,31,64,31,64,30,64,29,138,31,211,31,92,31,119,31,119,30,252,31,136,31,45,31,110,31,23,31,113,31,113,30,113,29,245,31,3,31,75,31,209,31,130,31,106,31,32,31,125,31,147,31,147,30,205,31,205,30,217,31,217,30,217,29,155,31,5,31,215,31,164,31,164,30,160,31,26,31,8,31,171,31,171,30,171,29,53,31,80,31,80,30,33,31,105,31,203,31,109,31,156,31,156,30,39,31,252,31,251,31,251,30,92,31,41,31,248,31,173,31,113,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
