-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_171 is
end project_tb_171;

architecture project_tb_arch_171 of project_tb_171 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 994;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,197,0,253,0,238,0,74,0,2,0,160,0,0,0,213,0,0,0,154,0,10,0,24,0,0,0,23,0,128,0,173,0,52,0,161,0,85,0,119,0,53,0,0,0,44,0,199,0,7,0,0,0,52,0,229,0,109,0,182,0,140,0,207,0,15,0,0,0,0,0,21,0,79,0,86,0,21,0,221,0,0,0,0,0,196,0,0,0,236,0,0,0,94,0,1,0,105,0,180,0,97,0,0,0,250,0,0,0,0,0,130,0,0,0,66,0,0,0,238,0,234,0,207,0,88,0,0,0,216,0,0,0,0,0,48,0,0,0,0,0,11,0,56,0,0,0,0,0,170,0,157,0,157,0,29,0,179,0,53,0,170,0,43,0,13,0,14,0,236,0,239,0,201,0,167,0,112,0,193,0,10,0,43,0,4,0,44,0,217,0,71,0,82,0,135,0,41,0,0,0,105,0,105,0,47,0,138,0,205,0,185,0,207,0,179,0,114,0,144,0,17,0,230,0,170,0,218,0,0,0,93,0,183,0,0,0,116,0,71,0,126,0,81,0,123,0,31,0,131,0,74,0,94,0,0,0,110,0,58,0,159,0,105,0,235,0,201,0,49,0,181,0,55,0,0,0,158,0,0,0,163,0,8,0,230,0,116,0,133,0,123,0,27,0,212,0,121,0,40,0,0,0,0,0,165,0,0,0,136,0,222,0,100,0,215,0,224,0,101,0,115,0,26,0,55,0,31,0,149,0,0,0,230,0,222,0,0,0,223,0,55,0,244,0,72,0,130,0,74,0,0,0,11,0,72,0,202,0,39,0,48,0,29,0,33,0,50,0,13,0,45,0,11,0,2,0,171,0,135,0,170,0,104,0,0,0,0,0,188,0,221,0,213,0,133,0,178,0,221,0,119,0,202,0,12,0,0,0,0,0,155,0,67,0,218,0,126,0,9,0,79,0,0,0,87,0,0,0,188,0,146,0,238,0,196,0,61,0,219,0,24,0,87,0,200,0,250,0,133,0,247,0,0,0,249,0,108,0,173,0,200,0,183,0,218,0,0,0,47,0,212,0,0,0,0,0,26,0,20,0,110,0,0,0,5,0,208,0,27,0,0,0,123,0,32,0,52,0,172,0,167,0,0,0,48,0,62,0,143,0,0,0,71,0,223,0,175,0,65,0,110,0,199,0,210,0,95,0,1,0,0,0,145,0,0,0,0,0,0,0,250,0,0,0,202,0,180,0,34,0,59,0,67,0,0,0,103,0,90,0,226,0,0,0,64,0,27,0,6,0,86,0,255,0,29,0,206,0,97,0,146,0,148,0,0,0,0,0,39,0,100,0,224,0,174,0,168,0,0,0,180,0,247,0,115,0,87,0,133,0,146,0,156,0,253,0,96,0,0,0,66,0,66,0,217,0,0,0,89,0,68,0,111,0,175,0,142,0,54,0,0,0,240,0,101,0,0,0,0,0,0,0,132,0,170,0,192,0,220,0,65,0,177,0,105,0,27,0,0,0,0,0,201,0,227,0,186,0,229,0,86,0,174,0,0,0,23,0,151,0,0,0,90,0,134,0,169,0,12,0,63,0,0,0,0,0,34,0,168,0,0,0,108,0,115,0,0,0,218,0,134,0,141,0,29,0,179,0,0,0,60,0,0,0,158,0,242,0,148,0,52,0,120,0,160,0,0,0,244,0,0,0,154,0,148,0,58,0,0,0,214,0,76,0,242,0,30,0,101,0,215,0,0,0,219,0,195,0,10,0,170,0,46,0,137,0,103,0,184,0,0,0,2,0,118,0,112,0,107,0,0,0,80,0,0,0,0,0,52,0,152,0,152,0,237,0,0,0,155,0,89,0,189,0,29,0,192,0,233,0,0,0,149,0,225,0,223,0,215,0,84,0,69,0,51,0,156,0,128,0,184,0,31,0,0,0,144,0,35,0,0,0,179,0,0,0,226,0,2,0,135,0,196,0,0,0,126,0,0,0,129,0,118,0,186,0,104,0,62,0,43,0,0,0,0,0,220,0,52,0,59,0,125,0,247,0,68,0,0,0,191,0,19,0,99,0,197,0,90,0,226,0,0,0,51,0,79,0,0,0,95,0,18,0,0,0,25,0,54,0,218,0,157,0,0,0,23,0,0,0,0,0,101,0,80,0,154,0,220,0,186,0,126,0,22,0,0,0,0,0,87,0,29,0,0,0,0,0,0,0,0,0,25,0,214,0,167,0,25,0,189,0,0,0,217,0,34,0,208,0,194,0,243,0,179,0,228,0,232,0,49,0,0,0,0,0,93,0,150,0,169,0,252,0,177,0,140,0,203,0,209,0,169,0,0,0,25,0,183,0,207,0,108,0,0,0,19,0,152,0,70,0,66,0,63,0,60,0,0,0,175,0,135,0,0,0,32,0,132,0,0,0,25,0,0,0,77,0,6,0,195,0,0,0,0,0,110,0,61,0,0,0,0,0,70,0,232,0,178,0,93,0,225,0,0,0,239,0,0,0,237,0,208,0,231,0,165,0,89,0,87,0,60,0,81,0,83,0,36,0,0,0,24,0,70,0,199,0,66,0,147,0,130,0,247,0,0,0,199,0,214,0,6,0,33,0,217,0,202,0,249,0,225,0,239,0,11,0,245,0,190,0,80,0,65,0,0,0,8,0,236,0,122,0,0,0,0,0,198,0,189,0,118,0,74,0,0,0,7,0,158,0,42,0,64,0,0,0,50,0,164,0,86,0,0,0,125,0,46,0,0,0,0,0,40,0,87,0,66,0,0,0,40,0,221,0,157,0,38,0,242,0,0,0,149,0,193,0,49,0,138,0,140,0,0,0,93,0,46,0,0,0,234,0,72,0,179,0,111,0,229,0,173,0,77,0,78,0,227,0,194,0,104,0,205,0,2,0,104,0,0,0,129,0,235,0,0,0,166,0,36,0,192,0,166,0,88,0,143,0,196,0,0,0,169,0,129,0,198,0,182,0,225,0,198,0,0,0,0,0,4,0,125,0,18,0,63,0,29,0,106,0,0,0,17,0,6,0,82,0,177,0,0,0,0,0,138,0,168,0,0,0,46,0,239,0,234,0,118,0,126,0,237,0,155,0,0,0,202,0,100,0,141,0,121,0,135,0,0,0,148,0,131,0,63,0,30,0,138,0,118,0,160,0,92,0,2,0,97,0,174,0,42,0,80,0,219,0,0,0,117,0,167,0,75,0,64,0,215,0,0,0,139,0,0,0,86,0,0,0,0,0,82,0,208,0,163,0,179,0,216,0,0,0,169,0,0,0,123,0,240,0,107,0,0,0,0,0,28,0,41,0,220,0,175,0,18,0,0,0,15,0,50,0,0,0,217,0,74,0,96,0,220,0,248,0,192,0,8,0,214,0,241,0,225,0,182,0,147,0,158,0,224,0,0,0,81,0,25,0,119,0,126,0,0,0,189,0,0,0,0,0,128,0,200,0,41,0,146,0,0,0,190,0,42,0,22,0,158,0,14,0,55,0,0,0,221,0,239,0,7,0,23,0,213,0,0,0,61,0,223,0,230,0,58,0,57,0,189,0,101,0,169,0,248,0,6,0,70,0,42,0,9,0,30,0,26,0,174,0,165,0,133,0,144,0,0,0,78,0,0,0,0,0,0,0,151,0,17,0,177,0,27,0,0,0,196,0,152,0,71,0,74,0,0,0,9,0,51,0,158,0,0,0,228,0,125,0,0,0,195,0,144,0,101,0,250,0,0,0,106,0,27,0,214,0,42,0,0,0,178,0,0,0,84,0,76,0,194,0,69,0,164,0,64,0,0,0,242,0,109,0,104,0,249,0,121,0,0,0,27,0,7,0,92,0,77,0,80,0,0,0,0,0,0,0,62,0,254,0,125,0,54,0,118,0,0,0,137,0,235,0,133,0,218,0,235,0,0,0,0,0,152,0,0,0,24,0,10,0,120,0,40,0,37,0,40,0,0,0,244,0,95,0,193,0,164,0,0,0,125,0,0,0,196,0,31,0,137,0,201,0,0,0,111,0,51,0,102,0,119,0,235,0,0,0,242,0,0,0,115,0,40,0,226,0,178,0,47,0,0,0,216,0,16,0,26,0,113,0,254,0,230,0,205,0,33,0,55,0,0,0,225,0,0,0,86,0,71,0,125,0,36,0,0,0,31,0,0,0,61,0,31,0,153,0,0,0,132,0,101,0,107,0,123,0,0,0,222,0,151,0,0,0,65,0,111,0,243,0,110,0,72,0,49,0,121,0,143,0,128,0,80,0,53,0,0,0,107,0,0,0,210,0,0,0,180,0,0,0,96,0,152,0,0,0,50,0,19,0,39,0,216,0,157,0,116,0,112,0,115,0,18,0,59,0,217,0,245,0,0,0,220,0,27,0,121,0,8,0,70,0,91,0,162,0,121,0,63,0,242,0,140,0,197,0,152,0,225,0,79,0,64,0,114,0,197,0,83,0,166,0,28,0,237,0);
signal scenario_full  : scenario_type := (0,0,197,31,253,31,238,31,74,31,2,31,160,31,160,30,213,31,213,30,154,31,10,31,24,31,24,30,23,31,128,31,173,31,52,31,161,31,85,31,119,31,53,31,53,30,44,31,199,31,7,31,7,30,52,31,229,31,109,31,182,31,140,31,207,31,15,31,15,30,15,29,21,31,79,31,86,31,21,31,221,31,221,30,221,29,196,31,196,30,236,31,236,30,94,31,1,31,105,31,180,31,97,31,97,30,250,31,250,30,250,29,130,31,130,30,66,31,66,30,238,31,234,31,207,31,88,31,88,30,216,31,216,30,216,29,48,31,48,30,48,29,11,31,56,31,56,30,56,29,170,31,157,31,157,31,29,31,179,31,53,31,170,31,43,31,13,31,14,31,236,31,239,31,201,31,167,31,112,31,193,31,10,31,43,31,4,31,44,31,217,31,71,31,82,31,135,31,41,31,41,30,105,31,105,31,47,31,138,31,205,31,185,31,207,31,179,31,114,31,144,31,17,31,230,31,170,31,218,31,218,30,93,31,183,31,183,30,116,31,71,31,126,31,81,31,123,31,31,31,131,31,74,31,94,31,94,30,110,31,58,31,159,31,105,31,235,31,201,31,49,31,181,31,55,31,55,30,158,31,158,30,163,31,8,31,230,31,116,31,133,31,123,31,27,31,212,31,121,31,40,31,40,30,40,29,165,31,165,30,136,31,222,31,100,31,215,31,224,31,101,31,115,31,26,31,55,31,31,31,149,31,149,30,230,31,222,31,222,30,223,31,55,31,244,31,72,31,130,31,74,31,74,30,11,31,72,31,202,31,39,31,48,31,29,31,33,31,50,31,13,31,45,31,11,31,2,31,171,31,135,31,170,31,104,31,104,30,104,29,188,31,221,31,213,31,133,31,178,31,221,31,119,31,202,31,12,31,12,30,12,29,155,31,67,31,218,31,126,31,9,31,79,31,79,30,87,31,87,30,188,31,146,31,238,31,196,31,61,31,219,31,24,31,87,31,200,31,250,31,133,31,247,31,247,30,249,31,108,31,173,31,200,31,183,31,218,31,218,30,47,31,212,31,212,30,212,29,26,31,20,31,110,31,110,30,5,31,208,31,27,31,27,30,123,31,32,31,52,31,172,31,167,31,167,30,48,31,62,31,143,31,143,30,71,31,223,31,175,31,65,31,110,31,199,31,210,31,95,31,1,31,1,30,145,31,145,30,145,29,145,28,250,31,250,30,202,31,180,31,34,31,59,31,67,31,67,30,103,31,90,31,226,31,226,30,64,31,27,31,6,31,86,31,255,31,29,31,206,31,97,31,146,31,148,31,148,30,148,29,39,31,100,31,224,31,174,31,168,31,168,30,180,31,247,31,115,31,87,31,133,31,146,31,156,31,253,31,96,31,96,30,66,31,66,31,217,31,217,30,89,31,68,31,111,31,175,31,142,31,54,31,54,30,240,31,101,31,101,30,101,29,101,28,132,31,170,31,192,31,220,31,65,31,177,31,105,31,27,31,27,30,27,29,201,31,227,31,186,31,229,31,86,31,174,31,174,30,23,31,151,31,151,30,90,31,134,31,169,31,12,31,63,31,63,30,63,29,34,31,168,31,168,30,108,31,115,31,115,30,218,31,134,31,141,31,29,31,179,31,179,30,60,31,60,30,158,31,242,31,148,31,52,31,120,31,160,31,160,30,244,31,244,30,154,31,148,31,58,31,58,30,214,31,76,31,242,31,30,31,101,31,215,31,215,30,219,31,195,31,10,31,170,31,46,31,137,31,103,31,184,31,184,30,2,31,118,31,112,31,107,31,107,30,80,31,80,30,80,29,52,31,152,31,152,31,237,31,237,30,155,31,89,31,189,31,29,31,192,31,233,31,233,30,149,31,225,31,223,31,215,31,84,31,69,31,51,31,156,31,128,31,184,31,31,31,31,30,144,31,35,31,35,30,179,31,179,30,226,31,2,31,135,31,196,31,196,30,126,31,126,30,129,31,118,31,186,31,104,31,62,31,43,31,43,30,43,29,220,31,52,31,59,31,125,31,247,31,68,31,68,30,191,31,19,31,99,31,197,31,90,31,226,31,226,30,51,31,79,31,79,30,95,31,18,31,18,30,25,31,54,31,218,31,157,31,157,30,23,31,23,30,23,29,101,31,80,31,154,31,220,31,186,31,126,31,22,31,22,30,22,29,87,31,29,31,29,30,29,29,29,28,29,27,25,31,214,31,167,31,25,31,189,31,189,30,217,31,34,31,208,31,194,31,243,31,179,31,228,31,232,31,49,31,49,30,49,29,93,31,150,31,169,31,252,31,177,31,140,31,203,31,209,31,169,31,169,30,25,31,183,31,207,31,108,31,108,30,19,31,152,31,70,31,66,31,63,31,60,31,60,30,175,31,135,31,135,30,32,31,132,31,132,30,25,31,25,30,77,31,6,31,195,31,195,30,195,29,110,31,61,31,61,30,61,29,70,31,232,31,178,31,93,31,225,31,225,30,239,31,239,30,237,31,208,31,231,31,165,31,89,31,87,31,60,31,81,31,83,31,36,31,36,30,24,31,70,31,199,31,66,31,147,31,130,31,247,31,247,30,199,31,214,31,6,31,33,31,217,31,202,31,249,31,225,31,239,31,11,31,245,31,190,31,80,31,65,31,65,30,8,31,236,31,122,31,122,30,122,29,198,31,189,31,118,31,74,31,74,30,7,31,158,31,42,31,64,31,64,30,50,31,164,31,86,31,86,30,125,31,46,31,46,30,46,29,40,31,87,31,66,31,66,30,40,31,221,31,157,31,38,31,242,31,242,30,149,31,193,31,49,31,138,31,140,31,140,30,93,31,46,31,46,30,234,31,72,31,179,31,111,31,229,31,173,31,77,31,78,31,227,31,194,31,104,31,205,31,2,31,104,31,104,30,129,31,235,31,235,30,166,31,36,31,192,31,166,31,88,31,143,31,196,31,196,30,169,31,129,31,198,31,182,31,225,31,198,31,198,30,198,29,4,31,125,31,18,31,63,31,29,31,106,31,106,30,17,31,6,31,82,31,177,31,177,30,177,29,138,31,168,31,168,30,46,31,239,31,234,31,118,31,126,31,237,31,155,31,155,30,202,31,100,31,141,31,121,31,135,31,135,30,148,31,131,31,63,31,30,31,138,31,118,31,160,31,92,31,2,31,97,31,174,31,42,31,80,31,219,31,219,30,117,31,167,31,75,31,64,31,215,31,215,30,139,31,139,30,86,31,86,30,86,29,82,31,208,31,163,31,179,31,216,31,216,30,169,31,169,30,123,31,240,31,107,31,107,30,107,29,28,31,41,31,220,31,175,31,18,31,18,30,15,31,50,31,50,30,217,31,74,31,96,31,220,31,248,31,192,31,8,31,214,31,241,31,225,31,182,31,147,31,158,31,224,31,224,30,81,31,25,31,119,31,126,31,126,30,189,31,189,30,189,29,128,31,200,31,41,31,146,31,146,30,190,31,42,31,22,31,158,31,14,31,55,31,55,30,221,31,239,31,7,31,23,31,213,31,213,30,61,31,223,31,230,31,58,31,57,31,189,31,101,31,169,31,248,31,6,31,70,31,42,31,9,31,30,31,26,31,174,31,165,31,133,31,144,31,144,30,78,31,78,30,78,29,78,28,151,31,17,31,177,31,27,31,27,30,196,31,152,31,71,31,74,31,74,30,9,31,51,31,158,31,158,30,228,31,125,31,125,30,195,31,144,31,101,31,250,31,250,30,106,31,27,31,214,31,42,31,42,30,178,31,178,30,84,31,76,31,194,31,69,31,164,31,64,31,64,30,242,31,109,31,104,31,249,31,121,31,121,30,27,31,7,31,92,31,77,31,80,31,80,30,80,29,80,28,62,31,254,31,125,31,54,31,118,31,118,30,137,31,235,31,133,31,218,31,235,31,235,30,235,29,152,31,152,30,24,31,10,31,120,31,40,31,37,31,40,31,40,30,244,31,95,31,193,31,164,31,164,30,125,31,125,30,196,31,31,31,137,31,201,31,201,30,111,31,51,31,102,31,119,31,235,31,235,30,242,31,242,30,115,31,40,31,226,31,178,31,47,31,47,30,216,31,16,31,26,31,113,31,254,31,230,31,205,31,33,31,55,31,55,30,225,31,225,30,86,31,71,31,125,31,36,31,36,30,31,31,31,30,61,31,31,31,153,31,153,30,132,31,101,31,107,31,123,31,123,30,222,31,151,31,151,30,65,31,111,31,243,31,110,31,72,31,49,31,121,31,143,31,128,31,80,31,53,31,53,30,107,31,107,30,210,31,210,30,180,31,180,30,96,31,152,31,152,30,50,31,19,31,39,31,216,31,157,31,116,31,112,31,115,31,18,31,59,31,217,31,245,31,245,30,220,31,27,31,121,31,8,31,70,31,91,31,162,31,121,31,63,31,242,31,140,31,197,31,152,31,225,31,79,31,64,31,114,31,197,31,83,31,166,31,28,31,237,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
