-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_359 is
end project_tb_359;

architecture project_tb_arch_359 of project_tb_359 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 312;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,152,0,87,0,0,0,187,0,53,0,100,0,197,0,213,0,59,0,57,0,138,0,157,0,180,0,177,0,0,0,215,0,141,0,0,0,115,0,0,0,178,0,161,0,21,0,102,0,203,0,150,0,61,0,172,0,4,0,63,0,21,0,108,0,24,0,0,0,60,0,0,0,7,0,22,0,0,0,127,0,49,0,254,0,2,0,174,0,0,0,98,0,153,0,155,0,157,0,0,0,201,0,190,0,183,0,50,0,218,0,112,0,69,0,193,0,25,0,0,0,175,0,16,0,0,0,27,0,0,0,166,0,24,0,36,0,0,0,113,0,0,0,0,0,227,0,0,0,63,0,73,0,77,0,153,0,99,0,44,0,155,0,45,0,210,0,56,0,154,0,121,0,0,0,87,0,0,0,110,0,131,0,200,0,218,0,102,0,7,0,174,0,0,0,0,0,188,0,172,0,182,0,95,0,162,0,115,0,222,0,0,0,0,0,19,0,171,0,141,0,97,0,0,0,255,0,191,0,52,0,14,0,237,0,88,0,20,0,52,0,79,0,115,0,11,0,113,0,82,0,0,0,78,0,61,0,233,0,44,0,255,0,220,0,127,0,95,0,16,0,8,0,110,0,0,0,0,0,150,0,0,0,0,0,77,0,0,0,130,0,40,0,0,0,198,0,169,0,9,0,199,0,30,0,91,0,85,0,120,0,4,0,65,0,169,0,0,0,70,0,125,0,0,0,151,0,136,0,203,0,44,0,194,0,192,0,0,0,161,0,26,0,131,0,64,0,214,0,96,0,47,0,172,0,168,0,172,0,124,0,253,0,196,0,79,0,110,0,0,0,154,0,175,0,0,0,0,0,0,0,194,0,194,0,50,0,144,0,183,0,163,0,57,0,231,0,20,0,197,0,235,0,215,0,224,0,7,0,112,0,98,0,222,0,200,0,71,0,35,0,185,0,138,0,0,0,238,0,114,0,137,0,0,0,0,0,47,0,51,0,210,0,88,0,19,0,3,0,88,0,238,0,126,0,57,0,0,0,0,0,134,0,12,0,104,0,0,0,0,0,0,0,236,0,82,0,198,0,73,0,1,0,188,0,2,0,248,0,133,0,27,0,78,0,35,0,222,0,0,0,219,0,159,0,116,0,0,0,0,0,194,0,139,0,96,0,205,0,89,0,0,0,11,0,76,0,0,0,10,0,237,0,0,0,0,0,12,0,41,0,148,0,0,0,0,0,144,0,0,0,32,0,46,0,107,0,239,0,0,0,147,0,12,0,205,0,0,0,62,0,159,0,0,0,187,0,0,0,0,0,117,0,12,0,176,0,106,0,175,0,81,0,44,0,44,0,168,0,96,0,15,0,0,0,123,0,111,0,121,0,12,0,10,0,203,0,0,0,61,0,186,0);
signal scenario_full  : scenario_type := (135,31,152,31,87,31,87,30,187,31,53,31,100,31,197,31,213,31,59,31,57,31,138,31,157,31,180,31,177,31,177,30,215,31,141,31,141,30,115,31,115,30,178,31,161,31,21,31,102,31,203,31,150,31,61,31,172,31,4,31,63,31,21,31,108,31,24,31,24,30,60,31,60,30,7,31,22,31,22,30,127,31,49,31,254,31,2,31,174,31,174,30,98,31,153,31,155,31,157,31,157,30,201,31,190,31,183,31,50,31,218,31,112,31,69,31,193,31,25,31,25,30,175,31,16,31,16,30,27,31,27,30,166,31,24,31,36,31,36,30,113,31,113,30,113,29,227,31,227,30,63,31,73,31,77,31,153,31,99,31,44,31,155,31,45,31,210,31,56,31,154,31,121,31,121,30,87,31,87,30,110,31,131,31,200,31,218,31,102,31,7,31,174,31,174,30,174,29,188,31,172,31,182,31,95,31,162,31,115,31,222,31,222,30,222,29,19,31,171,31,141,31,97,31,97,30,255,31,191,31,52,31,14,31,237,31,88,31,20,31,52,31,79,31,115,31,11,31,113,31,82,31,82,30,78,31,61,31,233,31,44,31,255,31,220,31,127,31,95,31,16,31,8,31,110,31,110,30,110,29,150,31,150,30,150,29,77,31,77,30,130,31,40,31,40,30,198,31,169,31,9,31,199,31,30,31,91,31,85,31,120,31,4,31,65,31,169,31,169,30,70,31,125,31,125,30,151,31,136,31,203,31,44,31,194,31,192,31,192,30,161,31,26,31,131,31,64,31,214,31,96,31,47,31,172,31,168,31,172,31,124,31,253,31,196,31,79,31,110,31,110,30,154,31,175,31,175,30,175,29,175,28,194,31,194,31,50,31,144,31,183,31,163,31,57,31,231,31,20,31,197,31,235,31,215,31,224,31,7,31,112,31,98,31,222,31,200,31,71,31,35,31,185,31,138,31,138,30,238,31,114,31,137,31,137,30,137,29,47,31,51,31,210,31,88,31,19,31,3,31,88,31,238,31,126,31,57,31,57,30,57,29,134,31,12,31,104,31,104,30,104,29,104,28,236,31,82,31,198,31,73,31,1,31,188,31,2,31,248,31,133,31,27,31,78,31,35,31,222,31,222,30,219,31,159,31,116,31,116,30,116,29,194,31,139,31,96,31,205,31,89,31,89,30,11,31,76,31,76,30,10,31,237,31,237,30,237,29,12,31,41,31,148,31,148,30,148,29,144,31,144,30,32,31,46,31,107,31,239,31,239,30,147,31,12,31,205,31,205,30,62,31,159,31,159,30,187,31,187,30,187,29,117,31,12,31,176,31,106,31,175,31,81,31,44,31,44,31,168,31,96,31,15,31,15,30,123,31,111,31,121,31,12,31,10,31,203,31,203,30,61,31,186,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
