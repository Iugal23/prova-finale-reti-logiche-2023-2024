-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_558 is
end project_tb_558;

architecture project_tb_arch_558 of project_tb_558 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 941;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (57,0,86,0,226,0,195,0,0,0,0,0,0,0,0,0,215,0,55,0,42,0,36,0,0,0,220,0,46,0,170,0,194,0,144,0,23,0,238,0,58,0,241,0,0,0,73,0,115,0,36,0,124,0,139,0,206,0,25,0,0,0,189,0,0,0,161,0,0,0,0,0,60,0,216,0,14,0,3,0,0,0,122,0,0,0,183,0,33,0,209,0,0,0,151,0,126,0,83,0,29,0,0,0,38,0,150,0,251,0,181,0,177,0,80,0,222,0,0,0,243,0,0,0,207,0,152,0,153,0,0,0,57,0,135,0,109,0,109,0,93,0,42,0,65,0,234,0,150,0,226,0,0,0,205,0,71,0,0,0,216,0,165,0,0,0,73,0,0,0,5,0,37,0,106,0,42,0,45,0,6,0,94,0,175,0,86,0,41,0,200,0,147,0,247,0,251,0,115,0,7,0,139,0,146,0,0,0,0,0,223,0,0,0,54,0,211,0,82,0,223,0,0,0,184,0,45,0,234,0,65,0,3,0,3,0,53,0,246,0,0,0,162,0,63,0,99,0,0,0,66,0,0,0,13,0,233,0,92,0,91,0,51,0,206,0,216,0,173,0,48,0,191,0,233,0,0,0,120,0,191,0,91,0,21,0,187,0,145,0,100,0,0,0,0,0,0,0,226,0,45,0,186,0,32,0,220,0,0,0,0,0,53,0,40,0,82,0,0,0,0,0,98,0,245,0,35,0,0,0,0,0,121,0,0,0,172,0,64,0,0,0,136,0,165,0,223,0,169,0,50,0,188,0,29,0,243,0,77,0,0,0,104,0,0,0,207,0,167,0,49,0,216,0,69,0,35,0,224,0,17,0,102,0,238,0,0,0,60,0,146,0,143,0,0,0,235,0,26,0,62,0,0,0,0,0,195,0,199,0,252,0,151,0,245,0,89,0,0,0,0,0,162,0,0,0,0,0,0,0,216,0,0,0,54,0,87,0,172,0,15,0,78,0,94,0,55,0,67,0,0,0,0,0,84,0,176,0,0,0,150,0,238,0,0,0,89,0,218,0,208,0,119,0,241,0,108,0,251,0,58,0,0,0,150,0,204,0,238,0,243,0,27,0,185,0,145,0,127,0,46,0,236,0,0,0,157,0,191,0,158,0,180,0,12,0,61,0,15,0,176,0,194,0,86,0,18,0,247,0,159,0,185,0,170,0,0,0,185,0,188,0,51,0,233,0,218,0,235,0,200,0,137,0,159,0,167,0,0,0,192,0,0,0,85,0,166,0,227,0,0,0,0,0,6,0,208,0,0,0,143,0,96,0,70,0,227,0,82,0,0,0,206,0,107,0,167,0,97,0,25,0,143,0,0,0,64,0,247,0,55,0,186,0,0,0,78,0,0,0,11,0,31,0,0,0,53,0,0,0,0,0,71,0,71,0,71,0,230,0,184,0,0,0,201,0,151,0,124,0,125,0,67,0,7,0,103,0,29,0,227,0,4,0,16,0,0,0,44,0,255,0,173,0,207,0,0,0,2,0,81,0,52,0,179,0,184,0,132,0,22,0,21,0,26,0,0,0,17,0,65,0,234,0,117,0,103,0,103,0,189,0,63,0,131,0,226,0,77,0,149,0,0,0,0,0,171,0,177,0,0,0,0,0,206,0,81,0,92,0,128,0,0,0,202,0,160,0,82,0,0,0,239,0,121,0,250,0,19,0,167,0,82,0,0,0,228,0,68,0,221,0,213,0,71,0,27,0,5,0,193,0,103,0,218,0,88,0,189,0,120,0,89,0,0,0,77,0,47,0,75,0,223,0,173,0,76,0,0,0,0,0,42,0,38,0,75,0,180,0,197,0,38,0,213,0,10,0,158,0,17,0,56,0,7,0,192,0,47,0,65,0,0,0,0,0,65,0,196,0,0,0,226,0,14,0,60,0,158,0,172,0,10,0,16,0,241,0,230,0,0,0,212,0,86,0,165,0,31,0,0,0,27,0,146,0,197,0,165,0,68,0,77,0,38,0,77,0,41,0,192,0,0,0,29,0,46,0,209,0,52,0,11,0,159,0,190,0,243,0,139,0,224,0,151,0,241,0,179,0,227,0,108,0,102,0,23,0,152,0,0,0,49,0,63,0,223,0,207,0,58,0,48,0,246,0,9,0,179,0,144,0,66,0,158,0,148,0,250,0,169,0,0,0,2,0,116,0,0,0,0,0,200,0,212,0,96,0,21,0,133,0,11,0,240,0,14,0,135,0,170,0,250,0,0,0,164,0,68,0,198,0,0,0,125,0,243,0,0,0,144,0,190,0,148,0,164,0,8,0,0,0,93,0,237,0,216,0,28,0,209,0,16,0,145,0,148,0,79,0,225,0,229,0,89,0,103,0,146,0,131,0,94,0,118,0,167,0,48,0,6,0,2,0,0,0,83,0,0,0,198,0,0,0,232,0,194,0,26,0,0,0,0,0,43,0,123,0,188,0,0,0,76,0,252,0,47,0,231,0,0,0,29,0,50,0,224,0,224,0,0,0,195,0,7,0,249,0,68,0,17,0,126,0,26,0,56,0,0,0,66,0,114,0,149,0,0,0,122,0,9,0,182,0,86,0,0,0,33,0,93,0,0,0,195,0,9,0,125,0,194,0,239,0,1,0,42,0,240,0,40,0,4,0,207,0,204,0,107,0,0,0,31,0,0,0,209,0,125,0,0,0,0,0,131,0,8,0,59,0,84,0,0,0,179,0,215,0,105,0,190,0,244,0,73,0,134,0,0,0,175,0,18,0,193,0,17,0,30,0,241,0,197,0,80,0,107,0,216,0,146,0,244,0,8,0,0,0,234,0,113,0,71,0,197,0,46,0,234,0,84,0,0,0,160,0,122,0,25,0,14,0,0,0,186,0,89,0,137,0,140,0,80,0,0,0,50,0,102,0,189,0,43,0,165,0,142,0,200,0,0,0,137,0,177,0,188,0,0,0,157,0,0,0,3,0,105,0,15,0,87,0,0,0,0,0,188,0,99,0,27,0,42,0,150,0,111,0,122,0,233,0,44,0,149,0,245,0,236,0,0,0,205,0,15,0,179,0,237,0,202,0,153,0,232,0,32,0,128,0,145,0,68,0,0,0,248,0,31,0,108,0,160,0,61,0,226,0,158,0,0,0,0,0,37,0,0,0,0,0,0,0,147,0,209,0,18,0,23,0,242,0,132,0,23,0,169,0,163,0,60,0,31,0,203,0,0,0,93,0,72,0,0,0,81,0,139,0,0,0,33,0,0,0,0,0,30,0,0,0,79,0,104,0,0,0,97,0,0,0,91,0,237,0,94,0,177,0,133,0,0,0,172,0,0,0,234,0,0,0,91,0,57,0,0,0,18,0,35,0,13,0,47,0,136,0,113,0,91,0,0,0,55,0,58,0,15,0,55,0,80,0,129,0,99,0,194,0,195,0,87,0,101,0,61,0,0,0,36,0,0,0,91,0,0,0,100,0,33,0,149,0,220,0,161,0,149,0,157,0,147,0,89,0,0,0,213,0,98,0,0,0,0,0,194,0,0,0,0,0,135,0,237,0,0,0,207,0,0,0,0,0,227,0,0,0,108,0,211,0,162,0,24,0,216,0,213,0,23,0,147,0,0,0,252,0,62,0,191,0,147,0,253,0,247,0,0,0,202,0,165,0,107,0,1,0,208,0,0,0,219,0,210,0,50,0,125,0,112,0,0,0,77,0,0,0,47,0,69,0,54,0,21,0,46,0,18,0,28,0,151,0,20,0,0,0,99,0,0,0,54,0,111,0,0,0,141,0,201,0,105,0,19,0,127,0,0,0,0,0,19,0,0,0,244,0,203,0,0,0,0,0,143,0,0,0,63,0,197,0,130,0,248,0,102,0,75,0,101,0,12,0,173,0,208,0,87,0,33,0,56,0,0,0,130,0,190,0,46,0,92,0,87,0,0,0,117,0,102,0,142,0,233,0,0,0,42,0,31,0,0,0,0,0,124,0,0,0,75,0,16,0,197,0,0,0,43,0,199,0,15,0,0,0,96,0,198,0,61,0,243,0,240,0,18,0,32,0,122,0,106,0,14,0,78,0,54,0,218,0,0,0,99,0,236,0,53,0,0,0,33,0,49,0,95,0,169,0,45,0,37,0,64,0,131,0,209,0,34,0,193,0,0,0,147,0,204,0,79,0,0,0,248,0,73,0,74,0,48,0,150,0,129,0,0,0,30,0,255,0,122,0);
signal scenario_full  : scenario_type := (57,31,86,31,226,31,195,31,195,30,195,29,195,28,195,27,215,31,55,31,42,31,36,31,36,30,220,31,46,31,170,31,194,31,144,31,23,31,238,31,58,31,241,31,241,30,73,31,115,31,36,31,124,31,139,31,206,31,25,31,25,30,189,31,189,30,161,31,161,30,161,29,60,31,216,31,14,31,3,31,3,30,122,31,122,30,183,31,33,31,209,31,209,30,151,31,126,31,83,31,29,31,29,30,38,31,150,31,251,31,181,31,177,31,80,31,222,31,222,30,243,31,243,30,207,31,152,31,153,31,153,30,57,31,135,31,109,31,109,31,93,31,42,31,65,31,234,31,150,31,226,31,226,30,205,31,71,31,71,30,216,31,165,31,165,30,73,31,73,30,5,31,37,31,106,31,42,31,45,31,6,31,94,31,175,31,86,31,41,31,200,31,147,31,247,31,251,31,115,31,7,31,139,31,146,31,146,30,146,29,223,31,223,30,54,31,211,31,82,31,223,31,223,30,184,31,45,31,234,31,65,31,3,31,3,31,53,31,246,31,246,30,162,31,63,31,99,31,99,30,66,31,66,30,13,31,233,31,92,31,91,31,51,31,206,31,216,31,173,31,48,31,191,31,233,31,233,30,120,31,191,31,91,31,21,31,187,31,145,31,100,31,100,30,100,29,100,28,226,31,45,31,186,31,32,31,220,31,220,30,220,29,53,31,40,31,82,31,82,30,82,29,98,31,245,31,35,31,35,30,35,29,121,31,121,30,172,31,64,31,64,30,136,31,165,31,223,31,169,31,50,31,188,31,29,31,243,31,77,31,77,30,104,31,104,30,207,31,167,31,49,31,216,31,69,31,35,31,224,31,17,31,102,31,238,31,238,30,60,31,146,31,143,31,143,30,235,31,26,31,62,31,62,30,62,29,195,31,199,31,252,31,151,31,245,31,89,31,89,30,89,29,162,31,162,30,162,29,162,28,216,31,216,30,54,31,87,31,172,31,15,31,78,31,94,31,55,31,67,31,67,30,67,29,84,31,176,31,176,30,150,31,238,31,238,30,89,31,218,31,208,31,119,31,241,31,108,31,251,31,58,31,58,30,150,31,204,31,238,31,243,31,27,31,185,31,145,31,127,31,46,31,236,31,236,30,157,31,191,31,158,31,180,31,12,31,61,31,15,31,176,31,194,31,86,31,18,31,247,31,159,31,185,31,170,31,170,30,185,31,188,31,51,31,233,31,218,31,235,31,200,31,137,31,159,31,167,31,167,30,192,31,192,30,85,31,166,31,227,31,227,30,227,29,6,31,208,31,208,30,143,31,96,31,70,31,227,31,82,31,82,30,206,31,107,31,167,31,97,31,25,31,143,31,143,30,64,31,247,31,55,31,186,31,186,30,78,31,78,30,11,31,31,31,31,30,53,31,53,30,53,29,71,31,71,31,71,31,230,31,184,31,184,30,201,31,151,31,124,31,125,31,67,31,7,31,103,31,29,31,227,31,4,31,16,31,16,30,44,31,255,31,173,31,207,31,207,30,2,31,81,31,52,31,179,31,184,31,132,31,22,31,21,31,26,31,26,30,17,31,65,31,234,31,117,31,103,31,103,31,189,31,63,31,131,31,226,31,77,31,149,31,149,30,149,29,171,31,177,31,177,30,177,29,206,31,81,31,92,31,128,31,128,30,202,31,160,31,82,31,82,30,239,31,121,31,250,31,19,31,167,31,82,31,82,30,228,31,68,31,221,31,213,31,71,31,27,31,5,31,193,31,103,31,218,31,88,31,189,31,120,31,89,31,89,30,77,31,47,31,75,31,223,31,173,31,76,31,76,30,76,29,42,31,38,31,75,31,180,31,197,31,38,31,213,31,10,31,158,31,17,31,56,31,7,31,192,31,47,31,65,31,65,30,65,29,65,31,196,31,196,30,226,31,14,31,60,31,158,31,172,31,10,31,16,31,241,31,230,31,230,30,212,31,86,31,165,31,31,31,31,30,27,31,146,31,197,31,165,31,68,31,77,31,38,31,77,31,41,31,192,31,192,30,29,31,46,31,209,31,52,31,11,31,159,31,190,31,243,31,139,31,224,31,151,31,241,31,179,31,227,31,108,31,102,31,23,31,152,31,152,30,49,31,63,31,223,31,207,31,58,31,48,31,246,31,9,31,179,31,144,31,66,31,158,31,148,31,250,31,169,31,169,30,2,31,116,31,116,30,116,29,200,31,212,31,96,31,21,31,133,31,11,31,240,31,14,31,135,31,170,31,250,31,250,30,164,31,68,31,198,31,198,30,125,31,243,31,243,30,144,31,190,31,148,31,164,31,8,31,8,30,93,31,237,31,216,31,28,31,209,31,16,31,145,31,148,31,79,31,225,31,229,31,89,31,103,31,146,31,131,31,94,31,118,31,167,31,48,31,6,31,2,31,2,30,83,31,83,30,198,31,198,30,232,31,194,31,26,31,26,30,26,29,43,31,123,31,188,31,188,30,76,31,252,31,47,31,231,31,231,30,29,31,50,31,224,31,224,31,224,30,195,31,7,31,249,31,68,31,17,31,126,31,26,31,56,31,56,30,66,31,114,31,149,31,149,30,122,31,9,31,182,31,86,31,86,30,33,31,93,31,93,30,195,31,9,31,125,31,194,31,239,31,1,31,42,31,240,31,40,31,4,31,207,31,204,31,107,31,107,30,31,31,31,30,209,31,125,31,125,30,125,29,131,31,8,31,59,31,84,31,84,30,179,31,215,31,105,31,190,31,244,31,73,31,134,31,134,30,175,31,18,31,193,31,17,31,30,31,241,31,197,31,80,31,107,31,216,31,146,31,244,31,8,31,8,30,234,31,113,31,71,31,197,31,46,31,234,31,84,31,84,30,160,31,122,31,25,31,14,31,14,30,186,31,89,31,137,31,140,31,80,31,80,30,50,31,102,31,189,31,43,31,165,31,142,31,200,31,200,30,137,31,177,31,188,31,188,30,157,31,157,30,3,31,105,31,15,31,87,31,87,30,87,29,188,31,99,31,27,31,42,31,150,31,111,31,122,31,233,31,44,31,149,31,245,31,236,31,236,30,205,31,15,31,179,31,237,31,202,31,153,31,232,31,32,31,128,31,145,31,68,31,68,30,248,31,31,31,108,31,160,31,61,31,226,31,158,31,158,30,158,29,37,31,37,30,37,29,37,28,147,31,209,31,18,31,23,31,242,31,132,31,23,31,169,31,163,31,60,31,31,31,203,31,203,30,93,31,72,31,72,30,81,31,139,31,139,30,33,31,33,30,33,29,30,31,30,30,79,31,104,31,104,30,97,31,97,30,91,31,237,31,94,31,177,31,133,31,133,30,172,31,172,30,234,31,234,30,91,31,57,31,57,30,18,31,35,31,13,31,47,31,136,31,113,31,91,31,91,30,55,31,58,31,15,31,55,31,80,31,129,31,99,31,194,31,195,31,87,31,101,31,61,31,61,30,36,31,36,30,91,31,91,30,100,31,33,31,149,31,220,31,161,31,149,31,157,31,147,31,89,31,89,30,213,31,98,31,98,30,98,29,194,31,194,30,194,29,135,31,237,31,237,30,207,31,207,30,207,29,227,31,227,30,108,31,211,31,162,31,24,31,216,31,213,31,23,31,147,31,147,30,252,31,62,31,191,31,147,31,253,31,247,31,247,30,202,31,165,31,107,31,1,31,208,31,208,30,219,31,210,31,50,31,125,31,112,31,112,30,77,31,77,30,47,31,69,31,54,31,21,31,46,31,18,31,28,31,151,31,20,31,20,30,99,31,99,30,54,31,111,31,111,30,141,31,201,31,105,31,19,31,127,31,127,30,127,29,19,31,19,30,244,31,203,31,203,30,203,29,143,31,143,30,63,31,197,31,130,31,248,31,102,31,75,31,101,31,12,31,173,31,208,31,87,31,33,31,56,31,56,30,130,31,190,31,46,31,92,31,87,31,87,30,117,31,102,31,142,31,233,31,233,30,42,31,31,31,31,30,31,29,124,31,124,30,75,31,16,31,197,31,197,30,43,31,199,31,15,31,15,30,96,31,198,31,61,31,243,31,240,31,18,31,32,31,122,31,106,31,14,31,78,31,54,31,218,31,218,30,99,31,236,31,53,31,53,30,33,31,49,31,95,31,169,31,45,31,37,31,64,31,131,31,209,31,34,31,193,31,193,30,147,31,204,31,79,31,79,30,248,31,73,31,74,31,48,31,150,31,129,31,129,30,30,31,255,31,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
