-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 795;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (210,0,252,0,88,0,183,0,192,0,177,0,124,0,0,0,0,0,189,0,94,0,0,0,0,0,242,0,199,0,0,0,158,0,116,0,0,0,0,0,81,0,0,0,109,0,0,0,222,0,255,0,0,0,0,0,32,0,0,0,254,0,18,0,0,0,177,0,252,0,12,0,0,0,227,0,94,0,148,0,9,0,189,0,29,0,0,0,184,0,253,0,227,0,213,0,106,0,101,0,0,0,0,0,22,0,253,0,83,0,194,0,53,0,185,0,0,0,184,0,162,0,179,0,71,0,126,0,46,0,33,0,56,0,0,0,226,0,120,0,18,0,249,0,0,0,230,0,0,0,197,0,33,0,0,0,0,0,68,0,165,0,34,0,227,0,137,0,182,0,236,0,0,0,0,0,124,0,153,0,223,0,133,0,130,0,224,0,194,0,239,0,254,0,113,0,123,0,244,0,0,0,15,0,254,0,133,0,192,0,140,0,0,0,13,0,212,0,103,0,237,0,37,0,0,0,216,0,0,0,114,0,97,0,166,0,0,0,110,0,170,0,73,0,15,0,0,0,31,0,37,0,120,0,0,0,166,0,0,0,119,0,254,0,154,0,174,0,118,0,234,0,58,0,0,0,169,0,35,0,201,0,230,0,82,0,141,0,0,0,196,0,39,0,0,0,0,0,0,0,114,0,0,0,47,0,0,0,65,0,54,0,157,0,245,0,181,0,0,0,16,0,178,0,137,0,144,0,175,0,157,0,104,0,114,0,0,0,189,0,97,0,243,0,116,0,246,0,84,0,0,0,66,0,152,0,87,0,52,0,104,0,218,0,165,0,102,0,88,0,172,0,188,0,21,0,182,0,190,0,206,0,209,0,193,0,0,0,176,0,0,0,205,0,144,0,54,0,148,0,163,0,78,0,167,0,96,0,22,0,68,0,220,0,244,0,39,0,65,0,212,0,89,0,0,0,68,0,30,0,90,0,236,0,198,0,67,0,49,0,184,0,33,0,0,0,0,0,0,0,15,0,0,0,126,0,29,0,0,0,0,0,110,0,51,0,237,0,195,0,158,0,159,0,129,0,0,0,174,0,248,0,73,0,0,0,134,0,249,0,130,0,20,0,24,0,196,0,0,0,0,0,145,0,92,0,79,0,196,0,133,0,142,0,146,0,95,0,27,0,205,0,30,0,232,0,144,0,0,0,22,0,155,0,0,0,50,0,161,0,0,0,80,0,161,0,100,0,0,0,193,0,156,0,0,0,0,0,36,0,197,0,198,0,235,0,236,0,143,0,0,0,143,0,0,0,180,0,0,0,238,0,165,0,173,0,81,0,198,0,89,0,230,0,217,0,44,0,76,0,0,0,141,0,0,0,73,0,159,0,115,0,146,0,229,0,176,0,206,0,84,0,73,0,33,0,202,0,36,0,2,0,234,0,0,0,224,0,16,0,84,0,147,0,29,0,225,0,176,0,0,0,0,0,228,0,157,0,144,0,0,0,109,0,9,0,0,0,148,0,96,0,157,0,113,0,166,0,210,0,136,0,0,0,100,0,151,0,31,0,0,0,84,0,169,0,0,0,59,0,233,0,0,0,158,0,213,0,0,0,166,0,0,0,157,0,155,0,209,0,3,0,188,0,198,0,50,0,13,0,73,0,230,0,0,0,214,0,223,0,205,0,102,0,241,0,81,0,105,0,207,0,26,0,108,0,88,0,22,0,104,0,91,0,0,0,237,0,160,0,28,0,197,0,174,0,0,0,0,0,202,0,237,0,0,0,0,0,80,0,152,0,0,0,159,0,71,0,215,0,0,0,155,0,184,0,160,0,98,0,0,0,0,0,206,0,94,0,223,0,0,0,8,0,181,0,247,0,0,0,71,0,191,0,168,0,156,0,152,0,250,0,0,0,5,0,249,0,46,0,239,0,135,0,83,0,209,0,0,0,129,0,64,0,219,0,129,0,70,0,66,0,111,0,252,0,217,0,0,0,163,0,171,0,205,0,141,0,5,0,232,0,0,0,74,0,7,0,182,0,68,0,100,0,207,0,172,0,158,0,165,0,159,0,0,0,25,0,187,0,123,0,1,0,0,0,164,0,209,0,173,0,229,0,141,0,85,0,165,0,145,0,105,0,165,0,107,0,0,0,144,0,0,0,104,0,36,0,24,0,146,0,0,0,93,0,10,0,192,0,0,0,120,0,15,0,184,0,205,0,171,0,76,0,0,0,94,0,7,0,88,0,29,0,6,0,0,0,42,0,42,0,0,0,0,0,95,0,142,0,235,0,114,0,148,0,78,0,60,0,130,0,143,0,77,0,0,0,229,0,4,0,0,0,72,0,122,0,0,0,171,0,135,0,0,0,169,0,0,0,67,0,145,0,238,0,217,0,0,0,22,0,15,0,148,0,187,0,61,0,0,0,0,0,122,0,36,0,61,0,0,0,18,0,0,0,217,0,46,0,114,0,184,0,0,0,0,0,0,0,31,0,114,0,130,0,31,0,0,0,197,0,0,0,94,0,60,0,100,0,197,0,0,0,0,0,0,0,242,0,106,0,0,0,0,0,57,0,34,0,19,0,250,0,25,0,0,0,35,0,89,0,0,0,195,0,96,0,42,0,130,0,78,0,0,0,220,0,70,0,0,0,229,0,169,0,113,0,77,0,199,0,247,0,57,0,26,0,34,0,0,0,235,0,172,0,217,0,22,0,16,0,0,0,0,0,122,0,221,0,124,0,0,0,153,0,0,0,0,0,194,0,209,0,0,0,0,0,6,0,246,0,50,0,0,0,99,0,115,0,235,0,95,0,153,0,72,0,166,0,1,0,235,0,0,0,87,0,201,0,85,0,79,0,13,0,0,0,0,0,221,0,135,0,185,0,0,0,31,0,34,0,167,0,0,0,151,0,79,0,86,0,58,0,136,0,202,0,141,0,85,0,93,0,51,0,0,0,5,0,69,0,50,0,20,0,188,0,114,0,0,0,149,0,51,0,173,0,208,0,0,0,104,0,48,0,0,0,92,0,62,0,16,0,183,0,227,0,82,0,240,0,46,0,137,0,218,0,204,0,56,0,80,0,99,0,65,0,204,0,156,0,214,0,161,0,70,0,164,0,6,0,208,0,80,0,0,0,0,0,145,0,147,0,254,0,211,0,0,0,44,0,202,0,31,0,0,0,16,0,244,0,140,0,134,0,46,0,245,0,0,0,187,0,237,0,0,0,36,0,206,0,104,0,152,0,143,0,0,0,130,0,0,0,48,0,86,0,0,0,154,0,97,0,32,0,227,0,1,0,21,0,168,0,6,0,0,0,241,0,72,0,53,0,0,0,0,0,248,0,155,0,176,0,217,0,0,0,98,0,83,0,225,0,206,0,204,0,60,0,0,0,154,0,37,0,133,0,68,0,0,0,166,0,213,0,15,0,182,0,190,0,57,0,30,0,44,0,0,0,111,0,121,0,169,0,231,0,0,0,181,0,202,0,87,0,0,0,81,0,196,0,80,0,234,0,27,0,251,0,0,0,0,0,70,0,0,0,190,0,0,0,205,0,4,0,62,0,0,0,0,0,42,0,178,0,195,0,212,0);
signal scenario_full  : scenario_type := (210,31,252,31,88,31,183,31,192,31,177,31,124,31,124,30,124,29,189,31,94,31,94,30,94,29,242,31,199,31,199,30,158,31,116,31,116,30,116,29,81,31,81,30,109,31,109,30,222,31,255,31,255,30,255,29,32,31,32,30,254,31,18,31,18,30,177,31,252,31,12,31,12,30,227,31,94,31,148,31,9,31,189,31,29,31,29,30,184,31,253,31,227,31,213,31,106,31,101,31,101,30,101,29,22,31,253,31,83,31,194,31,53,31,185,31,185,30,184,31,162,31,179,31,71,31,126,31,46,31,33,31,56,31,56,30,226,31,120,31,18,31,249,31,249,30,230,31,230,30,197,31,33,31,33,30,33,29,68,31,165,31,34,31,227,31,137,31,182,31,236,31,236,30,236,29,124,31,153,31,223,31,133,31,130,31,224,31,194,31,239,31,254,31,113,31,123,31,244,31,244,30,15,31,254,31,133,31,192,31,140,31,140,30,13,31,212,31,103,31,237,31,37,31,37,30,216,31,216,30,114,31,97,31,166,31,166,30,110,31,170,31,73,31,15,31,15,30,31,31,37,31,120,31,120,30,166,31,166,30,119,31,254,31,154,31,174,31,118,31,234,31,58,31,58,30,169,31,35,31,201,31,230,31,82,31,141,31,141,30,196,31,39,31,39,30,39,29,39,28,114,31,114,30,47,31,47,30,65,31,54,31,157,31,245,31,181,31,181,30,16,31,178,31,137,31,144,31,175,31,157,31,104,31,114,31,114,30,189,31,97,31,243,31,116,31,246,31,84,31,84,30,66,31,152,31,87,31,52,31,104,31,218,31,165,31,102,31,88,31,172,31,188,31,21,31,182,31,190,31,206,31,209,31,193,31,193,30,176,31,176,30,205,31,144,31,54,31,148,31,163,31,78,31,167,31,96,31,22,31,68,31,220,31,244,31,39,31,65,31,212,31,89,31,89,30,68,31,30,31,90,31,236,31,198,31,67,31,49,31,184,31,33,31,33,30,33,29,33,28,15,31,15,30,126,31,29,31,29,30,29,29,110,31,51,31,237,31,195,31,158,31,159,31,129,31,129,30,174,31,248,31,73,31,73,30,134,31,249,31,130,31,20,31,24,31,196,31,196,30,196,29,145,31,92,31,79,31,196,31,133,31,142,31,146,31,95,31,27,31,205,31,30,31,232,31,144,31,144,30,22,31,155,31,155,30,50,31,161,31,161,30,80,31,161,31,100,31,100,30,193,31,156,31,156,30,156,29,36,31,197,31,198,31,235,31,236,31,143,31,143,30,143,31,143,30,180,31,180,30,238,31,165,31,173,31,81,31,198,31,89,31,230,31,217,31,44,31,76,31,76,30,141,31,141,30,73,31,159,31,115,31,146,31,229,31,176,31,206,31,84,31,73,31,33,31,202,31,36,31,2,31,234,31,234,30,224,31,16,31,84,31,147,31,29,31,225,31,176,31,176,30,176,29,228,31,157,31,144,31,144,30,109,31,9,31,9,30,148,31,96,31,157,31,113,31,166,31,210,31,136,31,136,30,100,31,151,31,31,31,31,30,84,31,169,31,169,30,59,31,233,31,233,30,158,31,213,31,213,30,166,31,166,30,157,31,155,31,209,31,3,31,188,31,198,31,50,31,13,31,73,31,230,31,230,30,214,31,223,31,205,31,102,31,241,31,81,31,105,31,207,31,26,31,108,31,88,31,22,31,104,31,91,31,91,30,237,31,160,31,28,31,197,31,174,31,174,30,174,29,202,31,237,31,237,30,237,29,80,31,152,31,152,30,159,31,71,31,215,31,215,30,155,31,184,31,160,31,98,31,98,30,98,29,206,31,94,31,223,31,223,30,8,31,181,31,247,31,247,30,71,31,191,31,168,31,156,31,152,31,250,31,250,30,5,31,249,31,46,31,239,31,135,31,83,31,209,31,209,30,129,31,64,31,219,31,129,31,70,31,66,31,111,31,252,31,217,31,217,30,163,31,171,31,205,31,141,31,5,31,232,31,232,30,74,31,7,31,182,31,68,31,100,31,207,31,172,31,158,31,165,31,159,31,159,30,25,31,187,31,123,31,1,31,1,30,164,31,209,31,173,31,229,31,141,31,85,31,165,31,145,31,105,31,165,31,107,31,107,30,144,31,144,30,104,31,36,31,24,31,146,31,146,30,93,31,10,31,192,31,192,30,120,31,15,31,184,31,205,31,171,31,76,31,76,30,94,31,7,31,88,31,29,31,6,31,6,30,42,31,42,31,42,30,42,29,95,31,142,31,235,31,114,31,148,31,78,31,60,31,130,31,143,31,77,31,77,30,229,31,4,31,4,30,72,31,122,31,122,30,171,31,135,31,135,30,169,31,169,30,67,31,145,31,238,31,217,31,217,30,22,31,15,31,148,31,187,31,61,31,61,30,61,29,122,31,36,31,61,31,61,30,18,31,18,30,217,31,46,31,114,31,184,31,184,30,184,29,184,28,31,31,114,31,130,31,31,31,31,30,197,31,197,30,94,31,60,31,100,31,197,31,197,30,197,29,197,28,242,31,106,31,106,30,106,29,57,31,34,31,19,31,250,31,25,31,25,30,35,31,89,31,89,30,195,31,96,31,42,31,130,31,78,31,78,30,220,31,70,31,70,30,229,31,169,31,113,31,77,31,199,31,247,31,57,31,26,31,34,31,34,30,235,31,172,31,217,31,22,31,16,31,16,30,16,29,122,31,221,31,124,31,124,30,153,31,153,30,153,29,194,31,209,31,209,30,209,29,6,31,246,31,50,31,50,30,99,31,115,31,235,31,95,31,153,31,72,31,166,31,1,31,235,31,235,30,87,31,201,31,85,31,79,31,13,31,13,30,13,29,221,31,135,31,185,31,185,30,31,31,34,31,167,31,167,30,151,31,79,31,86,31,58,31,136,31,202,31,141,31,85,31,93,31,51,31,51,30,5,31,69,31,50,31,20,31,188,31,114,31,114,30,149,31,51,31,173,31,208,31,208,30,104,31,48,31,48,30,92,31,62,31,16,31,183,31,227,31,82,31,240,31,46,31,137,31,218,31,204,31,56,31,80,31,99,31,65,31,204,31,156,31,214,31,161,31,70,31,164,31,6,31,208,31,80,31,80,30,80,29,145,31,147,31,254,31,211,31,211,30,44,31,202,31,31,31,31,30,16,31,244,31,140,31,134,31,46,31,245,31,245,30,187,31,237,31,237,30,36,31,206,31,104,31,152,31,143,31,143,30,130,31,130,30,48,31,86,31,86,30,154,31,97,31,32,31,227,31,1,31,21,31,168,31,6,31,6,30,241,31,72,31,53,31,53,30,53,29,248,31,155,31,176,31,217,31,217,30,98,31,83,31,225,31,206,31,204,31,60,31,60,30,154,31,37,31,133,31,68,31,68,30,166,31,213,31,15,31,182,31,190,31,57,31,30,31,44,31,44,30,111,31,121,31,169,31,231,31,231,30,181,31,202,31,87,31,87,30,81,31,196,31,80,31,234,31,27,31,251,31,251,30,251,29,70,31,70,30,190,31,190,30,205,31,4,31,62,31,62,30,62,29,42,31,178,31,195,31,212,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
