-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 638;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (76,0,10,0,0,0,219,0,52,0,0,0,4,0,0,0,206,0,177,0,74,0,22,0,55,0,231,0,0,0,125,0,35,0,23,0,0,0,53,0,190,0,0,0,240,0,126,0,28,0,0,0,255,0,61,0,61,0,0,0,43,0,104,0,58,0,89,0,0,0,143,0,82,0,75,0,0,0,209,0,62,0,235,0,25,0,250,0,171,0,21,0,193,0,0,0,124,0,36,0,254,0,0,0,71,0,0,0,241,0,87,0,117,0,34,0,0,0,0,0,186,0,43,0,239,0,215,0,101,0,126,0,0,0,136,0,23,0,174,0,107,0,144,0,135,0,238,0,94,0,230,0,183,0,218,0,226,0,15,0,0,0,117,0,0,0,147,0,65,0,15,0,96,0,153,0,1,0,120,0,228,0,0,0,181,0,164,0,0,0,251,0,224,0,125,0,32,0,34,0,155,0,0,0,151,0,189,0,196,0,164,0,242,0,171,0,122,0,188,0,66,0,146,0,210,0,152,0,252,0,105,0,28,0,85,0,38,0,186,0,76,0,52,0,9,0,93,0,165,0,138,0,242,0,197,0,0,0,26,0,0,0,184,0,0,0,0,0,209,0,0,0,92,0,75,0,0,0,112,0,179,0,86,0,0,0,21,0,0,0,0,0,0,0,137,0,81,0,178,0,202,0,208,0,49,0,182,0,142,0,1,0,63,0,210,0,242,0,85,0,17,0,225,0,240,0,203,0,208,0,140,0,119,0,142,0,0,0,196,0,191,0,240,0,33,0,4,0,150,0,123,0,81,0,1,0,9,0,235,0,0,0,170,0,185,0,173,0,203,0,150,0,149,0,0,0,0,0,243,0,4,0,224,0,0,0,94,0,36,0,186,0,132,0,88,0,220,0,0,0,87,0,224,0,208,0,246,0,0,0,185,0,248,0,0,0,161,0,118,0,183,0,175,0,146,0,18,0,167,0,57,0,158,0,222,0,138,0,219,0,255,0,132,0,235,0,220,0,186,0,104,0,198,0,0,0,0,0,126,0,255,0,0,0,136,0,39,0,223,0,27,0,102,0,98,0,157,0,226,0,33,0,175,0,151,0,32,0,77,0,188,0,227,0,91,0,254,0,239,0,169,0,40,0,0,0,52,0,202,0,73,0,200,0,0,0,0,0,156,0,100,0,235,0,186,0,164,0,137,0,210,0,0,0,189,0,189,0,66,0,30,0,36,0,0,0,33,0,217,0,235,0,116,0,157,0,33,0,104,0,0,0,59,0,75,0,0,0,0,0,54,0,52,0,99,0,111,0,0,0,0,0,0,0,0,0,118,0,123,0,38,0,93,0,43,0,153,0,84,0,0,0,239,0,51,0,255,0,106,0,103,0,192,0,0,0,29,0,0,0,0,0,41,0,120,0,104,0,119,0,88,0,0,0,140,0,230,0,0,0,205,0,0,0,0,0,28,0,214,0,0,0,221,0,0,0,0,0,83,0,64,0,58,0,175,0,178,0,137,0,188,0,76,0,81,0,215,0,0,0,176,0,177,0,209,0,99,0,233,0,166,0,30,0,0,0,93,0,22,0,86,0,246,0,77,0,190,0,180,0,103,0,54,0,0,0,216,0,88,0,139,0,210,0,155,0,0,0,141,0,182,0,0,0,72,0,127,0,0,0,77,0,34,0,185,0,213,0,202,0,122,0,0,0,0,0,216,0,208,0,36,0,255,0,81,0,0,0,0,0,165,0,194,0,0,0,213,0,0,0,251,0,51,0,0,0,9,0,64,0,148,0,220,0,83,0,0,0,40,0,153,0,23,0,117,0,146,0,149,0,0,0,96,0,0,0,61,0,200,0,34,0,0,0,131,0,0,0,188,0,0,0,110,0,206,0,30,0,0,0,172,0,122,0,0,0,36,0,0,0,212,0,81,0,172,0,0,0,220,0,230,0,168,0,186,0,150,0,0,0,88,0,0,0,169,0,120,0,49,0,2,0,0,0,155,0,40,0,39,0,0,0,191,0,71,0,32,0,0,0,95,0,251,0,7,0,55,0,0,0,158,0,245,0,4,0,0,0,149,0,0,0,87,0,211,0,0,0,236,0,160,0,211,0,0,0,0,0,91,0,249,0,75,0,94,0,220,0,75,0,0,0,0,0,181,0,25,0,156,0,136,0,27,0,0,0,191,0,102,0,154,0,0,0,16,0,55,0,85,0,118,0,166,0,3,0,163,0,49,0,30,0,0,0,0,0,170,0,209,0,0,0,21,0,190,0,248,0,124,0,13,0,210,0,93,0,33,0,10,0,0,0,20,0,158,0,39,0,139,0,21,0,210,0,109,0,0,0,160,0,224,0,0,0,111,0,0,0,170,0,225,0,68,0,51,0,153,0,175,0,245,0,0,0,2,0,173,0,186,0,251,0,216,0,117,0,186,0,149,0,215,0,1,0,125,0,185,0,0,0,96,0,196,0,242,0,67,0,96,0,223,0,148,0,30,0,212,0,231,0,136,0,147,0,0,0,0,0,148,0,136,0,0,0,225,0,0,0,196,0,252,0,213,0,74,0,102,0,0,0,185,0,60,0,167,0,119,0,97,0,0,0,240,0,244,0,251,0,87,0,163,0,48,0,196,0,13,0,232,0,212,0,232,0,19,0,41,0,227,0,233,0,25,0,232,0,200,0,0,0,90,0,86,0,166,0,8,0,225,0,24,0,14,0,99,0,145,0,67,0,0,0,0,0,111,0,0,0,145,0,0,0,0,0,216,0,0,0,188,0,182,0,171,0,0,0,15,0,229,0,0,0,0,0,195,0,238,0,33,0,200,0,0,0,236,0,0,0,131,0,129,0,0,0,153,0,45,0,65,0,133,0,109,0,81,0);
signal scenario_full  : scenario_type := (76,31,10,31,10,30,219,31,52,31,52,30,4,31,4,30,206,31,177,31,74,31,22,31,55,31,231,31,231,30,125,31,35,31,23,31,23,30,53,31,190,31,190,30,240,31,126,31,28,31,28,30,255,31,61,31,61,31,61,30,43,31,104,31,58,31,89,31,89,30,143,31,82,31,75,31,75,30,209,31,62,31,235,31,25,31,250,31,171,31,21,31,193,31,193,30,124,31,36,31,254,31,254,30,71,31,71,30,241,31,87,31,117,31,34,31,34,30,34,29,186,31,43,31,239,31,215,31,101,31,126,31,126,30,136,31,23,31,174,31,107,31,144,31,135,31,238,31,94,31,230,31,183,31,218,31,226,31,15,31,15,30,117,31,117,30,147,31,65,31,15,31,96,31,153,31,1,31,120,31,228,31,228,30,181,31,164,31,164,30,251,31,224,31,125,31,32,31,34,31,155,31,155,30,151,31,189,31,196,31,164,31,242,31,171,31,122,31,188,31,66,31,146,31,210,31,152,31,252,31,105,31,28,31,85,31,38,31,186,31,76,31,52,31,9,31,93,31,165,31,138,31,242,31,197,31,197,30,26,31,26,30,184,31,184,30,184,29,209,31,209,30,92,31,75,31,75,30,112,31,179,31,86,31,86,30,21,31,21,30,21,29,21,28,137,31,81,31,178,31,202,31,208,31,49,31,182,31,142,31,1,31,63,31,210,31,242,31,85,31,17,31,225,31,240,31,203,31,208,31,140,31,119,31,142,31,142,30,196,31,191,31,240,31,33,31,4,31,150,31,123,31,81,31,1,31,9,31,235,31,235,30,170,31,185,31,173,31,203,31,150,31,149,31,149,30,149,29,243,31,4,31,224,31,224,30,94,31,36,31,186,31,132,31,88,31,220,31,220,30,87,31,224,31,208,31,246,31,246,30,185,31,248,31,248,30,161,31,118,31,183,31,175,31,146,31,18,31,167,31,57,31,158,31,222,31,138,31,219,31,255,31,132,31,235,31,220,31,186,31,104,31,198,31,198,30,198,29,126,31,255,31,255,30,136,31,39,31,223,31,27,31,102,31,98,31,157,31,226,31,33,31,175,31,151,31,32,31,77,31,188,31,227,31,91,31,254,31,239,31,169,31,40,31,40,30,52,31,202,31,73,31,200,31,200,30,200,29,156,31,100,31,235,31,186,31,164,31,137,31,210,31,210,30,189,31,189,31,66,31,30,31,36,31,36,30,33,31,217,31,235,31,116,31,157,31,33,31,104,31,104,30,59,31,75,31,75,30,75,29,54,31,52,31,99,31,111,31,111,30,111,29,111,28,111,27,118,31,123,31,38,31,93,31,43,31,153,31,84,31,84,30,239,31,51,31,255,31,106,31,103,31,192,31,192,30,29,31,29,30,29,29,41,31,120,31,104,31,119,31,88,31,88,30,140,31,230,31,230,30,205,31,205,30,205,29,28,31,214,31,214,30,221,31,221,30,221,29,83,31,64,31,58,31,175,31,178,31,137,31,188,31,76,31,81,31,215,31,215,30,176,31,177,31,209,31,99,31,233,31,166,31,30,31,30,30,93,31,22,31,86,31,246,31,77,31,190,31,180,31,103,31,54,31,54,30,216,31,88,31,139,31,210,31,155,31,155,30,141,31,182,31,182,30,72,31,127,31,127,30,77,31,34,31,185,31,213,31,202,31,122,31,122,30,122,29,216,31,208,31,36,31,255,31,81,31,81,30,81,29,165,31,194,31,194,30,213,31,213,30,251,31,51,31,51,30,9,31,64,31,148,31,220,31,83,31,83,30,40,31,153,31,23,31,117,31,146,31,149,31,149,30,96,31,96,30,61,31,200,31,34,31,34,30,131,31,131,30,188,31,188,30,110,31,206,31,30,31,30,30,172,31,122,31,122,30,36,31,36,30,212,31,81,31,172,31,172,30,220,31,230,31,168,31,186,31,150,31,150,30,88,31,88,30,169,31,120,31,49,31,2,31,2,30,155,31,40,31,39,31,39,30,191,31,71,31,32,31,32,30,95,31,251,31,7,31,55,31,55,30,158,31,245,31,4,31,4,30,149,31,149,30,87,31,211,31,211,30,236,31,160,31,211,31,211,30,211,29,91,31,249,31,75,31,94,31,220,31,75,31,75,30,75,29,181,31,25,31,156,31,136,31,27,31,27,30,191,31,102,31,154,31,154,30,16,31,55,31,85,31,118,31,166,31,3,31,163,31,49,31,30,31,30,30,30,29,170,31,209,31,209,30,21,31,190,31,248,31,124,31,13,31,210,31,93,31,33,31,10,31,10,30,20,31,158,31,39,31,139,31,21,31,210,31,109,31,109,30,160,31,224,31,224,30,111,31,111,30,170,31,225,31,68,31,51,31,153,31,175,31,245,31,245,30,2,31,173,31,186,31,251,31,216,31,117,31,186,31,149,31,215,31,1,31,125,31,185,31,185,30,96,31,196,31,242,31,67,31,96,31,223,31,148,31,30,31,212,31,231,31,136,31,147,31,147,30,147,29,148,31,136,31,136,30,225,31,225,30,196,31,252,31,213,31,74,31,102,31,102,30,185,31,60,31,167,31,119,31,97,31,97,30,240,31,244,31,251,31,87,31,163,31,48,31,196,31,13,31,232,31,212,31,232,31,19,31,41,31,227,31,233,31,25,31,232,31,200,31,200,30,90,31,86,31,166,31,8,31,225,31,24,31,14,31,99,31,145,31,67,31,67,30,67,29,111,31,111,30,145,31,145,30,145,29,216,31,216,30,188,31,182,31,171,31,171,30,15,31,229,31,229,30,229,29,195,31,238,31,33,31,200,31,200,30,236,31,236,30,131,31,129,31,129,30,153,31,45,31,65,31,133,31,109,31,81,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
