-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_838 is
end project_tb_838;

architecture project_tb_arch_838 of project_tb_838 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 721;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (151,0,98,0,135,0,233,0,0,0,0,0,61,0,177,0,172,0,136,0,54,0,62,0,134,0,244,0,93,0,193,0,137,0,94,0,0,0,0,0,168,0,70,0,202,0,174,0,0,0,168,0,0,0,0,0,45,0,67,0,118,0,108,0,137,0,133,0,55,0,167,0,0,0,0,0,100,0,0,0,228,0,83,0,223,0,5,0,0,0,0,0,143,0,90,0,0,0,95,0,212,0,44,0,130,0,233,0,219,0,160,0,145,0,98,0,105,0,151,0,123,0,168,0,115,0,0,0,132,0,66,0,159,0,0,0,235,0,134,0,0,0,0,0,91,0,3,0,0,0,53,0,221,0,168,0,29,0,150,0,5,0,0,0,0,0,0,0,131,0,0,0,0,0,0,0,205,0,43,0,0,0,71,0,94,0,101,0,191,0,203,0,157,0,0,0,0,0,220,0,7,0,157,0,0,0,184,0,0,0,249,0,213,0,134,0,22,0,194,0,56,0,224,0,0,0,0,0,255,0,179,0,0,0,113,0,186,0,35,0,132,0,255,0,141,0,160,0,86,0,0,0,118,0,230,0,0,0,162,0,0,0,0,0,149,0,125,0,0,0,238,0,60,0,206,0,215,0,13,0,84,0,0,0,138,0,0,0,235,0,237,0,236,0,46,0,205,0,4,0,0,0,199,0,27,0,0,0,244,0,185,0,71,0,167,0,80,0,186,0,0,0,0,0,78,0,0,0,0,0,205,0,73,0,157,0,125,0,10,0,180,0,75,0,0,0,0,0,222,0,62,0,82,0,156,0,0,0,0,0,201,0,0,0,0,0,82,0,0,0,0,0,0,0,112,0,0,0,0,0,195,0,2,0,248,0,223,0,123,0,0,0,2,0,27,0,57,0,145,0,47,0,128,0,0,0,239,0,243,0,150,0,194,0,0,0,234,0,39,0,0,0,144,0,66,0,146,0,0,0,112,0,210,0,0,0,250,0,204,0,217,0,82,0,136,0,0,0,0,0,147,0,147,0,158,0,131,0,49,0,136,0,189,0,192,0,237,0,183,0,50,0,125,0,227,0,94,0,0,0,136,0,28,0,197,0,0,0,225,0,14,0,6,0,38,0,67,0,87,0,156,0,130,0,32,0,0,0,99,0,101,0,235,0,73,0,248,0,117,0,0,0,0,0,180,0,119,0,5,0,185,0,0,0,101,0,49,0,101,0,207,0,247,0,187,0,0,0,234,0,103,0,145,0,0,0,40,0,157,0,104,0,0,0,160,0,243,0,169,0,91,0,191,0,169,0,219,0,165,0,71,0,118,0,0,0,95,0,122,0,19,0,255,0,210,0,144,0,177,0,143,0,0,0,252,0,247,0,115,0,0,0,158,0,171,0,120,0,0,0,0,0,223,0,32,0,61,0,6,0,0,0,20,0,0,0,42,0,0,0,30,0,0,0,120,0,62,0,0,0,240,0,87,0,129,0,0,0,37,0,143,0,0,0,180,0,156,0,11,0,93,0,136,0,227,0,151,0,89,0,10,0,180,0,244,0,157,0,202,0,192,0,218,0,226,0,35,0,31,0,0,0,173,0,0,0,104,0,106,0,53,0,99,0,248,0,228,0,151,0,96,0,68,0,214,0,112,0,186,0,0,0,140,0,0,0,239,0,0,0,0,0,228,0,208,0,0,0,134,0,238,0,94,0,20,0,0,0,0,0,0,0,0,0,187,0,0,0,0,0,196,0,187,0,136,0,0,0,26,0,0,0,0,0,44,0,147,0,91,0,215,0,8,0,212,0,0,0,41,0,11,0,111,0,226,0,0,0,0,0,0,0,0,0,0,0,224,0,0,0,151,0,0,0,96,0,253,0,191,0,49,0,101,0,141,0,0,0,0,0,37,0,150,0,244,0,32,0,11,0,34,0,138,0,8,0,229,0,86,0,102,0,168,0,17,0,0,0,15,0,45,0,122,0,86,0,65,0,0,0,157,0,221,0,96,0,78,0,31,0,60,0,152,0,48,0,136,0,120,0,62,0,23,0,204,0,59,0,191,0,50,0,0,0,118,0,9,0,23,0,65,0,21,0,0,0,37,0,11,0,132,0,229,0,197,0,143,0,0,0,187,0,113,0,161,0,149,0,27,0,206,0,82,0,78,0,23,0,47,0,42,0,110,0,202,0,223,0,0,0,151,0,54,0,66,0,97,0,250,0,0,0,16,0,0,0,197,0,107,0,128,0,118,0,0,0,0,0,46,0,185,0,170,0,163,0,6,0,82,0,103,0,24,0,84,0,188,0,60,0,67,0,67,0,184,0,212,0,58,0,253,0,87,0,155,0,182,0,145,0,0,0,64,0,155,0,135,0,183,0,155,0,185,0,0,0,2,0,0,0,82,0,115,0,53,0,142,0,97,0,175,0,0,0,197,0,2,0,10,0,0,0,189,0,99,0,150,0,254,0,0,0,36,0,75,0,214,0,92,0,198,0,93,0,176,0,0,0,27,0,234,0,248,0,71,0,186,0,47,0,40,0,0,0,247,0,240,0,207,0,158,0,103,0,121,0,245,0,0,0,16,0,152,0,30,0,4,0,45,0,0,0,98,0,126,0,115,0,138,0,141,0,200,0,193,0,0,0,10,0,0,0,117,0,0,0,105,0,249,0,0,0,137,0,44,0,126,0,184,0,60,0,223,0,18,0,30,0,109,0,0,0,189,0,84,0,201,0,188,0,7,0,50,0,154,0,3,0,190,0,238,0,31,0,0,0,151,0,0,0,247,0,121,0,162,0,137,0,153,0,189,0,196,0,218,0,88,0,185,0,20,0,0,0,70,0,42,0,90,0,235,0,0,0,173,0,179,0,0,0,76,0,119,0,165,0,0,0,118,0,9,0,17,0,164,0,14,0,137,0,88,0,135,0,0,0,222,0,202,0,230,0,253,0,163,0,165,0,103,0,0,0,182,0,0,0,10,0,194,0,227,0,53,0,187,0,102,0,5,0,153,0,237,0,219,0,209,0,128,0,0,0,0,0,0,0,0,0,3,0,181,0,118,0,224,0,92,0,0,0,139,0,0,0,97,0,144,0,85,0,140,0,241,0,125,0,142,0,171,0,0,0,152,0,119,0,120,0,99,0,209,0,242,0,97,0,227,0,72,0,204,0,0,0,197,0,250,0,5,0,0,0,0,0,122,0,183,0,3,0,195,0,0,0,88,0,0,0,183,0,143,0,203,0,164,0,175,0,181,0,199,0);
signal scenario_full  : scenario_type := (151,31,98,31,135,31,233,31,233,30,233,29,61,31,177,31,172,31,136,31,54,31,62,31,134,31,244,31,93,31,193,31,137,31,94,31,94,30,94,29,168,31,70,31,202,31,174,31,174,30,168,31,168,30,168,29,45,31,67,31,118,31,108,31,137,31,133,31,55,31,167,31,167,30,167,29,100,31,100,30,228,31,83,31,223,31,5,31,5,30,5,29,143,31,90,31,90,30,95,31,212,31,44,31,130,31,233,31,219,31,160,31,145,31,98,31,105,31,151,31,123,31,168,31,115,31,115,30,132,31,66,31,159,31,159,30,235,31,134,31,134,30,134,29,91,31,3,31,3,30,53,31,221,31,168,31,29,31,150,31,5,31,5,30,5,29,5,28,131,31,131,30,131,29,131,28,205,31,43,31,43,30,71,31,94,31,101,31,191,31,203,31,157,31,157,30,157,29,220,31,7,31,157,31,157,30,184,31,184,30,249,31,213,31,134,31,22,31,194,31,56,31,224,31,224,30,224,29,255,31,179,31,179,30,113,31,186,31,35,31,132,31,255,31,141,31,160,31,86,31,86,30,118,31,230,31,230,30,162,31,162,30,162,29,149,31,125,31,125,30,238,31,60,31,206,31,215,31,13,31,84,31,84,30,138,31,138,30,235,31,237,31,236,31,46,31,205,31,4,31,4,30,199,31,27,31,27,30,244,31,185,31,71,31,167,31,80,31,186,31,186,30,186,29,78,31,78,30,78,29,205,31,73,31,157,31,125,31,10,31,180,31,75,31,75,30,75,29,222,31,62,31,82,31,156,31,156,30,156,29,201,31,201,30,201,29,82,31,82,30,82,29,82,28,112,31,112,30,112,29,195,31,2,31,248,31,223,31,123,31,123,30,2,31,27,31,57,31,145,31,47,31,128,31,128,30,239,31,243,31,150,31,194,31,194,30,234,31,39,31,39,30,144,31,66,31,146,31,146,30,112,31,210,31,210,30,250,31,204,31,217,31,82,31,136,31,136,30,136,29,147,31,147,31,158,31,131,31,49,31,136,31,189,31,192,31,237,31,183,31,50,31,125,31,227,31,94,31,94,30,136,31,28,31,197,31,197,30,225,31,14,31,6,31,38,31,67,31,87,31,156,31,130,31,32,31,32,30,99,31,101,31,235,31,73,31,248,31,117,31,117,30,117,29,180,31,119,31,5,31,185,31,185,30,101,31,49,31,101,31,207,31,247,31,187,31,187,30,234,31,103,31,145,31,145,30,40,31,157,31,104,31,104,30,160,31,243,31,169,31,91,31,191,31,169,31,219,31,165,31,71,31,118,31,118,30,95,31,122,31,19,31,255,31,210,31,144,31,177,31,143,31,143,30,252,31,247,31,115,31,115,30,158,31,171,31,120,31,120,30,120,29,223,31,32,31,61,31,6,31,6,30,20,31,20,30,42,31,42,30,30,31,30,30,120,31,62,31,62,30,240,31,87,31,129,31,129,30,37,31,143,31,143,30,180,31,156,31,11,31,93,31,136,31,227,31,151,31,89,31,10,31,180,31,244,31,157,31,202,31,192,31,218,31,226,31,35,31,31,31,31,30,173,31,173,30,104,31,106,31,53,31,99,31,248,31,228,31,151,31,96,31,68,31,214,31,112,31,186,31,186,30,140,31,140,30,239,31,239,30,239,29,228,31,208,31,208,30,134,31,238,31,94,31,20,31,20,30,20,29,20,28,20,27,187,31,187,30,187,29,196,31,187,31,136,31,136,30,26,31,26,30,26,29,44,31,147,31,91,31,215,31,8,31,212,31,212,30,41,31,11,31,111,31,226,31,226,30,226,29,226,28,226,27,226,26,224,31,224,30,151,31,151,30,96,31,253,31,191,31,49,31,101,31,141,31,141,30,141,29,37,31,150,31,244,31,32,31,11,31,34,31,138,31,8,31,229,31,86,31,102,31,168,31,17,31,17,30,15,31,45,31,122,31,86,31,65,31,65,30,157,31,221,31,96,31,78,31,31,31,60,31,152,31,48,31,136,31,120,31,62,31,23,31,204,31,59,31,191,31,50,31,50,30,118,31,9,31,23,31,65,31,21,31,21,30,37,31,11,31,132,31,229,31,197,31,143,31,143,30,187,31,113,31,161,31,149,31,27,31,206,31,82,31,78,31,23,31,47,31,42,31,110,31,202,31,223,31,223,30,151,31,54,31,66,31,97,31,250,31,250,30,16,31,16,30,197,31,107,31,128,31,118,31,118,30,118,29,46,31,185,31,170,31,163,31,6,31,82,31,103,31,24,31,84,31,188,31,60,31,67,31,67,31,184,31,212,31,58,31,253,31,87,31,155,31,182,31,145,31,145,30,64,31,155,31,135,31,183,31,155,31,185,31,185,30,2,31,2,30,82,31,115,31,53,31,142,31,97,31,175,31,175,30,197,31,2,31,10,31,10,30,189,31,99,31,150,31,254,31,254,30,36,31,75,31,214,31,92,31,198,31,93,31,176,31,176,30,27,31,234,31,248,31,71,31,186,31,47,31,40,31,40,30,247,31,240,31,207,31,158,31,103,31,121,31,245,31,245,30,16,31,152,31,30,31,4,31,45,31,45,30,98,31,126,31,115,31,138,31,141,31,200,31,193,31,193,30,10,31,10,30,117,31,117,30,105,31,249,31,249,30,137,31,44,31,126,31,184,31,60,31,223,31,18,31,30,31,109,31,109,30,189,31,84,31,201,31,188,31,7,31,50,31,154,31,3,31,190,31,238,31,31,31,31,30,151,31,151,30,247,31,121,31,162,31,137,31,153,31,189,31,196,31,218,31,88,31,185,31,20,31,20,30,70,31,42,31,90,31,235,31,235,30,173,31,179,31,179,30,76,31,119,31,165,31,165,30,118,31,9,31,17,31,164,31,14,31,137,31,88,31,135,31,135,30,222,31,202,31,230,31,253,31,163,31,165,31,103,31,103,30,182,31,182,30,10,31,194,31,227,31,53,31,187,31,102,31,5,31,153,31,237,31,219,31,209,31,128,31,128,30,128,29,128,28,128,27,3,31,181,31,118,31,224,31,92,31,92,30,139,31,139,30,97,31,144,31,85,31,140,31,241,31,125,31,142,31,171,31,171,30,152,31,119,31,120,31,99,31,209,31,242,31,97,31,227,31,72,31,204,31,204,30,197,31,250,31,5,31,5,30,5,29,122,31,183,31,3,31,195,31,195,30,88,31,88,30,183,31,143,31,203,31,164,31,175,31,181,31,199,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
