-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_140 is
end project_tb_140;

architecture project_tb_arch_140 of project_tb_140 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 790;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,0,0,0,0,138,0,0,0,51,0,45,0,38,0,154,0,180,0,102,0,189,0,12,0,36,0,0,0,235,0,20,0,122,0,51,0,106,0,237,0,152,0,0,0,0,0,90,0,217,0,38,0,0,0,155,0,147,0,205,0,254,0,94,0,125,0,89,0,59,0,154,0,188,0,71,0,175,0,0,0,188,0,104,0,190,0,0,0,6,0,3,0,101,0,112,0,180,0,196,0,0,0,240,0,0,0,215,0,85,0,0,0,47,0,202,0,73,0,30,0,0,0,190,0,120,0,206,0,179,0,253,0,73,0,143,0,0,0,16,0,124,0,187,0,60,0,33,0,0,0,8,0,0,0,0,0,64,0,37,0,109,0,0,0,11,0,0,0,123,0,0,0,185,0,53,0,115,0,0,0,62,0,0,0,4,0,227,0,119,0,8,0,82,0,4,0,83,0,115,0,53,0,0,0,27,0,0,0,231,0,71,0,199,0,145,0,206,0,177,0,126,0,17,0,153,0,1,0,135,0,33,0,38,0,22,0,22,0,0,0,0,0,54,0,148,0,11,0,165,0,222,0,136,0,76,0,44,0,220,0,98,0,155,0,249,0,77,0,0,0,0,0,214,0,252,0,42,0,203,0,186,0,106,0,210,0,16,0,191,0,0,0,194,0,2,0,0,0,36,0,236,0,213,0,38,0,191,0,0,0,0,0,136,0,117,0,129,0,192,0,0,0,0,0,0,0,207,0,0,0,0,0,7,0,86,0,90,0,59,0,110,0,0,0,0,0,173,0,77,0,108,0,0,0,0,0,167,0,249,0,0,0,245,0,209,0,0,0,0,0,180,0,0,0,115,0,65,0,0,0,145,0,0,0,146,0,201,0,83,0,0,0,247,0,109,0,17,0,94,0,70,0,183,0,55,0,249,0,197,0,0,0,125,0,41,0,167,0,146,0,6,0,9,0,131,0,0,0,156,0,86,0,48,0,66,0,243,0,136,0,0,0,177,0,188,0,159,0,194,0,160,0,132,0,89,0,222,0,0,0,85,0,0,0,12,0,155,0,141,0,31,0,199,0,193,0,74,0,108,0,28,0,216,0,16,0,0,0,68,0,173,0,239,0,69,0,0,0,149,0,3,0,219,0,50,0,126,0,142,0,0,0,101,0,43,0,202,0,0,0,0,0,105,0,51,0,214,0,0,0,188,0,40,0,123,0,0,0,0,0,45,0,0,0,243,0,182,0,199,0,240,0,22,0,107,0,163,0,209,0,216,0,0,0,0,0,37,0,184,0,203,0,140,0,0,0,46,0,97,0,125,0,46,0,91,0,140,0,50,0,112,0,63,0,139,0,0,0,0,0,47,0,152,0,0,0,0,0,26,0,43,0,204,0,0,0,123,0,19,0,170,0,54,0,164,0,187,0,167,0,18,0,116,0,112,0,0,0,34,0,0,0,0,0,251,0,145,0,174,0,134,0,200,0,0,0,128,0,0,0,240,0,85,0,122,0,85,0,117,0,165,0,51,0,244,0,102,0,83,0,72,0,76,0,126,0,99,0,216,0,0,0,185,0,0,0,45,0,218,0,78,0,0,0,126,0,0,0,212,0,171,0,182,0,161,0,72,0,0,0,250,0,242,0,7,0,0,0,96,0,6,0,0,0,228,0,183,0,174,0,255,0,24,0,100,0,230,0,0,0,18,0,102,0,78,0,47,0,0,0,197,0,166,0,125,0,48,0,45,0,188,0,87,0,0,0,0,0,49,0,171,0,0,0,12,0,13,0,57,0,102,0,0,0,0,0,87,0,0,0,151,0,80,0,0,0,8,0,0,0,0,0,136,0,251,0,44,0,90,0,0,0,204,0,146,0,127,0,187,0,133,0,0,0,34,0,0,0,67,0,55,0,25,0,173,0,35,0,89,0,221,0,22,0,0,0,145,0,4,0,41,0,54,0,86,0,140,0,38,0,0,0,0,0,52,0,225,0,25,0,173,0,0,0,121,0,82,0,25,0,86,0,42,0,129,0,72,0,241,0,192,0,139,0,46,0,89,0,68,0,0,0,144,0,23,0,137,0,0,0,138,0,163,0,0,0,133,0,88,0,0,0,0,0,138,0,22,0,0,0,101,0,40,0,84,0,101,0,0,0,0,0,0,0,196,0,126,0,0,0,144,0,65,0,39,0,48,0,116,0,126,0,106,0,105,0,0,0,140,0,0,0,35,0,0,0,25,0,223,0,88,0,130,0,16,0,99,0,36,0,15,0,233,0,137,0,209,0,0,0,234,0,129,0,0,0,105,0,146,0,104,0,0,0,139,0,217,0,54,0,60,0,239,0,116,0,68,0,11,0,0,0,0,0,52,0,252,0,189,0,53,0,94,0,149,0,0,0,0,0,130,0,160,0,23,0,0,0,0,0,215,0,66,0,0,0,215,0,97,0,135,0,0,0,234,0,147,0,236,0,1,0,69,0,105,0,101,0,90,0,0,0,231,0,130,0,81,0,124,0,250,0,117,0,0,0,151,0,0,0,0,0,119,0,135,0,9,0,219,0,25,0,87,0,36,0,137,0,185,0,224,0,193,0,189,0,181,0,193,0,0,0,55,0,0,0,94,0,239,0,181,0,174,0,128,0,176,0,224,0,0,0,161,0,113,0,160,0,96,0,22,0,0,0,57,0,86,0,143,0,104,0,43,0,0,0,253,0,14,0,154,0,0,0,48,0,151,0,121,0,202,0,96,0,121,0,166,0,176,0,129,0,0,0,0,0,124,0,98,0,131,0,0,0,22,0,242,0,0,0,61,0,163,0,57,0,0,0,170,0,127,0,190,0,0,0,65,0,61,0,108,0,0,0,90,0,221,0,206,0,191,0,15,0,123,0,7,0,50,0,54,0,253,0,140,0,0,0,0,0,119,0,116,0,133,0,133,0,171,0,0,0,14,0,59,0,27,0,80,0,57,0,175,0,0,0,101,0,0,0,0,0,148,0,19,0,0,0,165,0,64,0,86,0,120,0,91,0,179,0,188,0,242,0,0,0,218,0,212,0,144,0,28,0,148,0,0,0,250,0,83,0,222,0,205,0,108,0,152,0,231,0,92,0,108,0,132,0,0,0,148,0,0,0,0,0,4,0,202,0,133,0,0,0,166,0,0,0,229,0,80,0,86,0,186,0,162,0,33,0,99,0,3,0,0,0,247,0,66,0,181,0,171,0,194,0,3,0,0,0,92,0,193,0,109,0,153,0,0,0,208,0,122,0,67,0,101,0,0,0,78,0,0,0,0,0,124,0,168,0,0,0,76,0,152,0,242,0,20,0,3,0,90,0,110,0,217,0,104,0,0,0,38,0,0,0,82,0,108,0,0,0,198,0,245,0,165,0,0,0,254,0,137,0,146,0,255,0,146,0,132,0,49,0,50,0,162,0,163,0,0,0,43,0,222,0,46,0,194,0,0,0,197,0,53,0,32,0,0,0,0,0,97,0,212,0,184,0,104,0,86,0,0,0,194,0,163,0,44,0,0,0,0,0,0,0,180,0,74,0,150,0,241,0,0,0,117,0);
signal scenario_full  : scenario_type := (36,31,36,30,36,29,138,31,138,30,51,31,45,31,38,31,154,31,180,31,102,31,189,31,12,31,36,31,36,30,235,31,20,31,122,31,51,31,106,31,237,31,152,31,152,30,152,29,90,31,217,31,38,31,38,30,155,31,147,31,205,31,254,31,94,31,125,31,89,31,59,31,154,31,188,31,71,31,175,31,175,30,188,31,104,31,190,31,190,30,6,31,3,31,101,31,112,31,180,31,196,31,196,30,240,31,240,30,215,31,85,31,85,30,47,31,202,31,73,31,30,31,30,30,190,31,120,31,206,31,179,31,253,31,73,31,143,31,143,30,16,31,124,31,187,31,60,31,33,31,33,30,8,31,8,30,8,29,64,31,37,31,109,31,109,30,11,31,11,30,123,31,123,30,185,31,53,31,115,31,115,30,62,31,62,30,4,31,227,31,119,31,8,31,82,31,4,31,83,31,115,31,53,31,53,30,27,31,27,30,231,31,71,31,199,31,145,31,206,31,177,31,126,31,17,31,153,31,1,31,135,31,33,31,38,31,22,31,22,31,22,30,22,29,54,31,148,31,11,31,165,31,222,31,136,31,76,31,44,31,220,31,98,31,155,31,249,31,77,31,77,30,77,29,214,31,252,31,42,31,203,31,186,31,106,31,210,31,16,31,191,31,191,30,194,31,2,31,2,30,36,31,236,31,213,31,38,31,191,31,191,30,191,29,136,31,117,31,129,31,192,31,192,30,192,29,192,28,207,31,207,30,207,29,7,31,86,31,90,31,59,31,110,31,110,30,110,29,173,31,77,31,108,31,108,30,108,29,167,31,249,31,249,30,245,31,209,31,209,30,209,29,180,31,180,30,115,31,65,31,65,30,145,31,145,30,146,31,201,31,83,31,83,30,247,31,109,31,17,31,94,31,70,31,183,31,55,31,249,31,197,31,197,30,125,31,41,31,167,31,146,31,6,31,9,31,131,31,131,30,156,31,86,31,48,31,66,31,243,31,136,31,136,30,177,31,188,31,159,31,194,31,160,31,132,31,89,31,222,31,222,30,85,31,85,30,12,31,155,31,141,31,31,31,199,31,193,31,74,31,108,31,28,31,216,31,16,31,16,30,68,31,173,31,239,31,69,31,69,30,149,31,3,31,219,31,50,31,126,31,142,31,142,30,101,31,43,31,202,31,202,30,202,29,105,31,51,31,214,31,214,30,188,31,40,31,123,31,123,30,123,29,45,31,45,30,243,31,182,31,199,31,240,31,22,31,107,31,163,31,209,31,216,31,216,30,216,29,37,31,184,31,203,31,140,31,140,30,46,31,97,31,125,31,46,31,91,31,140,31,50,31,112,31,63,31,139,31,139,30,139,29,47,31,152,31,152,30,152,29,26,31,43,31,204,31,204,30,123,31,19,31,170,31,54,31,164,31,187,31,167,31,18,31,116,31,112,31,112,30,34,31,34,30,34,29,251,31,145,31,174,31,134,31,200,31,200,30,128,31,128,30,240,31,85,31,122,31,85,31,117,31,165,31,51,31,244,31,102,31,83,31,72,31,76,31,126,31,99,31,216,31,216,30,185,31,185,30,45,31,218,31,78,31,78,30,126,31,126,30,212,31,171,31,182,31,161,31,72,31,72,30,250,31,242,31,7,31,7,30,96,31,6,31,6,30,228,31,183,31,174,31,255,31,24,31,100,31,230,31,230,30,18,31,102,31,78,31,47,31,47,30,197,31,166,31,125,31,48,31,45,31,188,31,87,31,87,30,87,29,49,31,171,31,171,30,12,31,13,31,57,31,102,31,102,30,102,29,87,31,87,30,151,31,80,31,80,30,8,31,8,30,8,29,136,31,251,31,44,31,90,31,90,30,204,31,146,31,127,31,187,31,133,31,133,30,34,31,34,30,67,31,55,31,25,31,173,31,35,31,89,31,221,31,22,31,22,30,145,31,4,31,41,31,54,31,86,31,140,31,38,31,38,30,38,29,52,31,225,31,25,31,173,31,173,30,121,31,82,31,25,31,86,31,42,31,129,31,72,31,241,31,192,31,139,31,46,31,89,31,68,31,68,30,144,31,23,31,137,31,137,30,138,31,163,31,163,30,133,31,88,31,88,30,88,29,138,31,22,31,22,30,101,31,40,31,84,31,101,31,101,30,101,29,101,28,196,31,126,31,126,30,144,31,65,31,39,31,48,31,116,31,126,31,106,31,105,31,105,30,140,31,140,30,35,31,35,30,25,31,223,31,88,31,130,31,16,31,99,31,36,31,15,31,233,31,137,31,209,31,209,30,234,31,129,31,129,30,105,31,146,31,104,31,104,30,139,31,217,31,54,31,60,31,239,31,116,31,68,31,11,31,11,30,11,29,52,31,252,31,189,31,53,31,94,31,149,31,149,30,149,29,130,31,160,31,23,31,23,30,23,29,215,31,66,31,66,30,215,31,97,31,135,31,135,30,234,31,147,31,236,31,1,31,69,31,105,31,101,31,90,31,90,30,231,31,130,31,81,31,124,31,250,31,117,31,117,30,151,31,151,30,151,29,119,31,135,31,9,31,219,31,25,31,87,31,36,31,137,31,185,31,224,31,193,31,189,31,181,31,193,31,193,30,55,31,55,30,94,31,239,31,181,31,174,31,128,31,176,31,224,31,224,30,161,31,113,31,160,31,96,31,22,31,22,30,57,31,86,31,143,31,104,31,43,31,43,30,253,31,14,31,154,31,154,30,48,31,151,31,121,31,202,31,96,31,121,31,166,31,176,31,129,31,129,30,129,29,124,31,98,31,131,31,131,30,22,31,242,31,242,30,61,31,163,31,57,31,57,30,170,31,127,31,190,31,190,30,65,31,61,31,108,31,108,30,90,31,221,31,206,31,191,31,15,31,123,31,7,31,50,31,54,31,253,31,140,31,140,30,140,29,119,31,116,31,133,31,133,31,171,31,171,30,14,31,59,31,27,31,80,31,57,31,175,31,175,30,101,31,101,30,101,29,148,31,19,31,19,30,165,31,64,31,86,31,120,31,91,31,179,31,188,31,242,31,242,30,218,31,212,31,144,31,28,31,148,31,148,30,250,31,83,31,222,31,205,31,108,31,152,31,231,31,92,31,108,31,132,31,132,30,148,31,148,30,148,29,4,31,202,31,133,31,133,30,166,31,166,30,229,31,80,31,86,31,186,31,162,31,33,31,99,31,3,31,3,30,247,31,66,31,181,31,171,31,194,31,3,31,3,30,92,31,193,31,109,31,153,31,153,30,208,31,122,31,67,31,101,31,101,30,78,31,78,30,78,29,124,31,168,31,168,30,76,31,152,31,242,31,20,31,3,31,90,31,110,31,217,31,104,31,104,30,38,31,38,30,82,31,108,31,108,30,198,31,245,31,165,31,165,30,254,31,137,31,146,31,255,31,146,31,132,31,49,31,50,31,162,31,163,31,163,30,43,31,222,31,46,31,194,31,194,30,197,31,53,31,32,31,32,30,32,29,97,31,212,31,184,31,104,31,86,31,86,30,194,31,163,31,44,31,44,30,44,29,44,28,180,31,74,31,150,31,241,31,241,30,117,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
