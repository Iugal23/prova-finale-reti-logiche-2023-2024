-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_372 is
end project_tb_372;

architecture project_tb_arch_372 of project_tb_372 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 324;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,146,0,112,0,143,0,40,0,79,0,28,0,190,0,63,0,0,0,0,0,162,0,0,0,37,0,32,0,28,0,0,0,207,0,76,0,0,0,252,0,203,0,0,0,177,0,0,0,0,0,184,0,0,0,237,0,0,0,14,0,249,0,143,0,205,0,159,0,0,0,0,0,89,0,156,0,14,0,130,0,0,0,5,0,38,0,175,0,241,0,0,0,0,0,181,0,134,0,165,0,204,0,85,0,0,0,232,0,0,0,89,0,101,0,225,0,95,0,201,0,0,0,185,0,50,0,0,0,0,0,111,0,93,0,3,0,73,0,0,0,13,0,33,0,56,0,0,0,208,0,245,0,87,0,0,0,64,0,68,0,180,0,135,0,237,0,110,0,116,0,241,0,40,0,143,0,190,0,46,0,0,0,0,0,0,0,132,0,1,0,229,0,214,0,92,0,162,0,133,0,204,0,173,0,0,0,92,0,20,0,0,0,127,0,58,0,236,0,28,0,240,0,231,0,0,0,100,0,204,0,155,0,60,0,138,0,75,0,43,0,125,0,16,0,88,0,0,0,227,0,215,0,80,0,115,0,99,0,13,0,141,0,0,0,142,0,125,0,248,0,174,0,8,0,25,0,60,0,240,0,178,0,211,0,89,0,95,0,161,0,253,0,0,0,31,0,0,0,0,0,0,0,54,0,139,0,0,0,173,0,154,0,118,0,250,0,0,0,11,0,0,0,130,0,17,0,83,0,161,0,0,0,252,0,0,0,72,0,2,0,241,0,162,0,177,0,163,0,61,0,98,0,111,0,0,0,2,0,0,0,155,0,0,0,197,0,243,0,161,0,138,0,234,0,203,0,225,0,114,0,102,0,216,0,16,0,207,0,191,0,186,0,255,0,57,0,5,0,43,0,227,0,68,0,122,0,118,0,86,0,236,0,80,0,101,0,0,0,0,0,239,0,0,0,26,0,105,0,230,0,63,0,172,0,0,0,92,0,82,0,159,0,10,0,11,0,198,0,153,0,0,0,222,0,0,0,192,0,125,0,102,0,104,0,243,0,0,0,136,0,255,0,206,0,126,0,154,0,103,0,0,0,204,0,0,0,182,0,4,0,64,0,114,0,226,0,77,0,0,0,110,0,161,0,11,0,172,0,0,0,0,0,236,0,205,0,116,0,198,0,222,0,60,0,78,0,44,0,0,0,25,0,115,0,0,0,60,0,78,0,243,0,105,0,0,0,76,0,11,0,0,0,134,0,149,0,197,0,255,0,136,0,240,0,159,0,107,0,121,0,0,0,32,0,251,0,0,0,75,0,112,0,92,0,95,0,167,0,123,0,37,0,67,0,123,0,122,0,209,0,67,0,78,0,48,0,122,0,120,0,120,0,103,0,0,0,0,0,247,0,239,0,15,0,0,0,38,0,244,0,0,0,205,0,0,0,48,0,48,0,51,0,146,0,221,0);
signal scenario_full  : scenario_type := (109,31,146,31,112,31,143,31,40,31,79,31,28,31,190,31,63,31,63,30,63,29,162,31,162,30,37,31,32,31,28,31,28,30,207,31,76,31,76,30,252,31,203,31,203,30,177,31,177,30,177,29,184,31,184,30,237,31,237,30,14,31,249,31,143,31,205,31,159,31,159,30,159,29,89,31,156,31,14,31,130,31,130,30,5,31,38,31,175,31,241,31,241,30,241,29,181,31,134,31,165,31,204,31,85,31,85,30,232,31,232,30,89,31,101,31,225,31,95,31,201,31,201,30,185,31,50,31,50,30,50,29,111,31,93,31,3,31,73,31,73,30,13,31,33,31,56,31,56,30,208,31,245,31,87,31,87,30,64,31,68,31,180,31,135,31,237,31,110,31,116,31,241,31,40,31,143,31,190,31,46,31,46,30,46,29,46,28,132,31,1,31,229,31,214,31,92,31,162,31,133,31,204,31,173,31,173,30,92,31,20,31,20,30,127,31,58,31,236,31,28,31,240,31,231,31,231,30,100,31,204,31,155,31,60,31,138,31,75,31,43,31,125,31,16,31,88,31,88,30,227,31,215,31,80,31,115,31,99,31,13,31,141,31,141,30,142,31,125,31,248,31,174,31,8,31,25,31,60,31,240,31,178,31,211,31,89,31,95,31,161,31,253,31,253,30,31,31,31,30,31,29,31,28,54,31,139,31,139,30,173,31,154,31,118,31,250,31,250,30,11,31,11,30,130,31,17,31,83,31,161,31,161,30,252,31,252,30,72,31,2,31,241,31,162,31,177,31,163,31,61,31,98,31,111,31,111,30,2,31,2,30,155,31,155,30,197,31,243,31,161,31,138,31,234,31,203,31,225,31,114,31,102,31,216,31,16,31,207,31,191,31,186,31,255,31,57,31,5,31,43,31,227,31,68,31,122,31,118,31,86,31,236,31,80,31,101,31,101,30,101,29,239,31,239,30,26,31,105,31,230,31,63,31,172,31,172,30,92,31,82,31,159,31,10,31,11,31,198,31,153,31,153,30,222,31,222,30,192,31,125,31,102,31,104,31,243,31,243,30,136,31,255,31,206,31,126,31,154,31,103,31,103,30,204,31,204,30,182,31,4,31,64,31,114,31,226,31,77,31,77,30,110,31,161,31,11,31,172,31,172,30,172,29,236,31,205,31,116,31,198,31,222,31,60,31,78,31,44,31,44,30,25,31,115,31,115,30,60,31,78,31,243,31,105,31,105,30,76,31,11,31,11,30,134,31,149,31,197,31,255,31,136,31,240,31,159,31,107,31,121,31,121,30,32,31,251,31,251,30,75,31,112,31,92,31,95,31,167,31,123,31,37,31,67,31,123,31,122,31,209,31,67,31,78,31,48,31,122,31,120,31,120,31,103,31,103,30,103,29,247,31,239,31,15,31,15,30,38,31,244,31,244,30,205,31,205,30,48,31,48,31,51,31,146,31,221,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
