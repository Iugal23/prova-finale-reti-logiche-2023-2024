-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_503 is
end project_tb_503;

architecture project_tb_arch_503 of project_tb_503 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 813;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,79,0,8,0,169,0,40,0,53,0,191,0,0,0,174,0,139,0,121,0,0,0,141,0,128,0,108,0,151,0,0,0,151,0,0,0,37,0,193,0,12,0,185,0,0,0,248,0,11,0,12,0,242,0,220,0,69,0,226,0,22,0,24,0,86,0,174,0,75,0,0,0,0,0,55,0,0,0,30,0,194,0,244,0,85,0,183,0,89,0,125,0,0,0,3,0,47,0,179,0,0,0,11,0,7,0,0,0,70,0,122,0,0,0,0,0,1,0,0,0,99,0,211,0,0,0,223,0,65,0,217,0,187,0,219,0,0,0,0,0,3,0,224,0,53,0,32,0,0,0,192,0,38,0,0,0,117,0,217,0,146,0,99,0,202,0,88,0,249,0,143,0,105,0,150,0,165,0,15,0,200,0,86,0,244,0,83,0,84,0,236,0,179,0,99,0,63,0,24,0,37,0,0,0,255,0,153,0,174,0,99,0,0,0,184,0,78,0,148,0,0,0,72,0,170,0,138,0,158,0,245,0,187,0,166,0,152,0,0,0,252,0,215,0,10,0,2,0,33,0,39,0,0,0,14,0,72,0,0,0,196,0,0,0,245,0,224,0,26,0,7,0,165,0,170,0,104,0,130,0,83,0,150,0,214,0,75,0,154,0,123,0,190,0,144,0,161,0,88,0,32,0,158,0,162,0,49,0,156,0,94,0,234,0,0,0,5,0,32,0,170,0,66,0,103,0,188,0,24,0,235,0,132,0,0,0,0,0,235,0,0,0,0,0,140,0,0,0,0,0,4,0,136,0,152,0,3,0,32,0,246,0,186,0,95,0,183,0,7,0,255,0,0,0,10,0,158,0,39,0,190,0,194,0,74,0,11,0,69,0,205,0,156,0,0,0,47,0,67,0,127,0,0,0,0,0,208,0,189,0,177,0,103,0,154,0,98,0,0,0,27,0,25,0,0,0,199,0,0,0,0,0,0,0,221,0,99,0,252,0,18,0,119,0,0,0,17,0,107,0,74,0,12,0,170,0,143,0,147,0,120,0,0,0,57,0,146,0,239,0,239,0,51,0,167,0,29,0,97,0,97,0,149,0,123,0,0,0,0,0,192,0,157,0,236,0,240,0,152,0,157,0,182,0,169,0,28,0,0,0,130,0,0,0,0,0,211,0,252,0,60,0,179,0,229,0,19,0,59,0,171,0,125,0,212,0,217,0,83,0,0,0,229,0,160,0,189,0,198,0,253,0,0,0,28,0,70,0,228,0,229,0,68,0,129,0,0,0,115,0,0,0,204,0,122,0,109,0,236,0,159,0,209,0,41,0,36,0,251,0,0,0,45,0,77,0,3,0,251,0,115,0,215,0,0,0,57,0,67,0,173,0,0,0,38,0,0,0,132,0,154,0,0,0,115,0,0,0,139,0,0,0,42,0,250,0,75,0,114,0,228,0,201,0,184,0,123,0,0,0,0,0,0,0,0,0,0,0,79,0,77,0,0,0,252,0,135,0,0,0,0,0,184,0,24,0,114,0,18,0,0,0,227,0,86,0,0,0,194,0,250,0,99,0,103,0,175,0,20,0,0,0,21,0,226,0,0,0,250,0,216,0,62,0,0,0,0,0,165,0,150,0,166,0,2,0,152,0,130,0,64,0,202,0,221,0,0,0,5,0,0,0,102,0,0,0,166,0,67,0,0,0,204,0,215,0,215,0,0,0,87,0,89,0,216,0,244,0,117,0,96,0,60,0,248,0,194,0,127,0,0,0,0,0,73,0,117,0,178,0,100,0,0,0,44,0,67,0,142,0,97,0,0,0,0,0,51,0,0,0,190,0,227,0,0,0,34,0,0,0,36,0,211,0,0,0,151,0,0,0,198,0,57,0,185,0,219,0,0,0,0,0,0,0,132,0,199,0,0,0,146,0,0,0,75,0,0,0,201,0,212,0,74,0,181,0,255,0,91,0,213,0,0,0,106,0,65,0,160,0,104,0,45,0,254,0,0,0,141,0,187,0,93,0,0,0,7,0,165,0,86,0,240,0,83,0,0,0,237,0,5,0,102,0,137,0,146,0,206,0,63,0,181,0,227,0,147,0,120,0,158,0,66,0,91,0,249,0,229,0,208,0,22,0,192,0,195,0,0,0,33,0,255,0,206,0,42,0,149,0,0,0,160,0,82,0,163,0,226,0,103,0,0,0,215,0,105,0,19,0,179,0,244,0,94,0,88,0,0,0,0,0,0,0,107,0,0,0,101,0,88,0,129,0,176,0,32,0,214,0,0,0,166,0,58,0,0,0,152,0,207,0,36,0,254,0,0,0,131,0,100,0,254,0,170,0,28,0,252,0,29,0,0,0,161,0,231,0,240,0,0,0,20,0,157,0,236,0,180,0,0,0,205,0,82,0,0,0,202,0,126,0,226,0,18,0,72,0,51,0,224,0,52,0,7,0,254,0,53,0,0,0,37,0,0,0,0,0,0,0,48,0,0,0,22,0,227,0,128,0,57,0,211,0,63,0,244,0,243,0,218,0,36,0,203,0,62,0,17,0,193,0,0,0,246,0,139,0,135,0,0,0,238,0,122,0,186,0,127,0,85,0,118,0,203,0,251,0,195,0,137,0,0,0,232,0,131,0,206,0,38,0,248,0,131,0,246,0,115,0,145,0,0,0,209,0,248,0,22,0,100,0,78,0,99,0,58,0,0,0,213,0,0,0,10,0,35,0,0,0,55,0,0,0,0,0,49,0,75,0,106,0,64,0,213,0,147,0,86,0,16,0,103,0,154,0,73,0,175,0,88,0,86,0,0,0,11,0,114,0,13,0,168,0,27,0,0,0,57,0,0,0,117,0,106,0,45,0,158,0,72,0,47,0,0,0,160,0,148,0,226,0,0,0,12,0,117,0,101,0,106,0,0,0,0,0,75,0,141,0,0,0,193,0,149,0,140,0,56,0,166,0,38,0,80,0,220,0,200,0,44,0,4,0,211,0,251,0,0,0,140,0,206,0,80,0,0,0,174,0,158,0,0,0,162,0,212,0,151,0,157,0,192,0,253,0,212,0,231,0,245,0,123,0,148,0,50,0,157,0,254,0,0,0,116,0,0,0,0,0,67,0,0,0,190,0,147,0,0,0,223,0,0,0,130,0,21,0,24,0,87,0,0,0,183,0,6,0,0,0,208,0,56,0,193,0,5,0,159,0,74,0,132,0,0,0,145,0,0,0,247,0,113,0,0,0,137,0,155,0,251,0,241,0,61,0,183,0,161,0,144,0,237,0,169,0,225,0,0,0,93,0,0,0,0,0,0,0,26,0,0,0,25,0,137,0,184,0,114,0,111,0,92,0,0,0,160,0,0,0,244,0,152,0,186,0,205,0,177,0,129,0,161,0,27,0,0,0,1,0,0,0,42,0,154,0,34,0,192,0,0,0,191,0,191,0,73,0,88,0,130,0,0,0,0,0,0,0,131,0,0,0,162,0,0,0,58,0,23,0,245,0,0,0,120,0,0,0,243,0,234,0,0,0,0,0,28,0,86,0,233,0,0,0,198,0,111,0,228,0,21,0,140,0,31,0,236,0,13,0,147,0,0,0,49,0,94,0,138,0,235,0,187,0,0,0,91,0,101,0,166,0,224,0,110,0,124,0,0,0,91,0,190,0);
signal scenario_full  : scenario_type := (1,31,79,31,8,31,169,31,40,31,53,31,191,31,191,30,174,31,139,31,121,31,121,30,141,31,128,31,108,31,151,31,151,30,151,31,151,30,37,31,193,31,12,31,185,31,185,30,248,31,11,31,12,31,242,31,220,31,69,31,226,31,22,31,24,31,86,31,174,31,75,31,75,30,75,29,55,31,55,30,30,31,194,31,244,31,85,31,183,31,89,31,125,31,125,30,3,31,47,31,179,31,179,30,11,31,7,31,7,30,70,31,122,31,122,30,122,29,1,31,1,30,99,31,211,31,211,30,223,31,65,31,217,31,187,31,219,31,219,30,219,29,3,31,224,31,53,31,32,31,32,30,192,31,38,31,38,30,117,31,217,31,146,31,99,31,202,31,88,31,249,31,143,31,105,31,150,31,165,31,15,31,200,31,86,31,244,31,83,31,84,31,236,31,179,31,99,31,63,31,24,31,37,31,37,30,255,31,153,31,174,31,99,31,99,30,184,31,78,31,148,31,148,30,72,31,170,31,138,31,158,31,245,31,187,31,166,31,152,31,152,30,252,31,215,31,10,31,2,31,33,31,39,31,39,30,14,31,72,31,72,30,196,31,196,30,245,31,224,31,26,31,7,31,165,31,170,31,104,31,130,31,83,31,150,31,214,31,75,31,154,31,123,31,190,31,144,31,161,31,88,31,32,31,158,31,162,31,49,31,156,31,94,31,234,31,234,30,5,31,32,31,170,31,66,31,103,31,188,31,24,31,235,31,132,31,132,30,132,29,235,31,235,30,235,29,140,31,140,30,140,29,4,31,136,31,152,31,3,31,32,31,246,31,186,31,95,31,183,31,7,31,255,31,255,30,10,31,158,31,39,31,190,31,194,31,74,31,11,31,69,31,205,31,156,31,156,30,47,31,67,31,127,31,127,30,127,29,208,31,189,31,177,31,103,31,154,31,98,31,98,30,27,31,25,31,25,30,199,31,199,30,199,29,199,28,221,31,99,31,252,31,18,31,119,31,119,30,17,31,107,31,74,31,12,31,170,31,143,31,147,31,120,31,120,30,57,31,146,31,239,31,239,31,51,31,167,31,29,31,97,31,97,31,149,31,123,31,123,30,123,29,192,31,157,31,236,31,240,31,152,31,157,31,182,31,169,31,28,31,28,30,130,31,130,30,130,29,211,31,252,31,60,31,179,31,229,31,19,31,59,31,171,31,125,31,212,31,217,31,83,31,83,30,229,31,160,31,189,31,198,31,253,31,253,30,28,31,70,31,228,31,229,31,68,31,129,31,129,30,115,31,115,30,204,31,122,31,109,31,236,31,159,31,209,31,41,31,36,31,251,31,251,30,45,31,77,31,3,31,251,31,115,31,215,31,215,30,57,31,67,31,173,31,173,30,38,31,38,30,132,31,154,31,154,30,115,31,115,30,139,31,139,30,42,31,250,31,75,31,114,31,228,31,201,31,184,31,123,31,123,30,123,29,123,28,123,27,123,26,79,31,77,31,77,30,252,31,135,31,135,30,135,29,184,31,24,31,114,31,18,31,18,30,227,31,86,31,86,30,194,31,250,31,99,31,103,31,175,31,20,31,20,30,21,31,226,31,226,30,250,31,216,31,62,31,62,30,62,29,165,31,150,31,166,31,2,31,152,31,130,31,64,31,202,31,221,31,221,30,5,31,5,30,102,31,102,30,166,31,67,31,67,30,204,31,215,31,215,31,215,30,87,31,89,31,216,31,244,31,117,31,96,31,60,31,248,31,194,31,127,31,127,30,127,29,73,31,117,31,178,31,100,31,100,30,44,31,67,31,142,31,97,31,97,30,97,29,51,31,51,30,190,31,227,31,227,30,34,31,34,30,36,31,211,31,211,30,151,31,151,30,198,31,57,31,185,31,219,31,219,30,219,29,219,28,132,31,199,31,199,30,146,31,146,30,75,31,75,30,201,31,212,31,74,31,181,31,255,31,91,31,213,31,213,30,106,31,65,31,160,31,104,31,45,31,254,31,254,30,141,31,187,31,93,31,93,30,7,31,165,31,86,31,240,31,83,31,83,30,237,31,5,31,102,31,137,31,146,31,206,31,63,31,181,31,227,31,147,31,120,31,158,31,66,31,91,31,249,31,229,31,208,31,22,31,192,31,195,31,195,30,33,31,255,31,206,31,42,31,149,31,149,30,160,31,82,31,163,31,226,31,103,31,103,30,215,31,105,31,19,31,179,31,244,31,94,31,88,31,88,30,88,29,88,28,107,31,107,30,101,31,88,31,129,31,176,31,32,31,214,31,214,30,166,31,58,31,58,30,152,31,207,31,36,31,254,31,254,30,131,31,100,31,254,31,170,31,28,31,252,31,29,31,29,30,161,31,231,31,240,31,240,30,20,31,157,31,236,31,180,31,180,30,205,31,82,31,82,30,202,31,126,31,226,31,18,31,72,31,51,31,224,31,52,31,7,31,254,31,53,31,53,30,37,31,37,30,37,29,37,28,48,31,48,30,22,31,227,31,128,31,57,31,211,31,63,31,244,31,243,31,218,31,36,31,203,31,62,31,17,31,193,31,193,30,246,31,139,31,135,31,135,30,238,31,122,31,186,31,127,31,85,31,118,31,203,31,251,31,195,31,137,31,137,30,232,31,131,31,206,31,38,31,248,31,131,31,246,31,115,31,145,31,145,30,209,31,248,31,22,31,100,31,78,31,99,31,58,31,58,30,213,31,213,30,10,31,35,31,35,30,55,31,55,30,55,29,49,31,75,31,106,31,64,31,213,31,147,31,86,31,16,31,103,31,154,31,73,31,175,31,88,31,86,31,86,30,11,31,114,31,13,31,168,31,27,31,27,30,57,31,57,30,117,31,106,31,45,31,158,31,72,31,47,31,47,30,160,31,148,31,226,31,226,30,12,31,117,31,101,31,106,31,106,30,106,29,75,31,141,31,141,30,193,31,149,31,140,31,56,31,166,31,38,31,80,31,220,31,200,31,44,31,4,31,211,31,251,31,251,30,140,31,206,31,80,31,80,30,174,31,158,31,158,30,162,31,212,31,151,31,157,31,192,31,253,31,212,31,231,31,245,31,123,31,148,31,50,31,157,31,254,31,254,30,116,31,116,30,116,29,67,31,67,30,190,31,147,31,147,30,223,31,223,30,130,31,21,31,24,31,87,31,87,30,183,31,6,31,6,30,208,31,56,31,193,31,5,31,159,31,74,31,132,31,132,30,145,31,145,30,247,31,113,31,113,30,137,31,155,31,251,31,241,31,61,31,183,31,161,31,144,31,237,31,169,31,225,31,225,30,93,31,93,30,93,29,93,28,26,31,26,30,25,31,137,31,184,31,114,31,111,31,92,31,92,30,160,31,160,30,244,31,152,31,186,31,205,31,177,31,129,31,161,31,27,31,27,30,1,31,1,30,42,31,154,31,34,31,192,31,192,30,191,31,191,31,73,31,88,31,130,31,130,30,130,29,130,28,131,31,131,30,162,31,162,30,58,31,23,31,245,31,245,30,120,31,120,30,243,31,234,31,234,30,234,29,28,31,86,31,233,31,233,30,198,31,111,31,228,31,21,31,140,31,31,31,236,31,13,31,147,31,147,30,49,31,94,31,138,31,235,31,187,31,187,30,91,31,101,31,166,31,224,31,110,31,124,31,124,30,91,31,190,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
