-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_830 is
end project_tb_830;

architecture project_tb_arch_830 of project_tb_830 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 778;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (242,0,0,0,0,0,167,0,0,0,246,0,17,0,238,0,50,0,232,0,60,0,205,0,63,0,134,0,91,0,18,0,150,0,222,0,0,0,141,0,1,0,156,0,37,0,0,0,31,0,136,0,54,0,0,0,140,0,17,0,0,0,0,0,224,0,66,0,157,0,250,0,206,0,120,0,29,0,188,0,20,0,169,0,0,0,102,0,141,0,45,0,12,0,0,0,249,0,92,0,0,0,255,0,70,0,233,0,234,0,47,0,199,0,152,0,193,0,121,0,83,0,173,0,0,0,68,0,0,0,0,0,22,0,144,0,90,0,149,0,218,0,232,0,0,0,184,0,0,0,226,0,0,0,181,0,255,0,82,0,72,0,57,0,13,0,214,0,64,0,166,0,80,0,195,0,98,0,16,0,217,0,74,0,163,0,108,0,0,0,231,0,63,0,0,0,13,0,142,0,0,0,0,0,0,0,86,0,153,0,0,0,174,0,57,0,0,0,0,0,146,0,184,0,152,0,245,0,5,0,16,0,181,0,0,0,75,0,242,0,0,0,252,0,29,0,18,0,185,0,23,0,190,0,172,0,87,0,207,0,164,0,210,0,248,0,46,0,132,0,129,0,0,0,100,0,20,0,204,0,0,0,4,0,0,0,226,0,0,0,27,0,24,0,195,0,0,0,0,0,253,0,236,0,148,0,0,0,51,0,18,0,60,0,181,0,152,0,238,0,218,0,0,0,204,0,0,0,48,0,19,0,158,0,0,0,20,0,138,0,105,0,233,0,161,0,7,0,153,0,222,0,29,0,45,0,234,0,0,0,91,0,0,0,203,0,183,0,172,0,34,0,0,0,0,0,0,0,34,0,157,0,54,0,0,0,155,0,164,0,46,0,233,0,0,0,0,0,66,0,19,0,0,0,0,0,0,0,0,0,0,0,0,0,62,0,0,0,131,0,0,0,0,0,130,0,78,0,6,0,168,0,124,0,194,0,179,0,255,0,224,0,0,0,0,0,255,0,136,0,158,0,80,0,82,0,243,0,47,0,0,0,21,0,42,0,0,0,82,0,147,0,180,0,0,0,32,0,138,0,26,0,223,0,59,0,0,0,203,0,47,0,148,0,35,0,240,0,74,0,181,0,233,0,229,0,84,0,229,0,140,0,159,0,60,0,88,0,137,0,158,0,150,0,204,0,252,0,189,0,187,0,0,0,23,0,0,0,189,0,215,0,0,0,22,0,195,0,30,0,60,0,0,0,0,0,189,0,152,0,25,0,14,0,0,0,99,0,59,0,16,0,158,0,105,0,221,0,97,0,83,0,43,0,122,0,0,0,66,0,66,0,33,0,52,0,192,0,0,0,88,0,69,0,155,0,163,0,126,0,134,0,253,0,182,0,243,0,0,0,0,0,71,0,192,0,110,0,147,0,103,0,194,0,0,0,0,0,48,0,168,0,0,0,225,0,188,0,157,0,0,0,0,0,135,0,100,0,225,0,5,0,179,0,32,0,202,0,89,0,125,0,0,0,0,0,0,0,171,0,125,0,114,0,178,0,161,0,43,0,53,0,123,0,83,0,54,0,0,0,191,0,26,0,57,0,153,0,228,0,77,0,16,0,69,0,0,0,93,0,7,0,156,0,76,0,211,0,0,0,161,0,184,0,47,0,0,0,97,0,59,0,243,0,0,0,0,0,189,0,146,0,231,0,173,0,58,0,78,0,0,0,0,0,0,0,79,0,156,0,119,0,1,0,144,0,218,0,66,0,113,0,19,0,68,0,56,0,135,0,170,0,8,0,162,0,248,0,0,0,0,0,183,0,34,0,0,0,146,0,233,0,0,0,205,0,91,0,0,0,42,0,0,0,129,0,0,0,153,0,180,0,49,0,12,0,39,0,226,0,102,0,72,0,40,0,0,0,182,0,214,0,145,0,0,0,86,0,34,0,164,0,16,0,0,0,204,0,104,0,251,0,196,0,60,0,102,0,208,0,231,0,163,0,215,0,143,0,19,0,122,0,0,0,187,0,117,0,95,0,114,0,0,0,42,0,74,0,140,0,157,0,157,0,126,0,128,0,92,0,0,0,242,0,47,0,0,0,90,0,67,0,70,0,237,0,0,0,0,0,54,0,225,0,198,0,186,0,23,0,0,0,71,0,0,0,225,0,243,0,172,0,28,0,74,0,101,0,111,0,168,0,12,0,223,0,21,0,178,0,139,0,143,0,58,0,69,0,97,0,56,0,113,0,0,0,243,0,98,0,0,0,213,0,0,0,75,0,108,0,0,0,36,0,31,0,34,0,58,0,0,0,213,0,205,0,53,0,213,0,252,0,238,0,239,0,212,0,231,0,240,0,123,0,151,0,121,0,114,0,1,0,162,0,0,0,0,0,91,0,247,0,0,0,0,0,1,0,0,0,43,0,129,0,148,0,0,0,0,0,0,0,6,0,0,0,252,0,100,0,152,0,218,0,163,0,216,0,76,0,0,0,214,0,62,0,173,0,149,0,34,0,166,0,195,0,21,0,214,0,26,0,27,0,85,0,192,0,109,0,175,0,0,0,0,0,110,0,0,0,185,0,0,0,0,0,218,0,171,0,0,0,225,0,247,0,0,0,0,0,0,0,224,0,46,0,0,0,154,0,0,0,159,0,0,0,165,0,153,0,0,0,231,0,222,0,166,0,197,0,126,0,20,0,155,0,0,0,27,0,0,0,128,0,0,0,201,0,170,0,11,0,18,0,221,0,101,0,117,0,14,0,235,0,50,0,194,0,116,0,41,0,103,0,78,0,0,0,151,0,0,0,164,0,0,0,123,0,233,0,230,0,113,0,120,0,153,0,0,0,254,0,136,0,101,0,31,0,249,0,0,0,0,0,239,0,0,0,210,0,211,0,76,0,54,0,0,0,110,0,31,0,3,0,154,0,0,0,0,0,154,0,31,0,15,0,83,0,0,0,109,0,140,0,0,0,60,0,87,0,4,0,12,0,129,0,0,0,0,0,0,0,127,0,60,0,67,0,154,0,0,0,140,0,164,0,85,0,94,0,96,0,28,0,0,0,10,0,0,0,198,0,0,0,0,0,54,0,131,0,98,0,85,0,213,0,77,0,0,0,249,0,202,0,168,0,25,0,187,0,93,0,0,0,34,0,167,0,143,0,86,0,0,0,102,0,150,0,0,0,107,0,191,0,30,0,255,0,0,0,78,0,144,0,220,0,44,0,0,0,241,0,37,0,164,0,34,0,0,0,0,0,0,0,231,0,0,0,0,0,31,0,238,0,144,0,88,0,184,0,123,0,200,0,101,0,207,0,155,0,182,0,140,0,0,0,128,0,213,0,0,0,55,0,136,0,0,0,38,0,0,0,35,0,0,0,248,0,82,0,0,0,118,0,161,0,134,0,20,0,146,0,81,0,0,0,16,0,95,0,0,0,196,0,196,0,157,0,29,0,153,0,212,0,228,0,157,0,63,0,98,0,84,0,38,0,13,0,33,0,201,0,0,0,108,0);
signal scenario_full  : scenario_type := (242,31,242,30,242,29,167,31,167,30,246,31,17,31,238,31,50,31,232,31,60,31,205,31,63,31,134,31,91,31,18,31,150,31,222,31,222,30,141,31,1,31,156,31,37,31,37,30,31,31,136,31,54,31,54,30,140,31,17,31,17,30,17,29,224,31,66,31,157,31,250,31,206,31,120,31,29,31,188,31,20,31,169,31,169,30,102,31,141,31,45,31,12,31,12,30,249,31,92,31,92,30,255,31,70,31,233,31,234,31,47,31,199,31,152,31,193,31,121,31,83,31,173,31,173,30,68,31,68,30,68,29,22,31,144,31,90,31,149,31,218,31,232,31,232,30,184,31,184,30,226,31,226,30,181,31,255,31,82,31,72,31,57,31,13,31,214,31,64,31,166,31,80,31,195,31,98,31,16,31,217,31,74,31,163,31,108,31,108,30,231,31,63,31,63,30,13,31,142,31,142,30,142,29,142,28,86,31,153,31,153,30,174,31,57,31,57,30,57,29,146,31,184,31,152,31,245,31,5,31,16,31,181,31,181,30,75,31,242,31,242,30,252,31,29,31,18,31,185,31,23,31,190,31,172,31,87,31,207,31,164,31,210,31,248,31,46,31,132,31,129,31,129,30,100,31,20,31,204,31,204,30,4,31,4,30,226,31,226,30,27,31,24,31,195,31,195,30,195,29,253,31,236,31,148,31,148,30,51,31,18,31,60,31,181,31,152,31,238,31,218,31,218,30,204,31,204,30,48,31,19,31,158,31,158,30,20,31,138,31,105,31,233,31,161,31,7,31,153,31,222,31,29,31,45,31,234,31,234,30,91,31,91,30,203,31,183,31,172,31,34,31,34,30,34,29,34,28,34,31,157,31,54,31,54,30,155,31,164,31,46,31,233,31,233,30,233,29,66,31,19,31,19,30,19,29,19,28,19,27,19,26,19,25,62,31,62,30,131,31,131,30,131,29,130,31,78,31,6,31,168,31,124,31,194,31,179,31,255,31,224,31,224,30,224,29,255,31,136,31,158,31,80,31,82,31,243,31,47,31,47,30,21,31,42,31,42,30,82,31,147,31,180,31,180,30,32,31,138,31,26,31,223,31,59,31,59,30,203,31,47,31,148,31,35,31,240,31,74,31,181,31,233,31,229,31,84,31,229,31,140,31,159,31,60,31,88,31,137,31,158,31,150,31,204,31,252,31,189,31,187,31,187,30,23,31,23,30,189,31,215,31,215,30,22,31,195,31,30,31,60,31,60,30,60,29,189,31,152,31,25,31,14,31,14,30,99,31,59,31,16,31,158,31,105,31,221,31,97,31,83,31,43,31,122,31,122,30,66,31,66,31,33,31,52,31,192,31,192,30,88,31,69,31,155,31,163,31,126,31,134,31,253,31,182,31,243,31,243,30,243,29,71,31,192,31,110,31,147,31,103,31,194,31,194,30,194,29,48,31,168,31,168,30,225,31,188,31,157,31,157,30,157,29,135,31,100,31,225,31,5,31,179,31,32,31,202,31,89,31,125,31,125,30,125,29,125,28,171,31,125,31,114,31,178,31,161,31,43,31,53,31,123,31,83,31,54,31,54,30,191,31,26,31,57,31,153,31,228,31,77,31,16,31,69,31,69,30,93,31,7,31,156,31,76,31,211,31,211,30,161,31,184,31,47,31,47,30,97,31,59,31,243,31,243,30,243,29,189,31,146,31,231,31,173,31,58,31,78,31,78,30,78,29,78,28,79,31,156,31,119,31,1,31,144,31,218,31,66,31,113,31,19,31,68,31,56,31,135,31,170,31,8,31,162,31,248,31,248,30,248,29,183,31,34,31,34,30,146,31,233,31,233,30,205,31,91,31,91,30,42,31,42,30,129,31,129,30,153,31,180,31,49,31,12,31,39,31,226,31,102,31,72,31,40,31,40,30,182,31,214,31,145,31,145,30,86,31,34,31,164,31,16,31,16,30,204,31,104,31,251,31,196,31,60,31,102,31,208,31,231,31,163,31,215,31,143,31,19,31,122,31,122,30,187,31,117,31,95,31,114,31,114,30,42,31,74,31,140,31,157,31,157,31,126,31,128,31,92,31,92,30,242,31,47,31,47,30,90,31,67,31,70,31,237,31,237,30,237,29,54,31,225,31,198,31,186,31,23,31,23,30,71,31,71,30,225,31,243,31,172,31,28,31,74,31,101,31,111,31,168,31,12,31,223,31,21,31,178,31,139,31,143,31,58,31,69,31,97,31,56,31,113,31,113,30,243,31,98,31,98,30,213,31,213,30,75,31,108,31,108,30,36,31,31,31,34,31,58,31,58,30,213,31,205,31,53,31,213,31,252,31,238,31,239,31,212,31,231,31,240,31,123,31,151,31,121,31,114,31,1,31,162,31,162,30,162,29,91,31,247,31,247,30,247,29,1,31,1,30,43,31,129,31,148,31,148,30,148,29,148,28,6,31,6,30,252,31,100,31,152,31,218,31,163,31,216,31,76,31,76,30,214,31,62,31,173,31,149,31,34,31,166,31,195,31,21,31,214,31,26,31,27,31,85,31,192,31,109,31,175,31,175,30,175,29,110,31,110,30,185,31,185,30,185,29,218,31,171,31,171,30,225,31,247,31,247,30,247,29,247,28,224,31,46,31,46,30,154,31,154,30,159,31,159,30,165,31,153,31,153,30,231,31,222,31,166,31,197,31,126,31,20,31,155,31,155,30,27,31,27,30,128,31,128,30,201,31,170,31,11,31,18,31,221,31,101,31,117,31,14,31,235,31,50,31,194,31,116,31,41,31,103,31,78,31,78,30,151,31,151,30,164,31,164,30,123,31,233,31,230,31,113,31,120,31,153,31,153,30,254,31,136,31,101,31,31,31,249,31,249,30,249,29,239,31,239,30,210,31,211,31,76,31,54,31,54,30,110,31,31,31,3,31,154,31,154,30,154,29,154,31,31,31,15,31,83,31,83,30,109,31,140,31,140,30,60,31,87,31,4,31,12,31,129,31,129,30,129,29,129,28,127,31,60,31,67,31,154,31,154,30,140,31,164,31,85,31,94,31,96,31,28,31,28,30,10,31,10,30,198,31,198,30,198,29,54,31,131,31,98,31,85,31,213,31,77,31,77,30,249,31,202,31,168,31,25,31,187,31,93,31,93,30,34,31,167,31,143,31,86,31,86,30,102,31,150,31,150,30,107,31,191,31,30,31,255,31,255,30,78,31,144,31,220,31,44,31,44,30,241,31,37,31,164,31,34,31,34,30,34,29,34,28,231,31,231,30,231,29,31,31,238,31,144,31,88,31,184,31,123,31,200,31,101,31,207,31,155,31,182,31,140,31,140,30,128,31,213,31,213,30,55,31,136,31,136,30,38,31,38,30,35,31,35,30,248,31,82,31,82,30,118,31,161,31,134,31,20,31,146,31,81,31,81,30,16,31,95,31,95,30,196,31,196,31,157,31,29,31,153,31,212,31,228,31,157,31,63,31,98,31,84,31,38,31,13,31,33,31,201,31,201,30,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
