-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_18 is
end project_tb_18;

architecture project_tb_arch_18 of project_tb_18 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 206;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (191,0,235,0,2,0,0,0,106,0,50,0,218,0,0,0,168,0,134,0,0,0,211,0,84,0,115,0,0,0,235,0,71,0,139,0,102,0,1,0,84,0,0,0,158,0,154,0,137,0,138,0,135,0,82,0,0,0,197,0,192,0,0,0,86,0,110,0,235,0,209,0,166,0,111,0,119,0,239,0,31,0,195,0,251,0,187,0,112,0,31,0,241,0,135,0,137,0,197,0,228,0,104,0,48,0,0,0,139,0,44,0,201,0,147,0,0,0,52,0,74,0,0,0,0,0,213,0,134,0,76,0,254,0,211,0,22,0,0,0,60,0,172,0,199,0,227,0,43,0,114,0,70,0,248,0,109,0,79,0,0,0,113,0,0,0,0,0,160,0,0,0,38,0,123,0,27,0,210,0,8,0,140,0,33,0,43,0,0,0,226,0,0,0,143,0,0,0,0,0,148,0,178,0,193,0,178,0,170,0,0,0,235,0,175,0,166,0,73,0,0,0,49,0,0,0,49,0,34,0,176,0,0,0,165,0,229,0,0,0,139,0,0,0,189,0,231,0,143,0,60,0,0,0,11,0,92,0,212,0,238,0,227,0,47,0,180,0,52,0,67,0,214,0,120,0,0,0,79,0,118,0,86,0,163,0,168,0,72,0,24,0,251,0,116,0,162,0,83,0,223,0,197,0,0,0,229,0,59,0,142,0,68,0,231,0,135,0,69,0,98,0,0,0,245,0,148,0,163,0,132,0,122,0,0,0,66,0,104,0,125,0,160,0,14,0,219,0,0,0,238,0,120,0,0,0,0,0,0,0,83,0,127,0,0,0,216,0,0,0,216,0,199,0,129,0,104,0,0,0,96,0,0,0,93,0,0,0,0,0,46,0,28,0,135,0,255,0,0,0,247,0,227,0,209,0,108,0,227,0,56,0);
signal scenario_full  : scenario_type := (191,31,235,31,2,31,2,30,106,31,50,31,218,31,218,30,168,31,134,31,134,30,211,31,84,31,115,31,115,30,235,31,71,31,139,31,102,31,1,31,84,31,84,30,158,31,154,31,137,31,138,31,135,31,82,31,82,30,197,31,192,31,192,30,86,31,110,31,235,31,209,31,166,31,111,31,119,31,239,31,31,31,195,31,251,31,187,31,112,31,31,31,241,31,135,31,137,31,197,31,228,31,104,31,48,31,48,30,139,31,44,31,201,31,147,31,147,30,52,31,74,31,74,30,74,29,213,31,134,31,76,31,254,31,211,31,22,31,22,30,60,31,172,31,199,31,227,31,43,31,114,31,70,31,248,31,109,31,79,31,79,30,113,31,113,30,113,29,160,31,160,30,38,31,123,31,27,31,210,31,8,31,140,31,33,31,43,31,43,30,226,31,226,30,143,31,143,30,143,29,148,31,178,31,193,31,178,31,170,31,170,30,235,31,175,31,166,31,73,31,73,30,49,31,49,30,49,31,34,31,176,31,176,30,165,31,229,31,229,30,139,31,139,30,189,31,231,31,143,31,60,31,60,30,11,31,92,31,212,31,238,31,227,31,47,31,180,31,52,31,67,31,214,31,120,31,120,30,79,31,118,31,86,31,163,31,168,31,72,31,24,31,251,31,116,31,162,31,83,31,223,31,197,31,197,30,229,31,59,31,142,31,68,31,231,31,135,31,69,31,98,31,98,30,245,31,148,31,163,31,132,31,122,31,122,30,66,31,104,31,125,31,160,31,14,31,219,31,219,30,238,31,120,31,120,30,120,29,120,28,83,31,127,31,127,30,216,31,216,30,216,31,199,31,129,31,104,31,104,30,96,31,96,30,93,31,93,30,93,29,46,31,28,31,135,31,255,31,255,30,247,31,227,31,209,31,108,31,227,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
