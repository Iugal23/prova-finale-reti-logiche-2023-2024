-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_907 is
end project_tb_907;

architecture project_tb_arch_907 of project_tb_907 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 194;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,25,0,177,0,62,0,221,0,125,0,207,0,0,0,141,0,106,0,89,0,0,0,78,0,0,0,0,0,70,0,234,0,52,0,62,0,196,0,47,0,210,0,87,0,0,0,250,0,231,0,123,0,148,0,226,0,234,0,80,0,0,0,83,0,0,0,54,0,100,0,156,0,87,0,56,0,54,0,0,0,69,0,85,0,42,0,211,0,0,0,172,0,195,0,25,0,0,0,230,0,77,0,215,0,118,0,246,0,76,0,27,0,249,0,145,0,224,0,43,0,239,0,86,0,56,0,0,0,226,0,159,0,254,0,14,0,137,0,143,0,45,0,16,0,216,0,241,0,90,0,168,0,0,0,0,0,74,0,1,0,101,0,131,0,32,0,251,0,77,0,198,0,243,0,48,0,57,0,222,0,215,0,162,0,26,0,0,0,192,0,27,0,51,0,77,0,23,0,127,0,248,0,109,0,0,0,238,0,149,0,138,0,0,0,134,0,74,0,32,0,49,0,214,0,72,0,0,0,85,0,103,0,144,0,52,0,59,0,149,0,182,0,91,0,183,0,0,0,68,0,231,0,0,0,51,0,0,0,43,0,23,0,8,0,8,0,0,0,14,0,191,0,0,0,54,0,0,0,139,0,81,0,0,0,101,0,150,0,11,0,141,0,244,0,236,0,63,0,156,0,228,0,129,0,115,0,0,0,148,0,13,0,70,0,238,0,74,0,166,0,50,0,66,0,0,0,34,0,126,0,6,0,235,0,137,0,100,0,15,0,112,0,245,0,75,0,188,0,232,0,0,0,26,0,149,0,13,0,0,0,41,0,32,0,242,0,61,0,240,0,214,0,29,0,16,0,129,0,252,0,88,0,207,0,72,0);
signal scenario_full  : scenario_type := (136,31,25,31,177,31,62,31,221,31,125,31,207,31,207,30,141,31,106,31,89,31,89,30,78,31,78,30,78,29,70,31,234,31,52,31,62,31,196,31,47,31,210,31,87,31,87,30,250,31,231,31,123,31,148,31,226,31,234,31,80,31,80,30,83,31,83,30,54,31,100,31,156,31,87,31,56,31,54,31,54,30,69,31,85,31,42,31,211,31,211,30,172,31,195,31,25,31,25,30,230,31,77,31,215,31,118,31,246,31,76,31,27,31,249,31,145,31,224,31,43,31,239,31,86,31,56,31,56,30,226,31,159,31,254,31,14,31,137,31,143,31,45,31,16,31,216,31,241,31,90,31,168,31,168,30,168,29,74,31,1,31,101,31,131,31,32,31,251,31,77,31,198,31,243,31,48,31,57,31,222,31,215,31,162,31,26,31,26,30,192,31,27,31,51,31,77,31,23,31,127,31,248,31,109,31,109,30,238,31,149,31,138,31,138,30,134,31,74,31,32,31,49,31,214,31,72,31,72,30,85,31,103,31,144,31,52,31,59,31,149,31,182,31,91,31,183,31,183,30,68,31,231,31,231,30,51,31,51,30,43,31,23,31,8,31,8,31,8,30,14,31,191,31,191,30,54,31,54,30,139,31,81,31,81,30,101,31,150,31,11,31,141,31,244,31,236,31,63,31,156,31,228,31,129,31,115,31,115,30,148,31,13,31,70,31,238,31,74,31,166,31,50,31,66,31,66,30,34,31,126,31,6,31,235,31,137,31,100,31,15,31,112,31,245,31,75,31,188,31,232,31,232,30,26,31,149,31,13,31,13,30,41,31,32,31,242,31,61,31,240,31,214,31,29,31,16,31,129,31,252,31,88,31,207,31,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
