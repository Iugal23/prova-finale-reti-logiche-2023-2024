-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_933 is
end project_tb_933;

architecture project_tb_arch_933 of project_tb_933 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 851;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,158,0,99,0,107,0,20,0,106,0,0,0,189,0,125,0,86,0,44,0,134,0,0,0,31,0,250,0,0,0,246,0,121,0,71,0,205,0,187,0,201,0,119,0,8,0,211,0,0,0,0,0,0,0,247,0,176,0,99,0,153,0,167,0,115,0,252,0,0,0,107,0,157,0,2,0,91,0,0,0,0,0,62,0,200,0,237,0,147,0,0,0,57,0,76,0,0,0,140,0,77,0,70,0,123,0,179,0,96,0,0,0,165,0,86,0,148,0,248,0,128,0,11,0,215,0,0,0,1,0,210,0,212,0,245,0,11,0,113,0,93,0,42,0,119,0,75,0,93,0,160,0,152,0,0,0,42,0,0,0,0,0,37,0,57,0,97,0,59,0,0,0,225,0,28,0,199,0,135,0,60,0,78,0,153,0,1,0,47,0,102,0,22,0,29,0,249,0,177,0,107,0,232,0,0,0,220,0,0,0,59,0,0,0,195,0,82,0,47,0,101,0,121,0,0,0,185,0,0,0,131,0,0,0,14,0,89,0,255,0,137,0,0,0,39,0,185,0,233,0,0,0,141,0,234,0,0,0,235,0,224,0,0,0,140,0,11,0,145,0,64,0,130,0,53,0,206,0,173,0,97,0,32,0,135,0,61,0,4,0,74,0,76,0,148,0,123,0,116,0,59,0,97,0,93,0,247,0,171,0,0,0,156,0,227,0,86,0,228,0,55,0,47,0,41,0,127,0,246,0,102,0,0,0,253,0,173,0,0,0,242,0,24,0,97,0,220,0,124,0,88,0,172,0,55,0,69,0,0,0,0,0,112,0,40,0,26,0,35,0,202,0,227,0,146,0,219,0,0,0,15,0,0,0,127,0,0,0,247,0,0,0,0,0,151,0,0,0,12,0,147,0,38,0,0,0,248,0,28,0,228,0,225,0,130,0,182,0,174,0,97,0,221,0,88,0,140,0,194,0,163,0,171,0,0,0,0,0,40,0,206,0,0,0,220,0,216,0,0,0,15,0,221,0,2,0,0,0,235,0,83,0,0,0,29,0,159,0,160,0,111,0,0,0,0,0,128,0,244,0,195,0,182,0,37,0,254,0,67,0,20,0,0,0,178,0,0,0,135,0,206,0,207,0,226,0,158,0,43,0,255,0,65,0,165,0,117,0,129,0,140,0,65,0,103,0,16,0,16,0,83,0,254,0,96,0,173,0,0,0,68,0,244,0,179,0,162,0,178,0,0,0,189,0,28,0,138,0,45,0,215,0,213,0,236,0,0,0,107,0,62,0,0,0,250,0,0,0,39,0,0,0,208,0,1,0,180,0,118,0,98,0,0,0,0,0,21,0,133,0,196,0,0,0,129,0,99,0,194,0,65,0,53,0,0,0,212,0,240,0,103,0,144,0,96,0,229,0,0,0,195,0,0,0,209,0,192,0,0,0,187,0,69,0,170,0,0,0,0,0,33,0,82,0,129,0,212,0,152,0,230,0,107,0,236,0,0,0,0,0,0,0,0,0,128,0,0,0,192,0,177,0,21,0,125,0,224,0,33,0,0,0,247,0,241,0,64,0,222,0,237,0,159,0,234,0,17,0,140,0,197,0,0,0,194,0,122,0,53,0,57,0,154,0,232,0,1,0,182,0,89,0,100,0,242,0,207,0,225,0,240,0,94,0,38,0,250,0,210,0,0,0,167,0,206,0,0,0,85,0,0,0,151,0,7,0,121,0,48,0,38,0,27,0,0,0,185,0,39,0,176,0,243,0,149,0,86,0,161,0,82,0,69,0,115,0,226,0,0,0,85,0,130,0,229,0,204,0,113,0,241,0,121,0,214,0,0,0,136,0,115,0,0,0,0,0,249,0,137,0,100,0,82,0,111,0,78,0,74,0,220,0,247,0,42,0,33,0,0,0,122,0,154,0,0,0,184,0,195,0,81,0,89,0,113,0,56,0,179,0,16,0,191,0,203,0,23,0,110,0,0,0,149,0,0,0,69,0,12,0,59,0,150,0,204,0,215,0,68,0,41,0,145,0,82,0,177,0,80,0,75,0,153,0,246,0,197,0,200,0,6,0,238,0,228,0,73,0,0,0,84,0,0,0,89,0,155,0,210,0,222,0,150,0,75,0,153,0,243,0,5,0,0,0,192,0,14,0,68,0,213,0,235,0,165,0,107,0,0,0,153,0,99,0,0,0,79,0,0,0,148,0,218,0,73,0,0,0,135,0,0,0,0,0,19,0,93,0,0,0,208,0,105,0,93,0,29,0,0,0,212,0,148,0,135,0,241,0,0,0,0,0,127,0,83,0,20,0,230,0,195,0,56,0,215,0,0,0,212,0,120,0,0,0,75,0,168,0,139,0,27,0,255,0,67,0,62,0,170,0,143,0,219,0,130,0,92,0,250,0,135,0,203,0,0,0,222,0,64,0,23,0,0,0,8,0,94,0,155,0,195,0,32,0,123,0,0,0,36,0,89,0,127,0,142,0,186,0,100,0,211,0,250,0,0,0,224,0,10,0,77,0,0,0,97,0,236,0,187,0,174,0,0,0,68,0,65,0,201,0,0,0,244,0,133,0,0,0,77,0,209,0,126,0,198,0,0,0,80,0,51,0,21,0,0,0,240,0,200,0,43,0,0,0,149,0,214,0,59,0,37,0,52,0,0,0,167,0,34,0,150,0,64,0,236,0,181,0,57,0,19,0,157,0,0,0,190,0,91,0,0,0,241,0,0,0,0,0,0,0,119,0,0,0,0,0,253,0,0,0,77,0,0,0,214,0,26,0,236,0,246,0,34,0,203,0,0,0,38,0,178,0,137,0,119,0,21,0,238,0,103,0,155,0,191,0,171,0,223,0,158,0,23,0,234,0,222,0,107,0,239,0,63,0,98,0,125,0,187,0,32,0,226,0,195,0,143,0,24,0,0,0,75,0,156,0,0,0,195,0,62,0,237,0,95,0,0,0,81,0,248,0,55,0,93,0,193,0,107,0,69,0,49,0,222,0,4,0,119,0,104,0,0,0,0,0,178,0,0,0,0,0,53,0,111,0,19,0,100,0,0,0,107,0,3,0,0,0,0,0,203,0,100,0,0,0,12,0,105,0,125,0,211,0,215,0,67,0,111,0,255,0,70,0,32,0,0,0,134,0,94,0,87,0,0,0,243,0,236,0,135,0,0,0,91,0,36,0,50,0,64,0,0,0,173,0,232,0,94,0,188,0,210,0,55,0,80,0,75,0,89,0,235,0,0,0,66,0,70,0,93,0,251,0,104,0,0,0,213,0,34,0,0,0,0,0,207,0,207,0,36,0,0,0,70,0,0,0,192,0,119,0,0,0,4,0,111,0,0,0,191,0,194,0,254,0,160,0,187,0,0,0,184,0,64,0,0,0,251,0,18,0,184,0,23,0,11,0,147,0,67,0,184,0,199,0,143,0,140,0,255,0,206,0,166,0,0,0,0,0,66,0,209,0,76,0,150,0,111,0,52,0,181,0,16,0,0,0,250,0,82,0,0,0,199,0,164,0,7,0,0,0,0,0,53,0,32,0,239,0,179,0,176,0,0,0,68,0,6,0,101,0,0,0,0,0,222,0,93,0,111,0,66,0,116,0,184,0,59,0,0,0,174,0,0,0,25,0,0,0,187,0,184,0,0,0,21,0,152,0,229,0,37,0,253,0,104,0,112,0,205,0,189,0,222,0,81,0,66,0,180,0,113,0,0,0,0,0,127,0,102,0,133,0,223,0,114,0,16,0,103,0,0,0,165,0,245,0,0,0,165,0,180,0,74,0,125,0,0,0,102,0,10,0,0,0,249,0,189,0);
signal scenario_full  : scenario_type := (245,31,158,31,99,31,107,31,20,31,106,31,106,30,189,31,125,31,86,31,44,31,134,31,134,30,31,31,250,31,250,30,246,31,121,31,71,31,205,31,187,31,201,31,119,31,8,31,211,31,211,30,211,29,211,28,247,31,176,31,99,31,153,31,167,31,115,31,252,31,252,30,107,31,157,31,2,31,91,31,91,30,91,29,62,31,200,31,237,31,147,31,147,30,57,31,76,31,76,30,140,31,77,31,70,31,123,31,179,31,96,31,96,30,165,31,86,31,148,31,248,31,128,31,11,31,215,31,215,30,1,31,210,31,212,31,245,31,11,31,113,31,93,31,42,31,119,31,75,31,93,31,160,31,152,31,152,30,42,31,42,30,42,29,37,31,57,31,97,31,59,31,59,30,225,31,28,31,199,31,135,31,60,31,78,31,153,31,1,31,47,31,102,31,22,31,29,31,249,31,177,31,107,31,232,31,232,30,220,31,220,30,59,31,59,30,195,31,82,31,47,31,101,31,121,31,121,30,185,31,185,30,131,31,131,30,14,31,89,31,255,31,137,31,137,30,39,31,185,31,233,31,233,30,141,31,234,31,234,30,235,31,224,31,224,30,140,31,11,31,145,31,64,31,130,31,53,31,206,31,173,31,97,31,32,31,135,31,61,31,4,31,74,31,76,31,148,31,123,31,116,31,59,31,97,31,93,31,247,31,171,31,171,30,156,31,227,31,86,31,228,31,55,31,47,31,41,31,127,31,246,31,102,31,102,30,253,31,173,31,173,30,242,31,24,31,97,31,220,31,124,31,88,31,172,31,55,31,69,31,69,30,69,29,112,31,40,31,26,31,35,31,202,31,227,31,146,31,219,31,219,30,15,31,15,30,127,31,127,30,247,31,247,30,247,29,151,31,151,30,12,31,147,31,38,31,38,30,248,31,28,31,228,31,225,31,130,31,182,31,174,31,97,31,221,31,88,31,140,31,194,31,163,31,171,31,171,30,171,29,40,31,206,31,206,30,220,31,216,31,216,30,15,31,221,31,2,31,2,30,235,31,83,31,83,30,29,31,159,31,160,31,111,31,111,30,111,29,128,31,244,31,195,31,182,31,37,31,254,31,67,31,20,31,20,30,178,31,178,30,135,31,206,31,207,31,226,31,158,31,43,31,255,31,65,31,165,31,117,31,129,31,140,31,65,31,103,31,16,31,16,31,83,31,254,31,96,31,173,31,173,30,68,31,244,31,179,31,162,31,178,31,178,30,189,31,28,31,138,31,45,31,215,31,213,31,236,31,236,30,107,31,62,31,62,30,250,31,250,30,39,31,39,30,208,31,1,31,180,31,118,31,98,31,98,30,98,29,21,31,133,31,196,31,196,30,129,31,99,31,194,31,65,31,53,31,53,30,212,31,240,31,103,31,144,31,96,31,229,31,229,30,195,31,195,30,209,31,192,31,192,30,187,31,69,31,170,31,170,30,170,29,33,31,82,31,129,31,212,31,152,31,230,31,107,31,236,31,236,30,236,29,236,28,236,27,128,31,128,30,192,31,177,31,21,31,125,31,224,31,33,31,33,30,247,31,241,31,64,31,222,31,237,31,159,31,234,31,17,31,140,31,197,31,197,30,194,31,122,31,53,31,57,31,154,31,232,31,1,31,182,31,89,31,100,31,242,31,207,31,225,31,240,31,94,31,38,31,250,31,210,31,210,30,167,31,206,31,206,30,85,31,85,30,151,31,7,31,121,31,48,31,38,31,27,31,27,30,185,31,39,31,176,31,243,31,149,31,86,31,161,31,82,31,69,31,115,31,226,31,226,30,85,31,130,31,229,31,204,31,113,31,241,31,121,31,214,31,214,30,136,31,115,31,115,30,115,29,249,31,137,31,100,31,82,31,111,31,78,31,74,31,220,31,247,31,42,31,33,31,33,30,122,31,154,31,154,30,184,31,195,31,81,31,89,31,113,31,56,31,179,31,16,31,191,31,203,31,23,31,110,31,110,30,149,31,149,30,69,31,12,31,59,31,150,31,204,31,215,31,68,31,41,31,145,31,82,31,177,31,80,31,75,31,153,31,246,31,197,31,200,31,6,31,238,31,228,31,73,31,73,30,84,31,84,30,89,31,155,31,210,31,222,31,150,31,75,31,153,31,243,31,5,31,5,30,192,31,14,31,68,31,213,31,235,31,165,31,107,31,107,30,153,31,99,31,99,30,79,31,79,30,148,31,218,31,73,31,73,30,135,31,135,30,135,29,19,31,93,31,93,30,208,31,105,31,93,31,29,31,29,30,212,31,148,31,135,31,241,31,241,30,241,29,127,31,83,31,20,31,230,31,195,31,56,31,215,31,215,30,212,31,120,31,120,30,75,31,168,31,139,31,27,31,255,31,67,31,62,31,170,31,143,31,219,31,130,31,92,31,250,31,135,31,203,31,203,30,222,31,64,31,23,31,23,30,8,31,94,31,155,31,195,31,32,31,123,31,123,30,36,31,89,31,127,31,142,31,186,31,100,31,211,31,250,31,250,30,224,31,10,31,77,31,77,30,97,31,236,31,187,31,174,31,174,30,68,31,65,31,201,31,201,30,244,31,133,31,133,30,77,31,209,31,126,31,198,31,198,30,80,31,51,31,21,31,21,30,240,31,200,31,43,31,43,30,149,31,214,31,59,31,37,31,52,31,52,30,167,31,34,31,150,31,64,31,236,31,181,31,57,31,19,31,157,31,157,30,190,31,91,31,91,30,241,31,241,30,241,29,241,28,119,31,119,30,119,29,253,31,253,30,77,31,77,30,214,31,26,31,236,31,246,31,34,31,203,31,203,30,38,31,178,31,137,31,119,31,21,31,238,31,103,31,155,31,191,31,171,31,223,31,158,31,23,31,234,31,222,31,107,31,239,31,63,31,98,31,125,31,187,31,32,31,226,31,195,31,143,31,24,31,24,30,75,31,156,31,156,30,195,31,62,31,237,31,95,31,95,30,81,31,248,31,55,31,93,31,193,31,107,31,69,31,49,31,222,31,4,31,119,31,104,31,104,30,104,29,178,31,178,30,178,29,53,31,111,31,19,31,100,31,100,30,107,31,3,31,3,30,3,29,203,31,100,31,100,30,12,31,105,31,125,31,211,31,215,31,67,31,111,31,255,31,70,31,32,31,32,30,134,31,94,31,87,31,87,30,243,31,236,31,135,31,135,30,91,31,36,31,50,31,64,31,64,30,173,31,232,31,94,31,188,31,210,31,55,31,80,31,75,31,89,31,235,31,235,30,66,31,70,31,93,31,251,31,104,31,104,30,213,31,34,31,34,30,34,29,207,31,207,31,36,31,36,30,70,31,70,30,192,31,119,31,119,30,4,31,111,31,111,30,191,31,194,31,254,31,160,31,187,31,187,30,184,31,64,31,64,30,251,31,18,31,184,31,23,31,11,31,147,31,67,31,184,31,199,31,143,31,140,31,255,31,206,31,166,31,166,30,166,29,66,31,209,31,76,31,150,31,111,31,52,31,181,31,16,31,16,30,250,31,82,31,82,30,199,31,164,31,7,31,7,30,7,29,53,31,32,31,239,31,179,31,176,31,176,30,68,31,6,31,101,31,101,30,101,29,222,31,93,31,111,31,66,31,116,31,184,31,59,31,59,30,174,31,174,30,25,31,25,30,187,31,184,31,184,30,21,31,152,31,229,31,37,31,253,31,104,31,112,31,205,31,189,31,222,31,81,31,66,31,180,31,113,31,113,30,113,29,127,31,102,31,133,31,223,31,114,31,16,31,103,31,103,30,165,31,245,31,245,30,165,31,180,31,74,31,125,31,125,30,102,31,10,31,10,30,249,31,189,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
