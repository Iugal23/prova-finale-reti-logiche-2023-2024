-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_856 is
end project_tb_856;

architecture project_tb_arch_856 of project_tb_856 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 345;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (204,0,172,0,94,0,58,0,24,0,149,0,104,0,113,0,11,0,241,0,248,0,157,0,178,0,26,0,76,0,75,0,0,0,243,0,53,0,250,0,0,0,159,0,34,0,166,0,0,0,9,0,84,0,138,0,251,0,82,0,62,0,61,0,214,0,102,0,185,0,139,0,108,0,73,0,145,0,0,0,249,0,115,0,252,0,158,0,119,0,97,0,116,0,89,0,72,0,0,0,201,0,0,0,183,0,234,0,50,0,0,0,0,0,197,0,39,0,41,0,230,0,105,0,145,0,199,0,27,0,240,0,73,0,162,0,165,0,0,0,0,0,165,0,231,0,44,0,227,0,143,0,36,0,112,0,180,0,0,0,0,0,25,0,0,0,43,0,84,0,106,0,52,0,0,0,121,0,209,0,129,0,189,0,29,0,88,0,130,0,44,0,4,0,77,0,0,0,169,0,141,0,93,0,178,0,115,0,106,0,89,0,15,0,156,0,128,0,167,0,235,0,100,0,0,0,0,0,180,0,129,0,254,0,0,0,52,0,0,0,240,0,203,0,10,0,239,0,239,0,161,0,114,0,71,0,84,0,235,0,114,0,0,0,126,0,0,0,38,0,0,0,136,0,20,0,82,0,40,0,80,0,245,0,187,0,239,0,31,0,36,0,0,0,218,0,192,0,0,0,0,0,0,0,52,0,126,0,72,0,197,0,77,0,0,0,76,0,115,0,170,0,63,0,67,0,0,0,154,0,65,0,234,0,164,0,249,0,229,0,18,0,186,0,230,0,16,0,54,0,190,0,13,0,92,0,13,0,115,0,79,0,42,0,253,0,57,0,135,0,33,0,180,0,30,0,206,0,0,0,15,0,0,0,0,0,0,0,158,0,159,0,86,0,172,0,195,0,249,0,243,0,0,0,0,0,169,0,15,0,93,0,128,0,0,0,53,0,0,0,0,0,58,0,0,0,174,0,189,0,102,0,48,0,234,0,72,0,186,0,0,0,0,0,141,0,0,0,0,0,67,0,30,0,0,0,91,0,117,0,107,0,194,0,63,0,50,0,28,0,85,0,0,0,213,0,129,0,36,0,59,0,0,0,31,0,0,0,0,0,153,0,0,0,0,0,135,0,225,0,0,0,9,0,0,0,0,0,12,0,15,0,172,0,69,0,156,0,107,0,76,0,0,0,26,0,223,0,142,0,66,0,22,0,206,0,129,0,81,0,0,0,0,0,238,0,154,0,0,0,188,0,247,0,80,0,135,0,115,0,34,0,136,0,0,0,117,0,251,0,236,0,97,0,58,0,0,0,0,0,0,0,176,0,98,0,204,0,20,0,193,0,0,0,86,0,222,0,79,0,7,0,225,0,47,0,186,0,40,0,133,0,188,0,217,0,56,0,27,0,211,0,118,0,239,0,38,0,161,0,0,0,151,0,0,0,143,0,143,0,97,0,48,0,34,0,17,0,15,0,147,0,253,0,110,0,90,0,230,0,143,0,157,0,0,0,35,0,24,0,195,0,0,0,73,0,248,0,146,0,7,0,0,0,65,0,157,0,118,0);
signal scenario_full  : scenario_type := (204,31,172,31,94,31,58,31,24,31,149,31,104,31,113,31,11,31,241,31,248,31,157,31,178,31,26,31,76,31,75,31,75,30,243,31,53,31,250,31,250,30,159,31,34,31,166,31,166,30,9,31,84,31,138,31,251,31,82,31,62,31,61,31,214,31,102,31,185,31,139,31,108,31,73,31,145,31,145,30,249,31,115,31,252,31,158,31,119,31,97,31,116,31,89,31,72,31,72,30,201,31,201,30,183,31,234,31,50,31,50,30,50,29,197,31,39,31,41,31,230,31,105,31,145,31,199,31,27,31,240,31,73,31,162,31,165,31,165,30,165,29,165,31,231,31,44,31,227,31,143,31,36,31,112,31,180,31,180,30,180,29,25,31,25,30,43,31,84,31,106,31,52,31,52,30,121,31,209,31,129,31,189,31,29,31,88,31,130,31,44,31,4,31,77,31,77,30,169,31,141,31,93,31,178,31,115,31,106,31,89,31,15,31,156,31,128,31,167,31,235,31,100,31,100,30,100,29,180,31,129,31,254,31,254,30,52,31,52,30,240,31,203,31,10,31,239,31,239,31,161,31,114,31,71,31,84,31,235,31,114,31,114,30,126,31,126,30,38,31,38,30,136,31,20,31,82,31,40,31,80,31,245,31,187,31,239,31,31,31,36,31,36,30,218,31,192,31,192,30,192,29,192,28,52,31,126,31,72,31,197,31,77,31,77,30,76,31,115,31,170,31,63,31,67,31,67,30,154,31,65,31,234,31,164,31,249,31,229,31,18,31,186,31,230,31,16,31,54,31,190,31,13,31,92,31,13,31,115,31,79,31,42,31,253,31,57,31,135,31,33,31,180,31,30,31,206,31,206,30,15,31,15,30,15,29,15,28,158,31,159,31,86,31,172,31,195,31,249,31,243,31,243,30,243,29,169,31,15,31,93,31,128,31,128,30,53,31,53,30,53,29,58,31,58,30,174,31,189,31,102,31,48,31,234,31,72,31,186,31,186,30,186,29,141,31,141,30,141,29,67,31,30,31,30,30,91,31,117,31,107,31,194,31,63,31,50,31,28,31,85,31,85,30,213,31,129,31,36,31,59,31,59,30,31,31,31,30,31,29,153,31,153,30,153,29,135,31,225,31,225,30,9,31,9,30,9,29,12,31,15,31,172,31,69,31,156,31,107,31,76,31,76,30,26,31,223,31,142,31,66,31,22,31,206,31,129,31,81,31,81,30,81,29,238,31,154,31,154,30,188,31,247,31,80,31,135,31,115,31,34,31,136,31,136,30,117,31,251,31,236,31,97,31,58,31,58,30,58,29,58,28,176,31,98,31,204,31,20,31,193,31,193,30,86,31,222,31,79,31,7,31,225,31,47,31,186,31,40,31,133,31,188,31,217,31,56,31,27,31,211,31,118,31,239,31,38,31,161,31,161,30,151,31,151,30,143,31,143,31,97,31,48,31,34,31,17,31,15,31,147,31,253,31,110,31,90,31,230,31,143,31,157,31,157,30,35,31,24,31,195,31,195,30,73,31,248,31,146,31,7,31,7,30,65,31,157,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
