-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 660;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,203,0,0,0,172,0,134,0,57,0,45,0,0,0,27,0,0,0,120,0,115,0,1,0,0,0,49,0,21,0,0,0,67,0,149,0,162,0,202,0,185,0,185,0,101,0,0,0,146,0,163,0,30,0,0,0,0,0,255,0,55,0,157,0,137,0,255,0,199,0,221,0,16,0,0,0,31,0,1,0,10,0,92,0,181,0,57,0,85,0,60,0,30,0,0,0,0,0,19,0,0,0,79,0,212,0,98,0,22,0,228,0,102,0,151,0,163,0,165,0,217,0,239,0,26,0,0,0,208,0,62,0,155,0,0,0,110,0,16,0,105,0,0,0,167,0,15,0,8,0,255,0,125,0,34,0,219,0,230,0,26,0,233,0,106,0,0,0,154,0,0,0,220,0,0,0,165,0,148,0,95,0,0,0,94,0,216,0,1,0,18,0,11,0,152,0,3,0,0,0,43,0,70,0,12,0,106,0,204,0,0,0,0,0,248,0,90,0,205,0,123,0,32,0,197,0,0,0,207,0,73,0,147,0,229,0,95,0,249,0,226,0,185,0,122,0,0,0,170,0,210,0,19,0,25,0,45,0,105,0,95,0,188,0,170,0,78,0,110,0,7,0,0,0,145,0,140,0,182,0,148,0,0,0,166,0,136,0,138,0,9,0,254,0,170,0,114,0,130,0,7,0,96,0,232,0,222,0,218,0,171,0,0,0,131,0,63,0,71,0,153,0,194,0,0,0,28,0,68,0,0,0,0,0,150,0,10,0,143,0,90,0,170,0,147,0,0,0,92,0,216,0,15,0,13,0,237,0,0,0,76,0,254,0,0,0,3,0,191,0,224,0,25,0,120,0,158,0,0,0,52,0,112,0,129,0,169,0,91,0,87,0,0,0,141,0,200,0,174,0,216,0,117,0,0,0,3,0,4,0,223,0,0,0,0,0,183,0,250,0,0,0,177,0,9,0,0,0,219,0,27,0,170,0,66,0,169,0,0,0,0,0,180,0,71,0,33,0,201,0,116,0,92,0,73,0,155,0,0,0,0,0,214,0,204,0,42,0,119,0,81,0,188,0,0,0,176,0,13,0,120,0,167,0,0,0,0,0,202,0,90,0,0,0,0,0,164,0,253,0,173,0,0,0,247,0,142,0,79,0,156,0,0,0,26,0,217,0,224,0,242,0,184,0,21,0,134,0,241,0,8,0,214,0,129,0,183,0,15,0,201,0,79,0,219,0,169,0,218,0,72,0,134,0,119,0,178,0,6,0,129,0,0,0,0,0,6,0,34,0,7,0,0,0,120,0,191,0,93,0,12,0,228,0,202,0,86,0,174,0,183,0,154,0,22,0,65,0,50,0,60,0,0,0,0,0,28,0,169,0,0,0,187,0,160,0,0,0,179,0,187,0,0,0,60,0,0,0,240,0,164,0,53,0,122,0,0,0,123,0,170,0,49,0,120,0,121,0,0,0,11,0,216,0,127,0,15,0,166,0,26,0,252,0,32,0,0,0,63,0,15,0,52,0,142,0,211,0,117,0,204,0,83,0,0,0,233,0,39,0,146,0,235,0,0,0,44,0,0,0,99,0,0,0,242,0,0,0,101,0,237,0,171,0,0,0,0,0,56,0,139,0,201,0,97,0,92,0,0,0,120,0,18,0,109,0,172,0,0,0,0,0,1,0,18,0,89,0,0,0,93,0,38,0,0,0,200,0,226,0,171,0,170,0,0,0,0,0,102,0,58,0,0,0,42,0,159,0,59,0,236,0,113,0,78,0,0,0,39,0,122,0,44,0,162,0,169,0,253,0,0,0,137,0,111,0,18,0,197,0,175,0,130,0,99,0,0,0,221,0,3,0,145,0,199,0,0,0,70,0,51,0,148,0,0,0,0,0,125,0,9,0,46,0,50,0,239,0,230,0,232,0,115,0,242,0,90,0,50,0,0,0,241,0,248,0,183,0,175,0,27,0,101,0,37,0,87,0,57,0,227,0,90,0,101,0,0,0,122,0,0,0,157,0,84,0,219,0,0,0,81,0,138,0,80,0,79,0,224,0,50,0,241,0,37,0,17,0,211,0,154,0,73,0,176,0,215,0,181,0,229,0,0,0,102,0,139,0,102,0,0,0,12,0,55,0,0,0,0,0,26,0,0,0,122,0,5,0,36,0,121,0,133,0,0,0,224,0,0,0,0,0,40,0,0,0,110,0,219,0,20,0,106,0,0,0,251,0,78,0,25,0,76,0,85,0,193,0,248,0,248,0,105,0,161,0,224,0,199,0,121,0,251,0,0,0,0,0,0,0,62,0,179,0,28,0,0,0,44,0,39,0,36,0,44,0,76,0,51,0,155,0,0,0,150,0,160,0,149,0,179,0,250,0,225,0,0,0,25,0,137,0,14,0,131,0,0,0,3,0,0,0,0,0,107,0,211,0,0,0,123,0,135,0,219,0,231,0,0,0,84,0,0,0,249,0,42,0,160,0,246,0,252,0,67,0,81,0,212,0,167,0,0,0,131,0,58,0,79,0,0,0,80,0,116,0,0,0,49,0,110,0,1,0,242,0,50,0,0,0,0,0,52,0,145,0,137,0,127,0,152,0,134,0,172,0,0,0,0,0,0,0,98,0,198,0,192,0,235,0,0,0,155,0,0,0,254,0,54,0,173,0,112,0,133,0,60,0,128,0,225,0,0,0,0,0,50,0,189,0,119,0,22,0,177,0,94,0,123,0,0,0,119,0,160,0,240,0,0,0,121,0,144,0,76,0,192,0,148,0,0,0,254,0,106,0,72,0,26,0,83,0,198,0,178,0,0,0,21,0,74,0,203,0,0,0,219,0,35,0,182,0,103,0,99,0,101,0,222,0,126,0,0,0,25,0,0,0,0,0,168,0,3,0,5,0,0,0,0,0,204,0,0,0,218,0,11,0,0,0,1,0,58,0,221,0,20,0,0,0,0,0,0,0,230,0,217,0);
signal scenario_full  : scenario_type := (0,0,203,31,203,30,172,31,134,31,57,31,45,31,45,30,27,31,27,30,120,31,115,31,1,31,1,30,49,31,21,31,21,30,67,31,149,31,162,31,202,31,185,31,185,31,101,31,101,30,146,31,163,31,30,31,30,30,30,29,255,31,55,31,157,31,137,31,255,31,199,31,221,31,16,31,16,30,31,31,1,31,10,31,92,31,181,31,57,31,85,31,60,31,30,31,30,30,30,29,19,31,19,30,79,31,212,31,98,31,22,31,228,31,102,31,151,31,163,31,165,31,217,31,239,31,26,31,26,30,208,31,62,31,155,31,155,30,110,31,16,31,105,31,105,30,167,31,15,31,8,31,255,31,125,31,34,31,219,31,230,31,26,31,233,31,106,31,106,30,154,31,154,30,220,31,220,30,165,31,148,31,95,31,95,30,94,31,216,31,1,31,18,31,11,31,152,31,3,31,3,30,43,31,70,31,12,31,106,31,204,31,204,30,204,29,248,31,90,31,205,31,123,31,32,31,197,31,197,30,207,31,73,31,147,31,229,31,95,31,249,31,226,31,185,31,122,31,122,30,170,31,210,31,19,31,25,31,45,31,105,31,95,31,188,31,170,31,78,31,110,31,7,31,7,30,145,31,140,31,182,31,148,31,148,30,166,31,136,31,138,31,9,31,254,31,170,31,114,31,130,31,7,31,96,31,232,31,222,31,218,31,171,31,171,30,131,31,63,31,71,31,153,31,194,31,194,30,28,31,68,31,68,30,68,29,150,31,10,31,143,31,90,31,170,31,147,31,147,30,92,31,216,31,15,31,13,31,237,31,237,30,76,31,254,31,254,30,3,31,191,31,224,31,25,31,120,31,158,31,158,30,52,31,112,31,129,31,169,31,91,31,87,31,87,30,141,31,200,31,174,31,216,31,117,31,117,30,3,31,4,31,223,31,223,30,223,29,183,31,250,31,250,30,177,31,9,31,9,30,219,31,27,31,170,31,66,31,169,31,169,30,169,29,180,31,71,31,33,31,201,31,116,31,92,31,73,31,155,31,155,30,155,29,214,31,204,31,42,31,119,31,81,31,188,31,188,30,176,31,13,31,120,31,167,31,167,30,167,29,202,31,90,31,90,30,90,29,164,31,253,31,173,31,173,30,247,31,142,31,79,31,156,31,156,30,26,31,217,31,224,31,242,31,184,31,21,31,134,31,241,31,8,31,214,31,129,31,183,31,15,31,201,31,79,31,219,31,169,31,218,31,72,31,134,31,119,31,178,31,6,31,129,31,129,30,129,29,6,31,34,31,7,31,7,30,120,31,191,31,93,31,12,31,228,31,202,31,86,31,174,31,183,31,154,31,22,31,65,31,50,31,60,31,60,30,60,29,28,31,169,31,169,30,187,31,160,31,160,30,179,31,187,31,187,30,60,31,60,30,240,31,164,31,53,31,122,31,122,30,123,31,170,31,49,31,120,31,121,31,121,30,11,31,216,31,127,31,15,31,166,31,26,31,252,31,32,31,32,30,63,31,15,31,52,31,142,31,211,31,117,31,204,31,83,31,83,30,233,31,39,31,146,31,235,31,235,30,44,31,44,30,99,31,99,30,242,31,242,30,101,31,237,31,171,31,171,30,171,29,56,31,139,31,201,31,97,31,92,31,92,30,120,31,18,31,109,31,172,31,172,30,172,29,1,31,18,31,89,31,89,30,93,31,38,31,38,30,200,31,226,31,171,31,170,31,170,30,170,29,102,31,58,31,58,30,42,31,159,31,59,31,236,31,113,31,78,31,78,30,39,31,122,31,44,31,162,31,169,31,253,31,253,30,137,31,111,31,18,31,197,31,175,31,130,31,99,31,99,30,221,31,3,31,145,31,199,31,199,30,70,31,51,31,148,31,148,30,148,29,125,31,9,31,46,31,50,31,239,31,230,31,232,31,115,31,242,31,90,31,50,31,50,30,241,31,248,31,183,31,175,31,27,31,101,31,37,31,87,31,57,31,227,31,90,31,101,31,101,30,122,31,122,30,157,31,84,31,219,31,219,30,81,31,138,31,80,31,79,31,224,31,50,31,241,31,37,31,17,31,211,31,154,31,73,31,176,31,215,31,181,31,229,31,229,30,102,31,139,31,102,31,102,30,12,31,55,31,55,30,55,29,26,31,26,30,122,31,5,31,36,31,121,31,133,31,133,30,224,31,224,30,224,29,40,31,40,30,110,31,219,31,20,31,106,31,106,30,251,31,78,31,25,31,76,31,85,31,193,31,248,31,248,31,105,31,161,31,224,31,199,31,121,31,251,31,251,30,251,29,251,28,62,31,179,31,28,31,28,30,44,31,39,31,36,31,44,31,76,31,51,31,155,31,155,30,150,31,160,31,149,31,179,31,250,31,225,31,225,30,25,31,137,31,14,31,131,31,131,30,3,31,3,30,3,29,107,31,211,31,211,30,123,31,135,31,219,31,231,31,231,30,84,31,84,30,249,31,42,31,160,31,246,31,252,31,67,31,81,31,212,31,167,31,167,30,131,31,58,31,79,31,79,30,80,31,116,31,116,30,49,31,110,31,1,31,242,31,50,31,50,30,50,29,52,31,145,31,137,31,127,31,152,31,134,31,172,31,172,30,172,29,172,28,98,31,198,31,192,31,235,31,235,30,155,31,155,30,254,31,54,31,173,31,112,31,133,31,60,31,128,31,225,31,225,30,225,29,50,31,189,31,119,31,22,31,177,31,94,31,123,31,123,30,119,31,160,31,240,31,240,30,121,31,144,31,76,31,192,31,148,31,148,30,254,31,106,31,72,31,26,31,83,31,198,31,178,31,178,30,21,31,74,31,203,31,203,30,219,31,35,31,182,31,103,31,99,31,101,31,222,31,126,31,126,30,25,31,25,30,25,29,168,31,3,31,5,31,5,30,5,29,204,31,204,30,218,31,11,31,11,30,1,31,58,31,221,31,20,31,20,30,20,29,20,28,230,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
