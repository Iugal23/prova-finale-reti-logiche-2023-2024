-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_479 is
end project_tb_479;

architecture project_tb_arch_479 of project_tb_479 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 776;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (111,0,0,0,145,0,0,0,86,0,235,0,37,0,137,0,4,0,0,0,160,0,145,0,149,0,0,0,226,0,0,0,97,0,175,0,0,0,0,0,0,0,0,0,176,0,158,0,128,0,126,0,5,0,72,0,253,0,0,0,0,0,0,0,0,0,109,0,196,0,0,0,0,0,90,0,25,0,202,0,125,0,107,0,207,0,158,0,31,0,241,0,0,0,240,0,0,0,65,0,111,0,252,0,0,0,161,0,113,0,192,0,0,0,113,0,186,0,11,0,130,0,105,0,136,0,24,0,233,0,53,0,122,0,192,0,204,0,201,0,166,0,103,0,194,0,62,0,254,0,21,0,0,0,74,0,0,0,0,0,68,0,228,0,239,0,179,0,17,0,4,0,138,0,0,0,0,0,163,0,194,0,166,0,95,0,1,0,0,0,133,0,0,0,202,0,0,0,171,0,34,0,0,0,14,0,0,0,207,0,143,0,0,0,0,0,58,0,215,0,0,0,46,0,42,0,184,0,249,0,100,0,159,0,0,0,233,0,232,0,76,0,217,0,86,0,235,0,38,0,1,0,159,0,237,0,0,0,216,0,129,0,119,0,198,0,0,0,65,0,68,0,0,0,213,0,17,0,42,0,0,0,0,0,194,0,0,0,89,0,30,0,252,0,77,0,62,0,0,0,199,0,0,0,136,0,181,0,44,0,147,0,0,0,119,0,118,0,221,0,57,0,185,0,185,0,5,0,77,0,196,0,5,0,102,0,92,0,100,0,0,0,0,0,47,0,44,0,43,0,132,0,55,0,59,0,51,0,0,0,254,0,55,0,70,0,140,0,37,0,0,0,227,0,182,0,120,0,250,0,192,0,16,0,238,0,182,0,0,0,0,0,0,0,75,0,3,0,0,0,18,0,144,0,14,0,205,0,253,0,89,0,95,0,129,0,233,0,251,0,44,0,236,0,0,0,159,0,69,0,150,0,0,0,23,0,187,0,218,0,113,0,0,0,244,0,110,0,28,0,0,0,0,0,165,0,0,0,12,0,189,0,97,0,1,0,0,0,100,0,14,0,10,0,37,0,228,0,197,0,163,0,0,0,137,0,0,0,84,0,49,0,0,0,0,0,78,0,160,0,39,0,0,0,239,0,120,0,124,0,216,0,57,0,92,0,88,0,197,0,64,0,110,0,0,0,138,0,77,0,70,0,132,0,167,0,120,0,0,0,121,0,0,0,116,0,189,0,141,0,0,0,247,0,22,0,155,0,0,0,161,0,116,0,0,0,223,0,184,0,83,0,179,0,0,0,138,0,116,0,92,0,0,0,87,0,127,0,148,0,212,0,58,0,223,0,50,0,237,0,38,0,223,0,130,0,149,0,115,0,99,0,202,0,232,0,51,0,118,0,172,0,80,0,0,0,49,0,65,0,35,0,197,0,0,0,191,0,238,0,138,0,0,0,255,0,55,0,0,0,0,0,147,0,127,0,45,0,252,0,0,0,201,0,208,0,218,0,91,0,122,0,39,0,253,0,133,0,0,0,44,0,200,0,147,0,115,0,87,0,20,0,18,0,120,0,72,0,0,0,181,0,223,0,57,0,72,0,0,0,163,0,113,0,199,0,174,0,51,0,187,0,246,0,20,0,57,0,0,0,19,0,77,0,0,0,0,0,0,0,51,0,108,0,106,0,5,0,0,0,67,0,161,0,0,0,171,0,66,0,0,0,90,0,216,0,158,0,208,0,49,0,252,0,136,0,0,0,5,0,102,0,0,0,0,0,217,0,90,0,176,0,196,0,132,0,253,0,236,0,149,0,219,0,0,0,0,0,248,0,165,0,180,0,49,0,132,0,3,0,2,0,24,0,25,0,245,0,5,0,253,0,81,0,110,0,254,0,249,0,113,0,38,0,135,0,164,0,132,0,50,0,98,0,85,0,33,0,84,0,192,0,54,0,0,0,120,0,243,0,0,0,87,0,50,0,0,0,221,0,0,0,77,0,155,0,197,0,53,0,240,0,70,0,196,0,236,0,253,0,237,0,0,0,209,0,0,0,74,0,145,0,89,0,34,0,223,0,78,0,41,0,0,0,19,0,100,0,211,0,254,0,24,0,8,0,94,0,125,0,0,0,84,0,93,0,14,0,0,0,95,0,71,0,8,0,189,0,183,0,199,0,117,0,203,0,189,0,101,0,0,0,136,0,94,0,67,0,0,0,109,0,189,0,4,0,15,0,186,0,203,0,121,0,18,0,0,0,0,0,86,0,0,0,0,0,243,0,0,0,76,0,139,0,241,0,168,0,154,0,214,0,135,0,0,0,153,0,0,0,28,0,0,0,74,0,122,0,107,0,140,0,146,0,108,0,207,0,244,0,51,0,148,0,0,0,131,0,30,0,57,0,251,0,183,0,144,0,242,0,213,0,147,0,111,0,93,0,21,0,222,0,101,0,46,0,0,0,247,0,188,0,165,0,246,0,153,0,129,0,138,0,49,0,6,0,171,0,214,0,76,0,116,0,159,0,181,0,94,0,159,0,66,0,69,0,0,0,56,0,211,0,0,0,102,0,0,0,171,0,153,0,249,0,208,0,104,0,0,0,198,0,0,0,0,0,213,0,0,0,179,0,0,0,33,0,88,0,183,0,199,0,0,0,121,0,125,0,203,0,19,0,156,0,110,0,5,0,190,0,196,0,0,0,228,0,167,0,254,0,150,0,139,0,54,0,72,0,96,0,0,0,176,0,173,0,0,0,109,0,145,0,0,0,0,0,155,0,29,0,165,0,200,0,0,0,0,0,36,0,138,0,112,0,44,0,112,0,210,0,233,0,50,0,238,0,189,0,172,0,147,0,0,0,0,0,96,0,141,0,57,0,0,0,204,0,230,0,87,0,0,0,242,0,189,0,25,0,181,0,28,0,239,0,139,0,208,0,141,0,0,0,56,0,172,0,228,0,238,0,0,0,177,0,203,0,0,0,29,0,209,0,122,0,46,0,53,0,130,0,34,0,128,0,246,0,0,0,164,0,231,0,27,0,88,0,81,0,87,0,59,0,241,0,25,0,0,0,0,0,22,0,10,0,0,0,191,0,25,0,6,0,131,0,242,0,41,0,82,0,0,0,212,0,97,0,236,0,185,0,154,0,82,0,0,0,176,0,92,0,76,0,122,0,180,0,201,0,236,0,24,0,152,0,42,0,21,0,194,0,194,0,173,0,179,0,236,0,0,0,123,0,6,0,243,0,64,0,10,0,0,0,91,0,80,0,109,0,0,0,163,0,33,0,225,0,244,0,210,0,140,0,79,0,0,0,157,0,34,0,105,0,41,0,251,0,180,0,0,0,114,0,157,0,254,0,120,0,0,0,120,0,97,0,8,0,0,0,90,0,47,0,28,0,60,0,82,0,152,0,18,0,212,0,1,0,120,0,189,0,135,0,167,0,146,0,0,0,93,0,249,0,151,0,84,0,96,0,0,0,215,0,0,0,46,0,235,0,72,0,0,0);
signal scenario_full  : scenario_type := (111,31,111,30,145,31,145,30,86,31,235,31,37,31,137,31,4,31,4,30,160,31,145,31,149,31,149,30,226,31,226,30,97,31,175,31,175,30,175,29,175,28,175,27,176,31,158,31,128,31,126,31,5,31,72,31,253,31,253,30,253,29,253,28,253,27,109,31,196,31,196,30,196,29,90,31,25,31,202,31,125,31,107,31,207,31,158,31,31,31,241,31,241,30,240,31,240,30,65,31,111,31,252,31,252,30,161,31,113,31,192,31,192,30,113,31,186,31,11,31,130,31,105,31,136,31,24,31,233,31,53,31,122,31,192,31,204,31,201,31,166,31,103,31,194,31,62,31,254,31,21,31,21,30,74,31,74,30,74,29,68,31,228,31,239,31,179,31,17,31,4,31,138,31,138,30,138,29,163,31,194,31,166,31,95,31,1,31,1,30,133,31,133,30,202,31,202,30,171,31,34,31,34,30,14,31,14,30,207,31,143,31,143,30,143,29,58,31,215,31,215,30,46,31,42,31,184,31,249,31,100,31,159,31,159,30,233,31,232,31,76,31,217,31,86,31,235,31,38,31,1,31,159,31,237,31,237,30,216,31,129,31,119,31,198,31,198,30,65,31,68,31,68,30,213,31,17,31,42,31,42,30,42,29,194,31,194,30,89,31,30,31,252,31,77,31,62,31,62,30,199,31,199,30,136,31,181,31,44,31,147,31,147,30,119,31,118,31,221,31,57,31,185,31,185,31,5,31,77,31,196,31,5,31,102,31,92,31,100,31,100,30,100,29,47,31,44,31,43,31,132,31,55,31,59,31,51,31,51,30,254,31,55,31,70,31,140,31,37,31,37,30,227,31,182,31,120,31,250,31,192,31,16,31,238,31,182,31,182,30,182,29,182,28,75,31,3,31,3,30,18,31,144,31,14,31,205,31,253,31,89,31,95,31,129,31,233,31,251,31,44,31,236,31,236,30,159,31,69,31,150,31,150,30,23,31,187,31,218,31,113,31,113,30,244,31,110,31,28,31,28,30,28,29,165,31,165,30,12,31,189,31,97,31,1,31,1,30,100,31,14,31,10,31,37,31,228,31,197,31,163,31,163,30,137,31,137,30,84,31,49,31,49,30,49,29,78,31,160,31,39,31,39,30,239,31,120,31,124,31,216,31,57,31,92,31,88,31,197,31,64,31,110,31,110,30,138,31,77,31,70,31,132,31,167,31,120,31,120,30,121,31,121,30,116,31,189,31,141,31,141,30,247,31,22,31,155,31,155,30,161,31,116,31,116,30,223,31,184,31,83,31,179,31,179,30,138,31,116,31,92,31,92,30,87,31,127,31,148,31,212,31,58,31,223,31,50,31,237,31,38,31,223,31,130,31,149,31,115,31,99,31,202,31,232,31,51,31,118,31,172,31,80,31,80,30,49,31,65,31,35,31,197,31,197,30,191,31,238,31,138,31,138,30,255,31,55,31,55,30,55,29,147,31,127,31,45,31,252,31,252,30,201,31,208,31,218,31,91,31,122,31,39,31,253,31,133,31,133,30,44,31,200,31,147,31,115,31,87,31,20,31,18,31,120,31,72,31,72,30,181,31,223,31,57,31,72,31,72,30,163,31,113,31,199,31,174,31,51,31,187,31,246,31,20,31,57,31,57,30,19,31,77,31,77,30,77,29,77,28,51,31,108,31,106,31,5,31,5,30,67,31,161,31,161,30,171,31,66,31,66,30,90,31,216,31,158,31,208,31,49,31,252,31,136,31,136,30,5,31,102,31,102,30,102,29,217,31,90,31,176,31,196,31,132,31,253,31,236,31,149,31,219,31,219,30,219,29,248,31,165,31,180,31,49,31,132,31,3,31,2,31,24,31,25,31,245,31,5,31,253,31,81,31,110,31,254,31,249,31,113,31,38,31,135,31,164,31,132,31,50,31,98,31,85,31,33,31,84,31,192,31,54,31,54,30,120,31,243,31,243,30,87,31,50,31,50,30,221,31,221,30,77,31,155,31,197,31,53,31,240,31,70,31,196,31,236,31,253,31,237,31,237,30,209,31,209,30,74,31,145,31,89,31,34,31,223,31,78,31,41,31,41,30,19,31,100,31,211,31,254,31,24,31,8,31,94,31,125,31,125,30,84,31,93,31,14,31,14,30,95,31,71,31,8,31,189,31,183,31,199,31,117,31,203,31,189,31,101,31,101,30,136,31,94,31,67,31,67,30,109,31,189,31,4,31,15,31,186,31,203,31,121,31,18,31,18,30,18,29,86,31,86,30,86,29,243,31,243,30,76,31,139,31,241,31,168,31,154,31,214,31,135,31,135,30,153,31,153,30,28,31,28,30,74,31,122,31,107,31,140,31,146,31,108,31,207,31,244,31,51,31,148,31,148,30,131,31,30,31,57,31,251,31,183,31,144,31,242,31,213,31,147,31,111,31,93,31,21,31,222,31,101,31,46,31,46,30,247,31,188,31,165,31,246,31,153,31,129,31,138,31,49,31,6,31,171,31,214,31,76,31,116,31,159,31,181,31,94,31,159,31,66,31,69,31,69,30,56,31,211,31,211,30,102,31,102,30,171,31,153,31,249,31,208,31,104,31,104,30,198,31,198,30,198,29,213,31,213,30,179,31,179,30,33,31,88,31,183,31,199,31,199,30,121,31,125,31,203,31,19,31,156,31,110,31,5,31,190,31,196,31,196,30,228,31,167,31,254,31,150,31,139,31,54,31,72,31,96,31,96,30,176,31,173,31,173,30,109,31,145,31,145,30,145,29,155,31,29,31,165,31,200,31,200,30,200,29,36,31,138,31,112,31,44,31,112,31,210,31,233,31,50,31,238,31,189,31,172,31,147,31,147,30,147,29,96,31,141,31,57,31,57,30,204,31,230,31,87,31,87,30,242,31,189,31,25,31,181,31,28,31,239,31,139,31,208,31,141,31,141,30,56,31,172,31,228,31,238,31,238,30,177,31,203,31,203,30,29,31,209,31,122,31,46,31,53,31,130,31,34,31,128,31,246,31,246,30,164,31,231,31,27,31,88,31,81,31,87,31,59,31,241,31,25,31,25,30,25,29,22,31,10,31,10,30,191,31,25,31,6,31,131,31,242,31,41,31,82,31,82,30,212,31,97,31,236,31,185,31,154,31,82,31,82,30,176,31,92,31,76,31,122,31,180,31,201,31,236,31,24,31,152,31,42,31,21,31,194,31,194,31,173,31,179,31,236,31,236,30,123,31,6,31,243,31,64,31,10,31,10,30,91,31,80,31,109,31,109,30,163,31,33,31,225,31,244,31,210,31,140,31,79,31,79,30,157,31,34,31,105,31,41,31,251,31,180,31,180,30,114,31,157,31,254,31,120,31,120,30,120,31,97,31,8,31,8,30,90,31,47,31,28,31,60,31,82,31,152,31,18,31,212,31,1,31,120,31,189,31,135,31,167,31,146,31,146,30,93,31,249,31,151,31,84,31,96,31,96,30,215,31,215,30,46,31,235,31,72,31,72,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
