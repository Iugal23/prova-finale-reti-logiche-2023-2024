-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 847;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,187,0,139,0,178,0,156,0,0,0,48,0,35,0,32,0,57,0,156,0,103,0,166,0,248,0,255,0,250,0,199,0,1,0,87,0,54,0,185,0,15,0,0,0,21,0,126,0,221,0,199,0,170,0,198,0,166,0,214,0,0,0,163,0,234,0,64,0,2,0,217,0,117,0,0,0,0,0,146,0,233,0,0,0,36,0,0,0,216,0,172,0,212,0,177,0,110,0,98,0,230,0,134,0,8,0,223,0,48,0,97,0,35,0,134,0,81,0,156,0,58,0,0,0,197,0,135,0,86,0,76,0,4,0,178,0,182,0,147,0,0,0,250,0,191,0,0,0,243,0,182,0,164,0,139,0,185,0,53,0,214,0,235,0,106,0,2,0,0,0,223,0,198,0,124,0,184,0,181,0,4,0,7,0,5,0,0,0,48,0,0,0,0,0,0,0,79,0,77,0,217,0,63,0,39,0,11,0,40,0,10,0,96,0,99,0,0,0,0,0,141,0,128,0,12,0,232,0,241,0,217,0,0,0,245,0,0,0,222,0,0,0,103,0,198,0,228,0,0,0,86,0,180,0,0,0,0,0,123,0,246,0,0,0,0,0,249,0,220,0,15,0,159,0,74,0,69,0,34,0,176,0,0,0,53,0,0,0,255,0,128,0,101,0,0,0,185,0,82,0,207,0,221,0,218,0,249,0,243,0,228,0,11,0,41,0,117,0,124,0,0,0,0,0,161,0,200,0,122,0,81,0,55,0,15,0,91,0,32,0,15,0,0,0,148,0,163,0,108,0,192,0,78,0,0,0,164,0,46,0,190,0,113,0,117,0,0,0,0,0,95,0,0,0,199,0,40,0,0,0,174,0,82,0,37,0,7,0,0,0,0,0,164,0,102,0,37,0,43,0,113,0,0,0,87,0,0,0,25,0,181,0,238,0,0,0,0,0,17,0,183,0,72,0,230,0,103,0,44,0,253,0,115,0,0,0,245,0,178,0,0,0,54,0,212,0,0,0,213,0,19,0,37,0,157,0,132,0,106,0,93,0,191,0,164,0,112,0,255,0,214,0,107,0,0,0,31,0,37,0,229,0,173,0,35,0,21,0,0,0,219,0,188,0,43,0,0,0,66,0,61,0,227,0,58,0,96,0,0,0,2,0,0,0,0,0,107,0,0,0,0,0,140,0,192,0,86,0,26,0,224,0,36,0,58,0,208,0,88,0,41,0,74,0,145,0,59,0,75,0,224,0,127,0,140,0,111,0,59,0,122,0,73,0,26,0,0,0,0,0,0,0,43,0,34,0,80,0,255,0,0,0,0,0,0,0,156,0,69,0,178,0,188,0,4,0,94,0,125,0,142,0,243,0,0,0,132,0,53,0,0,0,243,0,250,0,216,0,132,0,11,0,5,0,50,0,218,0,0,0,182,0,54,0,180,0,164,0,167,0,0,0,190,0,51,0,0,0,0,0,253,0,120,0,0,0,47,0,0,0,7,0,161,0,52,0,0,0,253,0,0,0,0,0,167,0,172,0,134,0,246,0,112,0,0,0,18,0,128,0,0,0,156,0,196,0,221,0,242,0,45,0,188,0,185,0,206,0,4,0,171,0,0,0,227,0,212,0,193,0,114,0,143,0,0,0,201,0,199,0,0,0,7,0,76,0,102,0,75,0,131,0,123,0,0,0,199,0,251,0,220,0,196,0,232,0,164,0,101,0,1,0,22,0,239,0,48,0,0,0,125,0,250,0,0,0,41,0,220,0,0,0,46,0,98,0,128,0,246,0,60,0,32,0,61,0,151,0,0,0,98,0,153,0,0,0,94,0,185,0,184,0,31,0,240,0,15,0,205,0,249,0,231,0,62,0,0,0,226,0,170,0,0,0,0,0,156,0,236,0,92,0,228,0,0,0,34,0,64,0,0,0,0,0,213,0,0,0,168,0,0,0,204,0,7,0,9,0,156,0,163,0,65,0,178,0,255,0,0,0,152,0,0,0,245,0,152,0,240,0,36,0,137,0,0,0,0,0,89,0,219,0,180,0,180,0,0,0,3,0,10,0,219,0,0,0,180,0,237,0,0,0,120,0,84,0,155,0,0,0,24,0,0,0,3,0,24,0,31,0,26,0,164,0,138,0,84,0,120,0,5,0,181,0,30,0,67,0,243,0,18,0,78,0,245,0,51,0,0,0,0,0,0,0,214,0,207,0,237,0,216,0,116,0,119,0,223,0,229,0,0,0,62,0,251,0,192,0,167,0,209,0,181,0,0,0,214,0,153,0,190,0,14,0,38,0,152,0,63,0,122,0,221,0,75,0,4,0,203,0,222,0,35,0,217,0,36,0,131,0,69,0,186,0,152,0,70,0,0,0,122,0,188,0,226,0,0,0,29,0,0,0,162,0,230,0,0,0,229,0,31,0,139,0,216,0,209,0,191,0,70,0,137,0,91,0,22,0,144,0,164,0,235,0,0,0,97,0,125,0,87,0,129,0,0,0,250,0,126,0,47,0,45,0,68,0,0,0,0,0,113,0,53,0,113,0,0,0,216,0,220,0,82,0,0,0,0,0,174,0,48,0,132,0,10,0,143,0,0,0,55,0,33,0,251,0,121,0,134,0,41,0,144,0,227,0,12,0,191,0,249,0,121,0,170,0,199,0,1,0,43,0,111,0,152,0,0,0,20,0,237,0,176,0,11,0,105,0,0,0,225,0,0,0,80,0,244,0,67,0,150,0,233,0,226,0,0,0,220,0,69,0,0,0,68,0,175,0,0,0,20,0,12,0,0,0,122,0,160,0,244,0,64,0,180,0,179,0,0,0,230,0,99,0,3,0,0,0,253,0,176,0,129,0,230,0,0,0,25,0,33,0,229,0,136,0,147,0,0,0,10,0,189,0,87,0,0,0,54,0,3,0,132,0,141,0,0,0,108,0,6,0,0,0,127,0,168,0,0,0,193,0,106,0,101,0,0,0,99,0,180,0,22,0,151,0,152,0,166,0,179,0,33,0,0,0,210,0,0,0,0,0,155,0,177,0,32,0,2,0,122,0,243,0,0,0,232,0,0,0,0,0,31,0,251,0,180,0,19,0,215,0,128,0,157,0,117,0,80,0,153,0,0,0,112,0,241,0,169,0,22,0,0,0,0,0,164,0,0,0,177,0,209,0,0,0,208,0,29,0,0,0,95,0,102,0,0,0,66,0,134,0,0,0,175,0,11,0,0,0,238,0,4,0,0,0,0,0,100,0,167,0,84,0,219,0,168,0,24,0,153,0,132,0,168,0,0,0,207,0,40,0,80,0,86,0,136,0,7,0,225,0,114,0,9,0,67,0,11,0,134,0,238,0,172,0,247,0,147,0,106,0,30,0,0,0,216,0,198,0,186,0,97,0,205,0,0,0,31,0,252,0,232,0,0,0,193,0,136,0,0,0,48,0,52,0,243,0,32,0,56,0,11,0,148,0,62,0,115,0,9,0,232,0,114,0,0,0,53,0,8,0,80,0,200,0,162,0,114,0,90,0,40,0,56,0,69,0,163,0,14,0,0,0,211,0,0,0,86,0,244,0,73,0,39,0,213,0,78,0,0,0,6,0,131,0,0,0,0,0,144,0,0,0,0,0,0,0,166,0,123,0,61,0,99,0,0,0,182,0,66,0,233,0,190,0,0,0,7,0,222,0,196,0,0,0,22,0,146,0,203,0,153,0,0,0,70,0,23,0,245,0,7,0,106,0,191,0,108,0,253,0,38,0,21,0,0,0,150,0,45,0,201,0,193,0,0,0,161,0,78,0,0,0,214,0,74,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,187,31,139,31,178,31,156,31,156,30,48,31,35,31,32,31,57,31,156,31,103,31,166,31,248,31,255,31,250,31,199,31,1,31,87,31,54,31,185,31,15,31,15,30,21,31,126,31,221,31,199,31,170,31,198,31,166,31,214,31,214,30,163,31,234,31,64,31,2,31,217,31,117,31,117,30,117,29,146,31,233,31,233,30,36,31,36,30,216,31,172,31,212,31,177,31,110,31,98,31,230,31,134,31,8,31,223,31,48,31,97,31,35,31,134,31,81,31,156,31,58,31,58,30,197,31,135,31,86,31,76,31,4,31,178,31,182,31,147,31,147,30,250,31,191,31,191,30,243,31,182,31,164,31,139,31,185,31,53,31,214,31,235,31,106,31,2,31,2,30,223,31,198,31,124,31,184,31,181,31,4,31,7,31,5,31,5,30,48,31,48,30,48,29,48,28,79,31,77,31,217,31,63,31,39,31,11,31,40,31,10,31,96,31,99,31,99,30,99,29,141,31,128,31,12,31,232,31,241,31,217,31,217,30,245,31,245,30,222,31,222,30,103,31,198,31,228,31,228,30,86,31,180,31,180,30,180,29,123,31,246,31,246,30,246,29,249,31,220,31,15,31,159,31,74,31,69,31,34,31,176,31,176,30,53,31,53,30,255,31,128,31,101,31,101,30,185,31,82,31,207,31,221,31,218,31,249,31,243,31,228,31,11,31,41,31,117,31,124,31,124,30,124,29,161,31,200,31,122,31,81,31,55,31,15,31,91,31,32,31,15,31,15,30,148,31,163,31,108,31,192,31,78,31,78,30,164,31,46,31,190,31,113,31,117,31,117,30,117,29,95,31,95,30,199,31,40,31,40,30,174,31,82,31,37,31,7,31,7,30,7,29,164,31,102,31,37,31,43,31,113,31,113,30,87,31,87,30,25,31,181,31,238,31,238,30,238,29,17,31,183,31,72,31,230,31,103,31,44,31,253,31,115,31,115,30,245,31,178,31,178,30,54,31,212,31,212,30,213,31,19,31,37,31,157,31,132,31,106,31,93,31,191,31,164,31,112,31,255,31,214,31,107,31,107,30,31,31,37,31,229,31,173,31,35,31,21,31,21,30,219,31,188,31,43,31,43,30,66,31,61,31,227,31,58,31,96,31,96,30,2,31,2,30,2,29,107,31,107,30,107,29,140,31,192,31,86,31,26,31,224,31,36,31,58,31,208,31,88,31,41,31,74,31,145,31,59,31,75,31,224,31,127,31,140,31,111,31,59,31,122,31,73,31,26,31,26,30,26,29,26,28,43,31,34,31,80,31,255,31,255,30,255,29,255,28,156,31,69,31,178,31,188,31,4,31,94,31,125,31,142,31,243,31,243,30,132,31,53,31,53,30,243,31,250,31,216,31,132,31,11,31,5,31,50,31,218,31,218,30,182,31,54,31,180,31,164,31,167,31,167,30,190,31,51,31,51,30,51,29,253,31,120,31,120,30,47,31,47,30,7,31,161,31,52,31,52,30,253,31,253,30,253,29,167,31,172,31,134,31,246,31,112,31,112,30,18,31,128,31,128,30,156,31,196,31,221,31,242,31,45,31,188,31,185,31,206,31,4,31,171,31,171,30,227,31,212,31,193,31,114,31,143,31,143,30,201,31,199,31,199,30,7,31,76,31,102,31,75,31,131,31,123,31,123,30,199,31,251,31,220,31,196,31,232,31,164,31,101,31,1,31,22,31,239,31,48,31,48,30,125,31,250,31,250,30,41,31,220,31,220,30,46,31,98,31,128,31,246,31,60,31,32,31,61,31,151,31,151,30,98,31,153,31,153,30,94,31,185,31,184,31,31,31,240,31,15,31,205,31,249,31,231,31,62,31,62,30,226,31,170,31,170,30,170,29,156,31,236,31,92,31,228,31,228,30,34,31,64,31,64,30,64,29,213,31,213,30,168,31,168,30,204,31,7,31,9,31,156,31,163,31,65,31,178,31,255,31,255,30,152,31,152,30,245,31,152,31,240,31,36,31,137,31,137,30,137,29,89,31,219,31,180,31,180,31,180,30,3,31,10,31,219,31,219,30,180,31,237,31,237,30,120,31,84,31,155,31,155,30,24,31,24,30,3,31,24,31,31,31,26,31,164,31,138,31,84,31,120,31,5,31,181,31,30,31,67,31,243,31,18,31,78,31,245,31,51,31,51,30,51,29,51,28,214,31,207,31,237,31,216,31,116,31,119,31,223,31,229,31,229,30,62,31,251,31,192,31,167,31,209,31,181,31,181,30,214,31,153,31,190,31,14,31,38,31,152,31,63,31,122,31,221,31,75,31,4,31,203,31,222,31,35,31,217,31,36,31,131,31,69,31,186,31,152,31,70,31,70,30,122,31,188,31,226,31,226,30,29,31,29,30,162,31,230,31,230,30,229,31,31,31,139,31,216,31,209,31,191,31,70,31,137,31,91,31,22,31,144,31,164,31,235,31,235,30,97,31,125,31,87,31,129,31,129,30,250,31,126,31,47,31,45,31,68,31,68,30,68,29,113,31,53,31,113,31,113,30,216,31,220,31,82,31,82,30,82,29,174,31,48,31,132,31,10,31,143,31,143,30,55,31,33,31,251,31,121,31,134,31,41,31,144,31,227,31,12,31,191,31,249,31,121,31,170,31,199,31,1,31,43,31,111,31,152,31,152,30,20,31,237,31,176,31,11,31,105,31,105,30,225,31,225,30,80,31,244,31,67,31,150,31,233,31,226,31,226,30,220,31,69,31,69,30,68,31,175,31,175,30,20,31,12,31,12,30,122,31,160,31,244,31,64,31,180,31,179,31,179,30,230,31,99,31,3,31,3,30,253,31,176,31,129,31,230,31,230,30,25,31,33,31,229,31,136,31,147,31,147,30,10,31,189,31,87,31,87,30,54,31,3,31,132,31,141,31,141,30,108,31,6,31,6,30,127,31,168,31,168,30,193,31,106,31,101,31,101,30,99,31,180,31,22,31,151,31,152,31,166,31,179,31,33,31,33,30,210,31,210,30,210,29,155,31,177,31,32,31,2,31,122,31,243,31,243,30,232,31,232,30,232,29,31,31,251,31,180,31,19,31,215,31,128,31,157,31,117,31,80,31,153,31,153,30,112,31,241,31,169,31,22,31,22,30,22,29,164,31,164,30,177,31,209,31,209,30,208,31,29,31,29,30,95,31,102,31,102,30,66,31,134,31,134,30,175,31,11,31,11,30,238,31,4,31,4,30,4,29,100,31,167,31,84,31,219,31,168,31,24,31,153,31,132,31,168,31,168,30,207,31,40,31,80,31,86,31,136,31,7,31,225,31,114,31,9,31,67,31,11,31,134,31,238,31,172,31,247,31,147,31,106,31,30,31,30,30,216,31,198,31,186,31,97,31,205,31,205,30,31,31,252,31,232,31,232,30,193,31,136,31,136,30,48,31,52,31,243,31,32,31,56,31,11,31,148,31,62,31,115,31,9,31,232,31,114,31,114,30,53,31,8,31,80,31,200,31,162,31,114,31,90,31,40,31,56,31,69,31,163,31,14,31,14,30,211,31,211,30,86,31,244,31,73,31,39,31,213,31,78,31,78,30,6,31,131,31,131,30,131,29,144,31,144,30,144,29,144,28,166,31,123,31,61,31,99,31,99,30,182,31,66,31,233,31,190,31,190,30,7,31,222,31,196,31,196,30,22,31,146,31,203,31,153,31,153,30,70,31,23,31,245,31,7,31,106,31,191,31,108,31,253,31,38,31,21,31,21,30,150,31,45,31,201,31,193,31,193,30,161,31,78,31,78,30,214,31,74,31,74,30,74,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
