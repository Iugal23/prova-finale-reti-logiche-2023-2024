-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_82 is
end project_tb_82;

architecture project_tb_arch_82 of project_tb_82 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 655;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,95,0,224,0,94,0,47,0,11,0,0,0,166,0,217,0,108,0,178,0,247,0,23,0,218,0,199,0,0,0,0,0,240,0,168,0,51,0,197,0,51,0,64,0,0,0,30,0,104,0,148,0,156,0,0,0,14,0,111,0,127,0,0,0,85,0,253,0,91,0,0,0,121,0,186,0,52,0,44,0,28,0,105,0,37,0,217,0,87,0,5,0,25,0,112,0,57,0,0,0,0,0,156,0,141,0,35,0,56,0,0,0,218,0,0,0,19,0,37,0,0,0,201,0,0,0,212,0,191,0,161,0,187,0,220,0,123,0,176,0,0,0,227,0,0,0,152,0,207,0,133,0,219,0,0,0,20,0,167,0,0,0,152,0,199,0,26,0,0,0,134,0,0,0,38,0,70,0,176,0,106,0,88,0,62,0,0,0,0,0,182,0,0,0,166,0,78,0,10,0,0,0,0,0,214,0,0,0,98,0,195,0,138,0,232,0,23,0,0,0,138,0,6,0,214,0,210,0,119,0,165,0,55,0,53,0,179,0,32,0,151,0,54,0,40,0,124,0,0,0,173,0,0,0,0,0,230,0,75,0,205,0,225,0,210,0,83,0,149,0,66,0,0,0,195,0,223,0,213,0,0,0,53,0,0,0,68,0,150,0,0,0,166,0,253,0,0,0,0,0,251,0,165,0,93,0,0,0,61,0,115,0,67,0,179,0,132,0,0,0,61,0,29,0,59,0,0,0,0,0,0,0,0,0,241,0,60,0,171,0,0,0,115,0,177,0,140,0,250,0,132,0,6,0,0,0,250,0,0,0,127,0,0,0,206,0,82,0,253,0,197,0,0,0,60,0,130,0,23,0,245,0,27,0,239,0,173,0,7,0,232,0,0,0,227,0,187,0,181,0,14,0,231,0,108,0,0,0,0,0,62,0,247,0,41,0,124,0,143,0,0,0,0,0,91,0,0,0,0,0,0,0,166,0,112,0,153,0,0,0,216,0,47,0,144,0,225,0,248,0,0,0,232,0,85,0,47,0,74,0,151,0,236,0,94,0,113,0,0,0,92,0,7,0,0,0,148,0,0,0,50,0,195,0,31,0,0,0,223,0,0,0,82,0,111,0,194,0,0,0,108,0,108,0,0,0,33,0,193,0,224,0,14,0,127,0,181,0,237,0,248,0,0,0,100,0,132,0,0,0,0,0,114,0,0,0,170,0,0,0,120,0,231,0,0,0,80,0,29,0,17,0,178,0,99,0,154,0,0,0,0,0,0,0,46,0,61,0,75,0,1,0,8,0,235,0,176,0,64,0,183,0,0,0,73,0,196,0,78,0,170,0,195,0,214,0,224,0,27,0,13,0,48,0,248,0,164,0,0,0,56,0,35,0,183,0,194,0,129,0,234,0,0,0,193,0,0,0,144,0,33,0,64,0,241,0,122,0,0,0,0,0,182,0,220,0,170,0,95,0,192,0,182,0,105,0,102,0,18,0,216,0,90,0,0,0,234,0,92,0,255,0,206,0,165,0,141,0,183,0,43,0,119,0,41,0,12,0,198,0,0,0,164,0,215,0,233,0,181,0,187,0,152,0,75,0,88,0,137,0,144,0,179,0,171,0,0,0,210,0,0,0,161,0,153,0,247,0,5,0,105,0,180,0,85,0,0,0,138,0,104,0,0,0,0,0,0,0,168,0,0,0,105,0,0,0,42,0,73,0,0,0,0,0,69,0,0,0,216,0,176,0,5,0,0,0,0,0,122,0,0,0,0,0,120,0,15,0,84,0,114,0,168,0,0,0,48,0,169,0,45,0,106,0,219,0,0,0,43,0,0,0,85,0,163,0,20,0,0,0,37,0,94,0,31,0,151,0,0,0,187,0,0,0,29,0,0,0,0,0,0,0,221,0,0,0,16,0,156,0,226,0,237,0,165,0,0,0,22,0,59,0,214,0,0,0,230,0,51,0,81,0,198,0,162,0,90,0,31,0,124,0,0,0,210,0,191,0,204,0,125,0,39,0,0,0,215,0,248,0,214,0,229,0,0,0,5,0,206,0,0,0,0,0,14,0,61,0,92,0,97,0,37,0,0,0,30,0,128,0,250,0,174,0,0,0,0,0,123,0,3,0,146,0,164,0,0,0,187,0,180,0,82,0,201,0,79,0,67,0,254,0,251,0,227,0,43,0,227,0,138,0,12,0,75,0,0,0,0,0,0,0,33,0,26,0,0,0,168,0,254,0,194,0,57,0,97,0,120,0,81,0,243,0,204,0,87,0,93,0,5,0,78,0,89,0,0,0,140,0,0,0,70,0,0,0,0,0,145,0,75,0,94,0,230,0,10,0,26,0,0,0,183,0,193,0,221,0,214,0,32,0,158,0,39,0,131,0,48,0,224,0,232,0,61,0,239,0,147,0,52,0,110,0,10,0,0,0,50,0,20,0,76,0,242,0,114,0,207,0,250,0,15,0,188,0,186,0,241,0,80,0,107,0,33,0,46,0,180,0,99,0,0,0,0,0,6,0,0,0,0,0,187,0,0,0,240,0,90,0,35,0,188,0,226,0,255,0,122,0,100,0,131,0,137,0,196,0,0,0,145,0,63,0,197,0,89,0,0,0,0,0,233,0,153,0,228,0,38,0,142,0,0,0,189,0,33,0,123,0,58,0,126,0,198,0,0,0,149,0,4,0,38,0,244,0,0,0,142,0,51,0,172,0,111,0,0,0,126,0,154,0,124,0,0,0,0,0,52,0,201,0,0,0,104,0,157,0,76,0,14,0,0,0,61,0,95,0,49,0,146,0,39,0,125,0,169,0,31,0,0,0,237,0,99,0,128,0,169,0,251,0,0,0,0,0,214,0,71,0,0,0,0,0,34,0,0,0,195,0,166,0,193,0,84,0,1,0,10,0,223,0,144,0,55,0,115,0,0,0,12,0,28,0,132,0);
signal scenario_full  : scenario_type := (0,0,0,0,95,31,224,31,94,31,47,31,11,31,11,30,166,31,217,31,108,31,178,31,247,31,23,31,218,31,199,31,199,30,199,29,240,31,168,31,51,31,197,31,51,31,64,31,64,30,30,31,104,31,148,31,156,31,156,30,14,31,111,31,127,31,127,30,85,31,253,31,91,31,91,30,121,31,186,31,52,31,44,31,28,31,105,31,37,31,217,31,87,31,5,31,25,31,112,31,57,31,57,30,57,29,156,31,141,31,35,31,56,31,56,30,218,31,218,30,19,31,37,31,37,30,201,31,201,30,212,31,191,31,161,31,187,31,220,31,123,31,176,31,176,30,227,31,227,30,152,31,207,31,133,31,219,31,219,30,20,31,167,31,167,30,152,31,199,31,26,31,26,30,134,31,134,30,38,31,70,31,176,31,106,31,88,31,62,31,62,30,62,29,182,31,182,30,166,31,78,31,10,31,10,30,10,29,214,31,214,30,98,31,195,31,138,31,232,31,23,31,23,30,138,31,6,31,214,31,210,31,119,31,165,31,55,31,53,31,179,31,32,31,151,31,54,31,40,31,124,31,124,30,173,31,173,30,173,29,230,31,75,31,205,31,225,31,210,31,83,31,149,31,66,31,66,30,195,31,223,31,213,31,213,30,53,31,53,30,68,31,150,31,150,30,166,31,253,31,253,30,253,29,251,31,165,31,93,31,93,30,61,31,115,31,67,31,179,31,132,31,132,30,61,31,29,31,59,31,59,30,59,29,59,28,59,27,241,31,60,31,171,31,171,30,115,31,177,31,140,31,250,31,132,31,6,31,6,30,250,31,250,30,127,31,127,30,206,31,82,31,253,31,197,31,197,30,60,31,130,31,23,31,245,31,27,31,239,31,173,31,7,31,232,31,232,30,227,31,187,31,181,31,14,31,231,31,108,31,108,30,108,29,62,31,247,31,41,31,124,31,143,31,143,30,143,29,91,31,91,30,91,29,91,28,166,31,112,31,153,31,153,30,216,31,47,31,144,31,225,31,248,31,248,30,232,31,85,31,47,31,74,31,151,31,236,31,94,31,113,31,113,30,92,31,7,31,7,30,148,31,148,30,50,31,195,31,31,31,31,30,223,31,223,30,82,31,111,31,194,31,194,30,108,31,108,31,108,30,33,31,193,31,224,31,14,31,127,31,181,31,237,31,248,31,248,30,100,31,132,31,132,30,132,29,114,31,114,30,170,31,170,30,120,31,231,31,231,30,80,31,29,31,17,31,178,31,99,31,154,31,154,30,154,29,154,28,46,31,61,31,75,31,1,31,8,31,235,31,176,31,64,31,183,31,183,30,73,31,196,31,78,31,170,31,195,31,214,31,224,31,27,31,13,31,48,31,248,31,164,31,164,30,56,31,35,31,183,31,194,31,129,31,234,31,234,30,193,31,193,30,144,31,33,31,64,31,241,31,122,31,122,30,122,29,182,31,220,31,170,31,95,31,192,31,182,31,105,31,102,31,18,31,216,31,90,31,90,30,234,31,92,31,255,31,206,31,165,31,141,31,183,31,43,31,119,31,41,31,12,31,198,31,198,30,164,31,215,31,233,31,181,31,187,31,152,31,75,31,88,31,137,31,144,31,179,31,171,31,171,30,210,31,210,30,161,31,153,31,247,31,5,31,105,31,180,31,85,31,85,30,138,31,104,31,104,30,104,29,104,28,168,31,168,30,105,31,105,30,42,31,73,31,73,30,73,29,69,31,69,30,216,31,176,31,5,31,5,30,5,29,122,31,122,30,122,29,120,31,15,31,84,31,114,31,168,31,168,30,48,31,169,31,45,31,106,31,219,31,219,30,43,31,43,30,85,31,163,31,20,31,20,30,37,31,94,31,31,31,151,31,151,30,187,31,187,30,29,31,29,30,29,29,29,28,221,31,221,30,16,31,156,31,226,31,237,31,165,31,165,30,22,31,59,31,214,31,214,30,230,31,51,31,81,31,198,31,162,31,90,31,31,31,124,31,124,30,210,31,191,31,204,31,125,31,39,31,39,30,215,31,248,31,214,31,229,31,229,30,5,31,206,31,206,30,206,29,14,31,61,31,92,31,97,31,37,31,37,30,30,31,128,31,250,31,174,31,174,30,174,29,123,31,3,31,146,31,164,31,164,30,187,31,180,31,82,31,201,31,79,31,67,31,254,31,251,31,227,31,43,31,227,31,138,31,12,31,75,31,75,30,75,29,75,28,33,31,26,31,26,30,168,31,254,31,194,31,57,31,97,31,120,31,81,31,243,31,204,31,87,31,93,31,5,31,78,31,89,31,89,30,140,31,140,30,70,31,70,30,70,29,145,31,75,31,94,31,230,31,10,31,26,31,26,30,183,31,193,31,221,31,214,31,32,31,158,31,39,31,131,31,48,31,224,31,232,31,61,31,239,31,147,31,52,31,110,31,10,31,10,30,50,31,20,31,76,31,242,31,114,31,207,31,250,31,15,31,188,31,186,31,241,31,80,31,107,31,33,31,46,31,180,31,99,31,99,30,99,29,6,31,6,30,6,29,187,31,187,30,240,31,90,31,35,31,188,31,226,31,255,31,122,31,100,31,131,31,137,31,196,31,196,30,145,31,63,31,197,31,89,31,89,30,89,29,233,31,153,31,228,31,38,31,142,31,142,30,189,31,33,31,123,31,58,31,126,31,198,31,198,30,149,31,4,31,38,31,244,31,244,30,142,31,51,31,172,31,111,31,111,30,126,31,154,31,124,31,124,30,124,29,52,31,201,31,201,30,104,31,157,31,76,31,14,31,14,30,61,31,95,31,49,31,146,31,39,31,125,31,169,31,31,31,31,30,237,31,99,31,128,31,169,31,251,31,251,30,251,29,214,31,71,31,71,30,71,29,34,31,34,30,195,31,166,31,193,31,84,31,1,31,10,31,223,31,144,31,55,31,115,31,115,30,12,31,28,31,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
