-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 663;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,14,0,0,0,0,0,24,0,231,0,212,0,0,0,0,0,93,0,100,0,216,0,0,0,0,0,0,0,0,0,240,0,175,0,75,0,190,0,198,0,208,0,155,0,7,0,224,0,33,0,223,0,0,0,173,0,127,0,0,0,106,0,166,0,159,0,54,0,88,0,254,0,0,0,0,0,6,0,45,0,212,0,0,0,219,0,214,0,0,0,243,0,138,0,77,0,99,0,195,0,138,0,248,0,41,0,45,0,0,0,196,0,46,0,115,0,111,0,11,0,0,0,43,0,246,0,236,0,40,0,74,0,0,0,244,0,230,0,223,0,180,0,0,0,171,0,170,0,67,0,102,0,3,0,71,0,35,0,124,0,245,0,0,0,0,0,198,0,76,0,202,0,204,0,0,0,117,0,73,0,0,0,150,0,159,0,0,0,117,0,0,0,79,0,52,0,239,0,239,0,112,0,160,0,70,0,228,0,113,0,153,0,36,0,194,0,33,0,120,0,79,0,241,0,247,0,172,0,134,0,55,0,178,0,14,0,175,0,0,0,243,0,110,0,164,0,248,0,8,0,194,0,0,0,0,0,32,0,251,0,162,0,0,0,78,0,245,0,13,0,27,0,208,0,0,0,41,0,0,0,48,0,169,0,152,0,180,0,79,0,0,0,0,0,144,0,101,0,60,0,227,0,72,0,70,0,0,0,208,0,0,0,111,0,189,0,143,0,167,0,0,0,155,0,0,0,50,0,0,0,207,0,247,0,220,0,156,0,160,0,207,0,100,0,254,0,94,0,180,0,185,0,208,0,139,0,0,0,0,0,80,0,18,0,54,0,236,0,0,0,46,0,44,0,208,0,155,0,109,0,226,0,97,0,218,0,0,0,228,0,179,0,1,0,253,0,0,0,0,0,182,0,159,0,217,0,243,0,0,0,147,0,181,0,234,0,53,0,111,0,0,0,158,0,225,0,0,0,78,0,205,0,64,0,0,0,144,0,252,0,200,0,131,0,135,0,177,0,205,0,102,0,195,0,177,0,219,0,227,0,53,0,147,0,42,0,56,0,123,0,220,0,84,0,216,0,211,0,0,0,130,0,60,0,0,0,231,0,40,0,0,0,65,0,56,0,233,0,205,0,0,0,65,0,168,0,131,0,181,0,32,0,52,0,47,0,58,0,224,0,18,0,0,0,0,0,237,0,0,0,83,0,93,0,80,0,234,0,118,0,124,0,61,0,0,0,91,0,93,0,0,0,174,0,195,0,105,0,0,0,53,0,167,0,122,0,20,0,239,0,149,0,202,0,3,0,69,0,233,0,46,0,176,0,91,0,40,0,81,0,0,0,27,0,179,0,160,0,251,0,0,0,151,0,101,0,165,0,134,0,0,0,64,0,252,0,96,0,109,0,206,0,53,0,199,0,117,0,202,0,201,0,163,0,31,0,63,0,22,0,111,0,195,0,206,0,125,0,239,0,34,0,153,0,0,0,168,0,107,0,96,0,24,0,165,0,129,0,81,0,0,0,6,0,156,0,103,0,0,0,137,0,88,0,229,0,0,0,0,0,0,0,69,0,143,0,70,0,42,0,0,0,133,0,212,0,112,0,222,0,0,0,228,0,0,0,37,0,0,0,71,0,69,0,187,0,8,0,101,0,0,0,0,0,18,0,0,0,48,0,86,0,225,0,129,0,124,0,98,0,79,0,26,0,1,0,178,0,0,0,70,0,104,0,161,0,0,0,230,0,192,0,220,0,0,0,236,0,0,0,116,0,0,0,94,0,9,0,202,0,215,0,10,0,116,0,0,0,44,0,0,0,129,0,117,0,85,0,219,0,0,0,121,0,110,0,130,0,0,0,0,0,164,0,211,0,160,0,0,0,0,0,0,0,97,0,109,0,34,0,163,0,43,0,193,0,0,0,0,0,111,0,0,0,187,0,17,0,253,0,54,0,25,0,74,0,146,0,0,0,44,0,138,0,25,0,214,0,146,0,40,0,0,0,193,0,65,0,68,0,0,0,57,0,78,0,193,0,0,0,249,0,64,0,46,0,63,0,0,0,243,0,121,0,224,0,125,0,150,0,26,0,188,0,27,0,0,0,213,0,186,0,147,0,0,0,0,0,0,0,176,0,154,0,0,0,1,0,119,0,0,0,197,0,88,0,210,0,40,0,8,0,0,0,0,0,0,0,213,0,226,0,91,0,117,0,86,0,212,0,170,0,229,0,219,0,158,0,0,0,0,0,48,0,79,0,22,0,36,0,122,0,33,0,39,0,184,0,237,0,57,0,110,0,0,0,28,0,118,0,0,0,103,0,227,0,130,0,4,0,0,0,75,0,78,0,12,0,0,0,223,0,147,0,148,0,207,0,0,0,226,0,241,0,245,0,14,0,181,0,55,0,209,0,126,0,64,0,29,0,0,0,0,0,170,0,132,0,158,0,94,0,0,0,9,0,0,0,242,0,100,0,167,0,234,0,70,0,231,0,0,0,213,0,0,0,24,0,0,0,27,0,53,0,0,0,162,0,92,0,14,0,174,0,72,0,216,0,139,0,0,0,222,0,0,0,238,0,162,0,71,0,142,0,12,0,206,0,0,0,223,0,23,0,144,0,105,0,199,0,89,0,0,0,205,0,55,0,104,0,187,0,191,0,80,0,139,0,229,0,190,0,18,0,163,0,0,0,0,0,70,0,167,0,39,0,60,0,177,0,232,0,171,0,119,0,212,0,74,0,0,0,177,0,0,0,176,0,0,0,34,0,84,0,0,0,106,0,138,0,73,0,166,0,177,0,172,0,75,0,1,0,102,0,0,0,0,0,131,0,91,0,83,0,247,0,12,0,113,0,0,0,251,0,0,0,113,0,150,0,53,0,77,0,215,0,72,0,40,0,43,0,152,0,126,0,63,0,49,0,221,0,55,0,0,0,81,0,60,0,150,0,224,0,78,0,199,0,0,0,132,0,49,0,99,0,64,0,138,0,68,0,164,0);
signal scenario_full  : scenario_type := (0,0,14,31,14,30,14,29,24,31,231,31,212,31,212,30,212,29,93,31,100,31,216,31,216,30,216,29,216,28,216,27,240,31,175,31,75,31,190,31,198,31,208,31,155,31,7,31,224,31,33,31,223,31,223,30,173,31,127,31,127,30,106,31,166,31,159,31,54,31,88,31,254,31,254,30,254,29,6,31,45,31,212,31,212,30,219,31,214,31,214,30,243,31,138,31,77,31,99,31,195,31,138,31,248,31,41,31,45,31,45,30,196,31,46,31,115,31,111,31,11,31,11,30,43,31,246,31,236,31,40,31,74,31,74,30,244,31,230,31,223,31,180,31,180,30,171,31,170,31,67,31,102,31,3,31,71,31,35,31,124,31,245,31,245,30,245,29,198,31,76,31,202,31,204,31,204,30,117,31,73,31,73,30,150,31,159,31,159,30,117,31,117,30,79,31,52,31,239,31,239,31,112,31,160,31,70,31,228,31,113,31,153,31,36,31,194,31,33,31,120,31,79,31,241,31,247,31,172,31,134,31,55,31,178,31,14,31,175,31,175,30,243,31,110,31,164,31,248,31,8,31,194,31,194,30,194,29,32,31,251,31,162,31,162,30,78,31,245,31,13,31,27,31,208,31,208,30,41,31,41,30,48,31,169,31,152,31,180,31,79,31,79,30,79,29,144,31,101,31,60,31,227,31,72,31,70,31,70,30,208,31,208,30,111,31,189,31,143,31,167,31,167,30,155,31,155,30,50,31,50,30,207,31,247,31,220,31,156,31,160,31,207,31,100,31,254,31,94,31,180,31,185,31,208,31,139,31,139,30,139,29,80,31,18,31,54,31,236,31,236,30,46,31,44,31,208,31,155,31,109,31,226,31,97,31,218,31,218,30,228,31,179,31,1,31,253,31,253,30,253,29,182,31,159,31,217,31,243,31,243,30,147,31,181,31,234,31,53,31,111,31,111,30,158,31,225,31,225,30,78,31,205,31,64,31,64,30,144,31,252,31,200,31,131,31,135,31,177,31,205,31,102,31,195,31,177,31,219,31,227,31,53,31,147,31,42,31,56,31,123,31,220,31,84,31,216,31,211,31,211,30,130,31,60,31,60,30,231,31,40,31,40,30,65,31,56,31,233,31,205,31,205,30,65,31,168,31,131,31,181,31,32,31,52,31,47,31,58,31,224,31,18,31,18,30,18,29,237,31,237,30,83,31,93,31,80,31,234,31,118,31,124,31,61,31,61,30,91,31,93,31,93,30,174,31,195,31,105,31,105,30,53,31,167,31,122,31,20,31,239,31,149,31,202,31,3,31,69,31,233,31,46,31,176,31,91,31,40,31,81,31,81,30,27,31,179,31,160,31,251,31,251,30,151,31,101,31,165,31,134,31,134,30,64,31,252,31,96,31,109,31,206,31,53,31,199,31,117,31,202,31,201,31,163,31,31,31,63,31,22,31,111,31,195,31,206,31,125,31,239,31,34,31,153,31,153,30,168,31,107,31,96,31,24,31,165,31,129,31,81,31,81,30,6,31,156,31,103,31,103,30,137,31,88,31,229,31,229,30,229,29,229,28,69,31,143,31,70,31,42,31,42,30,133,31,212,31,112,31,222,31,222,30,228,31,228,30,37,31,37,30,71,31,69,31,187,31,8,31,101,31,101,30,101,29,18,31,18,30,48,31,86,31,225,31,129,31,124,31,98,31,79,31,26,31,1,31,178,31,178,30,70,31,104,31,161,31,161,30,230,31,192,31,220,31,220,30,236,31,236,30,116,31,116,30,94,31,9,31,202,31,215,31,10,31,116,31,116,30,44,31,44,30,129,31,117,31,85,31,219,31,219,30,121,31,110,31,130,31,130,30,130,29,164,31,211,31,160,31,160,30,160,29,160,28,97,31,109,31,34,31,163,31,43,31,193,31,193,30,193,29,111,31,111,30,187,31,17,31,253,31,54,31,25,31,74,31,146,31,146,30,44,31,138,31,25,31,214,31,146,31,40,31,40,30,193,31,65,31,68,31,68,30,57,31,78,31,193,31,193,30,249,31,64,31,46,31,63,31,63,30,243,31,121,31,224,31,125,31,150,31,26,31,188,31,27,31,27,30,213,31,186,31,147,31,147,30,147,29,147,28,176,31,154,31,154,30,1,31,119,31,119,30,197,31,88,31,210,31,40,31,8,31,8,30,8,29,8,28,213,31,226,31,91,31,117,31,86,31,212,31,170,31,229,31,219,31,158,31,158,30,158,29,48,31,79,31,22,31,36,31,122,31,33,31,39,31,184,31,237,31,57,31,110,31,110,30,28,31,118,31,118,30,103,31,227,31,130,31,4,31,4,30,75,31,78,31,12,31,12,30,223,31,147,31,148,31,207,31,207,30,226,31,241,31,245,31,14,31,181,31,55,31,209,31,126,31,64,31,29,31,29,30,29,29,170,31,132,31,158,31,94,31,94,30,9,31,9,30,242,31,100,31,167,31,234,31,70,31,231,31,231,30,213,31,213,30,24,31,24,30,27,31,53,31,53,30,162,31,92,31,14,31,174,31,72,31,216,31,139,31,139,30,222,31,222,30,238,31,162,31,71,31,142,31,12,31,206,31,206,30,223,31,23,31,144,31,105,31,199,31,89,31,89,30,205,31,55,31,104,31,187,31,191,31,80,31,139,31,229,31,190,31,18,31,163,31,163,30,163,29,70,31,167,31,39,31,60,31,177,31,232,31,171,31,119,31,212,31,74,31,74,30,177,31,177,30,176,31,176,30,34,31,84,31,84,30,106,31,138,31,73,31,166,31,177,31,172,31,75,31,1,31,102,31,102,30,102,29,131,31,91,31,83,31,247,31,12,31,113,31,113,30,251,31,251,30,113,31,150,31,53,31,77,31,215,31,72,31,40,31,43,31,152,31,126,31,63,31,49,31,221,31,55,31,55,30,81,31,60,31,150,31,224,31,78,31,199,31,199,30,132,31,49,31,99,31,64,31,138,31,68,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
