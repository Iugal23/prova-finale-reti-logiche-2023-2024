-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_981 is
end project_tb_981;

architecture project_tb_arch_981 of project_tb_981 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 743;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (18,0,158,0,3,0,73,0,61,0,63,0,10,0,172,0,72,0,250,0,31,0,4,0,0,0,157,0,19,0,207,0,8,0,0,0,224,0,0,0,45,0,168,0,18,0,87,0,51,0,6,0,172,0,144,0,57,0,26,0,25,0,72,0,73,0,0,0,190,0,145,0,0,0,131,0,147,0,13,0,57,0,11,0,141,0,157,0,0,0,105,0,95,0,17,0,0,0,153,0,188,0,123,0,61,0,144,0,13,0,47,0,84,0,0,0,187,0,171,0,0,0,21,0,20,0,234,0,252,0,0,0,103,0,231,0,77,0,21,0,0,0,221,0,0,0,0,0,0,0,199,0,0,0,84,0,246,0,142,0,78,0,43,0,107,0,127,0,233,0,240,0,137,0,6,0,206,0,79,0,0,0,138,0,246,0,101,0,31,0,152,0,115,0,84,0,183,0,85,0,101,0,122,0,0,0,0,0,5,0,68,0,92,0,74,0,0,0,122,0,90,0,27,0,0,0,112,0,90,0,151,0,134,0,114,0,32,0,211,0,0,0,226,0,64,0,0,0,145,0,54,0,223,0,190,0,209,0,148,0,124,0,0,0,99,0,52,0,220,0,0,0,193,0,30,0,234,0,197,0,0,0,0,0,129,0,0,0,7,0,249,0,145,0,211,0,57,0,81,0,0,0,0,0,236,0,110,0,0,0,0,0,0,0,213,0,118,0,41,0,184,0,161,0,43,0,0,0,130,0,62,0,0,0,54,0,20,0,51,0,162,0,60,0,176,0,188,0,120,0,200,0,34,0,0,0,193,0,186,0,172,0,158,0,44,0,81,0,217,0,105,0,191,0,0,0,0,0,164,0,104,0,56,0,0,0,241,0,77,0,0,0,0,0,248,0,203,0,169,0,67,0,78,0,0,0,147,0,159,0,112,0,191,0,135,0,61,0,166,0,220,0,210,0,196,0,43,0,235,0,3,0,162,0,212,0,211,0,0,0,41,0,82,0,58,0,246,0,49,0,17,0,2,0,246,0,74,0,0,0,0,0,0,0,179,0,0,0,0,0,85,0,249,0,10,0,193,0,51,0,42,0,191,0,43,0,46,0,0,0,240,0,201,0,70,0,108,0,131,0,100,0,0,0,49,0,0,0,0,0,243,0,36,0,75,0,200,0,2,0,17,0,111,0,171,0,24,0,0,0,228,0,162,0,76,0,55,0,125,0,0,0,23,0,104,0,207,0,51,0,146,0,227,0,0,0,0,0,79,0,53,0,0,0,64,0,150,0,35,0,93,0,120,0,45,0,220,0,64,0,172,0,103,0,0,0,81,0,137,0,116,0,64,0,92,0,122,0,48,0,124,0,252,0,255,0,57,0,117,0,232,0,0,0,65,0,0,0,86,0,185,0,41,0,168,0,139,0,101,0,1,0,147,0,96,0,0,0,111,0,81,0,155,0,0,0,237,0,187,0,214,0,0,0,111,0,0,0,2,0,159,0,240,0,154,0,108,0,129,0,64,0,212,0,0,0,0,0,164,0,43,0,0,0,0,0,150,0,16,0,92,0,246,0,156,0,66,0,86,0,117,0,0,0,111,0,94,0,0,0,206,0,73,0,0,0,30,0,121,0,110,0,151,0,80,0,26,0,105,0,199,0,129,0,0,0,0,0,134,0,0,0,129,0,90,0,0,0,0,0,243,0,0,0,193,0,182,0,220,0,127,0,52,0,163,0,224,0,0,0,205,0,83,0,31,0,148,0,18,0,41,0,0,0,148,0,0,0,116,0,229,0,23,0,188,0,34,0,2,0,103,0,1,0,64,0,191,0,0,0,113,0,3,0,0,0,45,0,47,0,0,0,204,0,131,0,110,0,0,0,0,0,205,0,74,0,84,0,0,0,0,0,47,0,63,0,169,0,191,0,24,0,118,0,34,0,190,0,153,0,0,0,132,0,159,0,0,0,222,0,0,0,5,0,189,0,238,0,0,0,69,0,156,0,64,0,0,0,209,0,170,0,54,0,61,0,238,0,181,0,23,0,123,0,245,0,0,0,69,0,10,0,85,0,159,0,0,0,211,0,204,0,148,0,223,0,0,0,140,0,153,0,200,0,0,0,75,0,219,0,61,0,149,0,0,0,93,0,112,0,96,0,48,0,49,0,182,0,0,0,3,0,205,0,105,0,0,0,230,0,140,0,215,0,0,0,187,0,99,0,68,0,32,0,242,0,14,0,158,0,5,0,228,0,23,0,0,0,135,0,0,0,0,0,238,0,104,0,0,0,12,0,187,0,0,0,83,0,71,0,4,0,166,0,0,0,170,0,0,0,89,0,143,0,225,0,55,0,81,0,27,0,9,0,97,0,224,0,118,0,0,0,48,0,197,0,73,0,0,0,103,0,0,0,0,0,173,0,55,0,166,0,132,0,8,0,186,0,0,0,0,0,126,0,0,0,55,0,16,0,197,0,213,0,53,0,0,0,218,0,202,0,165,0,24,0,115,0,49,0,0,0,214,0,29,0,61,0,150,0,198,0,53,0,83,0,77,0,44,0,19,0,0,0,184,0,144,0,44,0,22,0,156,0,114,0,108,0,144,0,246,0,188,0,171,0,3,0,244,0,116,0,108,0,45,0,53,0,0,0,160,0,223,0,0,0,237,0,183,0,58,0,248,0,110,0,0,0,96,0,101,0,241,0,219,0,0,0,12,0,179,0,0,0,9,0,206,0,227,0,247,0,0,0,13,0,56,0,0,0,0,0,78,0,0,0,133,0,178,0,126,0,149,0,107,0,31,0,79,0,86,0,0,0,199,0,230,0,211,0,0,0,207,0,0,0,214,0,20,0,0,0,130,0,242,0,0,0,189,0,31,0,55,0,242,0,60,0,187,0,27,0,120,0,191,0,107,0,18,0,252,0,9,0,178,0,163,0,222,0,64,0,204,0,0,0,138,0,241,0,0,0,191,0,147,0,209,0,0,0,0,0,178,0,67,0,142,0,254,0,212,0,185,0,126,0,80,0,25,0,17,0,128,0,128,0,40,0,168,0,0,0,184,0,112,0,0,0,108,0,198,0,187,0,20,0,153,0,143,0,22,0,99,0,82,0,135,0,57,0,108,0,0,0,16,0,226,0,20,0,60,0,140,0,102,0,0,0,236,0,57,0,32,0,135,0,0,0,96,0,71,0,0,0,0,0,0,0,143,0,139,0,212,0,89,0,213,0,162,0,98,0,122,0,205,0,0,0,171,0,0,0,1,0,80,0,72,0,0,0,250,0,247,0,138,0,191,0,169,0,133,0,129,0,189,0,17,0,13,0,9,0,225,0,211,0,0,0,215,0,224,0,42,0,145,0);
signal scenario_full  : scenario_type := (18,31,158,31,3,31,73,31,61,31,63,31,10,31,172,31,72,31,250,31,31,31,4,31,4,30,157,31,19,31,207,31,8,31,8,30,224,31,224,30,45,31,168,31,18,31,87,31,51,31,6,31,172,31,144,31,57,31,26,31,25,31,72,31,73,31,73,30,190,31,145,31,145,30,131,31,147,31,13,31,57,31,11,31,141,31,157,31,157,30,105,31,95,31,17,31,17,30,153,31,188,31,123,31,61,31,144,31,13,31,47,31,84,31,84,30,187,31,171,31,171,30,21,31,20,31,234,31,252,31,252,30,103,31,231,31,77,31,21,31,21,30,221,31,221,30,221,29,221,28,199,31,199,30,84,31,246,31,142,31,78,31,43,31,107,31,127,31,233,31,240,31,137,31,6,31,206,31,79,31,79,30,138,31,246,31,101,31,31,31,152,31,115,31,84,31,183,31,85,31,101,31,122,31,122,30,122,29,5,31,68,31,92,31,74,31,74,30,122,31,90,31,27,31,27,30,112,31,90,31,151,31,134,31,114,31,32,31,211,31,211,30,226,31,64,31,64,30,145,31,54,31,223,31,190,31,209,31,148,31,124,31,124,30,99,31,52,31,220,31,220,30,193,31,30,31,234,31,197,31,197,30,197,29,129,31,129,30,7,31,249,31,145,31,211,31,57,31,81,31,81,30,81,29,236,31,110,31,110,30,110,29,110,28,213,31,118,31,41,31,184,31,161,31,43,31,43,30,130,31,62,31,62,30,54,31,20,31,51,31,162,31,60,31,176,31,188,31,120,31,200,31,34,31,34,30,193,31,186,31,172,31,158,31,44,31,81,31,217,31,105,31,191,31,191,30,191,29,164,31,104,31,56,31,56,30,241,31,77,31,77,30,77,29,248,31,203,31,169,31,67,31,78,31,78,30,147,31,159,31,112,31,191,31,135,31,61,31,166,31,220,31,210,31,196,31,43,31,235,31,3,31,162,31,212,31,211,31,211,30,41,31,82,31,58,31,246,31,49,31,17,31,2,31,246,31,74,31,74,30,74,29,74,28,179,31,179,30,179,29,85,31,249,31,10,31,193,31,51,31,42,31,191,31,43,31,46,31,46,30,240,31,201,31,70,31,108,31,131,31,100,31,100,30,49,31,49,30,49,29,243,31,36,31,75,31,200,31,2,31,17,31,111,31,171,31,24,31,24,30,228,31,162,31,76,31,55,31,125,31,125,30,23,31,104,31,207,31,51,31,146,31,227,31,227,30,227,29,79,31,53,31,53,30,64,31,150,31,35,31,93,31,120,31,45,31,220,31,64,31,172,31,103,31,103,30,81,31,137,31,116,31,64,31,92,31,122,31,48,31,124,31,252,31,255,31,57,31,117,31,232,31,232,30,65,31,65,30,86,31,185,31,41,31,168,31,139,31,101,31,1,31,147,31,96,31,96,30,111,31,81,31,155,31,155,30,237,31,187,31,214,31,214,30,111,31,111,30,2,31,159,31,240,31,154,31,108,31,129,31,64,31,212,31,212,30,212,29,164,31,43,31,43,30,43,29,150,31,16,31,92,31,246,31,156,31,66,31,86,31,117,31,117,30,111,31,94,31,94,30,206,31,73,31,73,30,30,31,121,31,110,31,151,31,80,31,26,31,105,31,199,31,129,31,129,30,129,29,134,31,134,30,129,31,90,31,90,30,90,29,243,31,243,30,193,31,182,31,220,31,127,31,52,31,163,31,224,31,224,30,205,31,83,31,31,31,148,31,18,31,41,31,41,30,148,31,148,30,116,31,229,31,23,31,188,31,34,31,2,31,103,31,1,31,64,31,191,31,191,30,113,31,3,31,3,30,45,31,47,31,47,30,204,31,131,31,110,31,110,30,110,29,205,31,74,31,84,31,84,30,84,29,47,31,63,31,169,31,191,31,24,31,118,31,34,31,190,31,153,31,153,30,132,31,159,31,159,30,222,31,222,30,5,31,189,31,238,31,238,30,69,31,156,31,64,31,64,30,209,31,170,31,54,31,61,31,238,31,181,31,23,31,123,31,245,31,245,30,69,31,10,31,85,31,159,31,159,30,211,31,204,31,148,31,223,31,223,30,140,31,153,31,200,31,200,30,75,31,219,31,61,31,149,31,149,30,93,31,112,31,96,31,48,31,49,31,182,31,182,30,3,31,205,31,105,31,105,30,230,31,140,31,215,31,215,30,187,31,99,31,68,31,32,31,242,31,14,31,158,31,5,31,228,31,23,31,23,30,135,31,135,30,135,29,238,31,104,31,104,30,12,31,187,31,187,30,83,31,71,31,4,31,166,31,166,30,170,31,170,30,89,31,143,31,225,31,55,31,81,31,27,31,9,31,97,31,224,31,118,31,118,30,48,31,197,31,73,31,73,30,103,31,103,30,103,29,173,31,55,31,166,31,132,31,8,31,186,31,186,30,186,29,126,31,126,30,55,31,16,31,197,31,213,31,53,31,53,30,218,31,202,31,165,31,24,31,115,31,49,31,49,30,214,31,29,31,61,31,150,31,198,31,53,31,83,31,77,31,44,31,19,31,19,30,184,31,144,31,44,31,22,31,156,31,114,31,108,31,144,31,246,31,188,31,171,31,3,31,244,31,116,31,108,31,45,31,53,31,53,30,160,31,223,31,223,30,237,31,183,31,58,31,248,31,110,31,110,30,96,31,101,31,241,31,219,31,219,30,12,31,179,31,179,30,9,31,206,31,227,31,247,31,247,30,13,31,56,31,56,30,56,29,78,31,78,30,133,31,178,31,126,31,149,31,107,31,31,31,79,31,86,31,86,30,199,31,230,31,211,31,211,30,207,31,207,30,214,31,20,31,20,30,130,31,242,31,242,30,189,31,31,31,55,31,242,31,60,31,187,31,27,31,120,31,191,31,107,31,18,31,252,31,9,31,178,31,163,31,222,31,64,31,204,31,204,30,138,31,241,31,241,30,191,31,147,31,209,31,209,30,209,29,178,31,67,31,142,31,254,31,212,31,185,31,126,31,80,31,25,31,17,31,128,31,128,31,40,31,168,31,168,30,184,31,112,31,112,30,108,31,198,31,187,31,20,31,153,31,143,31,22,31,99,31,82,31,135,31,57,31,108,31,108,30,16,31,226,31,20,31,60,31,140,31,102,31,102,30,236,31,57,31,32,31,135,31,135,30,96,31,71,31,71,30,71,29,71,28,143,31,139,31,212,31,89,31,213,31,162,31,98,31,122,31,205,31,205,30,171,31,171,30,1,31,80,31,72,31,72,30,250,31,247,31,138,31,191,31,169,31,133,31,129,31,189,31,17,31,13,31,9,31,225,31,211,31,211,30,215,31,224,31,42,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
