-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 174;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (58,0,64,0,54,0,195,0,202,0,0,0,22,0,0,0,196,0,138,0,140,0,8,0,0,0,176,0,109,0,94,0,0,0,57,0,0,0,163,0,29,0,142,0,234,0,35,0,46,0,174,0,115,0,233,0,0,0,235,0,196,0,0,0,0,0,31,0,226,0,104,0,180,0,0,0,135,0,169,0,160,0,65,0,161,0,126,0,18,0,104,0,245,0,137,0,5,0,72,0,0,0,0,0,0,0,111,0,244,0,99,0,19,0,128,0,176,0,141,0,131,0,67,0,4,0,175,0,224,0,222,0,63,0,16,0,71,0,197,0,162,0,157,0,142,0,0,0,55,0,241,0,140,0,0,0,14,0,165,0,0,0,0,0,17,0,231,0,224,0,73,0,114,0,92,0,248,0,26,0,222,0,23,0,79,0,99,0,11,0,103,0,112,0,206,0,0,0,205,0,53,0,113,0,149,0,177,0,22,0,0,0,89,0,44,0,148,0,120,0,102,0,232,0,194,0,255,0,15,0,173,0,127,0,0,0,0,0,44,0,0,0,18,0,166,0,14,0,165,0,1,0,227,0,97,0,173,0,0,0,237,0,165,0,86,0,66,0,25,0,0,0,94,0,247,0,80,0,148,0,0,0,16,0,2,0,100,0,148,0,190,0,106,0,0,0,163,0,89,0,214,0,190,0,28,0,57,0,30,0,0,0,188,0,66,0,198,0,79,0,154,0,222,0,104,0,0,0,72,0,147,0,153,0,204,0,0,0,120,0,70,0,218,0,76,0,56,0);
signal scenario_full  : scenario_type := (58,31,64,31,54,31,195,31,202,31,202,30,22,31,22,30,196,31,138,31,140,31,8,31,8,30,176,31,109,31,94,31,94,30,57,31,57,30,163,31,29,31,142,31,234,31,35,31,46,31,174,31,115,31,233,31,233,30,235,31,196,31,196,30,196,29,31,31,226,31,104,31,180,31,180,30,135,31,169,31,160,31,65,31,161,31,126,31,18,31,104,31,245,31,137,31,5,31,72,31,72,30,72,29,72,28,111,31,244,31,99,31,19,31,128,31,176,31,141,31,131,31,67,31,4,31,175,31,224,31,222,31,63,31,16,31,71,31,197,31,162,31,157,31,142,31,142,30,55,31,241,31,140,31,140,30,14,31,165,31,165,30,165,29,17,31,231,31,224,31,73,31,114,31,92,31,248,31,26,31,222,31,23,31,79,31,99,31,11,31,103,31,112,31,206,31,206,30,205,31,53,31,113,31,149,31,177,31,22,31,22,30,89,31,44,31,148,31,120,31,102,31,232,31,194,31,255,31,15,31,173,31,127,31,127,30,127,29,44,31,44,30,18,31,166,31,14,31,165,31,1,31,227,31,97,31,173,31,173,30,237,31,165,31,86,31,66,31,25,31,25,30,94,31,247,31,80,31,148,31,148,30,16,31,2,31,100,31,148,31,190,31,106,31,106,30,163,31,89,31,214,31,190,31,28,31,57,31,30,31,30,30,188,31,66,31,198,31,79,31,154,31,222,31,104,31,104,30,72,31,147,31,153,31,204,31,204,30,120,31,70,31,218,31,76,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
