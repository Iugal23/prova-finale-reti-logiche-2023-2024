-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 860;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (215,0,182,0,86,0,205,0,178,0,155,0,24,0,0,0,0,0,0,0,8,0,206,0,82,0,124,0,241,0,207,0,139,0,0,0,175,0,23,0,162,0,243,0,0,0,0,0,172,0,161,0,53,0,0,0,239,0,0,0,168,0,215,0,34,0,113,0,25,0,0,0,184,0,0,0,69,0,116,0,0,0,198,0,43,0,106,0,112,0,31,0,173,0,38,0,0,0,0,0,127,0,0,0,60,0,0,0,0,0,96,0,219,0,0,0,0,0,0,0,152,0,251,0,178,0,0,0,147,0,76,0,45,0,39,0,26,0,0,0,63,0,157,0,33,0,57,0,56,0,134,0,105,0,189,0,210,0,30,0,0,0,0,0,0,0,136,0,0,0,243,0,6,0,165,0,128,0,220,0,232,0,154,0,13,0,35,0,101,0,224,0,76,0,161,0,0,0,1,0,5,0,0,0,25,0,61,0,87,0,178,0,155,0,82,0,225,0,143,0,177,0,161,0,0,0,0,0,186,0,0,0,133,0,184,0,235,0,5,0,248,0,227,0,36,0,31,0,0,0,0,0,133,0,0,0,163,0,0,0,109,0,206,0,0,0,233,0,166,0,4,0,22,0,48,0,0,0,110,0,209,0,22,0,208,0,144,0,0,0,160,0,199,0,198,0,0,0,162,0,62,0,0,0,184,0,217,0,117,0,115,0,3,0,0,0,178,0,25,0,235,0,124,0,145,0,58,0,158,0,0,0,127,0,198,0,196,0,239,0,14,0,53,0,73,0,43,0,62,0,14,0,0,0,0,0,107,0,227,0,87,0,122,0,0,0,142,0,236,0,54,0,254,0,103,0,66,0,252,0,20,0,105,0,0,0,175,0,0,0,0,0,0,0,0,0,48,0,208,0,123,0,0,0,164,0,0,0,168,0,123,0,58,0,13,0,217,0,245,0,158,0,44,0,204,0,0,0,216,0,23,0,151,0,0,0,65,0,0,0,0,0,0,0,109,0,56,0,120,0,0,0,203,0,239,0,208,0,0,0,35,0,55,0,220,0,0,0,120,0,214,0,219,0,21,0,77,0,0,0,0,0,176,0,229,0,11,0,0,0,91,0,185,0,238,0,168,0,251,0,152,0,223,0,0,0,156,0,131,0,0,0,0,0,0,0,211,0,46,0,128,0,158,0,130,0,104,0,84,0,168,0,249,0,254,0,63,0,19,0,120,0,0,0,135,0,141,0,0,0,0,0,0,0,0,0,25,0,212,0,91,0,58,0,215,0,0,0,79,0,173,0,0,0,138,0,0,0,0,0,38,0,112,0,15,0,181,0,210,0,21,0,164,0,224,0,208,0,95,0,0,0,61,0,0,0,9,0,146,0,191,0,67,0,0,0,0,0,251,0,225,0,8,0,134,0,81,0,141,0,11,0,50,0,152,0,189,0,238,0,214,0,117,0,188,0,14,0,170,0,35,0,133,0,0,0,64,0,0,0,56,0,244,0,216,0,0,0,198,0,82,0,82,0,20,0,4,0,193,0,62,0,237,0,215,0,22,0,0,0,89,0,112,0,89,0,17,0,115,0,0,0,47,0,102,0,77,0,0,0,245,0,37,0,0,0,243,0,196,0,89,0,0,0,87,0,82,0,120,0,70,0,153,0,0,0,232,0,100,0,81,0,0,0,4,0,9,0,213,0,68,0,92,0,240,0,100,0,0,0,80,0,51,0,0,0,45,0,150,0,0,0,241,0,158,0,91,0,132,0,20,0,75,0,0,0,140,0,66,0,0,0,177,0,0,0,85,0,118,0,0,0,210,0,202,0,153,0,67,0,219,0,0,0,26,0,0,0,133,0,21,0,187,0,244,0,0,0,40,0,119,0,0,0,157,0,16,0,0,0,0,0,55,0,218,0,21,0,0,0,3,0,0,0,115,0,30,0,47,0,193,0,65,0,0,0,128,0,171,0,92,0,40,0,144,0,33,0,241,0,0,0,4,0,0,0,120,0,188,0,0,0,0,0,15,0,155,0,96,0,63,0,108,0,41,0,55,0,43,0,104,0,231,0,92,0,141,0,255,0,27,0,0,0,0,0,0,0,71,0,115,0,115,0,96,0,51,0,0,0,144,0,235,0,24,0,242,0,105,0,0,0,0,0,115,0,0,0,229,0,0,0,146,0,0,0,80,0,231,0,134,0,79,0,160,0,82,0,163,0,0,0,116,0,168,0,151,0,243,0,139,0,221,0,255,0,27,0,16,0,174,0,56,0,138,0,249,0,115,0,180,0,162,0,90,0,77,0,0,0,121,0,19,0,69,0,186,0,0,0,116,0,90,0,196,0,101,0,36,0,6,0,0,0,0,0,133,0,0,0,106,0,241,0,113,0,32,0,233,0,62,0,0,0,0,0,69,0,122,0,210,0,123,0,0,0,0,0,0,0,117,0,0,0,113,0,12,0,236,0,150,0,172,0,80,0,183,0,20,0,0,0,114,0,0,0,0,0,27,0,164,0,0,0,0,0,0,0,0,0,115,0,0,0,253,0,187,0,0,0,116,0,68,0,10,0,0,0,146,0,77,0,53,0,158,0,41,0,184,0,52,0,222,0,86,0,0,0,46,0,108,0,59,0,0,0,234,0,231,0,188,0,0,0,191,0,50,0,212,0,217,0,103,0,254,0,81,0,53,0,0,0,112,0,74,0,149,0,175,0,64,0,41,0,0,0,72,0,248,0,146,0,252,0,207,0,46,0,156,0,221,0,157,0,0,0,145,0,174,0,0,0,34,0,136,0,164,0,151,0,171,0,0,0,205,0,52,0,0,0,72,0,171,0,231,0,106,0,35,0,20,0,0,0,125,0,158,0,78,0,86,0,100,0,173,0,0,0,0,0,146,0,152,0,192,0,12,0,203,0,133,0,0,0,132,0,81,0,0,0,246,0,220,0,27,0,21,0,179,0,133,0,154,0,5,0,0,0,38,0,46,0,14,0,56,0,0,0,0,0,125,0,38,0,68,0,140,0,219,0,8,0,25,0,216,0,175,0,225,0,11,0,70,0,22,0,17,0,152,0,138,0,232,0,72,0,104,0,116,0,189,0,0,0,64,0,85,0,0,0,187,0,220,0,154,0,168,0,56,0,0,0,84,0,143,0,0,0,41,0,0,0,0,0,0,0,94,0,220,0,84,0,177,0,201,0,0,0,0,0,60,0,62,0,0,0,208,0,214,0,225,0,192,0,69,0,42,0,1,0,15,0,49,0,102,0,0,0,229,0,62,0,179,0,0,0,141,0,50,0,217,0,25,0,144,0,107,0,0,0,184,0,228,0,182,0,133,0,90,0,39,0,0,0,206,0,145,0,105,0,0,0,0,0,230,0,0,0,15,0,199,0,0,0,73,0,0,0,245,0,151,0,72,0,82,0,108,0,77,0,17,0,76,0,79,0,31,0,98,0,76,0,110,0,0,0,193,0,198,0,211,0,206,0,53,0,152,0,0,0,0,0,0,0,129,0,152,0,97,0,0,0,93,0,146,0,157,0,182,0,76,0,224,0,135,0,54,0,109,0,84,0,0,0,231,0,118,0,99,0,181,0,120,0,0,0,0,0,12,0,191,0,229,0,62,0,35,0,4,0,59,0,51,0,210,0,244,0,29,0,233,0,0,0,125,0,30,0,81,0,234,0,136,0,171,0,63,0,202,0,0,0,250,0,0,0,11,0,166,0,228,0,214,0,0,0,221,0,241,0,144,0,160,0,11,0,164,0,12,0,64,0,27,0,165,0,0,0,139,0,25,0,181,0,234,0,90,0,0,0,126,0,34,0,239,0,82,0,150,0,232,0,113,0,211,0,193,0,137,0,199,0,0,0,0,0,218,0,0,0);
signal scenario_full  : scenario_type := (215,31,182,31,86,31,205,31,178,31,155,31,24,31,24,30,24,29,24,28,8,31,206,31,82,31,124,31,241,31,207,31,139,31,139,30,175,31,23,31,162,31,243,31,243,30,243,29,172,31,161,31,53,31,53,30,239,31,239,30,168,31,215,31,34,31,113,31,25,31,25,30,184,31,184,30,69,31,116,31,116,30,198,31,43,31,106,31,112,31,31,31,173,31,38,31,38,30,38,29,127,31,127,30,60,31,60,30,60,29,96,31,219,31,219,30,219,29,219,28,152,31,251,31,178,31,178,30,147,31,76,31,45,31,39,31,26,31,26,30,63,31,157,31,33,31,57,31,56,31,134,31,105,31,189,31,210,31,30,31,30,30,30,29,30,28,136,31,136,30,243,31,6,31,165,31,128,31,220,31,232,31,154,31,13,31,35,31,101,31,224,31,76,31,161,31,161,30,1,31,5,31,5,30,25,31,61,31,87,31,178,31,155,31,82,31,225,31,143,31,177,31,161,31,161,30,161,29,186,31,186,30,133,31,184,31,235,31,5,31,248,31,227,31,36,31,31,31,31,30,31,29,133,31,133,30,163,31,163,30,109,31,206,31,206,30,233,31,166,31,4,31,22,31,48,31,48,30,110,31,209,31,22,31,208,31,144,31,144,30,160,31,199,31,198,31,198,30,162,31,62,31,62,30,184,31,217,31,117,31,115,31,3,31,3,30,178,31,25,31,235,31,124,31,145,31,58,31,158,31,158,30,127,31,198,31,196,31,239,31,14,31,53,31,73,31,43,31,62,31,14,31,14,30,14,29,107,31,227,31,87,31,122,31,122,30,142,31,236,31,54,31,254,31,103,31,66,31,252,31,20,31,105,31,105,30,175,31,175,30,175,29,175,28,175,27,48,31,208,31,123,31,123,30,164,31,164,30,168,31,123,31,58,31,13,31,217,31,245,31,158,31,44,31,204,31,204,30,216,31,23,31,151,31,151,30,65,31,65,30,65,29,65,28,109,31,56,31,120,31,120,30,203,31,239,31,208,31,208,30,35,31,55,31,220,31,220,30,120,31,214,31,219,31,21,31,77,31,77,30,77,29,176,31,229,31,11,31,11,30,91,31,185,31,238,31,168,31,251,31,152,31,223,31,223,30,156,31,131,31,131,30,131,29,131,28,211,31,46,31,128,31,158,31,130,31,104,31,84,31,168,31,249,31,254,31,63,31,19,31,120,31,120,30,135,31,141,31,141,30,141,29,141,28,141,27,25,31,212,31,91,31,58,31,215,31,215,30,79,31,173,31,173,30,138,31,138,30,138,29,38,31,112,31,15,31,181,31,210,31,21,31,164,31,224,31,208,31,95,31,95,30,61,31,61,30,9,31,146,31,191,31,67,31,67,30,67,29,251,31,225,31,8,31,134,31,81,31,141,31,11,31,50,31,152,31,189,31,238,31,214,31,117,31,188,31,14,31,170,31,35,31,133,31,133,30,64,31,64,30,56,31,244,31,216,31,216,30,198,31,82,31,82,31,20,31,4,31,193,31,62,31,237,31,215,31,22,31,22,30,89,31,112,31,89,31,17,31,115,31,115,30,47,31,102,31,77,31,77,30,245,31,37,31,37,30,243,31,196,31,89,31,89,30,87,31,82,31,120,31,70,31,153,31,153,30,232,31,100,31,81,31,81,30,4,31,9,31,213,31,68,31,92,31,240,31,100,31,100,30,80,31,51,31,51,30,45,31,150,31,150,30,241,31,158,31,91,31,132,31,20,31,75,31,75,30,140,31,66,31,66,30,177,31,177,30,85,31,118,31,118,30,210,31,202,31,153,31,67,31,219,31,219,30,26,31,26,30,133,31,21,31,187,31,244,31,244,30,40,31,119,31,119,30,157,31,16,31,16,30,16,29,55,31,218,31,21,31,21,30,3,31,3,30,115,31,30,31,47,31,193,31,65,31,65,30,128,31,171,31,92,31,40,31,144,31,33,31,241,31,241,30,4,31,4,30,120,31,188,31,188,30,188,29,15,31,155,31,96,31,63,31,108,31,41,31,55,31,43,31,104,31,231,31,92,31,141,31,255,31,27,31,27,30,27,29,27,28,71,31,115,31,115,31,96,31,51,31,51,30,144,31,235,31,24,31,242,31,105,31,105,30,105,29,115,31,115,30,229,31,229,30,146,31,146,30,80,31,231,31,134,31,79,31,160,31,82,31,163,31,163,30,116,31,168,31,151,31,243,31,139,31,221,31,255,31,27,31,16,31,174,31,56,31,138,31,249,31,115,31,180,31,162,31,90,31,77,31,77,30,121,31,19,31,69,31,186,31,186,30,116,31,90,31,196,31,101,31,36,31,6,31,6,30,6,29,133,31,133,30,106,31,241,31,113,31,32,31,233,31,62,31,62,30,62,29,69,31,122,31,210,31,123,31,123,30,123,29,123,28,117,31,117,30,113,31,12,31,236,31,150,31,172,31,80,31,183,31,20,31,20,30,114,31,114,30,114,29,27,31,164,31,164,30,164,29,164,28,164,27,115,31,115,30,253,31,187,31,187,30,116,31,68,31,10,31,10,30,146,31,77,31,53,31,158,31,41,31,184,31,52,31,222,31,86,31,86,30,46,31,108,31,59,31,59,30,234,31,231,31,188,31,188,30,191,31,50,31,212,31,217,31,103,31,254,31,81,31,53,31,53,30,112,31,74,31,149,31,175,31,64,31,41,31,41,30,72,31,248,31,146,31,252,31,207,31,46,31,156,31,221,31,157,31,157,30,145,31,174,31,174,30,34,31,136,31,164,31,151,31,171,31,171,30,205,31,52,31,52,30,72,31,171,31,231,31,106,31,35,31,20,31,20,30,125,31,158,31,78,31,86,31,100,31,173,31,173,30,173,29,146,31,152,31,192,31,12,31,203,31,133,31,133,30,132,31,81,31,81,30,246,31,220,31,27,31,21,31,179,31,133,31,154,31,5,31,5,30,38,31,46,31,14,31,56,31,56,30,56,29,125,31,38,31,68,31,140,31,219,31,8,31,25,31,216,31,175,31,225,31,11,31,70,31,22,31,17,31,152,31,138,31,232,31,72,31,104,31,116,31,189,31,189,30,64,31,85,31,85,30,187,31,220,31,154,31,168,31,56,31,56,30,84,31,143,31,143,30,41,31,41,30,41,29,41,28,94,31,220,31,84,31,177,31,201,31,201,30,201,29,60,31,62,31,62,30,208,31,214,31,225,31,192,31,69,31,42,31,1,31,15,31,49,31,102,31,102,30,229,31,62,31,179,31,179,30,141,31,50,31,217,31,25,31,144,31,107,31,107,30,184,31,228,31,182,31,133,31,90,31,39,31,39,30,206,31,145,31,105,31,105,30,105,29,230,31,230,30,15,31,199,31,199,30,73,31,73,30,245,31,151,31,72,31,82,31,108,31,77,31,17,31,76,31,79,31,31,31,98,31,76,31,110,31,110,30,193,31,198,31,211,31,206,31,53,31,152,31,152,30,152,29,152,28,129,31,152,31,97,31,97,30,93,31,146,31,157,31,182,31,76,31,224,31,135,31,54,31,109,31,84,31,84,30,231,31,118,31,99,31,181,31,120,31,120,30,120,29,12,31,191,31,229,31,62,31,35,31,4,31,59,31,51,31,210,31,244,31,29,31,233,31,233,30,125,31,30,31,81,31,234,31,136,31,171,31,63,31,202,31,202,30,250,31,250,30,11,31,166,31,228,31,214,31,214,30,221,31,241,31,144,31,160,31,11,31,164,31,12,31,64,31,27,31,165,31,165,30,139,31,25,31,181,31,234,31,90,31,90,30,126,31,34,31,239,31,82,31,150,31,232,31,113,31,211,31,193,31,137,31,199,31,199,30,199,29,218,31,218,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
