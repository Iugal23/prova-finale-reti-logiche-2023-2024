-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 155;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (170,0,100,0,132,0,213,0,0,0,195,0,0,0,220,0,212,0,86,0,34,0,0,0,177,0,24,0,22,0,84,0,212,0,87,0,197,0,5,0,0,0,76,0,192,0,194,0,95,0,64,0,44,0,14,0,39,0,135,0,221,0,247,0,0,0,0,0,0,0,87,0,161,0,153,0,0,0,183,0,0,0,0,0,0,0,195,0,8,0,212,0,95,0,76,0,46,0,41,0,208,0,0,0,193,0,139,0,116,0,108,0,135,0,128,0,30,0,250,0,187,0,120,0,163,0,107,0,0,0,62,0,0,0,190,0,38,0,109,0,220,0,41,0,125,0,215,0,131,0,108,0,130,0,244,0,0,0,223,0,214,0,173,0,9,0,109,0,178,0,172,0,196,0,220,0,190,0,0,0,20,0,107,0,241,0,218,0,158,0,127,0,106,0,235,0,0,0,42,0,43,0,148,0,160,0,46,0,0,0,212,0,183,0,167,0,0,0,10,0,0,0,75,0,169,0,131,0,76,0,129,0,225,0,37,0,71,0,116,0,0,0,153,0,62,0,127,0,240,0,55,0,186,0,28,0,188,0,255,0,61,0,39,0,0,0,112,0,151,0,217,0,11,0,207,0,0,0,0,0,17,0,165,0,60,0,167,0,232,0,0,0,231,0,63,0,110,0,92,0,255,0,1,0,137,0,14,0,220,0);
signal scenario_full  : scenario_type := (170,31,100,31,132,31,213,31,213,30,195,31,195,30,220,31,212,31,86,31,34,31,34,30,177,31,24,31,22,31,84,31,212,31,87,31,197,31,5,31,5,30,76,31,192,31,194,31,95,31,64,31,44,31,14,31,39,31,135,31,221,31,247,31,247,30,247,29,247,28,87,31,161,31,153,31,153,30,183,31,183,30,183,29,183,28,195,31,8,31,212,31,95,31,76,31,46,31,41,31,208,31,208,30,193,31,139,31,116,31,108,31,135,31,128,31,30,31,250,31,187,31,120,31,163,31,107,31,107,30,62,31,62,30,190,31,38,31,109,31,220,31,41,31,125,31,215,31,131,31,108,31,130,31,244,31,244,30,223,31,214,31,173,31,9,31,109,31,178,31,172,31,196,31,220,31,190,31,190,30,20,31,107,31,241,31,218,31,158,31,127,31,106,31,235,31,235,30,42,31,43,31,148,31,160,31,46,31,46,30,212,31,183,31,167,31,167,30,10,31,10,30,75,31,169,31,131,31,76,31,129,31,225,31,37,31,71,31,116,31,116,30,153,31,62,31,127,31,240,31,55,31,186,31,28,31,188,31,255,31,61,31,39,31,39,30,112,31,151,31,217,31,11,31,207,31,207,30,207,29,17,31,165,31,60,31,167,31,232,31,232,30,231,31,63,31,110,31,92,31,255,31,1,31,137,31,14,31,220,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
