-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 594;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (88,0,239,0,214,0,22,0,138,0,236,0,207,0,60,0,137,0,138,0,186,0,220,0,0,0,31,0,177,0,84,0,41,0,70,0,187,0,144,0,199,0,2,0,198,0,152,0,188,0,68,0,0,0,65,0,51,0,26,0,60,0,220,0,26,0,248,0,0,0,170,0,127,0,175,0,101,0,236,0,16,0,0,0,178,0,45,0,76,0,0,0,78,0,189,0,0,0,47,0,0,0,180,0,0,0,99,0,7,0,137,0,26,0,222,0,121,0,234,0,28,0,224,0,236,0,27,0,0,0,0,0,132,0,232,0,89,0,0,0,45,0,18,0,146,0,125,0,226,0,100,0,172,0,140,0,164,0,155,0,181,0,92,0,221,0,165,0,204,0,230,0,21,0,97,0,0,0,210,0,68,0,37,0,171,0,0,0,197,0,255,0,0,0,0,0,95,0,246,0,107,0,124,0,124,0,0,0,143,0,211,0,79,0,211,0,10,0,0,0,0,0,32,0,103,0,17,0,87,0,31,0,0,0,0,0,100,0,129,0,247,0,155,0,14,0,68,0,168,0,128,0,147,0,73,0,0,0,215,0,0,0,0,0,215,0,25,0,0,0,0,0,155,0,0,0,0,0,140,0,31,0,133,0,79,0,99,0,21,0,158,0,17,0,0,0,0,0,0,0,188,0,129,0,163,0,0,0,0,0,0,0,94,0,35,0,176,0,97,0,111,0,250,0,241,0,201,0,252,0,168,0,150,0,252,0,89,0,132,0,140,0,0,0,109,0,68,0,0,0,77,0,68,0,0,0,34,0,217,0,24,0,62,0,14,0,149,0,238,0,172,0,110,0,0,0,255,0,145,0,41,0,203,0,0,0,213,0,0,0,94,0,0,0,41,0,25,0,0,0,141,0,56,0,206,0,0,0,35,0,0,0,121,0,189,0,186,0,0,0,161,0,18,0,126,0,0,0,216,0,26,0,50,0,48,0,245,0,52,0,188,0,103,0,0,0,201,0,52,0,185,0,206,0,0,0,0,0,189,0,0,0,41,0,25,0,117,0,241,0,128,0,39,0,148,0,0,0,193,0,205,0,69,0,96,0,69,0,0,0,235,0,234,0,170,0,0,0,23,0,155,0,222,0,17,0,127,0,0,0,0,0,15,0,226,0,0,0,64,0,0,0,51,0,128,0,0,0,104,0,201,0,108,0,144,0,88,0,232,0,170,0,132,0,0,0,52,0,171,0,34,0,234,0,0,0,178,0,97,0,0,0,146,0,9,0,0,0,111,0,227,0,135,0,251,0,209,0,0,0,242,0,0,0,27,0,178,0,24,0,96,0,167,0,182,0,246,0,119,0,140,0,155,0,197,0,130,0,44,0,144,0,139,0,136,0,63,0,170,0,54,0,95,0,21,0,73,0,236,0,0,0,126,0,136,0,229,0,245,0,246,0,1,0,34,0,11,0,111,0,87,0,183,0,0,0,193,0,124,0,0,0,0,0,40,0,182,0,0,0,1,0,124,0,166,0,0,0,174,0,201,0,57,0,157,0,101,0,58,0,186,0,13,0,38,0,0,0,33,0,60,0,164,0,95,0,104,0,70,0,20,0,153,0,17,0,0,0,0,0,56,0,0,0,87,0,162,0,35,0,15,0,88,0,20,0,179,0,0,0,195,0,154,0,196,0,170,0,7,0,0,0,0,0,71,0,45,0,65,0,0,0,0,0,9,0,0,0,73,0,107,0,167,0,127,0,103,0,0,0,0,0,0,0,242,0,50,0,214,0,102,0,0,0,0,0,200,0,215,0,42,0,179,0,205,0,5,0,0,0,56,0,223,0,190,0,180,0,0,0,0,0,124,0,59,0,211,0,254,0,112,0,218,0,81,0,254,0,9,0,130,0,133,0,105,0,208,0,14,0,13,0,10,0,44,0,0,0,39,0,89,0,48,0,167,0,0,0,105,0,0,0,0,0,12,0,86,0,217,0,227,0,60,0,49,0,6,0,141,0,50,0,181,0,5,0,216,0,132,0,0,0,202,0,177,0,107,0,0,0,62,0,94,0,242,0,55,0,94,0,187,0,135,0,102,0,100,0,13,0,111,0,242,0,160,0,90,0,197,0,39,0,133,0,193,0,2,0,225,0,0,0,190,0,176,0,0,0,0,0,155,0,5,0,26,0,17,0,127,0,155,0,8,0,75,0,234,0,203,0,0,0,0,0,0,0,235,0,251,0,43,0,112,0,133,0,182,0,232,0,202,0,237,0,0,0,132,0,192,0,46,0,192,0,73,0,70,0,88,0,204,0,0,0,0,0,0,0,155,0,221,0,20,0,0,0,76,0,0,0,200,0,207,0,144,0,0,0,37,0,126,0,55,0,45,0,230,0,126,0,161,0,0,0,233,0,0,0,93,0,48,0,189,0,65,0,0,0,72,0,70,0,130,0,146,0,119,0,229,0,121,0,55,0,64,0,105,0,116,0,98,0,77,0,0,0,0,0,229,0,100,0,207,0,86,0,157,0,181,0,199,0,84,0,178,0,238,0,242,0,197,0,220,0,76,0,106,0,192,0,136,0,3,0,0,0,234,0,0,0,107,0,67,0,151,0,173,0,0,0,197,0,178,0,10,0,109,0,106,0,0,0,101,0,251,0,86,0,115,0,202,0,200,0,246,0,233,0);
signal scenario_full  : scenario_type := (88,31,239,31,214,31,22,31,138,31,236,31,207,31,60,31,137,31,138,31,186,31,220,31,220,30,31,31,177,31,84,31,41,31,70,31,187,31,144,31,199,31,2,31,198,31,152,31,188,31,68,31,68,30,65,31,51,31,26,31,60,31,220,31,26,31,248,31,248,30,170,31,127,31,175,31,101,31,236,31,16,31,16,30,178,31,45,31,76,31,76,30,78,31,189,31,189,30,47,31,47,30,180,31,180,30,99,31,7,31,137,31,26,31,222,31,121,31,234,31,28,31,224,31,236,31,27,31,27,30,27,29,132,31,232,31,89,31,89,30,45,31,18,31,146,31,125,31,226,31,100,31,172,31,140,31,164,31,155,31,181,31,92,31,221,31,165,31,204,31,230,31,21,31,97,31,97,30,210,31,68,31,37,31,171,31,171,30,197,31,255,31,255,30,255,29,95,31,246,31,107,31,124,31,124,31,124,30,143,31,211,31,79,31,211,31,10,31,10,30,10,29,32,31,103,31,17,31,87,31,31,31,31,30,31,29,100,31,129,31,247,31,155,31,14,31,68,31,168,31,128,31,147,31,73,31,73,30,215,31,215,30,215,29,215,31,25,31,25,30,25,29,155,31,155,30,155,29,140,31,31,31,133,31,79,31,99,31,21,31,158,31,17,31,17,30,17,29,17,28,188,31,129,31,163,31,163,30,163,29,163,28,94,31,35,31,176,31,97,31,111,31,250,31,241,31,201,31,252,31,168,31,150,31,252,31,89,31,132,31,140,31,140,30,109,31,68,31,68,30,77,31,68,31,68,30,34,31,217,31,24,31,62,31,14,31,149,31,238,31,172,31,110,31,110,30,255,31,145,31,41,31,203,31,203,30,213,31,213,30,94,31,94,30,41,31,25,31,25,30,141,31,56,31,206,31,206,30,35,31,35,30,121,31,189,31,186,31,186,30,161,31,18,31,126,31,126,30,216,31,26,31,50,31,48,31,245,31,52,31,188,31,103,31,103,30,201,31,52,31,185,31,206,31,206,30,206,29,189,31,189,30,41,31,25,31,117,31,241,31,128,31,39,31,148,31,148,30,193,31,205,31,69,31,96,31,69,31,69,30,235,31,234,31,170,31,170,30,23,31,155,31,222,31,17,31,127,31,127,30,127,29,15,31,226,31,226,30,64,31,64,30,51,31,128,31,128,30,104,31,201,31,108,31,144,31,88,31,232,31,170,31,132,31,132,30,52,31,171,31,34,31,234,31,234,30,178,31,97,31,97,30,146,31,9,31,9,30,111,31,227,31,135,31,251,31,209,31,209,30,242,31,242,30,27,31,178,31,24,31,96,31,167,31,182,31,246,31,119,31,140,31,155,31,197,31,130,31,44,31,144,31,139,31,136,31,63,31,170,31,54,31,95,31,21,31,73,31,236,31,236,30,126,31,136,31,229,31,245,31,246,31,1,31,34,31,11,31,111,31,87,31,183,31,183,30,193,31,124,31,124,30,124,29,40,31,182,31,182,30,1,31,124,31,166,31,166,30,174,31,201,31,57,31,157,31,101,31,58,31,186,31,13,31,38,31,38,30,33,31,60,31,164,31,95,31,104,31,70,31,20,31,153,31,17,31,17,30,17,29,56,31,56,30,87,31,162,31,35,31,15,31,88,31,20,31,179,31,179,30,195,31,154,31,196,31,170,31,7,31,7,30,7,29,71,31,45,31,65,31,65,30,65,29,9,31,9,30,73,31,107,31,167,31,127,31,103,31,103,30,103,29,103,28,242,31,50,31,214,31,102,31,102,30,102,29,200,31,215,31,42,31,179,31,205,31,5,31,5,30,56,31,223,31,190,31,180,31,180,30,180,29,124,31,59,31,211,31,254,31,112,31,218,31,81,31,254,31,9,31,130,31,133,31,105,31,208,31,14,31,13,31,10,31,44,31,44,30,39,31,89,31,48,31,167,31,167,30,105,31,105,30,105,29,12,31,86,31,217,31,227,31,60,31,49,31,6,31,141,31,50,31,181,31,5,31,216,31,132,31,132,30,202,31,177,31,107,31,107,30,62,31,94,31,242,31,55,31,94,31,187,31,135,31,102,31,100,31,13,31,111,31,242,31,160,31,90,31,197,31,39,31,133,31,193,31,2,31,225,31,225,30,190,31,176,31,176,30,176,29,155,31,5,31,26,31,17,31,127,31,155,31,8,31,75,31,234,31,203,31,203,30,203,29,203,28,235,31,251,31,43,31,112,31,133,31,182,31,232,31,202,31,237,31,237,30,132,31,192,31,46,31,192,31,73,31,70,31,88,31,204,31,204,30,204,29,204,28,155,31,221,31,20,31,20,30,76,31,76,30,200,31,207,31,144,31,144,30,37,31,126,31,55,31,45,31,230,31,126,31,161,31,161,30,233,31,233,30,93,31,48,31,189,31,65,31,65,30,72,31,70,31,130,31,146,31,119,31,229,31,121,31,55,31,64,31,105,31,116,31,98,31,77,31,77,30,77,29,229,31,100,31,207,31,86,31,157,31,181,31,199,31,84,31,178,31,238,31,242,31,197,31,220,31,76,31,106,31,192,31,136,31,3,31,3,30,234,31,234,30,107,31,67,31,151,31,173,31,173,30,197,31,178,31,10,31,109,31,106,31,106,30,101,31,251,31,86,31,115,31,202,31,200,31,246,31,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
