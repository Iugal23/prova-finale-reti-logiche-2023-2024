-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_824 is
end project_tb_824;

architecture project_tb_arch_824 of project_tb_824 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 726;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,22,0,103,0,202,0,16,0,0,0,6,0,0,0,183,0,4,0,63,0,0,0,157,0,237,0,198,0,72,0,132,0,229,0,0,0,142,0,255,0,203,0,0,0,0,0,0,0,221,0,143,0,0,0,60,0,18,0,49,0,4,0,216,0,235,0,151,0,0,0,0,0,131,0,217,0,127,0,0,0,206,0,0,0,244,0,204,0,146,0,82,0,96,0,200,0,0,0,0,0,222,0,212,0,47,0,0,0,244,0,107,0,0,0,27,0,0,0,101,0,156,0,0,0,0,0,76,0,104,0,0,0,0,0,48,0,249,0,38,0,74,0,120,0,63,0,40,0,93,0,100,0,97,0,109,0,0,0,7,0,49,0,77,0,72,0,72,0,15,0,24,0,0,0,61,0,194,0,0,0,45,0,0,0,249,0,3,0,161,0,102,0,81,0,38,0,0,0,130,0,0,0,127,0,202,0,5,0,170,0,0,0,93,0,217,0,153,0,0,0,0,0,16,0,0,0,163,0,88,0,0,0,116,0,147,0,181,0,75,0,170,0,1,0,51,0,0,0,92,0,251,0,0,0,199,0,91,0,169,0,0,0,215,0,0,0,224,0,191,0,16,0,228,0,0,0,0,0,182,0,183,0,13,0,135,0,152,0,44,0,34,0,71,0,0,0,155,0,33,0,37,0,152,0,19,0,54,0,64,0,188,0,1,0,163,0,0,0,161,0,0,0,69,0,0,0,146,0,170,0,245,0,189,0,215,0,91,0,0,0,201,0,0,0,111,0,73,0,0,0,248,0,0,0,0,0,106,0,62,0,2,0,141,0,132,0,206,0,149,0,21,0,88,0,219,0,238,0,0,0,142,0,26,0,47,0,230,0,202,0,85,0,0,0,119,0,198,0,230,0,241,0,182,0,0,0,216,0,12,0,85,0,4,0,140,0,229,0,200,0,0,0,215,0,0,0,30,0,239,0,110,0,0,0,80,0,224,0,0,0,76,0,14,0,0,0,172,0,0,0,167,0,5,0,155,0,0,0,91,0,49,0,0,0,90,0,131,0,224,0,234,0,188,0,72,0,140,0,119,0,205,0,15,0,0,0,40,0,0,0,194,0,164,0,55,0,144,0,10,0,80,0,0,0,52,0,0,0,0,0,187,0,0,0,55,0,182,0,181,0,195,0,229,0,255,0,0,0,112,0,0,0,0,0,0,0,148,0,82,0,112,0,0,0,166,0,21,0,203,0,103,0,129,0,43,0,38,0,191,0,17,0,107,0,20,0,1,0,193,0,215,0,135,0,100,0,251,0,191,0,0,0,58,0,47,0,213,0,0,0,134,0,114,0,1,0,251,0,0,0,99,0,0,0,198,0,189,0,167,0,160,0,53,0,0,0,0,0,59,0,158,0,211,0,90,0,20,0,35,0,0,0,136,0,5,0,244,0,0,0,25,0,140,0,201,0,177,0,36,0,0,0,24,0,0,0,18,0,104,0,0,0,58,0,66,0,120,0,29,0,235,0,95,0,0,0,228,0,95,0,0,0,13,0,89,0,28,0,113,0,72,0,103,0,36,0,196,0,225,0,66,0,0,0,131,0,92,0,163,0,108,0,63,0,140,0,144,0,39,0,49,0,153,0,240,0,201,0,0,0,0,0,36,0,0,0,113,0,97,0,123,0,205,0,45,0,0,0,40,0,59,0,135,0,203,0,11,0,255,0,42,0,141,0,0,0,83,0,58,0,212,0,0,0,185,0,127,0,195,0,81,0,108,0,0,0,70,0,175,0,0,0,43,0,218,0,18,0,140,0,0,0,63,0,249,0,74,0,178,0,56,0,178,0,186,0,195,0,162,0,92,0,0,0,176,0,144,0,240,0,0,0,93,0,72,0,171,0,40,0,0,0,0,0,54,0,74,0,219,0,141,0,86,0,151,0,82,0,98,0,163,0,27,0,41,0,15,0,73,0,0,0,0,0,4,0,214,0,20,0,115,0,177,0,105,0,4,0,3,0,73,0,46,0,142,0,66,0,0,0,0,0,70,0,93,0,78,0,75,0,65,0,0,0,209,0,0,0,140,0,23,0,226,0,89,0,115,0,0,0,208,0,0,0,231,0,124,0,222,0,100,0,80,0,183,0,29,0,237,0,52,0,108,0,96,0,0,0,114,0,22,0,0,0,191,0,179,0,162,0,149,0,19,0,232,0,59,0,131,0,183,0,120,0,98,0,215,0,126,0,37,0,182,0,238,0,213,0,218,0,136,0,0,0,0,0,0,0,235,0,117,0,55,0,190,0,237,0,227,0,0,0,0,0,13,0,198,0,199,0,0,0,0,0,25,0,2,0,12,0,0,0,52,0,9,0,170,0,0,0,248,0,175,0,0,0,226,0,112,0,20,0,44,0,231,0,196,0,161,0,219,0,233,0,129,0,205,0,170,0,0,0,86,0,236,0,75,0,159,0,119,0,13,0,77,0,158,0,23,0,200,0,0,0,154,0,190,0,0,0,79,0,7,0,167,0,0,0,186,0,131,0,226,0,117,0,88,0,46,0,0,0,12,0,44,0,81,0,84,0,38,0,181,0,176,0,47,0,120,0,207,0,170,0,254,0,75,0,153,0,35,0,111,0,237,0,25,0,153,0,74,0,0,0,69,0,168,0,5,0,148,0,47,0,0,0,0,0,100,0,237,0,67,0,44,0,235,0,36,0,84,0,0,0,0,0,149,0,185,0,123,0,0,0,201,0,0,0,0,0,182,0,0,0,134,0,252,0,0,0,101,0,223,0,89,0,175,0,0,0,3,0,0,0,214,0,0,0,0,0,74,0,193,0,203,0,150,0,247,0,182,0,0,0,144,0,37,0,0,0,193,0,251,0,46,0,0,0,237,0,191,0,12,0,225,0,16,0,0,0,153,0,194,0,0,0,160,0,210,0,0,0,202,0,207,0,34,0,81,0,80,0,0,0,0,0,2,0,219,0,204,0,0,0,193,0,96,0,46,0,188,0,0,0,102,0,65,0,0,0,226,0,0,0,92,0,0,0,100,0,203,0,202,0,176,0,213,0,150,0,36,0,154,0,90,0,202,0,0,0,136,0,45,0,15,0,0,0,185,0,63,0,238,0,0,0,53,0,0,0,201,0,207,0,217,0,236,0,123,0,94,0,166,0,15,0,72,0,0,0,96,0,0,0,156,0,120,0,51,0,7,0,0,0,161,0,247,0,4,0,254,0,230,0,0,0,110,0,14,0,14,0,188,0,0,0,87,0,79,0);
signal scenario_full  : scenario_type := (0,0,22,31,103,31,202,31,16,31,16,30,6,31,6,30,183,31,4,31,63,31,63,30,157,31,237,31,198,31,72,31,132,31,229,31,229,30,142,31,255,31,203,31,203,30,203,29,203,28,221,31,143,31,143,30,60,31,18,31,49,31,4,31,216,31,235,31,151,31,151,30,151,29,131,31,217,31,127,31,127,30,206,31,206,30,244,31,204,31,146,31,82,31,96,31,200,31,200,30,200,29,222,31,212,31,47,31,47,30,244,31,107,31,107,30,27,31,27,30,101,31,156,31,156,30,156,29,76,31,104,31,104,30,104,29,48,31,249,31,38,31,74,31,120,31,63,31,40,31,93,31,100,31,97,31,109,31,109,30,7,31,49,31,77,31,72,31,72,31,15,31,24,31,24,30,61,31,194,31,194,30,45,31,45,30,249,31,3,31,161,31,102,31,81,31,38,31,38,30,130,31,130,30,127,31,202,31,5,31,170,31,170,30,93,31,217,31,153,31,153,30,153,29,16,31,16,30,163,31,88,31,88,30,116,31,147,31,181,31,75,31,170,31,1,31,51,31,51,30,92,31,251,31,251,30,199,31,91,31,169,31,169,30,215,31,215,30,224,31,191,31,16,31,228,31,228,30,228,29,182,31,183,31,13,31,135,31,152,31,44,31,34,31,71,31,71,30,155,31,33,31,37,31,152,31,19,31,54,31,64,31,188,31,1,31,163,31,163,30,161,31,161,30,69,31,69,30,146,31,170,31,245,31,189,31,215,31,91,31,91,30,201,31,201,30,111,31,73,31,73,30,248,31,248,30,248,29,106,31,62,31,2,31,141,31,132,31,206,31,149,31,21,31,88,31,219,31,238,31,238,30,142,31,26,31,47,31,230,31,202,31,85,31,85,30,119,31,198,31,230,31,241,31,182,31,182,30,216,31,12,31,85,31,4,31,140,31,229,31,200,31,200,30,215,31,215,30,30,31,239,31,110,31,110,30,80,31,224,31,224,30,76,31,14,31,14,30,172,31,172,30,167,31,5,31,155,31,155,30,91,31,49,31,49,30,90,31,131,31,224,31,234,31,188,31,72,31,140,31,119,31,205,31,15,31,15,30,40,31,40,30,194,31,164,31,55,31,144,31,10,31,80,31,80,30,52,31,52,30,52,29,187,31,187,30,55,31,182,31,181,31,195,31,229,31,255,31,255,30,112,31,112,30,112,29,112,28,148,31,82,31,112,31,112,30,166,31,21,31,203,31,103,31,129,31,43,31,38,31,191,31,17,31,107,31,20,31,1,31,193,31,215,31,135,31,100,31,251,31,191,31,191,30,58,31,47,31,213,31,213,30,134,31,114,31,1,31,251,31,251,30,99,31,99,30,198,31,189,31,167,31,160,31,53,31,53,30,53,29,59,31,158,31,211,31,90,31,20,31,35,31,35,30,136,31,5,31,244,31,244,30,25,31,140,31,201,31,177,31,36,31,36,30,24,31,24,30,18,31,104,31,104,30,58,31,66,31,120,31,29,31,235,31,95,31,95,30,228,31,95,31,95,30,13,31,89,31,28,31,113,31,72,31,103,31,36,31,196,31,225,31,66,31,66,30,131,31,92,31,163,31,108,31,63,31,140,31,144,31,39,31,49,31,153,31,240,31,201,31,201,30,201,29,36,31,36,30,113,31,97,31,123,31,205,31,45,31,45,30,40,31,59,31,135,31,203,31,11,31,255,31,42,31,141,31,141,30,83,31,58,31,212,31,212,30,185,31,127,31,195,31,81,31,108,31,108,30,70,31,175,31,175,30,43,31,218,31,18,31,140,31,140,30,63,31,249,31,74,31,178,31,56,31,178,31,186,31,195,31,162,31,92,31,92,30,176,31,144,31,240,31,240,30,93,31,72,31,171,31,40,31,40,30,40,29,54,31,74,31,219,31,141,31,86,31,151,31,82,31,98,31,163,31,27,31,41,31,15,31,73,31,73,30,73,29,4,31,214,31,20,31,115,31,177,31,105,31,4,31,3,31,73,31,46,31,142,31,66,31,66,30,66,29,70,31,93,31,78,31,75,31,65,31,65,30,209,31,209,30,140,31,23,31,226,31,89,31,115,31,115,30,208,31,208,30,231,31,124,31,222,31,100,31,80,31,183,31,29,31,237,31,52,31,108,31,96,31,96,30,114,31,22,31,22,30,191,31,179,31,162,31,149,31,19,31,232,31,59,31,131,31,183,31,120,31,98,31,215,31,126,31,37,31,182,31,238,31,213,31,218,31,136,31,136,30,136,29,136,28,235,31,117,31,55,31,190,31,237,31,227,31,227,30,227,29,13,31,198,31,199,31,199,30,199,29,25,31,2,31,12,31,12,30,52,31,9,31,170,31,170,30,248,31,175,31,175,30,226,31,112,31,20,31,44,31,231,31,196,31,161,31,219,31,233,31,129,31,205,31,170,31,170,30,86,31,236,31,75,31,159,31,119,31,13,31,77,31,158,31,23,31,200,31,200,30,154,31,190,31,190,30,79,31,7,31,167,31,167,30,186,31,131,31,226,31,117,31,88,31,46,31,46,30,12,31,44,31,81,31,84,31,38,31,181,31,176,31,47,31,120,31,207,31,170,31,254,31,75,31,153,31,35,31,111,31,237,31,25,31,153,31,74,31,74,30,69,31,168,31,5,31,148,31,47,31,47,30,47,29,100,31,237,31,67,31,44,31,235,31,36,31,84,31,84,30,84,29,149,31,185,31,123,31,123,30,201,31,201,30,201,29,182,31,182,30,134,31,252,31,252,30,101,31,223,31,89,31,175,31,175,30,3,31,3,30,214,31,214,30,214,29,74,31,193,31,203,31,150,31,247,31,182,31,182,30,144,31,37,31,37,30,193,31,251,31,46,31,46,30,237,31,191,31,12,31,225,31,16,31,16,30,153,31,194,31,194,30,160,31,210,31,210,30,202,31,207,31,34,31,81,31,80,31,80,30,80,29,2,31,219,31,204,31,204,30,193,31,96,31,46,31,188,31,188,30,102,31,65,31,65,30,226,31,226,30,92,31,92,30,100,31,203,31,202,31,176,31,213,31,150,31,36,31,154,31,90,31,202,31,202,30,136,31,45,31,15,31,15,30,185,31,63,31,238,31,238,30,53,31,53,30,201,31,207,31,217,31,236,31,123,31,94,31,166,31,15,31,72,31,72,30,96,31,96,30,156,31,120,31,51,31,7,31,7,30,161,31,247,31,4,31,254,31,230,31,230,30,110,31,14,31,14,31,188,31,188,30,87,31,79,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
