-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 846;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,37,0,189,0,53,0,30,0,97,0,71,0,52,0,81,0,0,0,0,0,131,0,20,0,159,0,0,0,10,0,181,0,250,0,136,0,53,0,240,0,0,0,0,0,0,0,88,0,146,0,202,0,0,0,0,0,7,0,39,0,180,0,122,0,169,0,4,0,149,0,35,0,157,0,0,0,1,0,64,0,0,0,0,0,0,0,218,0,19,0,30,0,0,0,86,0,166,0,220,0,156,0,232,0,201,0,76,0,246,0,254,0,254,0,0,0,0,0,41,0,244,0,125,0,0,0,0,0,0,0,241,0,187,0,106,0,0,0,8,0,138,0,140,0,244,0,19,0,225,0,216,0,57,0,167,0,138,0,126,0,97,0,57,0,189,0,37,0,146,0,0,0,0,0,14,0,251,0,243,0,137,0,0,0,37,0,45,0,157,0,132,0,199,0,195,0,29,0,204,0,223,0,10,0,111,0,213,0,0,0,133,0,82,0,13,0,53,0,78,0,180,0,135,0,47,0,134,0,144,0,45,0,151,0,0,0,145,0,8,0,91,0,29,0,107,0,20,0,144,0,0,0,41,0,0,0,164,0,67,0,107,0,69,0,128,0,103,0,71,0,217,0,166,0,203,0,98,0,11,0,238,0,161,0,146,0,233,0,144,0,5,0,159,0,48,0,248,0,59,0,165,0,38,0,39,0,0,0,139,0,240,0,0,0,145,0,235,0,190,0,240,0,235,0,0,0,0,0,68,0,94,0,205,0,0,0,65,0,226,0,180,0,0,0,46,0,0,0,204,0,86,0,160,0,237,0,206,0,255,0,127,0,7,0,0,0,226,0,6,0,160,0,117,0,167,0,58,0,212,0,92,0,61,0,185,0,0,0,27,0,52,0,198,0,38,0,0,0,46,0,0,0,108,0,10,0,197,0,130,0,0,0,16,0,189,0,38,0,28,0,49,0,206,0,77,0,232,0,120,0,121,0,195,0,207,0,69,0,108,0,241,0,42,0,50,0,136,0,154,0,187,0,130,0,60,0,62,0,51,0,165,0,147,0,210,0,54,0,3,0,160,0,238,0,211,0,0,0,30,0,118,0,0,0,169,0,53,0,53,0,123,0,174,0,216,0,0,0,169,0,186,0,166,0,209,0,105,0,155,0,75,0,0,0,126,0,251,0,29,0,156,0,0,0,186,0,172,0,69,0,0,0,91,0,72,0,251,0,139,0,0,0,137,0,104,0,160,0,125,0,70,0,0,0,46,0,0,0,120,0,163,0,124,0,65,0,171,0,220,0,218,0,34,0,12,0,155,0,0,0,191,0,18,0,0,0,167,0,0,0,10,0,0,0,119,0,169,0,92,0,200,0,16,0,233,0,210,0,229,0,177,0,191,0,148,0,253,0,88,0,169,0,116,0,49,0,0,0,72,0,0,0,0,0,185,0,158,0,27,0,117,0,4,0,0,0,241,0,172,0,227,0,22,0,191,0,100,0,231,0,34,0,30,0,0,0,185,0,0,0,39,0,0,0,108,0,10,0,188,0,218,0,0,0,137,0,7,0,123,0,115,0,0,0,181,0,0,0,132,0,0,0,0,0,175,0,167,0,0,0,134,0,0,0,95,0,0,0,202,0,173,0,214,0,92,0,70,0,98,0,91,0,0,0,202,0,87,0,0,0,0,0,0,0,210,0,238,0,246,0,193,0,0,0,0,0,0,0,127,0,58,0,75,0,96,0,49,0,133,0,83,0,205,0,71,0,116,0,28,0,39,0,245,0,180,0,54,0,153,0,247,0,2,0,0,0,97,0,240,0,173,0,0,0,115,0,35,0,193,0,0,0,25,0,135,0,183,0,116,0,98,0,10,0,107,0,0,0,157,0,0,0,0,0,111,0,0,0,233,0,33,0,158,0,38,0,24,0,57,0,57,0,0,0,222,0,57,0,34,0,200,0,0,0,116,0,32,0,145,0,0,0,47,0,205,0,119,0,189,0,92,0,226,0,126,0,189,0,183,0,0,0,21,0,49,0,158,0,248,0,152,0,59,0,56,0,56,0,49,0,22,0,29,0,203,0,160,0,47,0,54,0,70,0,92,0,64,0,235,0,31,0,124,0,0,0,23,0,60,0,5,0,61,0,0,0,0,0,174,0,58,0,102,0,0,0,35,0,97,0,138,0,0,0,0,0,0,0,10,0,204,0,0,0,219,0,234,0,0,0,221,0,43,0,58,0,8,0,30,0,182,0,14,0,124,0,1,0,33,0,38,0,176,0,0,0,95,0,100,0,131,0,103,0,184,0,240,0,171,0,0,0,235,0,198,0,47,0,58,0,0,0,143,0,147,0,199,0,118,0,162,0,173,0,147,0,51,0,75,0,0,0,250,0,0,0,0,0,11,0,149,0,54,0,132,0,3,0,175,0,39,0,0,0,176,0,0,0,208,0,62,0,0,0,252,0,0,0,0,0,132,0,0,0,21,0,186,0,0,0,106,0,1,0,132,0,0,0,225,0,30,0,201,0,0,0,85,0,118,0,249,0,134,0,0,0,83,0,213,0,33,0,41,0,53,0,41,0,71,0,131,0,131,0,175,0,25,0,243,0,106,0,253,0,0,0,114,0,125,0,76,0,60,0,235,0,134,0,211,0,73,0,21,0,0,0,223,0,81,0,103,0,53,0,150,0,102,0,76,0,187,0,183,0,49,0,254,0,26,0,194,0,203,0,173,0,85,0,152,0,101,0,33,0,174,0,205,0,0,0,3,0,161,0,206,0,108,0,0,0,67,0,215,0,13,0,70,0,153,0,251,0,94,0,115,0,43,0,177,0,78,0,217,0,30,0,56,0,219,0,243,0,153,0,180,0,206,0,241,0,219,0,204,0,78,0,145,0,0,0,201,0,205,0,220,0,14,0,23,0,56,0,254,0,121,0,20,0,44,0,203,0,0,0,106,0,79,0,65,0,225,0,68,0,1,0,61,0,1,0,0,0,195,0,116,0,20,0,0,0,252,0,157,0,51,0,233,0,13,0,0,0,0,0,200,0,84,0,26,0,19,0,0,0,179,0,136,0,0,0,0,0,63,0,140,0,2,0,7,0,23,0,107,0,19,0,122,0,75,0,245,0,49,0,0,0,0,0,0,0,229,0,47,0,0,0,141,0,154,0,140,0,0,0,79,0,0,0,0,0,28,0,47,0,236,0,232,0,0,0,24,0,216,0,0,0,165,0,177,0,3,0,57,0,0,0,53,0,0,0,0,0,247,0,102,0,203,0,152,0,105,0,0,0,0,0,17,0,0,0,0,0,0,0,0,0,161,0,0,0,198,0,83,0,52,0,195,0,10,0,48,0,0,0,0,0,207,0,115,0,23,0,71,0,0,0,27,0,133,0,0,0,0,0,9,0,166,0,0,0,216,0,0,0,177,0,0,0,0,0,130,0,159,0,247,0,108,0,80,0,250,0,0,0,0,0,193,0,88,0,225,0,0,0,0,0,195,0,163,0,153,0,48,0,243,0,67,0,218,0,175,0,0,0,18,0,139,0,100,0,150,0,0,0,223,0,151,0,119,0,228,0,223,0,255,0,25,0,0,0,0,0,125,0,102,0,236,0,47,0,118,0,1,0,107,0,0,0,101,0,0,0,199,0,92,0,239,0,76,0,123,0,108,0,245,0,0,0,0,0,39,0,158,0,88,0,0,0,255,0,214,0,88,0,112,0,203,0,175,0,246,0,43,0,0,0,225,0,149,0,0,0,28,0,40,0,0,0,78,0,201,0,0,0,58,0,5,0,234,0,234,0,0,0,63,0,0,0,40,0);
signal scenario_full  : scenario_type := (0,0,37,31,189,31,53,31,30,31,97,31,71,31,52,31,81,31,81,30,81,29,131,31,20,31,159,31,159,30,10,31,181,31,250,31,136,31,53,31,240,31,240,30,240,29,240,28,88,31,146,31,202,31,202,30,202,29,7,31,39,31,180,31,122,31,169,31,4,31,149,31,35,31,157,31,157,30,1,31,64,31,64,30,64,29,64,28,218,31,19,31,30,31,30,30,86,31,166,31,220,31,156,31,232,31,201,31,76,31,246,31,254,31,254,31,254,30,254,29,41,31,244,31,125,31,125,30,125,29,125,28,241,31,187,31,106,31,106,30,8,31,138,31,140,31,244,31,19,31,225,31,216,31,57,31,167,31,138,31,126,31,97,31,57,31,189,31,37,31,146,31,146,30,146,29,14,31,251,31,243,31,137,31,137,30,37,31,45,31,157,31,132,31,199,31,195,31,29,31,204,31,223,31,10,31,111,31,213,31,213,30,133,31,82,31,13,31,53,31,78,31,180,31,135,31,47,31,134,31,144,31,45,31,151,31,151,30,145,31,8,31,91,31,29,31,107,31,20,31,144,31,144,30,41,31,41,30,164,31,67,31,107,31,69,31,128,31,103,31,71,31,217,31,166,31,203,31,98,31,11,31,238,31,161,31,146,31,233,31,144,31,5,31,159,31,48,31,248,31,59,31,165,31,38,31,39,31,39,30,139,31,240,31,240,30,145,31,235,31,190,31,240,31,235,31,235,30,235,29,68,31,94,31,205,31,205,30,65,31,226,31,180,31,180,30,46,31,46,30,204,31,86,31,160,31,237,31,206,31,255,31,127,31,7,31,7,30,226,31,6,31,160,31,117,31,167,31,58,31,212,31,92,31,61,31,185,31,185,30,27,31,52,31,198,31,38,31,38,30,46,31,46,30,108,31,10,31,197,31,130,31,130,30,16,31,189,31,38,31,28,31,49,31,206,31,77,31,232,31,120,31,121,31,195,31,207,31,69,31,108,31,241,31,42,31,50,31,136,31,154,31,187,31,130,31,60,31,62,31,51,31,165,31,147,31,210,31,54,31,3,31,160,31,238,31,211,31,211,30,30,31,118,31,118,30,169,31,53,31,53,31,123,31,174,31,216,31,216,30,169,31,186,31,166,31,209,31,105,31,155,31,75,31,75,30,126,31,251,31,29,31,156,31,156,30,186,31,172,31,69,31,69,30,91,31,72,31,251,31,139,31,139,30,137,31,104,31,160,31,125,31,70,31,70,30,46,31,46,30,120,31,163,31,124,31,65,31,171,31,220,31,218,31,34,31,12,31,155,31,155,30,191,31,18,31,18,30,167,31,167,30,10,31,10,30,119,31,169,31,92,31,200,31,16,31,233,31,210,31,229,31,177,31,191,31,148,31,253,31,88,31,169,31,116,31,49,31,49,30,72,31,72,30,72,29,185,31,158,31,27,31,117,31,4,31,4,30,241,31,172,31,227,31,22,31,191,31,100,31,231,31,34,31,30,31,30,30,185,31,185,30,39,31,39,30,108,31,10,31,188,31,218,31,218,30,137,31,7,31,123,31,115,31,115,30,181,31,181,30,132,31,132,30,132,29,175,31,167,31,167,30,134,31,134,30,95,31,95,30,202,31,173,31,214,31,92,31,70,31,98,31,91,31,91,30,202,31,87,31,87,30,87,29,87,28,210,31,238,31,246,31,193,31,193,30,193,29,193,28,127,31,58,31,75,31,96,31,49,31,133,31,83,31,205,31,71,31,116,31,28,31,39,31,245,31,180,31,54,31,153,31,247,31,2,31,2,30,97,31,240,31,173,31,173,30,115,31,35,31,193,31,193,30,25,31,135,31,183,31,116,31,98,31,10,31,107,31,107,30,157,31,157,30,157,29,111,31,111,30,233,31,33,31,158,31,38,31,24,31,57,31,57,31,57,30,222,31,57,31,34,31,200,31,200,30,116,31,32,31,145,31,145,30,47,31,205,31,119,31,189,31,92,31,226,31,126,31,189,31,183,31,183,30,21,31,49,31,158,31,248,31,152,31,59,31,56,31,56,31,49,31,22,31,29,31,203,31,160,31,47,31,54,31,70,31,92,31,64,31,235,31,31,31,124,31,124,30,23,31,60,31,5,31,61,31,61,30,61,29,174,31,58,31,102,31,102,30,35,31,97,31,138,31,138,30,138,29,138,28,10,31,204,31,204,30,219,31,234,31,234,30,221,31,43,31,58,31,8,31,30,31,182,31,14,31,124,31,1,31,33,31,38,31,176,31,176,30,95,31,100,31,131,31,103,31,184,31,240,31,171,31,171,30,235,31,198,31,47,31,58,31,58,30,143,31,147,31,199,31,118,31,162,31,173,31,147,31,51,31,75,31,75,30,250,31,250,30,250,29,11,31,149,31,54,31,132,31,3,31,175,31,39,31,39,30,176,31,176,30,208,31,62,31,62,30,252,31,252,30,252,29,132,31,132,30,21,31,186,31,186,30,106,31,1,31,132,31,132,30,225,31,30,31,201,31,201,30,85,31,118,31,249,31,134,31,134,30,83,31,213,31,33,31,41,31,53,31,41,31,71,31,131,31,131,31,175,31,25,31,243,31,106,31,253,31,253,30,114,31,125,31,76,31,60,31,235,31,134,31,211,31,73,31,21,31,21,30,223,31,81,31,103,31,53,31,150,31,102,31,76,31,187,31,183,31,49,31,254,31,26,31,194,31,203,31,173,31,85,31,152,31,101,31,33,31,174,31,205,31,205,30,3,31,161,31,206,31,108,31,108,30,67,31,215,31,13,31,70,31,153,31,251,31,94,31,115,31,43,31,177,31,78,31,217,31,30,31,56,31,219,31,243,31,153,31,180,31,206,31,241,31,219,31,204,31,78,31,145,31,145,30,201,31,205,31,220,31,14,31,23,31,56,31,254,31,121,31,20,31,44,31,203,31,203,30,106,31,79,31,65,31,225,31,68,31,1,31,61,31,1,31,1,30,195,31,116,31,20,31,20,30,252,31,157,31,51,31,233,31,13,31,13,30,13,29,200,31,84,31,26,31,19,31,19,30,179,31,136,31,136,30,136,29,63,31,140,31,2,31,7,31,23,31,107,31,19,31,122,31,75,31,245,31,49,31,49,30,49,29,49,28,229,31,47,31,47,30,141,31,154,31,140,31,140,30,79,31,79,30,79,29,28,31,47,31,236,31,232,31,232,30,24,31,216,31,216,30,165,31,177,31,3,31,57,31,57,30,53,31,53,30,53,29,247,31,102,31,203,31,152,31,105,31,105,30,105,29,17,31,17,30,17,29,17,28,17,27,161,31,161,30,198,31,83,31,52,31,195,31,10,31,48,31,48,30,48,29,207,31,115,31,23,31,71,31,71,30,27,31,133,31,133,30,133,29,9,31,166,31,166,30,216,31,216,30,177,31,177,30,177,29,130,31,159,31,247,31,108,31,80,31,250,31,250,30,250,29,193,31,88,31,225,31,225,30,225,29,195,31,163,31,153,31,48,31,243,31,67,31,218,31,175,31,175,30,18,31,139,31,100,31,150,31,150,30,223,31,151,31,119,31,228,31,223,31,255,31,25,31,25,30,25,29,125,31,102,31,236,31,47,31,118,31,1,31,107,31,107,30,101,31,101,30,199,31,92,31,239,31,76,31,123,31,108,31,245,31,245,30,245,29,39,31,158,31,88,31,88,30,255,31,214,31,88,31,112,31,203,31,175,31,246,31,43,31,43,30,225,31,149,31,149,30,28,31,40,31,40,30,78,31,201,31,201,30,58,31,5,31,234,31,234,31,234,30,63,31,63,30,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
