-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_550 is
end project_tb_550;

architecture project_tb_arch_550 of project_tb_550 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 290;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,125,0,198,0,7,0,250,0,39,0,0,0,32,0,3,0,0,0,55,0,186,0,23,0,123,0,154,0,0,0,8,0,19,0,135,0,30,0,0,0,230,0,161,0,38,0,0,0,141,0,0,0,249,0,111,0,153,0,140,0,178,0,161,0,214,0,171,0,0,0,151,0,42,0,108,0,157,0,0,0,0,0,99,0,28,0,254,0,195,0,75,0,0,0,56,0,0,0,0,0,0,0,45,0,0,0,130,0,0,0,10,0,171,0,88,0,237,0,0,0,31,0,123,0,176,0,150,0,212,0,0,0,16,0,199,0,0,0,255,0,235,0,193,0,2,0,215,0,0,0,107,0,74,0,223,0,223,0,70,0,225,0,52,0,0,0,18,0,58,0,181,0,179,0,0,0,0,0,255,0,29,0,0,0,0,0,0,0,202,0,61,0,212,0,188,0,0,0,0,0,0,0,210,0,0,0,90,0,69,0,0,0,253,0,0,0,67,0,14,0,135,0,0,0,114,0,188,0,174,0,48,0,0,0,38,0,46,0,167,0,132,0,0,0,75,0,104,0,42,0,0,0,67,0,93,0,238,0,0,0,158,0,50,0,182,0,204,0,125,0,239,0,42,0,61,0,44,0,0,0,50,0,0,0,167,0,159,0,61,0,235,0,70,0,197,0,250,0,60,0,139,0,130,0,0,0,0,0,7,0,0,0,8,0,122,0,10,0,160,0,11,0,45,0,209,0,81,0,43,0,11,0,224,0,102,0,236,0,0,0,0,0,9,0,64,0,221,0,70,0,242,0,200,0,85,0,28,0,194,0,0,0,42,0,0,0,217,0,11,0,76,0,91,0,67,0,71,0,108,0,149,0,219,0,0,0,207,0,125,0,184,0,31,0,14,0,0,0,206,0,190,0,73,0,0,0,33,0,0,0,32,0,16,0,247,0,22,0,25,0,0,0,147,0,129,0,194,0,166,0,190,0,30,0,238,0,27,0,85,0,192,0,0,0,107,0,166,0,205,0,97,0,0,0,0,0,243,0,79,0,41,0,214,0,23,0,0,0,254,0,143,0,73,0,123,0,45,0,0,0,192,0,0,0,152,0,217,0,57,0,214,0,154,0,129,0,0,0,3,0,106,0,231,0,172,0,54,0,11,0,97,0,0,0,249,0,0,0,219,0,150,0,36,0,178,0,33,0,4,0,0,0,50,0,221,0,48,0,188,0,0,0,0,0,0,0,185,0,0,0,0,0,0,0,0,0,255,0,232,0,102,0,169,0,69,0,3,0,126,0,31,0,94,0,81,0,0,0);
signal scenario_full  : scenario_type := (71,31,125,31,198,31,7,31,250,31,39,31,39,30,32,31,3,31,3,30,55,31,186,31,23,31,123,31,154,31,154,30,8,31,19,31,135,31,30,31,30,30,230,31,161,31,38,31,38,30,141,31,141,30,249,31,111,31,153,31,140,31,178,31,161,31,214,31,171,31,171,30,151,31,42,31,108,31,157,31,157,30,157,29,99,31,28,31,254,31,195,31,75,31,75,30,56,31,56,30,56,29,56,28,45,31,45,30,130,31,130,30,10,31,171,31,88,31,237,31,237,30,31,31,123,31,176,31,150,31,212,31,212,30,16,31,199,31,199,30,255,31,235,31,193,31,2,31,215,31,215,30,107,31,74,31,223,31,223,31,70,31,225,31,52,31,52,30,18,31,58,31,181,31,179,31,179,30,179,29,255,31,29,31,29,30,29,29,29,28,202,31,61,31,212,31,188,31,188,30,188,29,188,28,210,31,210,30,90,31,69,31,69,30,253,31,253,30,67,31,14,31,135,31,135,30,114,31,188,31,174,31,48,31,48,30,38,31,46,31,167,31,132,31,132,30,75,31,104,31,42,31,42,30,67,31,93,31,238,31,238,30,158,31,50,31,182,31,204,31,125,31,239,31,42,31,61,31,44,31,44,30,50,31,50,30,167,31,159,31,61,31,235,31,70,31,197,31,250,31,60,31,139,31,130,31,130,30,130,29,7,31,7,30,8,31,122,31,10,31,160,31,11,31,45,31,209,31,81,31,43,31,11,31,224,31,102,31,236,31,236,30,236,29,9,31,64,31,221,31,70,31,242,31,200,31,85,31,28,31,194,31,194,30,42,31,42,30,217,31,11,31,76,31,91,31,67,31,71,31,108,31,149,31,219,31,219,30,207,31,125,31,184,31,31,31,14,31,14,30,206,31,190,31,73,31,73,30,33,31,33,30,32,31,16,31,247,31,22,31,25,31,25,30,147,31,129,31,194,31,166,31,190,31,30,31,238,31,27,31,85,31,192,31,192,30,107,31,166,31,205,31,97,31,97,30,97,29,243,31,79,31,41,31,214,31,23,31,23,30,254,31,143,31,73,31,123,31,45,31,45,30,192,31,192,30,152,31,217,31,57,31,214,31,154,31,129,31,129,30,3,31,106,31,231,31,172,31,54,31,11,31,97,31,97,30,249,31,249,30,219,31,150,31,36,31,178,31,33,31,4,31,4,30,50,31,221,31,48,31,188,31,188,30,188,29,188,28,185,31,185,30,185,29,185,28,185,27,255,31,232,31,102,31,169,31,69,31,3,31,126,31,31,31,94,31,81,31,81,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
