-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 464;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (216,0,0,0,244,0,253,0,0,0,99,0,175,0,26,0,0,0,218,0,0,0,228,0,120,0,0,0,100,0,126,0,140,0,168,0,166,0,0,0,128,0,135,0,236,0,0,0,199,0,156,0,0,0,135,0,9,0,63,0,50,0,110,0,0,0,0,0,12,0,168,0,96,0,202,0,159,0,10,0,123,0,0,0,103,0,63,0,49,0,0,0,25,0,198,0,63,0,214,0,189,0,93,0,11,0,67,0,179,0,184,0,51,0,29,0,132,0,246,0,0,0,64,0,69,0,0,0,81,0,0,0,174,0,87,0,53,0,27,0,3,0,107,0,160,0,118,0,0,0,47,0,101,0,60,0,221,0,246,0,147,0,73,0,68,0,172,0,0,0,152,0,40,0,160,0,212,0,122,0,212,0,231,0,0,0,0,0,233,0,116,0,145,0,30,0,70,0,156,0,165,0,52,0,38,0,97,0,158,0,63,0,169,0,0,0,16,0,104,0,168,0,199,0,0,0,133,0,222,0,65,0,74,0,137,0,192,0,221,0,156,0,0,0,134,0,124,0,46,0,147,0,0,0,39,0,139,0,0,0,166,0,139,0,193,0,248,0,125,0,224,0,0,0,227,0,244,0,156,0,134,0,227,0,152,0,159,0,139,0,0,0,57,0,0,0,0,0,255,0,0,0,0,0,43,0,3,0,0,0,198,0,86,0,254,0,142,0,115,0,17,0,0,0,154,0,19,0,12,0,34,0,134,0,238,0,142,0,127,0,185,0,96,0,119,0,9,0,155,0,56,0,0,0,237,0,0,0,47,0,55,0,254,0,195,0,201,0,128,0,0,0,158,0,0,0,213,0,0,0,57,0,212,0,192,0,161,0,217,0,69,0,0,0,218,0,133,0,246,0,118,0,211,0,0,0,0,0,146,0,9,0,115,0,137,0,92,0,110,0,0,0,27,0,0,0,0,0,72,0,160,0,100,0,0,0,0,0,193,0,0,0,249,0,91,0,96,0,49,0,198,0,40,0,144,0,98,0,172,0,163,0,240,0,0,0,0,0,204,0,130,0,101,0,47,0,39,0,0,0,54,0,15,0,201,0,151,0,112,0,200,0,53,0,0,0,0,0,182,0,197,0,0,0,250,0,42,0,191,0,220,0,102,0,218,0,70,0,50,0,204,0,193,0,75,0,117,0,199,0,206,0,119,0,187,0,112,0,0,0,153,0,163,0,108,0,240,0,0,0,27,0,0,0,195,0,199,0,126,0,71,0,35,0,215,0,70,0,0,0,120,0,24,0,244,0,0,0,79,0,205,0,0,0,7,0,111,0,90,0,123,0,153,0,226,0,125,0,197,0,210,0,27,0,195,0,221,0,65,0,24,0,105,0,7,0,140,0,198,0,239,0,246,0,206,0,160,0,166,0,105,0,172,0,0,0,172,0,0,0,0,0,0,0,212,0,0,0,30,0,140,0,14,0,55,0,44,0,0,0,20,0,66,0,46,0,74,0,0,0,97,0,0,0,181,0,203,0,174,0,185,0,174,0,148,0,186,0,0,0,180,0,154,0,0,0,84,0,202,0,128,0,234,0,174,0,4,0,86,0,0,0,173,0,78,0,0,0,157,0,205,0,212,0,115,0,184,0,0,0,70,0,85,0,165,0,0,0,194,0,0,0,146,0,148,0,96,0,6,0,181,0,0,0,52,0,37,0,35,0,142,0,188,0,104,0,202,0,201,0,130,0,0,0,68,0,99,0,107,0,164,0,45,0,0,0,97,0,0,0,210,0,53,0,206,0,133,0,116,0,238,0,178,0,24,0,0,0,0,0,227,0,0,0,31,0,207,0,75,0,252,0,181,0,178,0,46,0,254,0,0,0,142,0,10,0,202,0,236,0,32,0,77,0,0,0,163,0,1,0,153,0,0,0,193,0,245,0,3,0,101,0,68,0,188,0,0,0,37,0,70,0,121,0,0,0,0,0,103,0,44,0,77,0,90,0,0,0,97,0,219,0,234,0,0,0,116,0,133,0,163,0,12,0,0,0,182,0,39,0,85,0,43,0,0,0,144,0,229,0,30,0,103,0,231,0,0,0);
signal scenario_full  : scenario_type := (216,31,216,30,244,31,253,31,253,30,99,31,175,31,26,31,26,30,218,31,218,30,228,31,120,31,120,30,100,31,126,31,140,31,168,31,166,31,166,30,128,31,135,31,236,31,236,30,199,31,156,31,156,30,135,31,9,31,63,31,50,31,110,31,110,30,110,29,12,31,168,31,96,31,202,31,159,31,10,31,123,31,123,30,103,31,63,31,49,31,49,30,25,31,198,31,63,31,214,31,189,31,93,31,11,31,67,31,179,31,184,31,51,31,29,31,132,31,246,31,246,30,64,31,69,31,69,30,81,31,81,30,174,31,87,31,53,31,27,31,3,31,107,31,160,31,118,31,118,30,47,31,101,31,60,31,221,31,246,31,147,31,73,31,68,31,172,31,172,30,152,31,40,31,160,31,212,31,122,31,212,31,231,31,231,30,231,29,233,31,116,31,145,31,30,31,70,31,156,31,165,31,52,31,38,31,97,31,158,31,63,31,169,31,169,30,16,31,104,31,168,31,199,31,199,30,133,31,222,31,65,31,74,31,137,31,192,31,221,31,156,31,156,30,134,31,124,31,46,31,147,31,147,30,39,31,139,31,139,30,166,31,139,31,193,31,248,31,125,31,224,31,224,30,227,31,244,31,156,31,134,31,227,31,152,31,159,31,139,31,139,30,57,31,57,30,57,29,255,31,255,30,255,29,43,31,3,31,3,30,198,31,86,31,254,31,142,31,115,31,17,31,17,30,154,31,19,31,12,31,34,31,134,31,238,31,142,31,127,31,185,31,96,31,119,31,9,31,155,31,56,31,56,30,237,31,237,30,47,31,55,31,254,31,195,31,201,31,128,31,128,30,158,31,158,30,213,31,213,30,57,31,212,31,192,31,161,31,217,31,69,31,69,30,218,31,133,31,246,31,118,31,211,31,211,30,211,29,146,31,9,31,115,31,137,31,92,31,110,31,110,30,27,31,27,30,27,29,72,31,160,31,100,31,100,30,100,29,193,31,193,30,249,31,91,31,96,31,49,31,198,31,40,31,144,31,98,31,172,31,163,31,240,31,240,30,240,29,204,31,130,31,101,31,47,31,39,31,39,30,54,31,15,31,201,31,151,31,112,31,200,31,53,31,53,30,53,29,182,31,197,31,197,30,250,31,42,31,191,31,220,31,102,31,218,31,70,31,50,31,204,31,193,31,75,31,117,31,199,31,206,31,119,31,187,31,112,31,112,30,153,31,163,31,108,31,240,31,240,30,27,31,27,30,195,31,199,31,126,31,71,31,35,31,215,31,70,31,70,30,120,31,24,31,244,31,244,30,79,31,205,31,205,30,7,31,111,31,90,31,123,31,153,31,226,31,125,31,197,31,210,31,27,31,195,31,221,31,65,31,24,31,105,31,7,31,140,31,198,31,239,31,246,31,206,31,160,31,166,31,105,31,172,31,172,30,172,31,172,30,172,29,172,28,212,31,212,30,30,31,140,31,14,31,55,31,44,31,44,30,20,31,66,31,46,31,74,31,74,30,97,31,97,30,181,31,203,31,174,31,185,31,174,31,148,31,186,31,186,30,180,31,154,31,154,30,84,31,202,31,128,31,234,31,174,31,4,31,86,31,86,30,173,31,78,31,78,30,157,31,205,31,212,31,115,31,184,31,184,30,70,31,85,31,165,31,165,30,194,31,194,30,146,31,148,31,96,31,6,31,181,31,181,30,52,31,37,31,35,31,142,31,188,31,104,31,202,31,201,31,130,31,130,30,68,31,99,31,107,31,164,31,45,31,45,30,97,31,97,30,210,31,53,31,206,31,133,31,116,31,238,31,178,31,24,31,24,30,24,29,227,31,227,30,31,31,207,31,75,31,252,31,181,31,178,31,46,31,254,31,254,30,142,31,10,31,202,31,236,31,32,31,77,31,77,30,163,31,1,31,153,31,153,30,193,31,245,31,3,31,101,31,68,31,188,31,188,30,37,31,70,31,121,31,121,30,121,29,103,31,44,31,77,31,90,31,90,30,97,31,219,31,234,31,234,30,116,31,133,31,163,31,12,31,12,30,182,31,39,31,85,31,43,31,43,30,144,31,229,31,30,31,103,31,231,31,231,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
