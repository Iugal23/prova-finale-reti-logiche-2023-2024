-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_202 is
end project_tb_202;

architecture project_tb_arch_202 of project_tb_202 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 947;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,0,0,10,0,0,0,221,0,59,0,253,0,0,0,112,0,98,0,54,0,47,0,218,0,43,0,189,0,82,0,98,0,224,0,189,0,136,0,89,0,246,0,5,0,79,0,219,0,0,0,19,0,69,0,3,0,0,0,117,0,0,0,5,0,0,0,119,0,97,0,164,0,223,0,4,0,0,0,215,0,6,0,255,0,75,0,127,0,18,0,0,0,0,0,39,0,0,0,37,0,20,0,0,0,33,0,150,0,129,0,0,0,88,0,0,0,0,0,191,0,86,0,196,0,73,0,201,0,235,0,188,0,164,0,0,0,127,0,249,0,65,0,0,0,36,0,0,0,124,0,0,0,226,0,112,0,18,0,202,0,186,0,255,0,57,0,0,0,0,0,204,0,250,0,29,0,169,0,35,0,134,0,56,0,151,0,177,0,0,0,228,0,115,0,153,0,51,0,40,0,239,0,0,0,63,0,216,0,0,0,1,0,187,0,204,0,4,0,229,0,64,0,0,0,93,0,158,0,60,0,138,0,134,0,7,0,82,0,0,0,137,0,0,0,0,0,33,0,99,0,0,0,0,0,75,0,53,0,225,0,0,0,204,0,171,0,77,0,153,0,29,0,162,0,48,0,248,0,19,0,82,0,151,0,218,0,0,0,138,0,183,0,151,0,72,0,82,0,213,0,203,0,23,0,251,0,27,0,70,0,211,0,186,0,227,0,0,0,0,0,85,0,165,0,48,0,120,0,228,0,125,0,0,0,249,0,235,0,0,0,0,0,201,0,49,0,189,0,128,0,190,0,194,0,252,0,126,0,255,0,17,0,0,0,0,0,114,0,169,0,154,0,151,0,173,0,0,0,12,0,41,0,119,0,0,0,219,0,178,0,14,0,7,0,10,0,33,0,221,0,18,0,120,0,26,0,166,0,130,0,120,0,57,0,153,0,162,0,129,0,126,0,79,0,0,0,0,0,192,0,0,0,57,0,0,0,0,0,99,0,6,0,229,0,173,0,45,0,0,0,201,0,161,0,197,0,0,0,0,0,12,0,15,0,0,0,107,0,109,0,176,0,196,0,152,0,0,0,80,0,252,0,107,0,190,0,183,0,0,0,170,0,90,0,78,0,11,0,170,0,184,0,0,0,220,0,114,0,237,0,40,0,0,0,213,0,168,0,37,0,149,0,255,0,212,0,63,0,146,0,23,0,0,0,0,0,249,0,33,0,0,0,0,0,173,0,0,0,135,0,0,0,249,0,78,0,213,0,130,0,79,0,221,0,0,0,67,0,248,0,15,0,16,0,0,0,42,0,161,0,220,0,0,0,198,0,0,0,0,0,135,0,110,0,142,0,77,0,145,0,189,0,190,0,50,0,0,0,131,0,0,0,5,0,166,0,17,0,77,0,44,0,200,0,0,0,106,0,77,0,40,0,62,0,217,0,255,0,172,0,202,0,121,0,125,0,55,0,20,0,0,0,156,0,224,0,0,0,98,0,0,0,0,0,203,0,116,0,140,0,42,0,168,0,155,0,168,0,104,0,24,0,66,0,0,0,4,0,167,0,122,0,188,0,9,0,131,0,26,0,0,0,11,0,55,0,98,0,156,0,172,0,0,0,143,0,201,0,159,0,57,0,0,0,97,0,28,0,167,0,71,0,0,0,0,0,213,0,78,0,0,0,0,0,101,0,53,0,51,0,174,0,36,0,48,0,97,0,150,0,211,0,0,0,0,0,162,0,7,0,235,0,0,0,103,0,121,0,3,0,223,0,218,0,35,0,168,0,0,0,0,0,127,0,230,0,127,0,163,0,81,0,94,0,33,0,0,0,100,0,70,0,170,0,86,0,109,0,95,0,190,0,188,0,0,0,81,0,0,0,88,0,175,0,7,0,162,0,174,0,113,0,245,0,4,0,150,0,133,0,153,0,23,0,77,0,108,0,25,0,76,0,76,0,81,0,28,0,0,0,57,0,71,0,171,0,0,0,107,0,106,0,117,0,138,0,204,0,146,0,201,0,14,0,90,0,143,0,209,0,0,0,46,0,51,0,187,0,112,0,56,0,182,0,73,0,165,0,239,0,255,0,0,0,163,0,39,0,58,0,225,0,194,0,56,0,70,0,161,0,75,0,108,0,204,0,0,0,41,0,30,0,25,0,74,0,30,0,131,0,0,0,88,0,12,0,107,0,145,0,86,0,245,0,48,0,234,0,196,0,236,0,246,0,0,0,254,0,112,0,0,0,0,0,101,0,84,0,52,0,100,0,181,0,149,0,0,0,53,0,204,0,0,0,233,0,107,0,221,0,84,0,197,0,18,0,0,0,0,0,67,0,177,0,54,0,139,0,11,0,171,0,24,0,62,0,28,0,125,0,0,0,27,0,41,0,73,0,170,0,157,0,98,0,19,0,173,0,0,0,95,0,100,0,22,0,0,0,29,0,234,0,47,0,10,0,179,0,241,0,11,0,0,0,198,0,31,0,0,0,35,0,0,0,32,0,70,0,74,0,112,0,45,0,60,0,70,0,20,0,0,0,75,0,0,0,125,0,24,0,0,0,168,0,0,0,11,0,163,0,125,0,140,0,0,0,177,0,98,0,173,0,135,0,205,0,230,0,21,0,63,0,0,0,236,0,107,0,0,0,24,0,71,0,180,0,150,0,18,0,144,0,243,0,230,0,247,0,58,0,198,0,52,0,0,0,38,0,126,0,113,0,26,0,235,0,183,0,179,0,120,0,221,0,187,0,127,0,86,0,211,0,122,0,106,0,199,0,0,0,77,0,144,0,10,0,146,0,115,0,162,0,50,0,127,0,116,0,201,0,205,0,0,0,129,0,0,0,68,0,108,0,0,0,0,0,251,0,22,0,0,0,105,0,91,0,179,0,86,0,16,0,180,0,166,0,80,0,49,0,239,0,73,0,197,0,118,0,252,0,206,0,126,0,248,0,180,0,31,0,13,0,67,0,162,0,0,0,220,0,54,0,59,0,234,0,59,0,250,0,74,0,0,0,94,0,44,0,85,0,179,0,87,0,107,0,0,0,39,0,52,0,0,0,0,0,97,0,86,0,249,0,172,0,33,0,0,0,179,0,0,0,154,0,137,0,112,0,66,0,33,0,108,0,0,0,0,0,245,0,229,0,79,0,255,0,224,0,65,0,133,0,91,0,66,0,206,0,116,0,68,0,29,0,105,0,24,0,99,0,51,0,0,0,226,0,137,0,120,0,161,0,6,0,203,0,189,0,0,0,0,0,98,0,52,0,212,0,221,0,46,0,166,0,0,0,51,0,0,0,0,0,0,0,0,0,25,0,139,0,161,0,27,0,55,0,241,0,31,0,0,0,39,0,119,0,0,0,187,0,212,0,186,0,224,0,255,0,134,0,21,0,85,0,25,0,146,0,79,0,62,0,203,0,255,0,0,0,23,0,158,0,161,0,23,0,0,0,0,0,97,0,26,0,190,0,0,0,211,0,80,0,0,0,189,0,210,0,226,0,174,0,67,0,127,0,0,0,182,0,0,0,166,0,0,0,175,0,65,0,89,0,245,0,5,0,0,0,102,0,8,0,248,0,0,0,251,0,20,0,0,0,7,0,220,0,0,0,88,0,44,0,142,0,18,0,247,0,175,0,70,0,21,0,242,0,0,0,163,0,99,0,5,0,56,0,209,0,0,0,1,0,0,0,125,0,112,0,0,0,160,0,182,0,212,0,224,0,181,0,121,0,0,0,34,0,30,0,0,0,77,0,0,0,209,0,96,0,145,0,199,0,61,0,167,0,0,0,0,0,239,0,169,0,112,0,0,0,72,0,2,0,104,0,255,0,58,0,0,0,74,0,159,0,150,0,67,0,89,0,149,0,33,0,230,0,113,0,248,0,0,0,62,0,174,0,103,0,8,0,70,0,155,0,34,0,1,0,252,0,54,0,249,0,126,0,46,0,2,0,23,0,0,0,0,0,45,0,4,0,163,0,51,0,0,0,31,0,52,0,40,0,170,0,65,0,90,0,173,0,249,0,234,0,138,0,0,0,0,0,69,0,115,0,119,0,0,0,118,0,187,0,247,0,0,0,85,0,0,0,0,0,0,0,0,0,28,0,84,0,0,0,25,0,145,0,0,0,179,0,114,0,0,0,174,0,118,0,5,0,0,0,153,0,179,0,9,0,0,0,179,0,176,0,107,0,46,0,0,0,246,0,0,0,120,0,122,0,100,0,168,0,99,0,8,0,0,0,172,0,233,0,235,0,220,0,212,0,253,0,205,0);
signal scenario_full  : scenario_type := (69,31,69,30,10,31,10,30,221,31,59,31,253,31,253,30,112,31,98,31,54,31,47,31,218,31,43,31,189,31,82,31,98,31,224,31,189,31,136,31,89,31,246,31,5,31,79,31,219,31,219,30,19,31,69,31,3,31,3,30,117,31,117,30,5,31,5,30,119,31,97,31,164,31,223,31,4,31,4,30,215,31,6,31,255,31,75,31,127,31,18,31,18,30,18,29,39,31,39,30,37,31,20,31,20,30,33,31,150,31,129,31,129,30,88,31,88,30,88,29,191,31,86,31,196,31,73,31,201,31,235,31,188,31,164,31,164,30,127,31,249,31,65,31,65,30,36,31,36,30,124,31,124,30,226,31,112,31,18,31,202,31,186,31,255,31,57,31,57,30,57,29,204,31,250,31,29,31,169,31,35,31,134,31,56,31,151,31,177,31,177,30,228,31,115,31,153,31,51,31,40,31,239,31,239,30,63,31,216,31,216,30,1,31,187,31,204,31,4,31,229,31,64,31,64,30,93,31,158,31,60,31,138,31,134,31,7,31,82,31,82,30,137,31,137,30,137,29,33,31,99,31,99,30,99,29,75,31,53,31,225,31,225,30,204,31,171,31,77,31,153,31,29,31,162,31,48,31,248,31,19,31,82,31,151,31,218,31,218,30,138,31,183,31,151,31,72,31,82,31,213,31,203,31,23,31,251,31,27,31,70,31,211,31,186,31,227,31,227,30,227,29,85,31,165,31,48,31,120,31,228,31,125,31,125,30,249,31,235,31,235,30,235,29,201,31,49,31,189,31,128,31,190,31,194,31,252,31,126,31,255,31,17,31,17,30,17,29,114,31,169,31,154,31,151,31,173,31,173,30,12,31,41,31,119,31,119,30,219,31,178,31,14,31,7,31,10,31,33,31,221,31,18,31,120,31,26,31,166,31,130,31,120,31,57,31,153,31,162,31,129,31,126,31,79,31,79,30,79,29,192,31,192,30,57,31,57,30,57,29,99,31,6,31,229,31,173,31,45,31,45,30,201,31,161,31,197,31,197,30,197,29,12,31,15,31,15,30,107,31,109,31,176,31,196,31,152,31,152,30,80,31,252,31,107,31,190,31,183,31,183,30,170,31,90,31,78,31,11,31,170,31,184,31,184,30,220,31,114,31,237,31,40,31,40,30,213,31,168,31,37,31,149,31,255,31,212,31,63,31,146,31,23,31,23,30,23,29,249,31,33,31,33,30,33,29,173,31,173,30,135,31,135,30,249,31,78,31,213,31,130,31,79,31,221,31,221,30,67,31,248,31,15,31,16,31,16,30,42,31,161,31,220,31,220,30,198,31,198,30,198,29,135,31,110,31,142,31,77,31,145,31,189,31,190,31,50,31,50,30,131,31,131,30,5,31,166,31,17,31,77,31,44,31,200,31,200,30,106,31,77,31,40,31,62,31,217,31,255,31,172,31,202,31,121,31,125,31,55,31,20,31,20,30,156,31,224,31,224,30,98,31,98,30,98,29,203,31,116,31,140,31,42,31,168,31,155,31,168,31,104,31,24,31,66,31,66,30,4,31,167,31,122,31,188,31,9,31,131,31,26,31,26,30,11,31,55,31,98,31,156,31,172,31,172,30,143,31,201,31,159,31,57,31,57,30,97,31,28,31,167,31,71,31,71,30,71,29,213,31,78,31,78,30,78,29,101,31,53,31,51,31,174,31,36,31,48,31,97,31,150,31,211,31,211,30,211,29,162,31,7,31,235,31,235,30,103,31,121,31,3,31,223,31,218,31,35,31,168,31,168,30,168,29,127,31,230,31,127,31,163,31,81,31,94,31,33,31,33,30,100,31,70,31,170,31,86,31,109,31,95,31,190,31,188,31,188,30,81,31,81,30,88,31,175,31,7,31,162,31,174,31,113,31,245,31,4,31,150,31,133,31,153,31,23,31,77,31,108,31,25,31,76,31,76,31,81,31,28,31,28,30,57,31,71,31,171,31,171,30,107,31,106,31,117,31,138,31,204,31,146,31,201,31,14,31,90,31,143,31,209,31,209,30,46,31,51,31,187,31,112,31,56,31,182,31,73,31,165,31,239,31,255,31,255,30,163,31,39,31,58,31,225,31,194,31,56,31,70,31,161,31,75,31,108,31,204,31,204,30,41,31,30,31,25,31,74,31,30,31,131,31,131,30,88,31,12,31,107,31,145,31,86,31,245,31,48,31,234,31,196,31,236,31,246,31,246,30,254,31,112,31,112,30,112,29,101,31,84,31,52,31,100,31,181,31,149,31,149,30,53,31,204,31,204,30,233,31,107,31,221,31,84,31,197,31,18,31,18,30,18,29,67,31,177,31,54,31,139,31,11,31,171,31,24,31,62,31,28,31,125,31,125,30,27,31,41,31,73,31,170,31,157,31,98,31,19,31,173,31,173,30,95,31,100,31,22,31,22,30,29,31,234,31,47,31,10,31,179,31,241,31,11,31,11,30,198,31,31,31,31,30,35,31,35,30,32,31,70,31,74,31,112,31,45,31,60,31,70,31,20,31,20,30,75,31,75,30,125,31,24,31,24,30,168,31,168,30,11,31,163,31,125,31,140,31,140,30,177,31,98,31,173,31,135,31,205,31,230,31,21,31,63,31,63,30,236,31,107,31,107,30,24,31,71,31,180,31,150,31,18,31,144,31,243,31,230,31,247,31,58,31,198,31,52,31,52,30,38,31,126,31,113,31,26,31,235,31,183,31,179,31,120,31,221,31,187,31,127,31,86,31,211,31,122,31,106,31,199,31,199,30,77,31,144,31,10,31,146,31,115,31,162,31,50,31,127,31,116,31,201,31,205,31,205,30,129,31,129,30,68,31,108,31,108,30,108,29,251,31,22,31,22,30,105,31,91,31,179,31,86,31,16,31,180,31,166,31,80,31,49,31,239,31,73,31,197,31,118,31,252,31,206,31,126,31,248,31,180,31,31,31,13,31,67,31,162,31,162,30,220,31,54,31,59,31,234,31,59,31,250,31,74,31,74,30,94,31,44,31,85,31,179,31,87,31,107,31,107,30,39,31,52,31,52,30,52,29,97,31,86,31,249,31,172,31,33,31,33,30,179,31,179,30,154,31,137,31,112,31,66,31,33,31,108,31,108,30,108,29,245,31,229,31,79,31,255,31,224,31,65,31,133,31,91,31,66,31,206,31,116,31,68,31,29,31,105,31,24,31,99,31,51,31,51,30,226,31,137,31,120,31,161,31,6,31,203,31,189,31,189,30,189,29,98,31,52,31,212,31,221,31,46,31,166,31,166,30,51,31,51,30,51,29,51,28,51,27,25,31,139,31,161,31,27,31,55,31,241,31,31,31,31,30,39,31,119,31,119,30,187,31,212,31,186,31,224,31,255,31,134,31,21,31,85,31,25,31,146,31,79,31,62,31,203,31,255,31,255,30,23,31,158,31,161,31,23,31,23,30,23,29,97,31,26,31,190,31,190,30,211,31,80,31,80,30,189,31,210,31,226,31,174,31,67,31,127,31,127,30,182,31,182,30,166,31,166,30,175,31,65,31,89,31,245,31,5,31,5,30,102,31,8,31,248,31,248,30,251,31,20,31,20,30,7,31,220,31,220,30,88,31,44,31,142,31,18,31,247,31,175,31,70,31,21,31,242,31,242,30,163,31,99,31,5,31,56,31,209,31,209,30,1,31,1,30,125,31,112,31,112,30,160,31,182,31,212,31,224,31,181,31,121,31,121,30,34,31,30,31,30,30,77,31,77,30,209,31,96,31,145,31,199,31,61,31,167,31,167,30,167,29,239,31,169,31,112,31,112,30,72,31,2,31,104,31,255,31,58,31,58,30,74,31,159,31,150,31,67,31,89,31,149,31,33,31,230,31,113,31,248,31,248,30,62,31,174,31,103,31,8,31,70,31,155,31,34,31,1,31,252,31,54,31,249,31,126,31,46,31,2,31,23,31,23,30,23,29,45,31,4,31,163,31,51,31,51,30,31,31,52,31,40,31,170,31,65,31,90,31,173,31,249,31,234,31,138,31,138,30,138,29,69,31,115,31,119,31,119,30,118,31,187,31,247,31,247,30,85,31,85,30,85,29,85,28,85,27,28,31,84,31,84,30,25,31,145,31,145,30,179,31,114,31,114,30,174,31,118,31,5,31,5,30,153,31,179,31,9,31,9,30,179,31,176,31,107,31,46,31,46,30,246,31,246,30,120,31,122,31,100,31,168,31,99,31,8,31,8,30,172,31,233,31,235,31,220,31,212,31,253,31,205,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
