-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 346;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (251,0,148,0,17,0,0,0,181,0,0,0,42,0,0,0,190,0,119,0,74,0,0,0,161,0,9,0,25,0,24,0,197,0,52,0,183,0,230,0,0,0,200,0,78,0,0,0,30,0,0,0,22,0,20,0,0,0,53,0,184,0,191,0,0,0,58,0,211,0,92,0,0,0,43,0,89,0,190,0,0,0,66,0,0,0,255,0,221,0,221,0,50,0,0,0,246,0,135,0,36,0,0,0,209,0,210,0,0,0,251,0,162,0,197,0,207,0,213,0,14,0,34,0,138,0,10,0,0,0,0,0,178,0,78,0,142,0,43,0,176,0,255,0,60,0,173,0,69,0,143,0,0,0,109,0,0,0,255,0,178,0,241,0,204,0,253,0,133,0,36,0,12,0,110,0,0,0,0,0,136,0,68,0,168,0,167,0,100,0,167,0,90,0,121,0,0,0,36,0,36,0,86,0,46,0,121,0,35,0,228,0,208,0,239,0,49,0,152,0,131,0,63,0,59,0,67,0,0,0,61,0,192,0,171,0,205,0,0,0,0,0,119,0,227,0,254,0,19,0,163,0,59,0,107,0,93,0,183,0,128,0,214,0,140,0,252,0,169,0,191,0,31,0,193,0,0,0,0,0,2,0,130,0,238,0,131,0,0,0,137,0,83,0,174,0,99,0,187,0,0,0,49,0,98,0,9,0,0,0,149,0,45,0,197,0,227,0,161,0,93,0,0,0,184,0,212,0,0,0,121,0,125,0,124,0,0,0,28,0,171,0,28,0,205,0,155,0,108,0,214,0,38,0,214,0,133,0,82,0,47,0,27,0,185,0,46,0,0,0,168,0,0,0,94,0,202,0,148,0,229,0,16,0,0,0,186,0,0,0,158,0,169,0,170,0,25,0,137,0,11,0,68,0,0,0,119,0,20,0,0,0,139,0,153,0,176,0,106,0,60,0,126,0,31,0,159,0,108,0,87,0,182,0,47,0,64,0,42,0,0,0,161,0,197,0,243,0,110,0,146,0,25,0,74,0,86,0,23,0,0,0,9,0,0,0,167,0,191,0,215,0,0,0,79,0,162,0,100,0,191,0,119,0,88,0,96,0,230,0,0,0,37,0,101,0,49,0,84,0,239,0,83,0,2,0,227,0,0,0,245,0,10,0,54,0,124,0,96,0,27,0,133,0,19,0,71,0,155,0,59,0,2,0,0,0,217,0,186,0,100,0,76,0,48,0,176,0,0,0,6,0,180,0,144,0,141,0,79,0,141,0,90,0,243,0,196,0,164,0,119,0,7,0,103,0,114,0,55,0,178,0,240,0,104,0,142,0,219,0,216,0,90,0,92,0,185,0,0,0,77,0,0,0,36,0,64,0,180,0,87,0,124,0,219,0,184,0,25,0,214,0,185,0,0,0,84,0,10,0,64,0,153,0,185,0,247,0,0,0,229,0,181,0,205,0,0,0,82,0,90,0,0,0,217,0,187,0,116,0,0,0,125,0,100,0,0,0,169,0,81,0,198,0,124,0,70,0,108,0,83,0,246,0,86,0,165,0,216,0,0,0);
signal scenario_full  : scenario_type := (251,31,148,31,17,31,17,30,181,31,181,30,42,31,42,30,190,31,119,31,74,31,74,30,161,31,9,31,25,31,24,31,197,31,52,31,183,31,230,31,230,30,200,31,78,31,78,30,30,31,30,30,22,31,20,31,20,30,53,31,184,31,191,31,191,30,58,31,211,31,92,31,92,30,43,31,89,31,190,31,190,30,66,31,66,30,255,31,221,31,221,31,50,31,50,30,246,31,135,31,36,31,36,30,209,31,210,31,210,30,251,31,162,31,197,31,207,31,213,31,14,31,34,31,138,31,10,31,10,30,10,29,178,31,78,31,142,31,43,31,176,31,255,31,60,31,173,31,69,31,143,31,143,30,109,31,109,30,255,31,178,31,241,31,204,31,253,31,133,31,36,31,12,31,110,31,110,30,110,29,136,31,68,31,168,31,167,31,100,31,167,31,90,31,121,31,121,30,36,31,36,31,86,31,46,31,121,31,35,31,228,31,208,31,239,31,49,31,152,31,131,31,63,31,59,31,67,31,67,30,61,31,192,31,171,31,205,31,205,30,205,29,119,31,227,31,254,31,19,31,163,31,59,31,107,31,93,31,183,31,128,31,214,31,140,31,252,31,169,31,191,31,31,31,193,31,193,30,193,29,2,31,130,31,238,31,131,31,131,30,137,31,83,31,174,31,99,31,187,31,187,30,49,31,98,31,9,31,9,30,149,31,45,31,197,31,227,31,161,31,93,31,93,30,184,31,212,31,212,30,121,31,125,31,124,31,124,30,28,31,171,31,28,31,205,31,155,31,108,31,214,31,38,31,214,31,133,31,82,31,47,31,27,31,185,31,46,31,46,30,168,31,168,30,94,31,202,31,148,31,229,31,16,31,16,30,186,31,186,30,158,31,169,31,170,31,25,31,137,31,11,31,68,31,68,30,119,31,20,31,20,30,139,31,153,31,176,31,106,31,60,31,126,31,31,31,159,31,108,31,87,31,182,31,47,31,64,31,42,31,42,30,161,31,197,31,243,31,110,31,146,31,25,31,74,31,86,31,23,31,23,30,9,31,9,30,167,31,191,31,215,31,215,30,79,31,162,31,100,31,191,31,119,31,88,31,96,31,230,31,230,30,37,31,101,31,49,31,84,31,239,31,83,31,2,31,227,31,227,30,245,31,10,31,54,31,124,31,96,31,27,31,133,31,19,31,71,31,155,31,59,31,2,31,2,30,217,31,186,31,100,31,76,31,48,31,176,31,176,30,6,31,180,31,144,31,141,31,79,31,141,31,90,31,243,31,196,31,164,31,119,31,7,31,103,31,114,31,55,31,178,31,240,31,104,31,142,31,219,31,216,31,90,31,92,31,185,31,185,30,77,31,77,30,36,31,64,31,180,31,87,31,124,31,219,31,184,31,25,31,214,31,185,31,185,30,84,31,10,31,64,31,153,31,185,31,247,31,247,30,229,31,181,31,205,31,205,30,82,31,90,31,90,30,217,31,187,31,116,31,116,30,125,31,100,31,100,30,169,31,81,31,198,31,124,31,70,31,108,31,83,31,246,31,86,31,165,31,216,31,216,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
