-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 181;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (204,0,0,0,0,0,0,0,140,0,112,0,165,0,216,0,107,0,172,0,124,0,14,0,236,0,172,0,67,0,183,0,0,0,167,0,96,0,0,0,137,0,204,0,134,0,86,0,0,0,208,0,247,0,34,0,178,0,0,0,148,0,123,0,130,0,199,0,105,0,249,0,251,0,53,0,188,0,165,0,253,0,46,0,224,0,0,0,155,0,134,0,38,0,123,0,252,0,146,0,47,0,183,0,174,0,245,0,0,0,252,0,106,0,0,0,205,0,46,0,28,0,164,0,226,0,88,0,48,0,58,0,178,0,133,0,216,0,27,0,0,0,133,0,249,0,8,0,0,0,0,0,244,0,107,0,0,0,16,0,0,0,0,0,0,0,24,0,0,0,43,0,240,0,189,0,222,0,0,0,14,0,0,0,60,0,0,0,81,0,74,0,217,0,28,0,184,0,140,0,245,0,146,0,237,0,118,0,216,0,154,0,151,0,0,0,0,0,205,0,0,0,38,0,75,0,184,0,0,0,48,0,145,0,197,0,141,0,139,0,133,0,56,0,112,0,243,0,217,0,248,0,213,0,62,0,0,0,246,0,0,0,194,0,54,0,32,0,212,0,109,0,197,0,171,0,147,0,211,0,179,0,86,0,25,0,48,0,0,0,210,0,254,0,0,0,102,0,221,0,105,0,0,0,0,0,212,0,8,0,0,0,242,0,0,0,16,0,49,0,105,0,19,0,191,0,32,0,122,0,214,0,20,0,0,0,53,0,124,0,0,0,160,0,116,0,0,0,204,0,199,0,250,0,42,0,0,0,115,0,253,0);
signal scenario_full  : scenario_type := (204,31,204,30,204,29,204,28,140,31,112,31,165,31,216,31,107,31,172,31,124,31,14,31,236,31,172,31,67,31,183,31,183,30,167,31,96,31,96,30,137,31,204,31,134,31,86,31,86,30,208,31,247,31,34,31,178,31,178,30,148,31,123,31,130,31,199,31,105,31,249,31,251,31,53,31,188,31,165,31,253,31,46,31,224,31,224,30,155,31,134,31,38,31,123,31,252,31,146,31,47,31,183,31,174,31,245,31,245,30,252,31,106,31,106,30,205,31,46,31,28,31,164,31,226,31,88,31,48,31,58,31,178,31,133,31,216,31,27,31,27,30,133,31,249,31,8,31,8,30,8,29,244,31,107,31,107,30,16,31,16,30,16,29,16,28,24,31,24,30,43,31,240,31,189,31,222,31,222,30,14,31,14,30,60,31,60,30,81,31,74,31,217,31,28,31,184,31,140,31,245,31,146,31,237,31,118,31,216,31,154,31,151,31,151,30,151,29,205,31,205,30,38,31,75,31,184,31,184,30,48,31,145,31,197,31,141,31,139,31,133,31,56,31,112,31,243,31,217,31,248,31,213,31,62,31,62,30,246,31,246,30,194,31,54,31,32,31,212,31,109,31,197,31,171,31,147,31,211,31,179,31,86,31,25,31,48,31,48,30,210,31,254,31,254,30,102,31,221,31,105,31,105,30,105,29,212,31,8,31,8,30,242,31,242,30,16,31,49,31,105,31,19,31,191,31,32,31,122,31,214,31,20,31,20,30,53,31,124,31,124,30,160,31,116,31,116,30,204,31,199,31,250,31,42,31,42,30,115,31,253,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
