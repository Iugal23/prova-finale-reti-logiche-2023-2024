-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 642;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (15,0,163,0,175,0,0,0,74,0,202,0,191,0,32,0,95,0,0,0,181,0,159,0,103,0,1,0,251,0,61,0,64,0,90,0,235,0,0,0,37,0,190,0,205,0,50,0,119,0,0,0,0,0,209,0,243,0,246,0,39,0,5,0,135,0,0,0,57,0,0,0,30,0,0,0,0,0,165,0,116,0,0,0,197,0,65,0,57,0,164,0,85,0,206,0,33,0,113,0,39,0,0,0,58,0,0,0,118,0,71,0,80,0,212,0,82,0,125,0,240,0,0,0,110,0,139,0,0,0,100,0,29,0,199,0,15,0,216,0,119,0,137,0,240,0,219,0,4,0,230,0,103,0,232,0,177,0,93,0,0,0,131,0,0,0,0,0,79,0,134,0,0,0,0,0,159,0,25,0,193,0,0,0,174,0,186,0,37,0,0,0,79,0,167,0,52,0,121,0,0,0,0,0,11,0,173,0,226,0,230,0,0,0,18,0,164,0,145,0,57,0,234,0,3,0,0,0,0,0,173,0,1,0,75,0,0,0,104,0,101,0,0,0,41,0,0,0,0,0,173,0,59,0,61,0,0,0,150,0,62,0,120,0,0,0,175,0,0,0,53,0,108,0,183,0,0,0,0,0,202,0,0,0,168,0,0,0,23,0,0,0,89,0,0,0,144,0,0,0,222,0,120,0,210,0,191,0,174,0,243,0,132,0,243,0,87,0,126,0,89,0,11,0,0,0,81,0,164,0,88,0,240,0,224,0,0,0,80,0,167,0,177,0,0,0,238,0,94,0,29,0,252,0,0,0,144,0,182,0,211,0,162,0,79,0,253,0,0,0,1,0,255,0,220,0,64,0,103,0,118,0,198,0,11,0,17,0,0,0,139,0,14,0,233,0,160,0,217,0,220,0,57,0,230,0,0,0,208,0,225,0,51,0,234,0,104,0,0,0,171,0,30,0,0,0,121,0,246,0,13,0,182,0,178,0,133,0,171,0,180,0,240,0,243,0,0,0,0,0,0,0,117,0,179,0,140,0,155,0,0,0,0,0,206,0,129,0,252,0,0,0,0,0,182,0,174,0,213,0,0,0,202,0,55,0,0,0,27,0,234,0,85,0,0,0,88,0,144,0,191,0,113,0,0,0,8,0,75,0,242,0,48,0,94,0,193,0,177,0,0,0,102,0,109,0,155,0,0,0,3,0,77,0,0,0,0,0,30,0,178,0,187,0,152,0,44,0,233,0,152,0,232,0,0,0,0,0,242,0,0,0,250,0,0,0,25,0,233,0,27,0,52,0,43,0,0,0,17,0,52,0,159,0,211,0,211,0,119,0,0,0,63,0,60,0,159,0,214,0,64,0,13,0,163,0,66,0,207,0,9,0,138,0,143,0,62,0,53,0,106,0,20,0,173,0,194,0,0,0,147,0,0,0,0,0,0,0,186,0,226,0,0,0,237,0,164,0,180,0,205,0,237,0,240,0,90,0,71,0,0,0,254,0,0,0,216,0,181,0,41,0,33,0,94,0,128,0,62,0,124,0,128,0,158,0,224,0,0,0,188,0,111,0,127,0,86,0,208,0,0,0,183,0,0,0,0,0,179,0,105,0,142,0,239,0,0,0,0,0,69,0,0,0,93,0,0,0,174,0,103,0,235,0,50,0,116,0,48,0,21,0,16,0,182,0,95,0,61,0,134,0,173,0,64,0,65,0,0,0,245,0,0,0,88,0,213,0,249,0,17,0,110,0,247,0,217,0,138,0,170,0,229,0,0,0,70,0,128,0,78,0,159,0,241,0,40,0,91,0,166,0,200,0,168,0,0,0,136,0,43,0,121,0,188,0,117,0,0,0,54,0,245,0,196,0,253,0,11,0,135,0,7,0,197,0,84,0,252,0,26,0,145,0,0,0,79,0,193,0,44,0,198,0,238,0,33,0,72,0,221,0,4,0,136,0,156,0,65,0,0,0,0,0,231,0,72,0,254,0,0,0,21,0,0,0,0,0,204,0,24,0,0,0,198,0,0,0,95,0,104,0,212,0,113,0,72,0,59,0,123,0,25,0,39,0,55,0,0,0,213,0,132,0,225,0,217,0,53,0,205,0,46,0,32,0,112,0,0,0,183,0,26,0,25,0,165,0,84,0,0,0,0,0,0,0,0,0,9,0,0,0,219,0,205,0,0,0,0,0,62,0,0,0,123,0,0,0,65,0,15,0,84,0,0,0,17,0,242,0,46,0,0,0,190,0,198,0,0,0,156,0,0,0,217,0,82,0,0,0,0,0,0,0,193,0,10,0,111,0,160,0,38,0,216,0,210,0,127,0,73,0,189,0,81,0,213,0,247,0,7,0,91,0,58,0,241,0,237,0,185,0,0,0,49,0,43,0,96,0,120,0,0,0,57,0,0,0,0,0,47,0,0,0,249,0,154,0,244,0,89,0,156,0,213,0,40,0,104,0,125,0,139,0,220,0,154,0,228,0,0,0,173,0,57,0,86,0,155,0,0,0,56,0,228,0,86,0,120,0,52,0,1,0,31,0,166,0,0,0,233,0,72,0,199,0,182,0,38,0,0,0,104,0,49,0,40,0,162,0,124,0,203,0,179,0,242,0,0,0,155,0,0,0,217,0,0,0,0,0,0,0,93,0,238,0,0,0,19,0,0,0,3,0,0,0,203,0,79,0,202,0,242,0,198,0,148,0,0,0,31,0,199,0,147,0,124,0,67,0,0,0,0,0,159,0,89,0,248,0,130,0,11,0,139,0,0,0,0,0,207,0,154,0,57,0,118,0,92,0,57,0,1,0,87,0,0,0,157,0,0,0,0,0,146,0,226,0,0,0,48,0,156,0,249,0,153,0,8,0,193,0,99,0,170,0,49,0,0,0,0,0,106,0);
signal scenario_full  : scenario_type := (15,31,163,31,175,31,175,30,74,31,202,31,191,31,32,31,95,31,95,30,181,31,159,31,103,31,1,31,251,31,61,31,64,31,90,31,235,31,235,30,37,31,190,31,205,31,50,31,119,31,119,30,119,29,209,31,243,31,246,31,39,31,5,31,135,31,135,30,57,31,57,30,30,31,30,30,30,29,165,31,116,31,116,30,197,31,65,31,57,31,164,31,85,31,206,31,33,31,113,31,39,31,39,30,58,31,58,30,118,31,71,31,80,31,212,31,82,31,125,31,240,31,240,30,110,31,139,31,139,30,100,31,29,31,199,31,15,31,216,31,119,31,137,31,240,31,219,31,4,31,230,31,103,31,232,31,177,31,93,31,93,30,131,31,131,30,131,29,79,31,134,31,134,30,134,29,159,31,25,31,193,31,193,30,174,31,186,31,37,31,37,30,79,31,167,31,52,31,121,31,121,30,121,29,11,31,173,31,226,31,230,31,230,30,18,31,164,31,145,31,57,31,234,31,3,31,3,30,3,29,173,31,1,31,75,31,75,30,104,31,101,31,101,30,41,31,41,30,41,29,173,31,59,31,61,31,61,30,150,31,62,31,120,31,120,30,175,31,175,30,53,31,108,31,183,31,183,30,183,29,202,31,202,30,168,31,168,30,23,31,23,30,89,31,89,30,144,31,144,30,222,31,120,31,210,31,191,31,174,31,243,31,132,31,243,31,87,31,126,31,89,31,11,31,11,30,81,31,164,31,88,31,240,31,224,31,224,30,80,31,167,31,177,31,177,30,238,31,94,31,29,31,252,31,252,30,144,31,182,31,211,31,162,31,79,31,253,31,253,30,1,31,255,31,220,31,64,31,103,31,118,31,198,31,11,31,17,31,17,30,139,31,14,31,233,31,160,31,217,31,220,31,57,31,230,31,230,30,208,31,225,31,51,31,234,31,104,31,104,30,171,31,30,31,30,30,121,31,246,31,13,31,182,31,178,31,133,31,171,31,180,31,240,31,243,31,243,30,243,29,243,28,117,31,179,31,140,31,155,31,155,30,155,29,206,31,129,31,252,31,252,30,252,29,182,31,174,31,213,31,213,30,202,31,55,31,55,30,27,31,234,31,85,31,85,30,88,31,144,31,191,31,113,31,113,30,8,31,75,31,242,31,48,31,94,31,193,31,177,31,177,30,102,31,109,31,155,31,155,30,3,31,77,31,77,30,77,29,30,31,178,31,187,31,152,31,44,31,233,31,152,31,232,31,232,30,232,29,242,31,242,30,250,31,250,30,25,31,233,31,27,31,52,31,43,31,43,30,17,31,52,31,159,31,211,31,211,31,119,31,119,30,63,31,60,31,159,31,214,31,64,31,13,31,163,31,66,31,207,31,9,31,138,31,143,31,62,31,53,31,106,31,20,31,173,31,194,31,194,30,147,31,147,30,147,29,147,28,186,31,226,31,226,30,237,31,164,31,180,31,205,31,237,31,240,31,90,31,71,31,71,30,254,31,254,30,216,31,181,31,41,31,33,31,94,31,128,31,62,31,124,31,128,31,158,31,224,31,224,30,188,31,111,31,127,31,86,31,208,31,208,30,183,31,183,30,183,29,179,31,105,31,142,31,239,31,239,30,239,29,69,31,69,30,93,31,93,30,174,31,103,31,235,31,50,31,116,31,48,31,21,31,16,31,182,31,95,31,61,31,134,31,173,31,64,31,65,31,65,30,245,31,245,30,88,31,213,31,249,31,17,31,110,31,247,31,217,31,138,31,170,31,229,31,229,30,70,31,128,31,78,31,159,31,241,31,40,31,91,31,166,31,200,31,168,31,168,30,136,31,43,31,121,31,188,31,117,31,117,30,54,31,245,31,196,31,253,31,11,31,135,31,7,31,197,31,84,31,252,31,26,31,145,31,145,30,79,31,193,31,44,31,198,31,238,31,33,31,72,31,221,31,4,31,136,31,156,31,65,31,65,30,65,29,231,31,72,31,254,31,254,30,21,31,21,30,21,29,204,31,24,31,24,30,198,31,198,30,95,31,104,31,212,31,113,31,72,31,59,31,123,31,25,31,39,31,55,31,55,30,213,31,132,31,225,31,217,31,53,31,205,31,46,31,32,31,112,31,112,30,183,31,26,31,25,31,165,31,84,31,84,30,84,29,84,28,84,27,9,31,9,30,219,31,205,31,205,30,205,29,62,31,62,30,123,31,123,30,65,31,15,31,84,31,84,30,17,31,242,31,46,31,46,30,190,31,198,31,198,30,156,31,156,30,217,31,82,31,82,30,82,29,82,28,193,31,10,31,111,31,160,31,38,31,216,31,210,31,127,31,73,31,189,31,81,31,213,31,247,31,7,31,91,31,58,31,241,31,237,31,185,31,185,30,49,31,43,31,96,31,120,31,120,30,57,31,57,30,57,29,47,31,47,30,249,31,154,31,244,31,89,31,156,31,213,31,40,31,104,31,125,31,139,31,220,31,154,31,228,31,228,30,173,31,57,31,86,31,155,31,155,30,56,31,228,31,86,31,120,31,52,31,1,31,31,31,166,31,166,30,233,31,72,31,199,31,182,31,38,31,38,30,104,31,49,31,40,31,162,31,124,31,203,31,179,31,242,31,242,30,155,31,155,30,217,31,217,30,217,29,217,28,93,31,238,31,238,30,19,31,19,30,3,31,3,30,203,31,79,31,202,31,242,31,198,31,148,31,148,30,31,31,199,31,147,31,124,31,67,31,67,30,67,29,159,31,89,31,248,31,130,31,11,31,139,31,139,30,139,29,207,31,154,31,57,31,118,31,92,31,57,31,1,31,87,31,87,30,157,31,157,30,157,29,146,31,226,31,226,30,48,31,156,31,249,31,153,31,8,31,193,31,99,31,170,31,49,31,49,30,49,29,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
