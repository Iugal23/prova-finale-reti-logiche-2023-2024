-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_197 is
end project_tb_197;

architecture project_tb_arch_197 of project_tb_197 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 879;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,64,0,208,0,86,0,0,0,138,0,0,0,84,0,221,0,29,0,190,0,26,0,30,0,120,0,0,0,48,0,88,0,182,0,4,0,172,0,237,0,229,0,101,0,140,0,240,0,53,0,0,0,162,0,206,0,0,0,0,0,0,0,60,0,69,0,250,0,88,0,28,0,37,0,43,0,196,0,20,0,18,0,133,0,101,0,236,0,221,0,12,0,218,0,0,0,171,0,210,0,26,0,110,0,0,0,205,0,0,0,179,0,106,0,0,0,93,0,253,0,216,0,0,0,179,0,23,0,6,0,233,0,56,0,104,0,0,0,150,0,109,0,78,0,91,0,6,0,5,0,83,0,0,0,219,0,0,0,61,0,40,0,210,0,219,0,165,0,60,0,0,0,225,0,42,0,243,0,50,0,103,0,0,0,163,0,201,0,207,0,0,0,84,0,155,0,253,0,164,0,41,0,141,0,0,0,53,0,135,0,0,0,83,0,0,0,32,0,150,0,153,0,0,0,0,0,0,0,69,0,0,0,192,0,68,0,202,0,0,0,0,0,45,0,239,0,238,0,199,0,1,0,203,0,0,0,62,0,0,0,235,0,27,0,0,0,0,0,0,0,99,0,191,0,140,0,10,0,199,0,0,0,246,0,116,0,202,0,135,0,0,0,0,0,174,0,0,0,139,0,78,0,248,0,102,0,199,0,64,0,89,0,251,0,176,0,234,0,46,0,187,0,250,0,118,0,57,0,183,0,132,0,245,0,255,0,131,0,83,0,0,0,67,0,180,0,44,0,91,0,248,0,128,0,89,0,245,0,211,0,171,0,29,0,226,0,237,0,235,0,237,0,115,0,105,0,98,0,220,0,96,0,101,0,113,0,193,0,152,0,166,0,40,0,0,0,109,0,0,0,198,0,199,0,0,0,49,0,161,0,148,0,207,0,0,0,246,0,39,0,77,0,84,0,77,0,103,0,251,0,22,0,0,0,74,0,80,0,62,0,238,0,6,0,68,0,0,0,230,0,163,0,243,0,249,0,246,0,176,0,74,0,44,0,66,0,196,0,215,0,166,0,240,0,0,0,0,0,230,0,123,0,164,0,114,0,0,0,193,0,0,0,128,0,75,0,238,0,113,0,143,0,90,0,184,0,94,0,200,0,91,0,0,0,247,0,51,0,0,0,131,0,184,0,121,0,133,0,151,0,2,0,0,0,240,0,106,0,248,0,105,0,127,0,43,0,166,0,0,0,213,0,45,0,0,0,68,0,177,0,137,0,62,0,108,0,194,0,166,0,134,0,135,0,245,0,101,0,0,0,118,0,168,0,0,0,0,0,169,0,217,0,0,0,27,0,161,0,1,0,101,0,0,0,165,0,233,0,140,0,37,0,77,0,90,0,200,0,69,0,85,0,83,0,0,0,0,0,119,0,147,0,167,0,0,0,182,0,221,0,190,0,123,0,83,0,151,0,15,0,0,0,196,0,204,0,80,0,70,0,249,0,0,0,86,0,0,0,0,0,111,0,187,0,228,0,0,0,248,0,71,0,240,0,41,0,143,0,201,0,238,0,108,0,0,0,0,0,148,0,0,0,36,0,44,0,41,0,125,0,73,0,101,0,42,0,197,0,113,0,255,0,220,0,158,0,0,0,213,0,46,0,119,0,73,0,0,0,0,0,109,0,80,0,15,0,0,0,215,0,0,0,0,0,0,0,111,0,71,0,20,0,112,0,0,0,60,0,16,0,232,0,202,0,0,0,0,0,50,0,139,0,0,0,75,0,0,0,247,0,190,0,132,0,132,0,224,0,20,0,173,0,236,0,22,0,0,0,214,0,29,0,29,0,125,0,55,0,126,0,175,0,39,0,199,0,17,0,245,0,138,0,79,0,134,0,59,0,129,0,0,0,122,0,0,0,141,0,112,0,145,0,0,0,233,0,0,0,0,0,0,0,1,0,251,0,134,0,65,0,87,0,99,0,192,0,0,0,137,0,20,0,51,0,197,0,120,0,61,0,60,0,85,0,233,0,230,0,243,0,107,0,84,0,139,0,0,0,201,0,45,0,132,0,129,0,194,0,0,0,130,0,41,0,5,0,191,0,98,0,0,0,145,0,212,0,0,0,0,0,57,0,255,0,85,0,94,0,194,0,0,0,60,0,32,0,20,0,149,0,0,0,184,0,132,0,204,0,215,0,70,0,136,0,0,0,7,0,33,0,64,0,149,0,206,0,82,0,179,0,185,0,0,0,0,0,225,0,62,0,142,0,131,0,210,0,234,0,245,0,0,0,148,0,0,0,149,0,36,0,0,0,254,0,132,0,200,0,241,0,0,0,187,0,47,0,0,0,51,0,0,0,94,0,0,0,196,0,141,0,194,0,0,0,0,0,0,0,0,0,0,0,0,0,201,0,0,0,104,0,40,0,172,0,134,0,229,0,82,0,218,0,68,0,0,0,169,0,40,0,105,0,89,0,98,0,195,0,150,0,226,0,0,0,141,0,254,0,78,0,220,0,86,0,206,0,90,0,0,0,47,0,0,0,82,0,173,0,178,0,150,0,223,0,57,0,115,0,0,0,127,0,10,0,12,0,0,0,80,0,244,0,0,0,65,0,88,0,224,0,201,0,10,0,15,0,235,0,218,0,0,0,0,0,149,0,57,0,0,0,0,0,0,0,83,0,86,0,102,0,51,0,96,0,236,0,0,0,0,0,139,0,229,0,0,0,32,0,0,0,90,0,27,0,50,0,0,0,62,0,191,0,124,0,52,0,157,0,189,0,136,0,236,0,0,0,184,0,91,0,0,0,0,0,159,0,0,0,13,0,163,0,124,0,0,0,12,0,0,0,54,0,107,0,54,0,156,0,0,0,0,0,0,0,28,0,24,0,252,0,120,0,206,0,0,0,0,0,99,0,77,0,95,0,227,0,193,0,65,0,126,0,40,0,18,0,228,0,34,0,169,0,0,0,209,0,156,0,0,0,142,0,41,0,179,0,65,0,222,0,7,0,165,0,113,0,159,0,236,0,150,0,195,0,0,0,5,0,140,0,70,0,26,0,158,0,52,0,17,0,98,0,243,0,66,0,154,0,0,0,115,0,152,0,47,0,0,0,150,0,136,0,0,0,0,0,2,0,166,0,116,0,152,0,186,0,141,0,131,0,124,0,71,0,223,0,4,0,120,0,2,0,225,0,246,0,208,0,172,0,237,0,193,0,31,0,0,0,107,0,122,0,126,0,226,0,168,0,152,0,99,0,0,0,216,0,183,0,0,0,0,0,70,0,251,0,254,0,56,0,0,0,0,0,51,0,98,0,220,0,0,0,62,0,230,0,0,0,105,0,29,0,105,0,0,0,71,0,0,0,188,0,0,0,157,0,69,0,71,0,181,0,0,0,144,0,151,0,173,0,135,0,93,0,203,0,25,0,152,0,115,0,252,0,179,0,87,0,195,0,136,0,92,0,0,0,162,0,0,0,58,0,3,0,116,0,3,0,168,0,62,0,194,0,140,0,234,0,35,0,36,0,234,0,75,0,103,0,253,0,0,0,101,0,58,0,0,0,113,0,223,0,171,0,0,0,93,0,63,0,117,0,182,0,255,0,130,0,11,0,98,0,184,0,222,0,44,0,129,0,39,0,206,0,123,0,43,0,201,0,103,0,199,0,216,0,138,0,134,0,137,0,28,0,15,0,64,0,122,0,216,0,0,0,119,0,73,0,31,0,110,0,132,0,178,0,0,0,31,0,28,0,57,0,166,0,107,0,50,0,132,0,117,0,168,0,43,0,0,0,233,0,254,0,155,0,134,0,25,0,36,0,147,0,0,0,3,0,113,0,0,0,223,0,205,0,0,0,190,0,0,0,254,0,92,0,0,0,0,0,238,0,79,0,221,0,134,0,106,0,0,0,0,0,0,0,18,0,234,0,125,0,58,0,175,0,187,0,12,0,233,0,44,0);
signal scenario_full  : scenario_type := (0,0,0,0,64,31,208,31,86,31,86,30,138,31,138,30,84,31,221,31,29,31,190,31,26,31,30,31,120,31,120,30,48,31,88,31,182,31,4,31,172,31,237,31,229,31,101,31,140,31,240,31,53,31,53,30,162,31,206,31,206,30,206,29,206,28,60,31,69,31,250,31,88,31,28,31,37,31,43,31,196,31,20,31,18,31,133,31,101,31,236,31,221,31,12,31,218,31,218,30,171,31,210,31,26,31,110,31,110,30,205,31,205,30,179,31,106,31,106,30,93,31,253,31,216,31,216,30,179,31,23,31,6,31,233,31,56,31,104,31,104,30,150,31,109,31,78,31,91,31,6,31,5,31,83,31,83,30,219,31,219,30,61,31,40,31,210,31,219,31,165,31,60,31,60,30,225,31,42,31,243,31,50,31,103,31,103,30,163,31,201,31,207,31,207,30,84,31,155,31,253,31,164,31,41,31,141,31,141,30,53,31,135,31,135,30,83,31,83,30,32,31,150,31,153,31,153,30,153,29,153,28,69,31,69,30,192,31,68,31,202,31,202,30,202,29,45,31,239,31,238,31,199,31,1,31,203,31,203,30,62,31,62,30,235,31,27,31,27,30,27,29,27,28,99,31,191,31,140,31,10,31,199,31,199,30,246,31,116,31,202,31,135,31,135,30,135,29,174,31,174,30,139,31,78,31,248,31,102,31,199,31,64,31,89,31,251,31,176,31,234,31,46,31,187,31,250,31,118,31,57,31,183,31,132,31,245,31,255,31,131,31,83,31,83,30,67,31,180,31,44,31,91,31,248,31,128,31,89,31,245,31,211,31,171,31,29,31,226,31,237,31,235,31,237,31,115,31,105,31,98,31,220,31,96,31,101,31,113,31,193,31,152,31,166,31,40,31,40,30,109,31,109,30,198,31,199,31,199,30,49,31,161,31,148,31,207,31,207,30,246,31,39,31,77,31,84,31,77,31,103,31,251,31,22,31,22,30,74,31,80,31,62,31,238,31,6,31,68,31,68,30,230,31,163,31,243,31,249,31,246,31,176,31,74,31,44,31,66,31,196,31,215,31,166,31,240,31,240,30,240,29,230,31,123,31,164,31,114,31,114,30,193,31,193,30,128,31,75,31,238,31,113,31,143,31,90,31,184,31,94,31,200,31,91,31,91,30,247,31,51,31,51,30,131,31,184,31,121,31,133,31,151,31,2,31,2,30,240,31,106,31,248,31,105,31,127,31,43,31,166,31,166,30,213,31,45,31,45,30,68,31,177,31,137,31,62,31,108,31,194,31,166,31,134,31,135,31,245,31,101,31,101,30,118,31,168,31,168,30,168,29,169,31,217,31,217,30,27,31,161,31,1,31,101,31,101,30,165,31,233,31,140,31,37,31,77,31,90,31,200,31,69,31,85,31,83,31,83,30,83,29,119,31,147,31,167,31,167,30,182,31,221,31,190,31,123,31,83,31,151,31,15,31,15,30,196,31,204,31,80,31,70,31,249,31,249,30,86,31,86,30,86,29,111,31,187,31,228,31,228,30,248,31,71,31,240,31,41,31,143,31,201,31,238,31,108,31,108,30,108,29,148,31,148,30,36,31,44,31,41,31,125,31,73,31,101,31,42,31,197,31,113,31,255,31,220,31,158,31,158,30,213,31,46,31,119,31,73,31,73,30,73,29,109,31,80,31,15,31,15,30,215,31,215,30,215,29,215,28,111,31,71,31,20,31,112,31,112,30,60,31,16,31,232,31,202,31,202,30,202,29,50,31,139,31,139,30,75,31,75,30,247,31,190,31,132,31,132,31,224,31,20,31,173,31,236,31,22,31,22,30,214,31,29,31,29,31,125,31,55,31,126,31,175,31,39,31,199,31,17,31,245,31,138,31,79,31,134,31,59,31,129,31,129,30,122,31,122,30,141,31,112,31,145,31,145,30,233,31,233,30,233,29,233,28,1,31,251,31,134,31,65,31,87,31,99,31,192,31,192,30,137,31,20,31,51,31,197,31,120,31,61,31,60,31,85,31,233,31,230,31,243,31,107,31,84,31,139,31,139,30,201,31,45,31,132,31,129,31,194,31,194,30,130,31,41,31,5,31,191,31,98,31,98,30,145,31,212,31,212,30,212,29,57,31,255,31,85,31,94,31,194,31,194,30,60,31,32,31,20,31,149,31,149,30,184,31,132,31,204,31,215,31,70,31,136,31,136,30,7,31,33,31,64,31,149,31,206,31,82,31,179,31,185,31,185,30,185,29,225,31,62,31,142,31,131,31,210,31,234,31,245,31,245,30,148,31,148,30,149,31,36,31,36,30,254,31,132,31,200,31,241,31,241,30,187,31,47,31,47,30,51,31,51,30,94,31,94,30,196,31,141,31,194,31,194,30,194,29,194,28,194,27,194,26,194,25,201,31,201,30,104,31,40,31,172,31,134,31,229,31,82,31,218,31,68,31,68,30,169,31,40,31,105,31,89,31,98,31,195,31,150,31,226,31,226,30,141,31,254,31,78,31,220,31,86,31,206,31,90,31,90,30,47,31,47,30,82,31,173,31,178,31,150,31,223,31,57,31,115,31,115,30,127,31,10,31,12,31,12,30,80,31,244,31,244,30,65,31,88,31,224,31,201,31,10,31,15,31,235,31,218,31,218,30,218,29,149,31,57,31,57,30,57,29,57,28,83,31,86,31,102,31,51,31,96,31,236,31,236,30,236,29,139,31,229,31,229,30,32,31,32,30,90,31,27,31,50,31,50,30,62,31,191,31,124,31,52,31,157,31,189,31,136,31,236,31,236,30,184,31,91,31,91,30,91,29,159,31,159,30,13,31,163,31,124,31,124,30,12,31,12,30,54,31,107,31,54,31,156,31,156,30,156,29,156,28,28,31,24,31,252,31,120,31,206,31,206,30,206,29,99,31,77,31,95,31,227,31,193,31,65,31,126,31,40,31,18,31,228,31,34,31,169,31,169,30,209,31,156,31,156,30,142,31,41,31,179,31,65,31,222,31,7,31,165,31,113,31,159,31,236,31,150,31,195,31,195,30,5,31,140,31,70,31,26,31,158,31,52,31,17,31,98,31,243,31,66,31,154,31,154,30,115,31,152,31,47,31,47,30,150,31,136,31,136,30,136,29,2,31,166,31,116,31,152,31,186,31,141,31,131,31,124,31,71,31,223,31,4,31,120,31,2,31,225,31,246,31,208,31,172,31,237,31,193,31,31,31,31,30,107,31,122,31,126,31,226,31,168,31,152,31,99,31,99,30,216,31,183,31,183,30,183,29,70,31,251,31,254,31,56,31,56,30,56,29,51,31,98,31,220,31,220,30,62,31,230,31,230,30,105,31,29,31,105,31,105,30,71,31,71,30,188,31,188,30,157,31,69,31,71,31,181,31,181,30,144,31,151,31,173,31,135,31,93,31,203,31,25,31,152,31,115,31,252,31,179,31,87,31,195,31,136,31,92,31,92,30,162,31,162,30,58,31,3,31,116,31,3,31,168,31,62,31,194,31,140,31,234,31,35,31,36,31,234,31,75,31,103,31,253,31,253,30,101,31,58,31,58,30,113,31,223,31,171,31,171,30,93,31,63,31,117,31,182,31,255,31,130,31,11,31,98,31,184,31,222,31,44,31,129,31,39,31,206,31,123,31,43,31,201,31,103,31,199,31,216,31,138,31,134,31,137,31,28,31,15,31,64,31,122,31,216,31,216,30,119,31,73,31,31,31,110,31,132,31,178,31,178,30,31,31,28,31,57,31,166,31,107,31,50,31,132,31,117,31,168,31,43,31,43,30,233,31,254,31,155,31,134,31,25,31,36,31,147,31,147,30,3,31,113,31,113,30,223,31,205,31,205,30,190,31,190,30,254,31,92,31,92,30,92,29,238,31,79,31,221,31,134,31,106,31,106,30,106,29,106,28,18,31,234,31,125,31,58,31,175,31,187,31,12,31,233,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
