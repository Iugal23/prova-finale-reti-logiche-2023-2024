-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_781 is
end project_tb_781;

architecture project_tb_arch_781 of project_tb_781 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 148;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,215,0,0,0,80,0,0,0,0,0,113,0,102,0,235,0,163,0,0,0,133,0,188,0,197,0,109,0,0,0,47,0,0,0,154,0,212,0,51,0,0,0,14,0,225,0,247,0,96,0,127,0,201,0,254,0,145,0,151,0,191,0,136,0,188,0,13,0,175,0,235,0,0,0,0,0,0,0,194,0,64,0,0,0,239,0,159,0,254,0,156,0,37,0,0,0,9,0,71,0,13,0,213,0,75,0,0,0,209,0,37,0,252,0,220,0,224,0,42,0,32,0,67,0,131,0,195,0,239,0,246,0,5,0,30,0,31,0,113,0,91,0,201,0,0,0,0,0,18,0,229,0,0,0,169,0,0,0,0,0,7,0,208,0,40,0,233,0,0,0,0,0,0,0,133,0,0,0,165,0,72,0,81,0,178,0,145,0,84,0,0,0,223,0,0,0,0,0,95,0,212,0,124,0,32,0,81,0,94,0,0,0,63,0,78,0,119,0,135,0,140,0,190,0,0,0,90,0,55,0,25,0,117,0,101,0,214,0,80,0,207,0,231,0,194,0,129,0,126,0,0,0,0,0,248,0,0,0,0,0,58,0,194,0,253,0,108,0,92,0,182,0,64,0,76,0,179,0,105,0,125,0,241,0,46,0,44,0,107,0,144,0,168,0);
signal scenario_full  : scenario_type := (0,0,215,31,215,30,80,31,80,30,80,29,113,31,102,31,235,31,163,31,163,30,133,31,188,31,197,31,109,31,109,30,47,31,47,30,154,31,212,31,51,31,51,30,14,31,225,31,247,31,96,31,127,31,201,31,254,31,145,31,151,31,191,31,136,31,188,31,13,31,175,31,235,31,235,30,235,29,235,28,194,31,64,31,64,30,239,31,159,31,254,31,156,31,37,31,37,30,9,31,71,31,13,31,213,31,75,31,75,30,209,31,37,31,252,31,220,31,224,31,42,31,32,31,67,31,131,31,195,31,239,31,246,31,5,31,30,31,31,31,113,31,91,31,201,31,201,30,201,29,18,31,229,31,229,30,169,31,169,30,169,29,7,31,208,31,40,31,233,31,233,30,233,29,233,28,133,31,133,30,165,31,72,31,81,31,178,31,145,31,84,31,84,30,223,31,223,30,223,29,95,31,212,31,124,31,32,31,81,31,94,31,94,30,63,31,78,31,119,31,135,31,140,31,190,31,190,30,90,31,55,31,25,31,117,31,101,31,214,31,80,31,207,31,231,31,194,31,129,31,126,31,126,30,126,29,248,31,248,30,248,29,58,31,194,31,253,31,108,31,92,31,182,31,64,31,76,31,179,31,105,31,125,31,241,31,46,31,44,31,107,31,144,31,168,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
