-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 240;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (28,0,0,0,114,0,226,0,64,0,91,0,19,0,52,0,222,0,0,0,0,0,89,0,107,0,124,0,0,0,178,0,173,0,229,0,78,0,0,0,54,0,179,0,181,0,120,0,171,0,250,0,97,0,192,0,56,0,73,0,22,0,17,0,168,0,222,0,173,0,165,0,117,0,49,0,94,0,132,0,173,0,97,0,0,0,187,0,10,0,101,0,134,0,121,0,0,0,139,0,0,0,146,0,0,0,71,0,193,0,136,0,254,0,62,0,0,0,189,0,0,0,6,0,10,0,67,0,29,0,0,0,40,0,218,0,64,0,0,0,224,0,69,0,171,0,5,0,81,0,17,0,28,0,24,0,0,0,0,0,121,0,170,0,235,0,18,0,107,0,144,0,195,0,130,0,195,0,90,0,0,0,141,0,108,0,0,0,132,0,0,0,146,0,0,0,211,0,41,0,204,0,4,0,50,0,17,0,0,0,58,0,66,0,52,0,0,0,0,0,56,0,23,0,19,0,36,0,0,0,147,0,218,0,0,0,0,0,0,0,31,0,0,0,204,0,2,0,153,0,220,0,0,0,146,0,0,0,208,0,237,0,253,0,0,0,45,0,0,0,151,0,88,0,114,0,241,0,231,0,0,0,13,0,131,0,25,0,166,0,0,0,0,0,184,0,201,0,249,0,224,0,121,0,0,0,0,0,48,0,167,0,223,0,224,0,243,0,204,0,166,0,19,0,103,0,212,0,0,0,217,0,0,0,128,0,0,0,76,0,152,0,100,0,18,0,168,0,251,0,200,0,157,0,100,0,202,0,0,0,188,0,0,0,19,0,0,0,0,0,0,0,61,0,214,0,186,0,4,0,0,0,127,0,178,0,55,0,129,0,210,0,86,0,0,0,197,0,237,0,32,0,18,0,125,0,187,0,201,0,95,0,0,0,132,0,38,0,25,0,0,0,112,0,0,0,232,0,71,0,95,0,254,0,192,0,6,0,92,0,129,0,143,0,80,0,0,0,123,0,91,0,250,0,8,0,206,0,102,0,99,0,140,0,154,0,114,0,76,0,161,0,153,0,149,0,0,0,0,0);
signal scenario_full  : scenario_type := (28,31,28,30,114,31,226,31,64,31,91,31,19,31,52,31,222,31,222,30,222,29,89,31,107,31,124,31,124,30,178,31,173,31,229,31,78,31,78,30,54,31,179,31,181,31,120,31,171,31,250,31,97,31,192,31,56,31,73,31,22,31,17,31,168,31,222,31,173,31,165,31,117,31,49,31,94,31,132,31,173,31,97,31,97,30,187,31,10,31,101,31,134,31,121,31,121,30,139,31,139,30,146,31,146,30,71,31,193,31,136,31,254,31,62,31,62,30,189,31,189,30,6,31,10,31,67,31,29,31,29,30,40,31,218,31,64,31,64,30,224,31,69,31,171,31,5,31,81,31,17,31,28,31,24,31,24,30,24,29,121,31,170,31,235,31,18,31,107,31,144,31,195,31,130,31,195,31,90,31,90,30,141,31,108,31,108,30,132,31,132,30,146,31,146,30,211,31,41,31,204,31,4,31,50,31,17,31,17,30,58,31,66,31,52,31,52,30,52,29,56,31,23,31,19,31,36,31,36,30,147,31,218,31,218,30,218,29,218,28,31,31,31,30,204,31,2,31,153,31,220,31,220,30,146,31,146,30,208,31,237,31,253,31,253,30,45,31,45,30,151,31,88,31,114,31,241,31,231,31,231,30,13,31,131,31,25,31,166,31,166,30,166,29,184,31,201,31,249,31,224,31,121,31,121,30,121,29,48,31,167,31,223,31,224,31,243,31,204,31,166,31,19,31,103,31,212,31,212,30,217,31,217,30,128,31,128,30,76,31,152,31,100,31,18,31,168,31,251,31,200,31,157,31,100,31,202,31,202,30,188,31,188,30,19,31,19,30,19,29,19,28,61,31,214,31,186,31,4,31,4,30,127,31,178,31,55,31,129,31,210,31,86,31,86,30,197,31,237,31,32,31,18,31,125,31,187,31,201,31,95,31,95,30,132,31,38,31,25,31,25,30,112,31,112,30,232,31,71,31,95,31,254,31,192,31,6,31,92,31,129,31,143,31,80,31,80,30,123,31,91,31,250,31,8,31,206,31,102,31,99,31,140,31,154,31,114,31,76,31,161,31,153,31,149,31,149,30,149,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
