-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 771;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,35,0,0,0,0,0,0,0,8,0,195,0,237,0,0,0,39,0,55,0,7,0,8,0,211,0,141,0,0,0,115,0,0,0,143,0,206,0,173,0,210,0,9,0,33,0,29,0,216,0,38,0,0,0,0,0,30,0,240,0,82,0,179,0,92,0,137,0,255,0,138,0,92,0,236,0,116,0,96,0,0,0,0,0,99,0,0,0,146,0,5,0,173,0,238,0,255,0,43,0,159,0,55,0,210,0,158,0,0,0,0,0,237,0,86,0,89,0,117,0,0,0,141,0,8,0,90,0,0,0,108,0,132,0,0,0,119,0,145,0,159,0,70,0,37,0,42,0,132,0,142,0,0,0,49,0,91,0,0,0,80,0,225,0,103,0,195,0,0,0,70,0,104,0,0,0,0,0,248,0,148,0,38,0,0,0,206,0,0,0,115,0,107,0,0,0,186,0,222,0,60,0,185,0,36,0,0,0,142,0,182,0,0,0,0,0,197,0,222,0,65,0,135,0,253,0,66,0,0,0,3,0,195,0,145,0,0,0,0,0,65,0,43,0,5,0,238,0,173,0,154,0,0,0,62,0,142,0,0,0,235,0,236,0,13,0,248,0,174,0,0,0,85,0,79,0,133,0,0,0,147,0,88,0,29,0,0,0,0,0,28,0,133,0,0,0,0,0,247,0,0,0,0,0,246,0,106,0,174,0,22,0,168,0,122,0,0,0,208,0,0,0,45,0,117,0,0,0,22,0,229,0,245,0,0,0,61,0,93,0,67,0,117,0,0,0,93,0,0,0,171,0,25,0,33,0,77,0,214,0,95,0,0,0,247,0,0,0,127,0,0,0,12,0,117,0,162,0,211,0,43,0,0,0,66,0,73,0,61,0,231,0,244,0,19,0,202,0,63,0,92,0,245,0,0,0,191,0,217,0,193,0,171,0,129,0,59,0,49,0,138,0,118,0,35,0,185,0,182,0,0,0,172,0,0,0,115,0,62,0,147,0,0,0,244,0,173,0,186,0,214,0,0,0,69,0,224,0,190,0,61,0,0,0,178,0,0,0,0,0,153,0,125,0,1,0,0,0,18,0,154,0,73,0,26,0,48,0,118,0,79,0,165,0,14,0,103,0,251,0,85,0,0,0,53,0,191,0,249,0,142,0,0,0,125,0,124,0,66,0,21,0,223,0,105,0,242,0,99,0,216,0,167,0,156,0,108,0,101,0,187,0,0,0,226,0,14,0,195,0,249,0,0,0,81,0,0,0,97,0,166,0,111,0,225,0,48,0,119,0,98,0,176,0,91,0,58,0,84,0,198,0,168,0,72,0,14,0,108,0,29,0,1,0,239,0,28,0,14,0,190,0,112,0,0,0,159,0,79,0,0,0,244,0,0,0,4,0,73,0,117,0,70,0,2,0,156,0,102,0,0,0,209,0,194,0,218,0,0,0,0,0,0,0,24,0,229,0,107,0,49,0,93,0,151,0,100,0,88,0,158,0,84,0,0,0,70,0,93,0,221,0,76,0,223,0,111,0,170,0,99,0,39,0,212,0,134,0,99,0,55,0,102,0,153,0,0,0,240,0,207,0,13,0,233,0,0,0,0,0,203,0,191,0,219,0,168,0,72,0,0,0,214,0,0,0,0,0,0,0,170,0,220,0,164,0,0,0,0,0,115,0,134,0,0,0,151,0,189,0,52,0,0,0,214,0,241,0,132,0,0,0,135,0,40,0,0,0,198,0,176,0,0,0,112,0,10,0,2,0,96,0,157,0,55,0,123,0,31,0,160,0,170,0,135,0,0,0,0,0,220,0,51,0,49,0,0,0,105,0,42,0,79,0,221,0,1,0,189,0,229,0,254,0,0,0,0,0,78,0,72,0,68,0,3,0,85,0,72,0,83,0,220,0,191,0,42,0,35,0,185,0,153,0,168,0,198,0,0,0,211,0,189,0,137,0,0,0,50,0,190,0,0,0,46,0,165,0,98,0,134,0,42,0,123,0,222,0,0,0,242,0,107,0,195,0,216,0,236,0,0,0,30,0,34,0,2,0,173,0,237,0,0,0,5,0,162,0,179,0,49,0,0,0,49,0,24,0,87,0,38,0,70,0,0,0,235,0,0,0,19,0,12,0,73,0,0,0,6,0,16,0,0,0,0,0,0,0,197,0,252,0,145,0,0,0,170,0,137,0,0,0,0,0,8,0,101,0,197,0,174,0,0,0,179,0,0,0,59,0,76,0,151,0,197,0,51,0,191,0,0,0,240,0,229,0,74,0,0,0,215,0,61,0,0,0,244,0,0,0,90,0,2,0,0,0,189,0,135,0,21,0,214,0,228,0,172,0,72,0,180,0,240,0,47,0,0,0,165,0,0,0,0,0,17,0,190,0,160,0,86,0,239,0,61,0,183,0,208,0,194,0,72,0,155,0,69,0,217,0,0,0,3,0,61,0,160,0,126,0,100,0,192,0,72,0,184,0,132,0,56,0,188,0,255,0,43,0,61,0,187,0,120,0,44,0,0,0,184,0,2,0,0,0,241,0,253,0,68,0,0,0,0,0,62,0,89,0,0,0,220,0,224,0,20,0,0,0,183,0,144,0,250,0,127,0,114,0,0,0,233,0,167,0,142,0,119,0,165,0,108,0,0,0,24,0,213,0,215,0,54,0,92,0,0,0,247,0,128,0,32,0,0,0,138,0,56,0,21,0,78,0,0,0,0,0,67,0,37,0,68,0,69,0,0,0,116,0,83,0,68,0,247,0,93,0,169,0,215,0,67,0,132,0,220,0,251,0,186,0,127,0,32,0,0,0,134,0,126,0,239,0,188,0,160,0,54,0,221,0,0,0,59,0,0,0,192,0,204,0,0,0,41,0,15,0,0,0,0,0,19,0,171,0,0,0,237,0,0,0,183,0,78,0,129,0,0,0,0,0,0,0,193,0,33,0,9,0,183,0,32,0,243,0,75,0,0,0,64,0,0,0,150,0,152,0,40,0,46,0,189,0,132,0,242,0,0,0,0,0,16,0,136,0,55,0,231,0,72,0,129,0,29,0,0,0,57,0,57,0,194,0,204,0,176,0,73,0,130,0,130,0,222,0,0,0,103,0,141,0,91,0,0,0,236,0,0,0,84,0,120,0,0,0,15,0,9,0,0,0,145,0,104,0,0,0,120,0,248,0,190,0,32,0,180,0,95,0,0,0,77,0,0,0,221,0,82,0,21,0,245,0,252,0,136,0,213,0,10,0,187,0,0,0,44,0,6,0,16,0,208,0,0,0,160,0,3,0,0,0,227,0,197,0,37,0,0,0,61,0,22,0,125,0,0,0,98,0,141,0,156,0,245,0,111,0,8,0,206,0,242,0,44,0,45,0,121,0,212,0,0,0,42,0,57,0,0,0,137,0,0,0,114,0,0,0,43,0,155,0,116,0,55,0,205,0,153,0,0,0,223,0,57,0,203,0,56,0,0,0);
signal scenario_full  : scenario_type := (0,0,35,31,35,30,35,29,35,28,8,31,195,31,237,31,237,30,39,31,55,31,7,31,8,31,211,31,141,31,141,30,115,31,115,30,143,31,206,31,173,31,210,31,9,31,33,31,29,31,216,31,38,31,38,30,38,29,30,31,240,31,82,31,179,31,92,31,137,31,255,31,138,31,92,31,236,31,116,31,96,31,96,30,96,29,99,31,99,30,146,31,5,31,173,31,238,31,255,31,43,31,159,31,55,31,210,31,158,31,158,30,158,29,237,31,86,31,89,31,117,31,117,30,141,31,8,31,90,31,90,30,108,31,132,31,132,30,119,31,145,31,159,31,70,31,37,31,42,31,132,31,142,31,142,30,49,31,91,31,91,30,80,31,225,31,103,31,195,31,195,30,70,31,104,31,104,30,104,29,248,31,148,31,38,31,38,30,206,31,206,30,115,31,107,31,107,30,186,31,222,31,60,31,185,31,36,31,36,30,142,31,182,31,182,30,182,29,197,31,222,31,65,31,135,31,253,31,66,31,66,30,3,31,195,31,145,31,145,30,145,29,65,31,43,31,5,31,238,31,173,31,154,31,154,30,62,31,142,31,142,30,235,31,236,31,13,31,248,31,174,31,174,30,85,31,79,31,133,31,133,30,147,31,88,31,29,31,29,30,29,29,28,31,133,31,133,30,133,29,247,31,247,30,247,29,246,31,106,31,174,31,22,31,168,31,122,31,122,30,208,31,208,30,45,31,117,31,117,30,22,31,229,31,245,31,245,30,61,31,93,31,67,31,117,31,117,30,93,31,93,30,171,31,25,31,33,31,77,31,214,31,95,31,95,30,247,31,247,30,127,31,127,30,12,31,117,31,162,31,211,31,43,31,43,30,66,31,73,31,61,31,231,31,244,31,19,31,202,31,63,31,92,31,245,31,245,30,191,31,217,31,193,31,171,31,129,31,59,31,49,31,138,31,118,31,35,31,185,31,182,31,182,30,172,31,172,30,115,31,62,31,147,31,147,30,244,31,173,31,186,31,214,31,214,30,69,31,224,31,190,31,61,31,61,30,178,31,178,30,178,29,153,31,125,31,1,31,1,30,18,31,154,31,73,31,26,31,48,31,118,31,79,31,165,31,14,31,103,31,251,31,85,31,85,30,53,31,191,31,249,31,142,31,142,30,125,31,124,31,66,31,21,31,223,31,105,31,242,31,99,31,216,31,167,31,156,31,108,31,101,31,187,31,187,30,226,31,14,31,195,31,249,31,249,30,81,31,81,30,97,31,166,31,111,31,225,31,48,31,119,31,98,31,176,31,91,31,58,31,84,31,198,31,168,31,72,31,14,31,108,31,29,31,1,31,239,31,28,31,14,31,190,31,112,31,112,30,159,31,79,31,79,30,244,31,244,30,4,31,73,31,117,31,70,31,2,31,156,31,102,31,102,30,209,31,194,31,218,31,218,30,218,29,218,28,24,31,229,31,107,31,49,31,93,31,151,31,100,31,88,31,158,31,84,31,84,30,70,31,93,31,221,31,76,31,223,31,111,31,170,31,99,31,39,31,212,31,134,31,99,31,55,31,102,31,153,31,153,30,240,31,207,31,13,31,233,31,233,30,233,29,203,31,191,31,219,31,168,31,72,31,72,30,214,31,214,30,214,29,214,28,170,31,220,31,164,31,164,30,164,29,115,31,134,31,134,30,151,31,189,31,52,31,52,30,214,31,241,31,132,31,132,30,135,31,40,31,40,30,198,31,176,31,176,30,112,31,10,31,2,31,96,31,157,31,55,31,123,31,31,31,160,31,170,31,135,31,135,30,135,29,220,31,51,31,49,31,49,30,105,31,42,31,79,31,221,31,1,31,189,31,229,31,254,31,254,30,254,29,78,31,72,31,68,31,3,31,85,31,72,31,83,31,220,31,191,31,42,31,35,31,185,31,153,31,168,31,198,31,198,30,211,31,189,31,137,31,137,30,50,31,190,31,190,30,46,31,165,31,98,31,134,31,42,31,123,31,222,31,222,30,242,31,107,31,195,31,216,31,236,31,236,30,30,31,34,31,2,31,173,31,237,31,237,30,5,31,162,31,179,31,49,31,49,30,49,31,24,31,87,31,38,31,70,31,70,30,235,31,235,30,19,31,12,31,73,31,73,30,6,31,16,31,16,30,16,29,16,28,197,31,252,31,145,31,145,30,170,31,137,31,137,30,137,29,8,31,101,31,197,31,174,31,174,30,179,31,179,30,59,31,76,31,151,31,197,31,51,31,191,31,191,30,240,31,229,31,74,31,74,30,215,31,61,31,61,30,244,31,244,30,90,31,2,31,2,30,189,31,135,31,21,31,214,31,228,31,172,31,72,31,180,31,240,31,47,31,47,30,165,31,165,30,165,29,17,31,190,31,160,31,86,31,239,31,61,31,183,31,208,31,194,31,72,31,155,31,69,31,217,31,217,30,3,31,61,31,160,31,126,31,100,31,192,31,72,31,184,31,132,31,56,31,188,31,255,31,43,31,61,31,187,31,120,31,44,31,44,30,184,31,2,31,2,30,241,31,253,31,68,31,68,30,68,29,62,31,89,31,89,30,220,31,224,31,20,31,20,30,183,31,144,31,250,31,127,31,114,31,114,30,233,31,167,31,142,31,119,31,165,31,108,31,108,30,24,31,213,31,215,31,54,31,92,31,92,30,247,31,128,31,32,31,32,30,138,31,56,31,21,31,78,31,78,30,78,29,67,31,37,31,68,31,69,31,69,30,116,31,83,31,68,31,247,31,93,31,169,31,215,31,67,31,132,31,220,31,251,31,186,31,127,31,32,31,32,30,134,31,126,31,239,31,188,31,160,31,54,31,221,31,221,30,59,31,59,30,192,31,204,31,204,30,41,31,15,31,15,30,15,29,19,31,171,31,171,30,237,31,237,30,183,31,78,31,129,31,129,30,129,29,129,28,193,31,33,31,9,31,183,31,32,31,243,31,75,31,75,30,64,31,64,30,150,31,152,31,40,31,46,31,189,31,132,31,242,31,242,30,242,29,16,31,136,31,55,31,231,31,72,31,129,31,29,31,29,30,57,31,57,31,194,31,204,31,176,31,73,31,130,31,130,31,222,31,222,30,103,31,141,31,91,31,91,30,236,31,236,30,84,31,120,31,120,30,15,31,9,31,9,30,145,31,104,31,104,30,120,31,248,31,190,31,32,31,180,31,95,31,95,30,77,31,77,30,221,31,82,31,21,31,245,31,252,31,136,31,213,31,10,31,187,31,187,30,44,31,6,31,16,31,208,31,208,30,160,31,3,31,3,30,227,31,197,31,37,31,37,30,61,31,22,31,125,31,125,30,98,31,141,31,156,31,245,31,111,31,8,31,206,31,242,31,44,31,45,31,121,31,212,31,212,30,42,31,57,31,57,30,137,31,137,30,114,31,114,30,43,31,155,31,116,31,55,31,205,31,153,31,153,30,223,31,57,31,203,31,56,31,56,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
