-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 686;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,152,0,235,0,141,0,76,0,29,0,114,0,220,0,47,0,34,0,27,0,214,0,22,0,246,0,162,0,0,0,12,0,0,0,191,0,0,0,0,0,149,0,93,0,31,0,177,0,185,0,100,0,28,0,221,0,63,0,204,0,74,0,9,0,140,0,155,0,97,0,0,0,90,0,220,0,221,0,125,0,126,0,18,0,154,0,0,0,62,0,43,0,213,0,100,0,29,0,0,0,159,0,0,0,47,0,159,0,52,0,112,0,0,0,0,0,240,0,70,0,181,0,38,0,160,0,241,0,248,0,0,0,31,0,240,0,152,0,200,0,252,0,234,0,165,0,144,0,185,0,0,0,0,0,187,0,39,0,77,0,24,0,232,0,19,0,250,0,169,0,152,0,37,0,252,0,117,0,188,0,0,0,212,0,0,0,40,0,0,0,0,0,67,0,0,0,22,0,143,0,121,0,0,0,218,0,134,0,96,0,137,0,192,0,205,0,168,0,255,0,201,0,134,0,135,0,98,0,19,0,226,0,0,0,169,0,181,0,159,0,246,0,198,0,124,0,0,0,168,0,43,0,93,0,58,0,0,0,85,0,165,0,46,0,135,0,0,0,0,0,155,0,140,0,2,0,197,0,186,0,178,0,0,0,0,0,204,0,95,0,240,0,213,0,0,0,2,0,166,0,137,0,45,0,0,0,222,0,119,0,189,0,195,0,13,0,19,0,234,0,206,0,0,0,171,0,37,0,0,0,158,0,223,0,112,0,178,0,155,0,0,0,109,0,247,0,0,0,46,0,220,0,0,0,3,0,145,0,15,0,255,0,242,0,193,0,244,0,125,0,205,0,51,0,45,0,19,0,66,0,160,0,92,0,0,0,250,0,0,0,51,0,101,0,141,0,66,0,0,0,0,0,170,0,1,0,169,0,83,0,239,0,127,0,0,0,0,0,125,0,112,0,19,0,254,0,0,0,7,0,196,0,83,0,0,0,128,0,0,0,141,0,91,0,0,0,116,0,89,0,78,0,137,0,0,0,0,0,232,0,186,0,198,0,111,0,0,0,21,0,247,0,150,0,124,0,164,0,216,0,0,0,207,0,86,0,68,0,0,0,85,0,84,0,19,0,251,0,0,0,0,0,172,0,240,0,0,0,0,0,0,0,138,0,172,0,252,0,75,0,159,0,0,0,249,0,0,0,0,0,173,0,245,0,8,0,36,0,118,0,173,0,86,0,31,0,151,0,134,0,64,0,137,0,62,0,91,0,131,0,184,0,179,0,196,0,0,0,0,0,189,0,0,0,215,0,0,0,134,0,24,0,0,0,0,0,62,0,177,0,96,0,168,0,126,0,237,0,126,0,50,0,209,0,109,0,198,0,0,0,164,0,210,0,253,0,30,0,227,0,0,0,191,0,60,0,0,0,112,0,0,0,198,0,189,0,0,0,128,0,157,0,210,0,56,0,185,0,0,0,182,0,34,0,0,0,121,0,246,0,215,0,122,0,222,0,0,0,112,0,0,0,145,0,0,0,13,0,0,0,199,0,72,0,205,0,168,0,37,0,204,0,97,0,158,0,0,0,0,0,118,0,104,0,18,0,86,0,67,0,0,0,150,0,13,0,236,0,193,0,32,0,158,0,227,0,36,0,0,0,47,0,88,0,61,0,67,0,198,0,118,0,166,0,168,0,34,0,35,0,0,0,0,0,33,0,0,0,33,0,151,0,211,0,84,0,183,0,0,0,0,0,194,0,34,0,191,0,98,0,147,0,124,0,185,0,56,0,32,0,107,0,235,0,97,0,118,0,128,0,194,0,0,0,178,0,93,0,150,0,243,0,33,0,54,0,227,0,142,0,209,0,19,0,112,0,0,0,2,0,87,0,234,0,0,0,176,0,14,0,89,0,96,0,0,0,0,0,222,0,176,0,0,0,97,0,90,0,202,0,29,0,250,0,54,0,72,0,166,0,191,0,238,0,0,0,0,0,199,0,206,0,75,0,207,0,148,0,20,0,247,0,197,0,0,0,0,0,31,0,0,0,207,0,157,0,100,0,150,0,95,0,0,0,137,0,87,0,80,0,10,0,120,0,129,0,246,0,75,0,107,0,15,0,56,0,255,0,9,0,254,0,187,0,210,0,0,0,250,0,0,0,250,0,153,0,145,0,0,0,137,0,56,0,0,0,71,0,235,0,63,0,0,0,0,0,191,0,232,0,245,0,36,0,32,0,103,0,3,0,139,0,0,0,18,0,243,0,189,0,103,0,0,0,52,0,0,0,137,0,0,0,39,0,0,0,124,0,165,0,90,0,63,0,31,0,26,0,235,0,189,0,248,0,0,0,250,0,7,0,158,0,168,0,105,0,105,0,0,0,145,0,68,0,30,0,57,0,225,0,0,0,0,0,0,0,80,0,127,0,136,0,200,0,10,0,178,0,125,0,115,0,53,0,135,0,0,0,129,0,44,0,61,0,65,0,38,0,0,0,62,0,0,0,116,0,133,0,245,0,0,0,0,0,163,0,99,0,0,0,51,0,18,0,0,0,46,0,89,0,138,0,87,0,249,0,75,0,0,0,238,0,147,0,47,0,234,0,118,0,220,0,165,0,216,0,213,0,27,0,116,0,126,0,70,0,0,0,140,0,0,0,84,0,17,0,0,0,220,0,243,0,117,0,115,0,0,0,250,0,215,0,92,0,138,0,201,0,0,0,123,0,0,0,180,0,183,0,80,0,12,0,62,0,0,0,44,0,84,0,0,0,33,0,135,0,0,0,120,0,3,0,0,0,194,0,22,0,150,0,0,0,0,0,170,0,0,0,99,0,0,0,0,0,0,0,248,0,240,0,176,0,224,0,145,0,253,0,106,0,11,0,78,0,30,0,142,0,111,0,64,0,0,0,0,0,73,0,0,0,231,0,129,0,211,0,209,0,27,0,39,0,76,0,0,0,230,0,205,0,78,0,137,0,57,0,125,0,122,0,187,0,1,0,0,0,106,0,146,0,122,0,205,0,70,0,35,0,0,0,0,0,16,0,94,0,16,0,0,0,98,0,0,0,0,0,0,0,99,0,0,0,104,0,251,0,147,0);
signal scenario_full  : scenario_type := (0,0,0,0,152,31,235,31,141,31,76,31,29,31,114,31,220,31,47,31,34,31,27,31,214,31,22,31,246,31,162,31,162,30,12,31,12,30,191,31,191,30,191,29,149,31,93,31,31,31,177,31,185,31,100,31,28,31,221,31,63,31,204,31,74,31,9,31,140,31,155,31,97,31,97,30,90,31,220,31,221,31,125,31,126,31,18,31,154,31,154,30,62,31,43,31,213,31,100,31,29,31,29,30,159,31,159,30,47,31,159,31,52,31,112,31,112,30,112,29,240,31,70,31,181,31,38,31,160,31,241,31,248,31,248,30,31,31,240,31,152,31,200,31,252,31,234,31,165,31,144,31,185,31,185,30,185,29,187,31,39,31,77,31,24,31,232,31,19,31,250,31,169,31,152,31,37,31,252,31,117,31,188,31,188,30,212,31,212,30,40,31,40,30,40,29,67,31,67,30,22,31,143,31,121,31,121,30,218,31,134,31,96,31,137,31,192,31,205,31,168,31,255,31,201,31,134,31,135,31,98,31,19,31,226,31,226,30,169,31,181,31,159,31,246,31,198,31,124,31,124,30,168,31,43,31,93,31,58,31,58,30,85,31,165,31,46,31,135,31,135,30,135,29,155,31,140,31,2,31,197,31,186,31,178,31,178,30,178,29,204,31,95,31,240,31,213,31,213,30,2,31,166,31,137,31,45,31,45,30,222,31,119,31,189,31,195,31,13,31,19,31,234,31,206,31,206,30,171,31,37,31,37,30,158,31,223,31,112,31,178,31,155,31,155,30,109,31,247,31,247,30,46,31,220,31,220,30,3,31,145,31,15,31,255,31,242,31,193,31,244,31,125,31,205,31,51,31,45,31,19,31,66,31,160,31,92,31,92,30,250,31,250,30,51,31,101,31,141,31,66,31,66,30,66,29,170,31,1,31,169,31,83,31,239,31,127,31,127,30,127,29,125,31,112,31,19,31,254,31,254,30,7,31,196,31,83,31,83,30,128,31,128,30,141,31,91,31,91,30,116,31,89,31,78,31,137,31,137,30,137,29,232,31,186,31,198,31,111,31,111,30,21,31,247,31,150,31,124,31,164,31,216,31,216,30,207,31,86,31,68,31,68,30,85,31,84,31,19,31,251,31,251,30,251,29,172,31,240,31,240,30,240,29,240,28,138,31,172,31,252,31,75,31,159,31,159,30,249,31,249,30,249,29,173,31,245,31,8,31,36,31,118,31,173,31,86,31,31,31,151,31,134,31,64,31,137,31,62,31,91,31,131,31,184,31,179,31,196,31,196,30,196,29,189,31,189,30,215,31,215,30,134,31,24,31,24,30,24,29,62,31,177,31,96,31,168,31,126,31,237,31,126,31,50,31,209,31,109,31,198,31,198,30,164,31,210,31,253,31,30,31,227,31,227,30,191,31,60,31,60,30,112,31,112,30,198,31,189,31,189,30,128,31,157,31,210,31,56,31,185,31,185,30,182,31,34,31,34,30,121,31,246,31,215,31,122,31,222,31,222,30,112,31,112,30,145,31,145,30,13,31,13,30,199,31,72,31,205,31,168,31,37,31,204,31,97,31,158,31,158,30,158,29,118,31,104,31,18,31,86,31,67,31,67,30,150,31,13,31,236,31,193,31,32,31,158,31,227,31,36,31,36,30,47,31,88,31,61,31,67,31,198,31,118,31,166,31,168,31,34,31,35,31,35,30,35,29,33,31,33,30,33,31,151,31,211,31,84,31,183,31,183,30,183,29,194,31,34,31,191,31,98,31,147,31,124,31,185,31,56,31,32,31,107,31,235,31,97,31,118,31,128,31,194,31,194,30,178,31,93,31,150,31,243,31,33,31,54,31,227,31,142,31,209,31,19,31,112,31,112,30,2,31,87,31,234,31,234,30,176,31,14,31,89,31,96,31,96,30,96,29,222,31,176,31,176,30,97,31,90,31,202,31,29,31,250,31,54,31,72,31,166,31,191,31,238,31,238,30,238,29,199,31,206,31,75,31,207,31,148,31,20,31,247,31,197,31,197,30,197,29,31,31,31,30,207,31,157,31,100,31,150,31,95,31,95,30,137,31,87,31,80,31,10,31,120,31,129,31,246,31,75,31,107,31,15,31,56,31,255,31,9,31,254,31,187,31,210,31,210,30,250,31,250,30,250,31,153,31,145,31,145,30,137,31,56,31,56,30,71,31,235,31,63,31,63,30,63,29,191,31,232,31,245,31,36,31,32,31,103,31,3,31,139,31,139,30,18,31,243,31,189,31,103,31,103,30,52,31,52,30,137,31,137,30,39,31,39,30,124,31,165,31,90,31,63,31,31,31,26,31,235,31,189,31,248,31,248,30,250,31,7,31,158,31,168,31,105,31,105,31,105,30,145,31,68,31,30,31,57,31,225,31,225,30,225,29,225,28,80,31,127,31,136,31,200,31,10,31,178,31,125,31,115,31,53,31,135,31,135,30,129,31,44,31,61,31,65,31,38,31,38,30,62,31,62,30,116,31,133,31,245,31,245,30,245,29,163,31,99,31,99,30,51,31,18,31,18,30,46,31,89,31,138,31,87,31,249,31,75,31,75,30,238,31,147,31,47,31,234,31,118,31,220,31,165,31,216,31,213,31,27,31,116,31,126,31,70,31,70,30,140,31,140,30,84,31,17,31,17,30,220,31,243,31,117,31,115,31,115,30,250,31,215,31,92,31,138,31,201,31,201,30,123,31,123,30,180,31,183,31,80,31,12,31,62,31,62,30,44,31,84,31,84,30,33,31,135,31,135,30,120,31,3,31,3,30,194,31,22,31,150,31,150,30,150,29,170,31,170,30,99,31,99,30,99,29,99,28,248,31,240,31,176,31,224,31,145,31,253,31,106,31,11,31,78,31,30,31,142,31,111,31,64,31,64,30,64,29,73,31,73,30,231,31,129,31,211,31,209,31,27,31,39,31,76,31,76,30,230,31,205,31,78,31,137,31,57,31,125,31,122,31,187,31,1,31,1,30,106,31,146,31,122,31,205,31,70,31,35,31,35,30,35,29,16,31,94,31,16,31,16,30,98,31,98,30,98,29,98,28,99,31,99,30,104,31,251,31,147,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
