-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_125 is
end project_tb_125;

architecture project_tb_arch_125 of project_tb_125 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 521;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (108,0,175,0,0,0,77,0,157,0,0,0,0,0,36,0,21,0,1,0,0,0,196,0,193,0,172,0,157,0,86,0,135,0,131,0,2,0,219,0,36,0,0,0,31,0,237,0,137,0,118,0,236,0,0,0,255,0,0,0,0,0,183,0,22,0,0,0,0,0,0,0,140,0,41,0,192,0,135,0,96,0,184,0,0,0,140,0,0,0,108,0,0,0,221,0,2,0,90,0,184,0,191,0,98,0,51,0,209,0,201,0,104,0,0,0,138,0,14,0,198,0,19,0,139,0,119,0,131,0,39,0,108,0,72,0,0,0,159,0,27,0,0,0,137,0,0,0,0,0,0,0,26,0,181,0,37,0,150,0,217,0,0,0,98,0,0,0,0,0,19,0,201,0,83,0,0,0,138,0,68,0,93,0,213,0,102,0,96,0,40,0,0,0,249,0,0,0,139,0,95,0,0,0,191,0,0,0,0,0,240,0,12,0,62,0,0,0,102,0,174,0,0,0,0,0,0,0,165,0,52,0,57,0,147,0,90,0,125,0,108,0,33,0,95,0,212,0,54,0,146,0,42,0,0,0,153,0,0,0,242,0,3,0,69,0,63,0,73,0,168,0,0,0,0,0,156,0,236,0,0,0,0,0,68,0,19,0,69,0,23,0,58,0,166,0,79,0,244,0,34,0,125,0,14,0,202,0,22,0,0,0,182,0,155,0,161,0,0,0,170,0,160,0,11,0,20,0,178,0,128,0,0,0,129,0,209,0,32,0,120,0,196,0,0,0,204,0,0,0,53,0,0,0,76,0,116,0,122,0,84,0,202,0,140,0,111,0,0,0,64,0,220,0,13,0,0,0,108,0,182,0,0,0,154,0,182,0,226,0,203,0,109,0,253,0,82,0,114,0,113,0,239,0,72,0,22,0,154,0,254,0,96,0,122,0,62,0,210,0,174,0,174,0,131,0,0,0,67,0,229,0,232,0,191,0,142,0,178,0,79,0,0,0,24,0,115,0,191,0,224,0,0,0,172,0,195,0,68,0,110,0,0,0,253,0,119,0,241,0,172,0,161,0,103,0,0,0,135,0,176,0,249,0,25,0,59,0,107,0,176,0,8,0,179,0,106,0,0,0,158,0,2,0,103,0,15,0,47,0,125,0,0,0,26,0,227,0,128,0,0,0,0,0,137,0,255,0,108,0,237,0,250,0,0,0,73,0,163,0,86,0,0,0,0,0,188,0,25,0,0,0,0,0,172,0,125,0,58,0,147,0,168,0,106,0,82,0,0,0,142,0,0,0,89,0,56,0,64,0,16,0,0,0,146,0,191,0,145,0,46,0,228,0,0,0,0,0,172,0,179,0,212,0,252,0,0,0,90,0,165,0,44,0,180,0,185,0,246,0,210,0,212,0,211,0,228,0,0,0,0,0,43,0,202,0,203,0,0,0,115,0,231,0,5,0,0,0,0,0,0,0,78,0,250,0,217,0,16,0,93,0,0,0,191,0,0,0,6,0,0,0,248,0,231,0,186,0,225,0,254,0,250,0,179,0,137,0,221,0,61,0,77,0,20,0,0,0,251,0,185,0,114,0,27,0,0,0,181,0,216,0,49,0,180,0,133,0,78,0,157,0,224,0,24,0,0,0,162,0,39,0,0,0,8,0,107,0,112,0,10,0,227,0,0,0,3,0,20,0,122,0,216,0,82,0,22,0,249,0,0,0,0,0,0,0,161,0,245,0,0,0,245,0,54,0,167,0,0,0,0,0,0,0,161,0,212,0,0,0,114,0,127,0,0,0,0,0,239,0,13,0,196,0,0,0,252,0,70,0,86,0,10,0,0,0,0,0,244,0,74,0,241,0,165,0,207,0,160,0,239,0,0,0,0,0,37,0,223,0,217,0,7,0,0,0,28,0,251,0,189,0,0,0,131,0,70,0,150,0,35,0,163,0,195,0,202,0,197,0,45,0,172,0,101,0,144,0,2,0,150,0,40,0,0,0,0,0,218,0,0,0,145,0,0,0,56,0,157,0,0,0,0,0,102,0,0,0,94,0,0,0,227,0,5,0,239,0,0,0,155,0,233,0,228,0,0,0,204,0,0,0,0,0,0,0,0,0,61,0,18,0,15,0,0,0,255,0,0,0,20,0,198,0,17,0,231,0,110,0,214,0,62,0,88,0,158,0,5,0,0,0,2,0,66,0,232,0,135,0,41,0,22,0,63,0,251,0,96,0,94,0,0,0,45,0,139,0,0,0,0,0,233,0,146,0,138,0,0,0,0,0,174,0,48,0,222,0,176,0,113,0,134,0,0,0,185,0,96,0,235,0,246,0,215,0,185,0,237,0,240,0);
signal scenario_full  : scenario_type := (108,31,175,31,175,30,77,31,157,31,157,30,157,29,36,31,21,31,1,31,1,30,196,31,193,31,172,31,157,31,86,31,135,31,131,31,2,31,219,31,36,31,36,30,31,31,237,31,137,31,118,31,236,31,236,30,255,31,255,30,255,29,183,31,22,31,22,30,22,29,22,28,140,31,41,31,192,31,135,31,96,31,184,31,184,30,140,31,140,30,108,31,108,30,221,31,2,31,90,31,184,31,191,31,98,31,51,31,209,31,201,31,104,31,104,30,138,31,14,31,198,31,19,31,139,31,119,31,131,31,39,31,108,31,72,31,72,30,159,31,27,31,27,30,137,31,137,30,137,29,137,28,26,31,181,31,37,31,150,31,217,31,217,30,98,31,98,30,98,29,19,31,201,31,83,31,83,30,138,31,68,31,93,31,213,31,102,31,96,31,40,31,40,30,249,31,249,30,139,31,95,31,95,30,191,31,191,30,191,29,240,31,12,31,62,31,62,30,102,31,174,31,174,30,174,29,174,28,165,31,52,31,57,31,147,31,90,31,125,31,108,31,33,31,95,31,212,31,54,31,146,31,42,31,42,30,153,31,153,30,242,31,3,31,69,31,63,31,73,31,168,31,168,30,168,29,156,31,236,31,236,30,236,29,68,31,19,31,69,31,23,31,58,31,166,31,79,31,244,31,34,31,125,31,14,31,202,31,22,31,22,30,182,31,155,31,161,31,161,30,170,31,160,31,11,31,20,31,178,31,128,31,128,30,129,31,209,31,32,31,120,31,196,31,196,30,204,31,204,30,53,31,53,30,76,31,116,31,122,31,84,31,202,31,140,31,111,31,111,30,64,31,220,31,13,31,13,30,108,31,182,31,182,30,154,31,182,31,226,31,203,31,109,31,253,31,82,31,114,31,113,31,239,31,72,31,22,31,154,31,254,31,96,31,122,31,62,31,210,31,174,31,174,31,131,31,131,30,67,31,229,31,232,31,191,31,142,31,178,31,79,31,79,30,24,31,115,31,191,31,224,31,224,30,172,31,195,31,68,31,110,31,110,30,253,31,119,31,241,31,172,31,161,31,103,31,103,30,135,31,176,31,249,31,25,31,59,31,107,31,176,31,8,31,179,31,106,31,106,30,158,31,2,31,103,31,15,31,47,31,125,31,125,30,26,31,227,31,128,31,128,30,128,29,137,31,255,31,108,31,237,31,250,31,250,30,73,31,163,31,86,31,86,30,86,29,188,31,25,31,25,30,25,29,172,31,125,31,58,31,147,31,168,31,106,31,82,31,82,30,142,31,142,30,89,31,56,31,64,31,16,31,16,30,146,31,191,31,145,31,46,31,228,31,228,30,228,29,172,31,179,31,212,31,252,31,252,30,90,31,165,31,44,31,180,31,185,31,246,31,210,31,212,31,211,31,228,31,228,30,228,29,43,31,202,31,203,31,203,30,115,31,231,31,5,31,5,30,5,29,5,28,78,31,250,31,217,31,16,31,93,31,93,30,191,31,191,30,6,31,6,30,248,31,231,31,186,31,225,31,254,31,250,31,179,31,137,31,221,31,61,31,77,31,20,31,20,30,251,31,185,31,114,31,27,31,27,30,181,31,216,31,49,31,180,31,133,31,78,31,157,31,224,31,24,31,24,30,162,31,39,31,39,30,8,31,107,31,112,31,10,31,227,31,227,30,3,31,20,31,122,31,216,31,82,31,22,31,249,31,249,30,249,29,249,28,161,31,245,31,245,30,245,31,54,31,167,31,167,30,167,29,167,28,161,31,212,31,212,30,114,31,127,31,127,30,127,29,239,31,13,31,196,31,196,30,252,31,70,31,86,31,10,31,10,30,10,29,244,31,74,31,241,31,165,31,207,31,160,31,239,31,239,30,239,29,37,31,223,31,217,31,7,31,7,30,28,31,251,31,189,31,189,30,131,31,70,31,150,31,35,31,163,31,195,31,202,31,197,31,45,31,172,31,101,31,144,31,2,31,150,31,40,31,40,30,40,29,218,31,218,30,145,31,145,30,56,31,157,31,157,30,157,29,102,31,102,30,94,31,94,30,227,31,5,31,239,31,239,30,155,31,233,31,228,31,228,30,204,31,204,30,204,29,204,28,204,27,61,31,18,31,15,31,15,30,255,31,255,30,20,31,198,31,17,31,231,31,110,31,214,31,62,31,88,31,158,31,5,31,5,30,2,31,66,31,232,31,135,31,41,31,22,31,63,31,251,31,96,31,94,31,94,30,45,31,139,31,139,30,139,29,233,31,146,31,138,31,138,30,138,29,174,31,48,31,222,31,176,31,113,31,134,31,134,30,185,31,96,31,235,31,246,31,215,31,185,31,237,31,240,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
