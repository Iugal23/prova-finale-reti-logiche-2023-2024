-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_808 is
end project_tb_808;

architecture project_tb_arch_808 of project_tb_808 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 837;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (39,0,0,0,239,0,30,0,0,0,156,0,0,0,0,0,183,0,0,0,111,0,0,0,168,0,240,0,79,0,106,0,109,0,229,0,0,0,239,0,154,0,0,0,3,0,184,0,244,0,105,0,71,0,30,0,180,0,211,0,58,0,125,0,87,0,106,0,71,0,153,0,84,0,105,0,9,0,40,0,0,0,182,0,197,0,154,0,193,0,151,0,191,0,102,0,24,0,203,0,240,0,56,0,10,0,0,0,35,0,216,0,40,0,85,0,0,0,32,0,172,0,202,0,0,0,0,0,179,0,0,0,112,0,0,0,31,0,20,0,35,0,159,0,118,0,253,0,253,0,249,0,224,0,0,0,145,0,166,0,0,0,0,0,163,0,90,0,163,0,113,0,42,0,175,0,0,0,0,0,0,0,42,0,63,0,0,0,0,0,31,0,215,0,173,0,33,0,177,0,90,0,118,0,18,0,21,0,243,0,0,0,13,0,123,0,204,0,234,0,0,0,229,0,0,0,104,0,87,0,0,0,10,0,67,0,43,0,0,0,50,0,0,0,162,0,0,0,166,0,254,0,31,0,227,0,0,0,207,0,234,0,95,0,72,0,233,0,207,0,209,0,50,0,192,0,0,0,0,0,0,0,142,0,0,0,19,0,81,0,68,0,0,0,253,0,124,0,0,0,0,0,173,0,251,0,233,0,0,0,161,0,0,0,68,0,234,0,0,0,77,0,0,0,159,0,161,0,210,0,0,0,110,0,0,0,120,0,93,0,12,0,253,0,111,0,217,0,137,0,229,0,0,0,0,0,43,0,0,0,69,0,156,0,219,0,59,0,0,0,0,0,160,0,40,0,193,0,240,0,8,0,0,0,100,0,103,0,37,0,212,0,215,0,212,0,132,0,32,0,70,0,80,0,150,0,91,0,56,0,68,0,45,0,0,0,211,0,130,0,0,0,0,0,47,0,0,0,4,0,166,0,242,0,30,0,39,0,230,0,158,0,3,0,0,0,162,0,72,0,176,0,203,0,18,0,127,0,0,0,0,0,202,0,42,0,198,0,231,0,39,0,0,0,0,0,169,0,191,0,165,0,24,0,178,0,104,0,55,0,241,0,81,0,110,0,154,0,133,0,0,0,28,0,145,0,206,0,110,0,240,0,0,0,172,0,31,0,37,0,0,0,84,0,0,0,136,0,0,0,142,0,103,0,121,0,37,0,101,0,0,0,118,0,0,0,213,0,105,0,138,0,30,0,125,0,112,0,60,0,12,0,153,0,179,0,0,0,207,0,182,0,81,0,136,0,178,0,0,0,113,0,0,0,7,0,51,0,0,0,73,0,25,0,187,0,234,0,0,0,0,0,166,0,11,0,24,0,0,0,191,0,127,0,0,0,48,0,0,0,32,0,232,0,245,0,89,0,91,0,83,0,47,0,191,0,103,0,191,0,150,0,186,0,171,0,116,0,117,0,25,0,112,0,156,0,34,0,141,0,9,0,89,0,20,0,124,0,230,0,195,0,48,0,163,0,0,0,117,0,250,0,200,0,0,0,0,0,11,0,0,0,220,0,171,0,49,0,229,0,0,0,158,0,0,0,0,0,24,0,31,0,117,0,255,0,0,0,98,0,189,0,55,0,104,0,0,0,65,0,55,0,173,0,0,0,103,0,0,0,106,0,211,0,187,0,172,0,163,0,126,0,132,0,80,0,0,0,170,0,50,0,75,0,137,0,209,0,132,0,0,0,208,0,42,0,57,0,102,0,47,0,170,0,88,0,0,0,0,0,132,0,0,0,241,0,214,0,0,0,199,0,120,0,204,0,215,0,52,0,0,0,78,0,48,0,218,0,152,0,0,0,0,0,234,0,65,0,94,0,146,0,222,0,0,0,73,0,192,0,4,0,0,0,0,0,128,0,230,0,207,0,0,0,43,0,167,0,56,0,231,0,239,0,31,0,145,0,110,0,172,0,235,0,88,0,0,0,207,0,0,0,239,0,111,0,56,0,234,0,226,0,185,0,84,0,41,0,0,0,148,0,127,0,160,0,0,0,64,0,65,0,221,0,164,0,243,0,221,0,0,0,132,0,9,0,236,0,32,0,139,0,23,0,0,0,228,0,171,0,169,0,0,0,145,0,207,0,77,0,0,0,195,0,195,0,88,0,216,0,70,0,150,0,198,0,5,0,0,0,172,0,0,0,91,0,0,0,188,0,189,0,60,0,184,0,80,0,0,0,139,0,0,0,0,0,0,0,124,0,0,0,251,0,15,0,172,0,114,0,143,0,117,0,247,0,143,0,94,0,0,0,152,0,217,0,241,0,3,0,0,0,129,0,0,0,229,0,118,0,0,0,113,0,65,0,0,0,53,0,136,0,56,0,0,0,0,0,228,0,0,0,33,0,0,0,0,0,0,0,35,0,8,0,138,0,244,0,239,0,22,0,85,0,244,0,6,0,187,0,67,0,174,0,220,0,159,0,0,0,171,0,14,0,66,0,0,0,202,0,59,0,208,0,230,0,150,0,197,0,44,0,225,0,95,0,10,0,38,0,8,0,186,0,170,0,0,0,0,0,0,0,0,0,151,0,121,0,135,0,4,0,22,0,69,0,180,0,210,0,254,0,99,0,185,0,105,0,19,0,184,0,245,0,0,0,141,0,0,0,0,0,78,0,172,0,91,0,0,0,19,0,152,0,135,0,91,0,109,0,84,0,249,0,120,0,94,0,199,0,101,0,26,0,240,0,0,0,0,0,1,0,142,0,172,0,0,0,0,0,0,0,206,0,107,0,226,0,210,0,221,0,17,0,211,0,251,0,111,0,114,0,0,0,19,0,0,0,0,0,87,0,173,0,117,0,145,0,6,0,12,0,61,0,0,0,97,0,97,0,66,0,0,0,102,0,110,0,58,0,160,0,174,0,0,0,0,0,153,0,219,0,0,0,26,0,17,0,217,0,215,0,200,0,0,0,50,0,0,0,194,0,40,0,253,0,104,0,14,0,0,0,159,0,57,0,179,0,250,0,0,0,21,0,107,0,68,0,155,0,191,0,210,0,234,0,179,0,84,0,62,0,228,0,202,0,144,0,165,0,50,0,133,0,0,0,148,0,0,0,0,0,210,0,68,0,33,0,49,0,200,0,0,0,133,0,0,0,210,0,0,0,148,0,2,0,45,0,0,0,0,0,103,0,236,0,167,0,0,0,255,0,71,0,0,0,78,0,75,0,0,0,50,0,191,0,28,0,79,0,117,0,214,0,196,0,154,0,72,0,191,0,227,0,134,0,102,0,205,0,204,0,0,0,192,0,17,0,165,0,30,0,122,0,0,0,171,0,170,0,225,0,0,0,0,0,78,0,26,0,13,0,105,0,0,0,62,0,72,0,35,0,135,0,102,0,193,0,129,0,214,0,62,0,32,0,41,0,217,0,9,0,126,0,159,0,134,0,202,0,54,0,0,0,115,0,235,0,0,0,12,0,210,0,248,0,85,0,14,0,51,0,199,0,137,0,156,0,88,0,82,0,248,0,59,0,138,0,1,0,111,0,233,0,95,0,218,0,0,0,100,0,122,0,181,0,134,0,17,0,185,0,46,0,237,0,0,0,39,0,164,0,61,0,215,0,37,0,44,0,129,0,10,0,239,0,86,0,27,0,143,0,14,0,20,0,0,0,0,0,212,0,235,0,128,0,129,0,0,0,241,0,168,0,0,0,194,0,206,0,156,0,0,0,12,0,33,0,81,0,183,0,240,0,253,0,132,0,14,0,9,0,0,0);
signal scenario_full  : scenario_type := (39,31,39,30,239,31,30,31,30,30,156,31,156,30,156,29,183,31,183,30,111,31,111,30,168,31,240,31,79,31,106,31,109,31,229,31,229,30,239,31,154,31,154,30,3,31,184,31,244,31,105,31,71,31,30,31,180,31,211,31,58,31,125,31,87,31,106,31,71,31,153,31,84,31,105,31,9,31,40,31,40,30,182,31,197,31,154,31,193,31,151,31,191,31,102,31,24,31,203,31,240,31,56,31,10,31,10,30,35,31,216,31,40,31,85,31,85,30,32,31,172,31,202,31,202,30,202,29,179,31,179,30,112,31,112,30,31,31,20,31,35,31,159,31,118,31,253,31,253,31,249,31,224,31,224,30,145,31,166,31,166,30,166,29,163,31,90,31,163,31,113,31,42,31,175,31,175,30,175,29,175,28,42,31,63,31,63,30,63,29,31,31,215,31,173,31,33,31,177,31,90,31,118,31,18,31,21,31,243,31,243,30,13,31,123,31,204,31,234,31,234,30,229,31,229,30,104,31,87,31,87,30,10,31,67,31,43,31,43,30,50,31,50,30,162,31,162,30,166,31,254,31,31,31,227,31,227,30,207,31,234,31,95,31,72,31,233,31,207,31,209,31,50,31,192,31,192,30,192,29,192,28,142,31,142,30,19,31,81,31,68,31,68,30,253,31,124,31,124,30,124,29,173,31,251,31,233,31,233,30,161,31,161,30,68,31,234,31,234,30,77,31,77,30,159,31,161,31,210,31,210,30,110,31,110,30,120,31,93,31,12,31,253,31,111,31,217,31,137,31,229,31,229,30,229,29,43,31,43,30,69,31,156,31,219,31,59,31,59,30,59,29,160,31,40,31,193,31,240,31,8,31,8,30,100,31,103,31,37,31,212,31,215,31,212,31,132,31,32,31,70,31,80,31,150,31,91,31,56,31,68,31,45,31,45,30,211,31,130,31,130,30,130,29,47,31,47,30,4,31,166,31,242,31,30,31,39,31,230,31,158,31,3,31,3,30,162,31,72,31,176,31,203,31,18,31,127,31,127,30,127,29,202,31,42,31,198,31,231,31,39,31,39,30,39,29,169,31,191,31,165,31,24,31,178,31,104,31,55,31,241,31,81,31,110,31,154,31,133,31,133,30,28,31,145,31,206,31,110,31,240,31,240,30,172,31,31,31,37,31,37,30,84,31,84,30,136,31,136,30,142,31,103,31,121,31,37,31,101,31,101,30,118,31,118,30,213,31,105,31,138,31,30,31,125,31,112,31,60,31,12,31,153,31,179,31,179,30,207,31,182,31,81,31,136,31,178,31,178,30,113,31,113,30,7,31,51,31,51,30,73,31,25,31,187,31,234,31,234,30,234,29,166,31,11,31,24,31,24,30,191,31,127,31,127,30,48,31,48,30,32,31,232,31,245,31,89,31,91,31,83,31,47,31,191,31,103,31,191,31,150,31,186,31,171,31,116,31,117,31,25,31,112,31,156,31,34,31,141,31,9,31,89,31,20,31,124,31,230,31,195,31,48,31,163,31,163,30,117,31,250,31,200,31,200,30,200,29,11,31,11,30,220,31,171,31,49,31,229,31,229,30,158,31,158,30,158,29,24,31,31,31,117,31,255,31,255,30,98,31,189,31,55,31,104,31,104,30,65,31,55,31,173,31,173,30,103,31,103,30,106,31,211,31,187,31,172,31,163,31,126,31,132,31,80,31,80,30,170,31,50,31,75,31,137,31,209,31,132,31,132,30,208,31,42,31,57,31,102,31,47,31,170,31,88,31,88,30,88,29,132,31,132,30,241,31,214,31,214,30,199,31,120,31,204,31,215,31,52,31,52,30,78,31,48,31,218,31,152,31,152,30,152,29,234,31,65,31,94,31,146,31,222,31,222,30,73,31,192,31,4,31,4,30,4,29,128,31,230,31,207,31,207,30,43,31,167,31,56,31,231,31,239,31,31,31,145,31,110,31,172,31,235,31,88,31,88,30,207,31,207,30,239,31,111,31,56,31,234,31,226,31,185,31,84,31,41,31,41,30,148,31,127,31,160,31,160,30,64,31,65,31,221,31,164,31,243,31,221,31,221,30,132,31,9,31,236,31,32,31,139,31,23,31,23,30,228,31,171,31,169,31,169,30,145,31,207,31,77,31,77,30,195,31,195,31,88,31,216,31,70,31,150,31,198,31,5,31,5,30,172,31,172,30,91,31,91,30,188,31,189,31,60,31,184,31,80,31,80,30,139,31,139,30,139,29,139,28,124,31,124,30,251,31,15,31,172,31,114,31,143,31,117,31,247,31,143,31,94,31,94,30,152,31,217,31,241,31,3,31,3,30,129,31,129,30,229,31,118,31,118,30,113,31,65,31,65,30,53,31,136,31,56,31,56,30,56,29,228,31,228,30,33,31,33,30,33,29,33,28,35,31,8,31,138,31,244,31,239,31,22,31,85,31,244,31,6,31,187,31,67,31,174,31,220,31,159,31,159,30,171,31,14,31,66,31,66,30,202,31,59,31,208,31,230,31,150,31,197,31,44,31,225,31,95,31,10,31,38,31,8,31,186,31,170,31,170,30,170,29,170,28,170,27,151,31,121,31,135,31,4,31,22,31,69,31,180,31,210,31,254,31,99,31,185,31,105,31,19,31,184,31,245,31,245,30,141,31,141,30,141,29,78,31,172,31,91,31,91,30,19,31,152,31,135,31,91,31,109,31,84,31,249,31,120,31,94,31,199,31,101,31,26,31,240,31,240,30,240,29,1,31,142,31,172,31,172,30,172,29,172,28,206,31,107,31,226,31,210,31,221,31,17,31,211,31,251,31,111,31,114,31,114,30,19,31,19,30,19,29,87,31,173,31,117,31,145,31,6,31,12,31,61,31,61,30,97,31,97,31,66,31,66,30,102,31,110,31,58,31,160,31,174,31,174,30,174,29,153,31,219,31,219,30,26,31,17,31,217,31,215,31,200,31,200,30,50,31,50,30,194,31,40,31,253,31,104,31,14,31,14,30,159,31,57,31,179,31,250,31,250,30,21,31,107,31,68,31,155,31,191,31,210,31,234,31,179,31,84,31,62,31,228,31,202,31,144,31,165,31,50,31,133,31,133,30,148,31,148,30,148,29,210,31,68,31,33,31,49,31,200,31,200,30,133,31,133,30,210,31,210,30,148,31,2,31,45,31,45,30,45,29,103,31,236,31,167,31,167,30,255,31,71,31,71,30,78,31,75,31,75,30,50,31,191,31,28,31,79,31,117,31,214,31,196,31,154,31,72,31,191,31,227,31,134,31,102,31,205,31,204,31,204,30,192,31,17,31,165,31,30,31,122,31,122,30,171,31,170,31,225,31,225,30,225,29,78,31,26,31,13,31,105,31,105,30,62,31,72,31,35,31,135,31,102,31,193,31,129,31,214,31,62,31,32,31,41,31,217,31,9,31,126,31,159,31,134,31,202,31,54,31,54,30,115,31,235,31,235,30,12,31,210,31,248,31,85,31,14,31,51,31,199,31,137,31,156,31,88,31,82,31,248,31,59,31,138,31,1,31,111,31,233,31,95,31,218,31,218,30,100,31,122,31,181,31,134,31,17,31,185,31,46,31,237,31,237,30,39,31,164,31,61,31,215,31,37,31,44,31,129,31,10,31,239,31,86,31,27,31,143,31,14,31,20,31,20,30,20,29,212,31,235,31,128,31,129,31,129,30,241,31,168,31,168,30,194,31,206,31,156,31,156,30,12,31,33,31,81,31,183,31,240,31,253,31,132,31,14,31,9,31,9,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
