-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_656 is
end project_tb_656;

architecture project_tb_arch_656 of project_tb_656 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 755;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,0,0,95,0,166,0,0,0,0,0,242,0,90,0,73,0,167,0,29,0,244,0,178,0,222,0,0,0,139,0,75,0,101,0,0,0,128,0,89,0,118,0,17,0,39,0,162,0,7,0,156,0,0,0,0,0,123,0,169,0,32,0,6,0,12,0,145,0,183,0,130,0,220,0,38,0,114,0,41,0,130,0,0,0,126,0,0,0,166,0,99,0,0,0,9,0,250,0,155,0,92,0,189,0,231,0,0,0,247,0,0,0,176,0,95,0,19,0,156,0,197,0,0,0,239,0,121,0,0,0,74,0,107,0,144,0,252,0,0,0,156,0,221,0,154,0,207,0,33,0,23,0,16,0,0,0,84,0,10,0,0,0,27,0,195,0,0,0,8,0,0,0,0,0,133,0,0,0,163,0,47,0,173,0,11,0,50,0,141,0,11,0,0,0,0,0,18,0,165,0,133,0,46,0,0,0,66,0,197,0,22,0,79,0,65,0,225,0,0,0,0,0,0,0,0,0,226,0,124,0,67,0,148,0,0,0,209,0,0,0,0,0,83,0,192,0,171,0,175,0,0,0,104,0,233,0,30,0,209,0,0,0,7,0,245,0,0,0,204,0,64,0,81,0,36,0,21,0,8,0,182,0,0,0,105,0,97,0,39,0,139,0,0,0,0,0,105,0,13,0,212,0,63,0,12,0,0,0,241,0,72,0,41,0,0,0,222,0,0,0,39,0,122,0,255,0,255,0,0,0,170,0,162,0,47,0,0,0,103,0,144,0,163,0,112,0,142,0,154,0,184,0,38,0,0,0,0,0,44,0,5,0,0,0,251,0,209,0,91,0,136,0,98,0,0,0,0,0,218,0,71,0,72,0,0,0,200,0,138,0,77,0,165,0,67,0,0,0,157,0,57,0,65,0,37,0,32,0,0,0,190,0,0,0,0,0,0,0,0,0,41,0,116,0,174,0,0,0,163,0,244,0,0,0,166,0,18,0,29,0,126,0,90,0,186,0,0,0,90,0,108,0,0,0,174,0,245,0,102,0,72,0,176,0,77,0,39,0,224,0,223,0,225,0,168,0,0,0,6,0,142,0,92,0,0,0,55,0,0,0,0,0,110,0,0,0,243,0,243,0,182,0,184,0,204,0,173,0,67,0,218,0,159,0,36,0,207,0,131,0,46,0,0,0,0,0,190,0,134,0,0,0,0,0,0,0,54,0,218,0,62,0,0,0,220,0,0,0,0,0,116,0,126,0,154,0,116,0,5,0,47,0,111,0,66,0,0,0,63,0,111,0,32,0,136,0,74,0,232,0,189,0,139,0,41,0,24,0,232,0,59,0,59,0,48,0,106,0,90,0,18,0,210,0,69,0,113,0,96,0,120,0,0,0,73,0,0,0,135,0,95,0,2,0,226,0,246,0,104,0,172,0,149,0,116,0,176,0,215,0,58,0,183,0,195,0,0,0,49,0,58,0,0,0,52,0,55,0,193,0,0,0,138,0,15,0,75,0,223,0,164,0,208,0,13,0,175,0,211,0,114,0,76,0,16,0,215,0,158,0,189,0,99,0,130,0,0,0,43,0,48,0,102,0,125,0,229,0,191,0,113,0,0,0,0,0,142,0,25,0,201,0,194,0,172,0,0,0,210,0,21,0,0,0,235,0,151,0,157,0,148,0,24,0,0,0,156,0,136,0,39,0,0,0,0,0,209,0,0,0,180,0,237,0,192,0,222,0,88,0,192,0,0,0,0,0,0,0,188,0,27,0,67,0,232,0,75,0,54,0,14,0,163,0,6,0,245,0,186,0,0,0,183,0,216,0,33,0,0,0,89,0,122,0,0,0,0,0,217,0,171,0,213,0,119,0,0,0,252,0,5,0,108,0,88,0,155,0,104,0,44,0,40,0,66,0,242,0,25,0,119,0,121,0,12,0,191,0,69,0,0,0,138,0,162,0,69,0,204,0,59,0,0,0,34,0,195,0,22,0,0,0,202,0,178,0,0,0,165,0,196,0,242,0,59,0,0,0,0,0,204,0,8,0,96,0,200,0,0,0,70,0,211,0,104,0,0,0,143,0,8,0,0,0,157,0,226,0,187,0,73,0,41,0,101,0,129,0,0,0,0,0,126,0,24,0,88,0,128,0,77,0,250,0,114,0,130,0,54,0,69,0,0,0,91,0,0,0,124,0,245,0,75,0,49,0,57,0,12,0,85,0,215,0,239,0,44,0,230,0,204,0,230,0,142,0,42,0,183,0,164,0,227,0,98,0,141,0,92,0,42,0,2,0,26,0,131,0,0,0,81,0,26,0,151,0,0,0,154,0,0,0,132,0,85,0,0,0,0,0,44,0,10,0,197,0,197,0,123,0,58,0,82,0,163,0,31,0,39,0,60,0,2,0,0,0,0,0,51,0,189,0,33,0,31,0,164,0,148,0,136,0,130,0,168,0,59,0,60,0,190,0,15,0,0,0,17,0,81,0,84,0,164,0,144,0,88,0,75,0,25,0,23,0,211,0,132,0,15,0,188,0,0,0,229,0,215,0,74,0,154,0,0,0,181,0,191,0,0,0,251,0,222,0,106,0,132,0,196,0,66,0,207,0,0,0,191,0,160,0,141,0,18,0,220,0,250,0,112,0,99,0,0,0,234,0,158,0,255,0,128,0,0,0,238,0,141,0,8,0,231,0,90,0,248,0,245,0,38,0,48,0,180,0,229,0,95,0,0,0,182,0,133,0,28,0,153,0,148,0,207,0,161,0,185,0,0,0,3,0,146,0,26,0,15,0,45,0,156,0,246,0,178,0,0,0,38,0,199,0,39,0,254,0,196,0,160,0,93,0,21,0,216,0,44,0,85,0,196,0,134,0,211,0,106,0,219,0,190,0,0,0,53,0,172,0,0,0,85,0,3,0,0,0,32,0,0,0,0,0,124,0,190,0,107,0,70,0,73,0,228,0,83,0,208,0,0,0,214,0,220,0,86,0,30,0,182,0,214,0,182,0,166,0,70,0,94,0,39,0,58,0,239,0,200,0,16,0,194,0,211,0,108,0,61,0,22,0,175,0,171,0,60,0,68,0,250,0,0,0,52,0,58,0,60,0,134,0,245,0,125,0,94,0,167,0,74,0,0,0,171,0,0,0,0,0,13,0,37,0,84,0,0,0,155,0,55,0,168,0,212,0,32,0,143,0,218,0,181,0,0,0,254,0,114,0,238,0,52,0,199,0,241,0,8,0,138,0,104,0,121,0,21,0,46,0,0,0,213,0,0,0,51,0,8,0,54,0,31,0,211,0,164,0,204,0,92,0,0,0,125,0,182,0,90,0,205,0,0,0,39,0,0,0,184,0,0,0,156,0,155,0,172,0,24,0,0,0,83,0,65,0,194,0,48,0,12,0);
signal scenario_full  : scenario_type := (68,31,68,30,95,31,166,31,166,30,166,29,242,31,90,31,73,31,167,31,29,31,244,31,178,31,222,31,222,30,139,31,75,31,101,31,101,30,128,31,89,31,118,31,17,31,39,31,162,31,7,31,156,31,156,30,156,29,123,31,169,31,32,31,6,31,12,31,145,31,183,31,130,31,220,31,38,31,114,31,41,31,130,31,130,30,126,31,126,30,166,31,99,31,99,30,9,31,250,31,155,31,92,31,189,31,231,31,231,30,247,31,247,30,176,31,95,31,19,31,156,31,197,31,197,30,239,31,121,31,121,30,74,31,107,31,144,31,252,31,252,30,156,31,221,31,154,31,207,31,33,31,23,31,16,31,16,30,84,31,10,31,10,30,27,31,195,31,195,30,8,31,8,30,8,29,133,31,133,30,163,31,47,31,173,31,11,31,50,31,141,31,11,31,11,30,11,29,18,31,165,31,133,31,46,31,46,30,66,31,197,31,22,31,79,31,65,31,225,31,225,30,225,29,225,28,225,27,226,31,124,31,67,31,148,31,148,30,209,31,209,30,209,29,83,31,192,31,171,31,175,31,175,30,104,31,233,31,30,31,209,31,209,30,7,31,245,31,245,30,204,31,64,31,81,31,36,31,21,31,8,31,182,31,182,30,105,31,97,31,39,31,139,31,139,30,139,29,105,31,13,31,212,31,63,31,12,31,12,30,241,31,72,31,41,31,41,30,222,31,222,30,39,31,122,31,255,31,255,31,255,30,170,31,162,31,47,31,47,30,103,31,144,31,163,31,112,31,142,31,154,31,184,31,38,31,38,30,38,29,44,31,5,31,5,30,251,31,209,31,91,31,136,31,98,31,98,30,98,29,218,31,71,31,72,31,72,30,200,31,138,31,77,31,165,31,67,31,67,30,157,31,57,31,65,31,37,31,32,31,32,30,190,31,190,30,190,29,190,28,190,27,41,31,116,31,174,31,174,30,163,31,244,31,244,30,166,31,18,31,29,31,126,31,90,31,186,31,186,30,90,31,108,31,108,30,174,31,245,31,102,31,72,31,176,31,77,31,39,31,224,31,223,31,225,31,168,31,168,30,6,31,142,31,92,31,92,30,55,31,55,30,55,29,110,31,110,30,243,31,243,31,182,31,184,31,204,31,173,31,67,31,218,31,159,31,36,31,207,31,131,31,46,31,46,30,46,29,190,31,134,31,134,30,134,29,134,28,54,31,218,31,62,31,62,30,220,31,220,30,220,29,116,31,126,31,154,31,116,31,5,31,47,31,111,31,66,31,66,30,63,31,111,31,32,31,136,31,74,31,232,31,189,31,139,31,41,31,24,31,232,31,59,31,59,31,48,31,106,31,90,31,18,31,210,31,69,31,113,31,96,31,120,31,120,30,73,31,73,30,135,31,95,31,2,31,226,31,246,31,104,31,172,31,149,31,116,31,176,31,215,31,58,31,183,31,195,31,195,30,49,31,58,31,58,30,52,31,55,31,193,31,193,30,138,31,15,31,75,31,223,31,164,31,208,31,13,31,175,31,211,31,114,31,76,31,16,31,215,31,158,31,189,31,99,31,130,31,130,30,43,31,48,31,102,31,125,31,229,31,191,31,113,31,113,30,113,29,142,31,25,31,201,31,194,31,172,31,172,30,210,31,21,31,21,30,235,31,151,31,157,31,148,31,24,31,24,30,156,31,136,31,39,31,39,30,39,29,209,31,209,30,180,31,237,31,192,31,222,31,88,31,192,31,192,30,192,29,192,28,188,31,27,31,67,31,232,31,75,31,54,31,14,31,163,31,6,31,245,31,186,31,186,30,183,31,216,31,33,31,33,30,89,31,122,31,122,30,122,29,217,31,171,31,213,31,119,31,119,30,252,31,5,31,108,31,88,31,155,31,104,31,44,31,40,31,66,31,242,31,25,31,119,31,121,31,12,31,191,31,69,31,69,30,138,31,162,31,69,31,204,31,59,31,59,30,34,31,195,31,22,31,22,30,202,31,178,31,178,30,165,31,196,31,242,31,59,31,59,30,59,29,204,31,8,31,96,31,200,31,200,30,70,31,211,31,104,31,104,30,143,31,8,31,8,30,157,31,226,31,187,31,73,31,41,31,101,31,129,31,129,30,129,29,126,31,24,31,88,31,128,31,77,31,250,31,114,31,130,31,54,31,69,31,69,30,91,31,91,30,124,31,245,31,75,31,49,31,57,31,12,31,85,31,215,31,239,31,44,31,230,31,204,31,230,31,142,31,42,31,183,31,164,31,227,31,98,31,141,31,92,31,42,31,2,31,26,31,131,31,131,30,81,31,26,31,151,31,151,30,154,31,154,30,132,31,85,31,85,30,85,29,44,31,10,31,197,31,197,31,123,31,58,31,82,31,163,31,31,31,39,31,60,31,2,31,2,30,2,29,51,31,189,31,33,31,31,31,164,31,148,31,136,31,130,31,168,31,59,31,60,31,190,31,15,31,15,30,17,31,81,31,84,31,164,31,144,31,88,31,75,31,25,31,23,31,211,31,132,31,15,31,188,31,188,30,229,31,215,31,74,31,154,31,154,30,181,31,191,31,191,30,251,31,222,31,106,31,132,31,196,31,66,31,207,31,207,30,191,31,160,31,141,31,18,31,220,31,250,31,112,31,99,31,99,30,234,31,158,31,255,31,128,31,128,30,238,31,141,31,8,31,231,31,90,31,248,31,245,31,38,31,48,31,180,31,229,31,95,31,95,30,182,31,133,31,28,31,153,31,148,31,207,31,161,31,185,31,185,30,3,31,146,31,26,31,15,31,45,31,156,31,246,31,178,31,178,30,38,31,199,31,39,31,254,31,196,31,160,31,93,31,21,31,216,31,44,31,85,31,196,31,134,31,211,31,106,31,219,31,190,31,190,30,53,31,172,31,172,30,85,31,3,31,3,30,32,31,32,30,32,29,124,31,190,31,107,31,70,31,73,31,228,31,83,31,208,31,208,30,214,31,220,31,86,31,30,31,182,31,214,31,182,31,166,31,70,31,94,31,39,31,58,31,239,31,200,31,16,31,194,31,211,31,108,31,61,31,22,31,175,31,171,31,60,31,68,31,250,31,250,30,52,31,58,31,60,31,134,31,245,31,125,31,94,31,167,31,74,31,74,30,171,31,171,30,171,29,13,31,37,31,84,31,84,30,155,31,55,31,168,31,212,31,32,31,143,31,218,31,181,31,181,30,254,31,114,31,238,31,52,31,199,31,241,31,8,31,138,31,104,31,121,31,21,31,46,31,46,30,213,31,213,30,51,31,8,31,54,31,31,31,211,31,164,31,204,31,92,31,92,30,125,31,182,31,90,31,205,31,205,30,39,31,39,30,184,31,184,30,156,31,155,31,172,31,24,31,24,30,83,31,65,31,194,31,48,31,12,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
