-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_833 is
end project_tb_833;

architecture project_tb_arch_833 of project_tb_833 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 460;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (187,0,178,0,132,0,45,0,65,0,90,0,7,0,183,0,28,0,91,0,0,0,193,0,6,0,112,0,55,0,32,0,111,0,0,0,0,0,0,0,0,0,30,0,56,0,83,0,32,0,229,0,124,0,79,0,40,0,204,0,9,0,229,0,95,0,203,0,5,0,0,0,98,0,0,0,0,0,17,0,73,0,36,0,0,0,46,0,145,0,6,0,115,0,237,0,51,0,178,0,93,0,61,0,198,0,95,0,243,0,96,0,121,0,0,0,119,0,229,0,217,0,128,0,80,0,67,0,0,0,200,0,0,0,0,0,226,0,0,0,193,0,225,0,20,0,28,0,21,0,138,0,92,0,1,0,78,0,13,0,0,0,0,0,26,0,133,0,221,0,35,0,0,0,185,0,9,0,244,0,171,0,0,0,223,0,45,0,61,0,202,0,67,0,52,0,188,0,233,0,86,0,80,0,36,0,117,0,211,0,211,0,197,0,245,0,83,0,0,0,135,0,190,0,26,0,0,0,186,0,170,0,0,0,72,0,176,0,151,0,0,0,0,0,245,0,0,0,0,0,0,0,0,0,36,0,102,0,73,0,163,0,113,0,0,0,110,0,112,0,168,0,36,0,192,0,199,0,167,0,206,0,0,0,203,0,226,0,0,0,225,0,124,0,143,0,161,0,7,0,169,0,244,0,194,0,0,0,112,0,81,0,0,0,104,0,194,0,89,0,196,0,222,0,0,0,120,0,14,0,66,0,104,0,17,0,149,0,0,0,190,0,148,0,0,0,87,0,250,0,205,0,0,0,62,0,20,0,142,0,69,0,74,0,208,0,61,0,0,0,0,0,203,0,179,0,223,0,56,0,48,0,0,0,89,0,12,0,192,0,58,0,86,0,201,0,15,0,0,0,0,0,246,0,100,0,63,0,0,0,0,0,0,0,71,0,109,0,53,0,45,0,144,0,155,0,0,0,0,0,238,0,86,0,237,0,119,0,217,0,0,0,186,0,0,0,26,0,87,0,230,0,251,0,196,0,56,0,253,0,22,0,23,0,86,0,14,0,186,0,103,0,0,0,0,0,164,0,137,0,0,0,0,0,172,0,47,0,97,0,138,0,21,0,29,0,207,0,161,0,251,0,180,0,232,0,220,0,208,0,90,0,219,0,116,0,249,0,0,0,37,0,38,0,20,0,232,0,249,0,118,0,203,0,162,0,93,0,0,0,174,0,205,0,202,0,32,0,0,0,0,0,9,0,195,0,0,0,214,0,177,0,121,0,116,0,0,0,193,0,0,0,189,0,219,0,75,0,124,0,156,0,116,0,0,0,19,0,177,0,20,0,89,0,0,0,183,0,84,0,251,0,192,0,45,0,36,0,0,0,150,0,169,0,0,0,0,0,50,0,250,0,148,0,104,0,0,0,162,0,101,0,54,0,242,0,252,0,184,0,0,0,22,0,0,0,34,0,166,0,190,0,0,0,200,0,0,0,125,0,111,0,4,0,96,0,46,0,140,0,125,0,155,0,253,0,0,0,0,0,156,0,187,0,124,0,59,0,7,0,234,0,167,0,48,0,149,0,255,0,82,0,211,0,126,0,44,0,95,0,25,0,15,0,41,0,0,0,0,0,0,0,241,0,223,0,29,0,209,0,152,0,149,0,178,0,26,0,174,0,189,0,224,0,91,0,0,0,0,0,45,0,29,0,46,0,20,0,0,0,4,0,9,0,0,0,214,0,249,0,0,0,0,0,0,0,99,0,27,0,161,0,120,0,29,0,101,0,0,0,120,0,0,0,2,0,0,0,188,0,0,0,172,0,239,0,141,0,120,0,22,0,176,0,10,0,115,0,26,0,129,0,209,0,110,0,0,0,128,0,95,0,0,0,0,0,125,0,19,0,34,0,201,0,215,0,248,0,53,0,88,0,183,0,90,0,0,0,0,0,0,0,38,0,192,0,11,0,169,0,36,0,0,0,146,0,0,0,183,0,0,0,4,0,133,0,230,0,50,0,82,0,188,0,76,0,187,0,169,0,23,0,38,0,0,0,204,0,93,0,0,0,1,0,150,0,154,0,0,0);
signal scenario_full  : scenario_type := (187,31,178,31,132,31,45,31,65,31,90,31,7,31,183,31,28,31,91,31,91,30,193,31,6,31,112,31,55,31,32,31,111,31,111,30,111,29,111,28,111,27,30,31,56,31,83,31,32,31,229,31,124,31,79,31,40,31,204,31,9,31,229,31,95,31,203,31,5,31,5,30,98,31,98,30,98,29,17,31,73,31,36,31,36,30,46,31,145,31,6,31,115,31,237,31,51,31,178,31,93,31,61,31,198,31,95,31,243,31,96,31,121,31,121,30,119,31,229,31,217,31,128,31,80,31,67,31,67,30,200,31,200,30,200,29,226,31,226,30,193,31,225,31,20,31,28,31,21,31,138,31,92,31,1,31,78,31,13,31,13,30,13,29,26,31,133,31,221,31,35,31,35,30,185,31,9,31,244,31,171,31,171,30,223,31,45,31,61,31,202,31,67,31,52,31,188,31,233,31,86,31,80,31,36,31,117,31,211,31,211,31,197,31,245,31,83,31,83,30,135,31,190,31,26,31,26,30,186,31,170,31,170,30,72,31,176,31,151,31,151,30,151,29,245,31,245,30,245,29,245,28,245,27,36,31,102,31,73,31,163,31,113,31,113,30,110,31,112,31,168,31,36,31,192,31,199,31,167,31,206,31,206,30,203,31,226,31,226,30,225,31,124,31,143,31,161,31,7,31,169,31,244,31,194,31,194,30,112,31,81,31,81,30,104,31,194,31,89,31,196,31,222,31,222,30,120,31,14,31,66,31,104,31,17,31,149,31,149,30,190,31,148,31,148,30,87,31,250,31,205,31,205,30,62,31,20,31,142,31,69,31,74,31,208,31,61,31,61,30,61,29,203,31,179,31,223,31,56,31,48,31,48,30,89,31,12,31,192,31,58,31,86,31,201,31,15,31,15,30,15,29,246,31,100,31,63,31,63,30,63,29,63,28,71,31,109,31,53,31,45,31,144,31,155,31,155,30,155,29,238,31,86,31,237,31,119,31,217,31,217,30,186,31,186,30,26,31,87,31,230,31,251,31,196,31,56,31,253,31,22,31,23,31,86,31,14,31,186,31,103,31,103,30,103,29,164,31,137,31,137,30,137,29,172,31,47,31,97,31,138,31,21,31,29,31,207,31,161,31,251,31,180,31,232,31,220,31,208,31,90,31,219,31,116,31,249,31,249,30,37,31,38,31,20,31,232,31,249,31,118,31,203,31,162,31,93,31,93,30,174,31,205,31,202,31,32,31,32,30,32,29,9,31,195,31,195,30,214,31,177,31,121,31,116,31,116,30,193,31,193,30,189,31,219,31,75,31,124,31,156,31,116,31,116,30,19,31,177,31,20,31,89,31,89,30,183,31,84,31,251,31,192,31,45,31,36,31,36,30,150,31,169,31,169,30,169,29,50,31,250,31,148,31,104,31,104,30,162,31,101,31,54,31,242,31,252,31,184,31,184,30,22,31,22,30,34,31,166,31,190,31,190,30,200,31,200,30,125,31,111,31,4,31,96,31,46,31,140,31,125,31,155,31,253,31,253,30,253,29,156,31,187,31,124,31,59,31,7,31,234,31,167,31,48,31,149,31,255,31,82,31,211,31,126,31,44,31,95,31,25,31,15,31,41,31,41,30,41,29,41,28,241,31,223,31,29,31,209,31,152,31,149,31,178,31,26,31,174,31,189,31,224,31,91,31,91,30,91,29,45,31,29,31,46,31,20,31,20,30,4,31,9,31,9,30,214,31,249,31,249,30,249,29,249,28,99,31,27,31,161,31,120,31,29,31,101,31,101,30,120,31,120,30,2,31,2,30,188,31,188,30,172,31,239,31,141,31,120,31,22,31,176,31,10,31,115,31,26,31,129,31,209,31,110,31,110,30,128,31,95,31,95,30,95,29,125,31,19,31,34,31,201,31,215,31,248,31,53,31,88,31,183,31,90,31,90,30,90,29,90,28,38,31,192,31,11,31,169,31,36,31,36,30,146,31,146,30,183,31,183,30,4,31,133,31,230,31,50,31,82,31,188,31,76,31,187,31,169,31,23,31,38,31,38,30,204,31,93,31,93,30,1,31,150,31,154,31,154,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
