-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 297;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,82,0,247,0,75,0,245,0,0,0,35,0,148,0,158,0,165,0,0,0,58,0,36,0,228,0,1,0,0,0,218,0,43,0,0,0,30,0,67,0,111,0,235,0,0,0,192,0,197,0,0,0,127,0,0,0,18,0,15,0,27,0,1,0,197,0,159,0,41,0,106,0,120,0,104,0,0,0,216,0,177,0,0,0,27,0,88,0,39,0,222,0,196,0,31,0,75,0,218,0,178,0,79,0,8,0,142,0,0,0,202,0,239,0,14,0,126,0,13,0,0,0,179,0,118,0,239,0,211,0,122,0,142,0,161,0,134,0,0,0,49,0,0,0,145,0,144,0,250,0,14,0,24,0,0,0,0,0,219,0,37,0,222,0,155,0,45,0,137,0,169,0,104,0,0,0,135,0,223,0,242,0,158,0,0,0,242,0,119,0,253,0,0,0,194,0,202,0,0,0,42,0,0,0,119,0,209,0,43,0,149,0,45,0,216,0,103,0,114,0,59,0,250,0,153,0,0,0,88,0,0,0,35,0,255,0,144,0,0,0,189,0,0,0,98,0,255,0,74,0,217,0,239,0,190,0,121,0,234,0,0,0,110,0,0,0,186,0,252,0,108,0,0,0,106,0,52,0,161,0,59,0,98,0,49,0,152,0,166,0,138,0,55,0,180,0,0,0,166,0,109,0,143,0,0,0,136,0,125,0,45,0,196,0,171,0,169,0,0,0,119,0,48,0,93,0,43,0,162,0,145,0,24,0,180,0,7,0,148,0,146,0,81,0,114,0,202,0,241,0,88,0,206,0,255,0,33,0,0,0,0,0,101,0,11,0,0,0,163,0,191,0,128,0,7,0,186,0,89,0,0,0,17,0,26,0,32,0,142,0,0,0,173,0,0,0,89,0,0,0,104,0,54,0,0,0,188,0,60,0,0,0,60,0,108,0,0,0,0,0,172,0,109,0,5,0,13,0,89,0,235,0,199,0,157,0,19,0,180,0,0,0,165,0,254,0,0,0,0,0,182,0,210,0,80,0,101,0,0,0,138,0,10,0,246,0,5,0,0,0,68,0,90,0,46,0,185,0,239,0,140,0,19,0,80,0,0,0,209,0,101,0,0,0,0,0,255,0,142,0,139,0,201,0,154,0,125,0,249,0,167,0,117,0,5,0,204,0,45,0,0,0,156,0,142,0,222,0,163,0,104,0,175,0,0,0,115,0,171,0,0,0,179,0,85,0,94,0,83,0,174,0,53,0,0,0,0,0,0,0,76,0,127,0,0,0,29,0,64,0,47,0,130,0,254,0,136,0,224,0,254,0,107,0,185,0,0,0,0,0,26,0);
signal scenario_full  : scenario_type := (0,0,82,31,247,31,75,31,245,31,245,30,35,31,148,31,158,31,165,31,165,30,58,31,36,31,228,31,1,31,1,30,218,31,43,31,43,30,30,31,67,31,111,31,235,31,235,30,192,31,197,31,197,30,127,31,127,30,18,31,15,31,27,31,1,31,197,31,159,31,41,31,106,31,120,31,104,31,104,30,216,31,177,31,177,30,27,31,88,31,39,31,222,31,196,31,31,31,75,31,218,31,178,31,79,31,8,31,142,31,142,30,202,31,239,31,14,31,126,31,13,31,13,30,179,31,118,31,239,31,211,31,122,31,142,31,161,31,134,31,134,30,49,31,49,30,145,31,144,31,250,31,14,31,24,31,24,30,24,29,219,31,37,31,222,31,155,31,45,31,137,31,169,31,104,31,104,30,135,31,223,31,242,31,158,31,158,30,242,31,119,31,253,31,253,30,194,31,202,31,202,30,42,31,42,30,119,31,209,31,43,31,149,31,45,31,216,31,103,31,114,31,59,31,250,31,153,31,153,30,88,31,88,30,35,31,255,31,144,31,144,30,189,31,189,30,98,31,255,31,74,31,217,31,239,31,190,31,121,31,234,31,234,30,110,31,110,30,186,31,252,31,108,31,108,30,106,31,52,31,161,31,59,31,98,31,49,31,152,31,166,31,138,31,55,31,180,31,180,30,166,31,109,31,143,31,143,30,136,31,125,31,45,31,196,31,171,31,169,31,169,30,119,31,48,31,93,31,43,31,162,31,145,31,24,31,180,31,7,31,148,31,146,31,81,31,114,31,202,31,241,31,88,31,206,31,255,31,33,31,33,30,33,29,101,31,11,31,11,30,163,31,191,31,128,31,7,31,186,31,89,31,89,30,17,31,26,31,32,31,142,31,142,30,173,31,173,30,89,31,89,30,104,31,54,31,54,30,188,31,60,31,60,30,60,31,108,31,108,30,108,29,172,31,109,31,5,31,13,31,89,31,235,31,199,31,157,31,19,31,180,31,180,30,165,31,254,31,254,30,254,29,182,31,210,31,80,31,101,31,101,30,138,31,10,31,246,31,5,31,5,30,68,31,90,31,46,31,185,31,239,31,140,31,19,31,80,31,80,30,209,31,101,31,101,30,101,29,255,31,142,31,139,31,201,31,154,31,125,31,249,31,167,31,117,31,5,31,204,31,45,31,45,30,156,31,142,31,222,31,163,31,104,31,175,31,175,30,115,31,171,31,171,30,179,31,85,31,94,31,83,31,174,31,53,31,53,30,53,29,53,28,76,31,127,31,127,30,29,31,64,31,47,31,130,31,254,31,136,31,224,31,254,31,107,31,185,31,185,30,185,29,26,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
