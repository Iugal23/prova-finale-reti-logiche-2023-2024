-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_896 is
end project_tb_896;

architecture project_tb_arch_896 of project_tb_896 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 658;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (99,0,245,0,154,0,0,0,0,0,0,0,127,0,231,0,32,0,190,0,215,0,0,0,85,0,192,0,140,0,192,0,148,0,15,0,0,0,0,0,208,0,151,0,161,0,0,0,181,0,64,0,29,0,31,0,73,0,0,0,62,0,226,0,22,0,228,0,101,0,145,0,120,0,98,0,221,0,15,0,0,0,47,0,10,0,163,0,14,0,54,0,247,0,0,0,0,0,81,0,137,0,62,0,55,0,192,0,223,0,0,0,92,0,0,0,201,0,0,0,121,0,250,0,233,0,193,0,68,0,73,0,90,0,66,0,12,0,125,0,0,0,82,0,55,0,250,0,0,0,113,0,231,0,119,0,155,0,49,0,119,0,91,0,73,0,54,0,0,0,0,0,148,0,210,0,34,0,148,0,57,0,0,0,0,0,144,0,143,0,148,0,0,0,0,0,199,0,207,0,214,0,103,0,46,0,7,0,0,0,15,0,0,0,0,0,182,0,58,0,206,0,131,0,104,0,103,0,0,0,28,0,160,0,86,0,17,0,190,0,147,0,181,0,113,0,235,0,0,0,141,0,0,0,94,0,88,0,164,0,121,0,0,0,8,0,235,0,0,0,0,0,0,0,91,0,0,0,129,0,46,0,250,0,232,0,22,0,150,0,150,0,7,0,208,0,139,0,175,0,192,0,0,0,63,0,204,0,65,0,0,0,72,0,67,0,0,0,78,0,228,0,81,0,212,0,162,0,0,0,61,0,0,0,242,0,154,0,43,0,78,0,151,0,0,0,31,0,23,0,225,0,94,0,0,0,122,0,55,0,208,0,0,0,0,0,219,0,83,0,72,0,142,0,110,0,89,0,0,0,0,0,118,0,0,0,0,0,0,0,38,0,98,0,55,0,225,0,95,0,202,0,16,0,0,0,136,0,216,0,0,0,49,0,0,0,60,0,115,0,108,0,115,0,0,0,0,0,12,0,0,0,135,0,115,0,248,0,236,0,207,0,0,0,118,0,187,0,127,0,134,0,160,0,101,0,217,0,80,0,212,0,232,0,0,0,47,0,39,0,89,0,235,0,223,0,0,0,0,0,179,0,129,0,254,0,207,0,0,0,125,0,0,0,109,0,138,0,236,0,164,0,160,0,0,0,36,0,145,0,197,0,36,0,212,0,197,0,94,0,91,0,237,0,56,0,106,0,91,0,141,0,231,0,206,0,0,0,150,0,187,0,179,0,160,0,0,0,222,0,175,0,0,0,101,0,84,0,40,0,0,0,72,0,0,0,245,0,118,0,0,0,149,0,0,0,149,0,193,0,0,0,163,0,25,0,223,0,64,0,40,0,227,0,0,0,144,0,8,0,171,0,124,0,0,0,196,0,117,0,0,0,0,0,115,0,37,0,183,0,63,0,161,0,175,0,77,0,138,0,18,0,0,0,90,0,9,0,11,0,232,0,0,0,241,0,158,0,144,0,45,0,38,0,151,0,0,0,77,0,163,0,85,0,0,0,0,0,0,0,132,0,91,0,0,0,220,0,148,0,115,0,105,0,69,0,2,0,129,0,138,0,249,0,0,0,141,0,148,0,128,0,35,0,218,0,183,0,23,0,115,0,136,0,0,0,129,0,58,0,0,0,120,0,141,0,90,0,136,0,85,0,29,0,100,0,111,0,95,0,72,0,154,0,102,0,0,0,0,0,126,0,0,0,207,0,39,0,95,0,0,0,52,0,0,0,215,0,160,0,251,0,244,0,202,0,242,0,32,0,194,0,233,0,203,0,220,0,230,0,164,0,84,0,13,0,142,0,177,0,0,0,63,0,199,0,0,0,157,0,74,0,0,0,0,0,204,0,79,0,59,0,0,0,199,0,14,0,0,0,216,0,222,0,41,0,69,0,89,0,0,0,0,0,25,0,15,0,238,0,108,0,52,0,0,0,54,0,0,0,241,0,18,0,35,0,236,0,12,0,23,0,0,0,254,0,64,0,133,0,0,0,0,0,131,0,91,0,243,0,245,0,136,0,0,0,213,0,225,0,0,0,164,0,224,0,226,0,64,0,132,0,100,0,105,0,208,0,86,0,0,0,95,0,50,0,0,0,62,0,0,0,99,0,150,0,186,0,146,0,69,0,184,0,25,0,0,0,34,0,91,0,255,0,54,0,236,0,222,0,90,0,0,0,0,0,177,0,9,0,247,0,110,0,0,0,246,0,0,0,136,0,119,0,211,0,95,0,164,0,0,0,0,0,57,0,29,0,84,0,185,0,115,0,44,0,0,0,0,0,92,0,153,0,149,0,125,0,29,0,0,0,37,0,79,0,160,0,0,0,0,0,23,0,217,0,0,0,52,0,52,0,255,0,48,0,75,0,253,0,173,0,0,0,97,0,240,0,87,0,160,0,0,0,182,0,45,0,237,0,241,0,0,0,11,0,221,0,150,0,104,0,6,0,0,0,168,0,124,0,121,0,172,0,135,0,56,0,231,0,248,0,183,0,47,0,93,0,197,0,242,0,0,0,0,0,0,0,85,0,0,0,79,0,0,0,121,0,242,0,218,0,184,0,90,0,85,0,113,0,0,0,190,0,3,0,226,0,121,0,249,0,37,0,204,0,55,0,147,0,166,0,211,0,0,0,162,0,94,0,30,0,0,0,28,0,43,0,140,0,166,0,0,0,235,0,64,0,115,0,229,0,214,0,151,0,39,0,0,0,119,0,89,0,70,0,220,0,0,0,0,0,0,0,179,0,136,0,41,0,205,0,168,0,223,0,218,0,80,0,233,0,147,0,182,0,166,0,174,0,36,0,180,0,9,0,0,0,216,0,179,0,0,0,0,0,171,0,76,0,13,0,87,0,0,0,0,0,153,0,164,0,0,0,0,0,221,0,92,0,136,0,39,0,68,0,0,0,14,0,209,0,75,0,135,0,181,0,66,0,0,0,0,0,164,0,49,0,144,0,0,0,33,0,57,0);
signal scenario_full  : scenario_type := (99,31,245,31,154,31,154,30,154,29,154,28,127,31,231,31,32,31,190,31,215,31,215,30,85,31,192,31,140,31,192,31,148,31,15,31,15,30,15,29,208,31,151,31,161,31,161,30,181,31,64,31,29,31,31,31,73,31,73,30,62,31,226,31,22,31,228,31,101,31,145,31,120,31,98,31,221,31,15,31,15,30,47,31,10,31,163,31,14,31,54,31,247,31,247,30,247,29,81,31,137,31,62,31,55,31,192,31,223,31,223,30,92,31,92,30,201,31,201,30,121,31,250,31,233,31,193,31,68,31,73,31,90,31,66,31,12,31,125,31,125,30,82,31,55,31,250,31,250,30,113,31,231,31,119,31,155,31,49,31,119,31,91,31,73,31,54,31,54,30,54,29,148,31,210,31,34,31,148,31,57,31,57,30,57,29,144,31,143,31,148,31,148,30,148,29,199,31,207,31,214,31,103,31,46,31,7,31,7,30,15,31,15,30,15,29,182,31,58,31,206,31,131,31,104,31,103,31,103,30,28,31,160,31,86,31,17,31,190,31,147,31,181,31,113,31,235,31,235,30,141,31,141,30,94,31,88,31,164,31,121,31,121,30,8,31,235,31,235,30,235,29,235,28,91,31,91,30,129,31,46,31,250,31,232,31,22,31,150,31,150,31,7,31,208,31,139,31,175,31,192,31,192,30,63,31,204,31,65,31,65,30,72,31,67,31,67,30,78,31,228,31,81,31,212,31,162,31,162,30,61,31,61,30,242,31,154,31,43,31,78,31,151,31,151,30,31,31,23,31,225,31,94,31,94,30,122,31,55,31,208,31,208,30,208,29,219,31,83,31,72,31,142,31,110,31,89,31,89,30,89,29,118,31,118,30,118,29,118,28,38,31,98,31,55,31,225,31,95,31,202,31,16,31,16,30,136,31,216,31,216,30,49,31,49,30,60,31,115,31,108,31,115,31,115,30,115,29,12,31,12,30,135,31,115,31,248,31,236,31,207,31,207,30,118,31,187,31,127,31,134,31,160,31,101,31,217,31,80,31,212,31,232,31,232,30,47,31,39,31,89,31,235,31,223,31,223,30,223,29,179,31,129,31,254,31,207,31,207,30,125,31,125,30,109,31,138,31,236,31,164,31,160,31,160,30,36,31,145,31,197,31,36,31,212,31,197,31,94,31,91,31,237,31,56,31,106,31,91,31,141,31,231,31,206,31,206,30,150,31,187,31,179,31,160,31,160,30,222,31,175,31,175,30,101,31,84,31,40,31,40,30,72,31,72,30,245,31,118,31,118,30,149,31,149,30,149,31,193,31,193,30,163,31,25,31,223,31,64,31,40,31,227,31,227,30,144,31,8,31,171,31,124,31,124,30,196,31,117,31,117,30,117,29,115,31,37,31,183,31,63,31,161,31,175,31,77,31,138,31,18,31,18,30,90,31,9,31,11,31,232,31,232,30,241,31,158,31,144,31,45,31,38,31,151,31,151,30,77,31,163,31,85,31,85,30,85,29,85,28,132,31,91,31,91,30,220,31,148,31,115,31,105,31,69,31,2,31,129,31,138,31,249,31,249,30,141,31,148,31,128,31,35,31,218,31,183,31,23,31,115,31,136,31,136,30,129,31,58,31,58,30,120,31,141,31,90,31,136,31,85,31,29,31,100,31,111,31,95,31,72,31,154,31,102,31,102,30,102,29,126,31,126,30,207,31,39,31,95,31,95,30,52,31,52,30,215,31,160,31,251,31,244,31,202,31,242,31,32,31,194,31,233,31,203,31,220,31,230,31,164,31,84,31,13,31,142,31,177,31,177,30,63,31,199,31,199,30,157,31,74,31,74,30,74,29,204,31,79,31,59,31,59,30,199,31,14,31,14,30,216,31,222,31,41,31,69,31,89,31,89,30,89,29,25,31,15,31,238,31,108,31,52,31,52,30,54,31,54,30,241,31,18,31,35,31,236,31,12,31,23,31,23,30,254,31,64,31,133,31,133,30,133,29,131,31,91,31,243,31,245,31,136,31,136,30,213,31,225,31,225,30,164,31,224,31,226,31,64,31,132,31,100,31,105,31,208,31,86,31,86,30,95,31,50,31,50,30,62,31,62,30,99,31,150,31,186,31,146,31,69,31,184,31,25,31,25,30,34,31,91,31,255,31,54,31,236,31,222,31,90,31,90,30,90,29,177,31,9,31,247,31,110,31,110,30,246,31,246,30,136,31,119,31,211,31,95,31,164,31,164,30,164,29,57,31,29,31,84,31,185,31,115,31,44,31,44,30,44,29,92,31,153,31,149,31,125,31,29,31,29,30,37,31,79,31,160,31,160,30,160,29,23,31,217,31,217,30,52,31,52,31,255,31,48,31,75,31,253,31,173,31,173,30,97,31,240,31,87,31,160,31,160,30,182,31,45,31,237,31,241,31,241,30,11,31,221,31,150,31,104,31,6,31,6,30,168,31,124,31,121,31,172,31,135,31,56,31,231,31,248,31,183,31,47,31,93,31,197,31,242,31,242,30,242,29,242,28,85,31,85,30,79,31,79,30,121,31,242,31,218,31,184,31,90,31,85,31,113,31,113,30,190,31,3,31,226,31,121,31,249,31,37,31,204,31,55,31,147,31,166,31,211,31,211,30,162,31,94,31,30,31,30,30,28,31,43,31,140,31,166,31,166,30,235,31,64,31,115,31,229,31,214,31,151,31,39,31,39,30,119,31,89,31,70,31,220,31,220,30,220,29,220,28,179,31,136,31,41,31,205,31,168,31,223,31,218,31,80,31,233,31,147,31,182,31,166,31,174,31,36,31,180,31,9,31,9,30,216,31,179,31,179,30,179,29,171,31,76,31,13,31,87,31,87,30,87,29,153,31,164,31,164,30,164,29,221,31,92,31,136,31,39,31,68,31,68,30,14,31,209,31,75,31,135,31,181,31,66,31,66,30,66,29,164,31,49,31,144,31,144,30,33,31,57,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
