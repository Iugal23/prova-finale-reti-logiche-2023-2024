-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_2 is
end project_tb_2;

architecture project_tb_arch_2 of project_tb_2 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 792;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (220,0,214,0,51,0,200,0,46,0,210,0,201,0,236,0,9,0,47,0,124,0,0,0,41,0,21,0,206,0,52,0,0,0,73,0,0,0,0,0,213,0,8,0,124,0,0,0,0,0,0,0,12,0,0,0,108,0,0,0,132,0,82,0,87,0,0,0,57,0,187,0,154,0,56,0,80,0,111,0,180,0,0,0,168,0,147,0,112,0,249,0,116,0,0,0,255,0,248,0,0,0,187,0,132,0,138,0,93,0,24,0,96,0,0,0,93,0,82,0,6,0,195,0,230,0,0,0,41,0,0,0,0,0,166,0,153,0,153,0,0,0,253,0,0,0,227,0,198,0,0,0,0,0,6,0,221,0,155,0,206,0,216,0,163,0,122,0,124,0,79,0,19,0,206,0,0,0,167,0,175,0,234,0,239,0,0,0,194,0,0,0,221,0,0,0,0,0,128,0,23,0,141,0,0,0,254,0,215,0,135,0,93,0,215,0,0,0,21,0,166,0,0,0,134,0,9,0,174,0,204,0,73,0,94,0,245,0,150,0,0,0,119,0,207,0,30,0,204,0,50,0,206,0,0,0,0,0,84,0,197,0,189,0,167,0,51,0,226,0,170,0,187,0,222,0,0,0,0,0,198,0,28,0,85,0,246,0,89,0,90,0,212,0,45,0,11,0,239,0,86,0,61,0,0,0,197,0,115,0,0,0,94,0,179,0,169,0,244,0,57,0,0,0,28,0,49,0,0,0,93,0,145,0,10,0,120,0,214,0,9,0,217,0,134,0,97,0,61,0,20,0,100,0,118,0,213,0,218,0,117,0,58,0,2,0,191,0,247,0,34,0,81,0,86,0,96,0,234,0,42,0,174,0,23,0,140,0,213,0,176,0,204,0,6,0,97,0,16,0,9,0,163,0,83,0,199,0,61,0,39,0,0,0,145,0,161,0,14,0,1,0,95,0,0,0,214,0,229,0,164,0,234,0,16,0,164,0,48,0,80,0,0,0,98,0,123,0,75,0,0,0,32,0,79,0,101,0,4,0,7,0,189,0,1,0,33,0,135,0,219,0,178,0,226,0,172,0,0,0,67,0,244,0,247,0,190,0,9,0,0,0,110,0,48,0,0,0,160,0,95,0,0,0,0,0,59,0,69,0,240,0,155,0,81,0,151,0,0,0,0,0,232,0,154,0,139,0,0,0,0,0,103,0,0,0,78,0,128,0,78,0,66,0,130,0,55,0,37,0,70,0,219,0,17,0,238,0,216,0,124,0,133,0,214,0,167,0,0,0,210,0,16,0,63,0,248,0,220,0,0,0,82,0,0,0,0,0,40,0,81,0,197,0,0,0,144,0,36,0,69,0,232,0,102,0,229,0,0,0,0,0,32,0,251,0,234,0,94,0,96,0,204,0,205,0,154,0,218,0,250,0,32,0,230,0,0,0,250,0,43,0,0,0,187,0,0,0,243,0,211,0,169,0,22,0,177,0,186,0,0,0,52,0,29,0,0,0,142,0,1,0,0,0,48,0,49,0,118,0,248,0,0,0,118,0,0,0,203,0,149,0,86,0,252,0,97,0,218,0,177,0,149,0,69,0,0,0,98,0,115,0,201,0,18,0,156,0,28,0,179,0,130,0,201,0,73,0,130,0,206,0,21,0,142,0,174,0,50,0,148,0,89,0,214,0,76,0,0,0,0,0,147,0,181,0,0,0,151,0,104,0,150,0,138,0,59,0,103,0,134,0,0,0,212,0,5,0,61,0,21,0,162,0,130,0,237,0,0,0,222,0,24,0,56,0,231,0,115,0,115,0,0,0,250,0,0,0,9,0,247,0,75,0,43,0,0,0,23,0,66,0,247,0,145,0,196,0,203,0,14,0,210,0,90,0,64,0,149,0,69,0,230,0,0,0,0,0,236,0,112,0,112,0,122,0,196,0,204,0,58,0,0,0,102,0,40,0,75,0,168,0,35,0,52,0,43,0,0,0,251,0,0,0,153,0,0,0,0,0,49,0,19,0,158,0,100,0,0,0,26,0,116,0,0,0,74,0,222,0,207,0,14,0,175,0,93,0,131,0,164,0,93,0,0,0,0,0,198,0,166,0,83,0,89,0,76,0,0,0,0,0,9,0,0,0,62,0,0,0,213,0,234,0,37,0,155,0,128,0,249,0,0,0,178,0,0,0,7,0,0,0,176,0,0,0,0,0,176,0,93,0,115,0,126,0,197,0,50,0,0,0,193,0,114,0,146,0,19,0,119,0,245,0,24,0,117,0,93,0,0,0,92,0,157,0,0,0,0,0,185,0,121,0,96,0,202,0,34,0,204,0,0,0,95,0,0,0,133,0,207,0,56,0,122,0,154,0,223,0,117,0,171,0,0,0,0,0,0,0,0,0,39,0,205,0,206,0,78,0,172,0,28,0,213,0,144,0,0,0,16,0,130,0,12,0,0,0,87,0,26,0,168,0,223,0,212,0,24,0,218,0,0,0,0,0,0,0,229,0,215,0,244,0,44,0,56,0,82,0,195,0,0,0,212,0,222,0,0,0,134,0,113,0,17,0,121,0,12,0,0,0,50,0,0,0,142,0,169,0,240,0,131,0,217,0,41,0,163,0,60,0,155,0,202,0,33,0,0,0,0,0,138,0,88,0,0,0,74,0,0,0,138,0,173,0,72,0,239,0,33,0,213,0,97,0,79,0,63,0,41,0,0,0,204,0,196,0,190,0,0,0,115,0,191,0,31,0,0,0,213,0,178,0,80,0,163,0,171,0,213,0,122,0,197,0,139,0,178,0,42,0,112,0,0,0,26,0,190,0,0,0,0,0,216,0,156,0,0,0,106,0,159,0,99,0,151,0,84,0,0,0,53,0,88,0,126,0,77,0,59,0,110,0,0,0,82,0,0,0,0,0,80,0,115,0,228,0,209,0,0,0,118,0,0,0,15,0,127,0,111,0,206,0,118,0,254,0,116,0,61,0,0,0,162,0,112,0,95,0,94,0,0,0,20,0,0,0,98,0,0,0,42,0,215,0,101,0,159,0,74,0,0,0,89,0,143,0,174,0,131,0,240,0,0,0,14,0,0,0,176,0,191,0,211,0,147,0,201,0,145,0,63,0,235,0,121,0,92,0,197,0,191,0,176,0,63,0,0,0,16,0,139,0,145,0,101,0,0,0,247,0,184,0,8,0,54,0,128,0,0,0,0,0,210,0,196,0,149,0,241,0,54,0,227,0,0,0,195,0,7,0,161,0,19,0,48,0,184,0,0,0,0,0,253,0,168,0,14,0,89,0,27,0,160,0,159,0,34,0,209,0,102,0,155,0,190,0,168,0,108,0,0,0,37,0,180,0,0,0,83,0,80,0,227,0,224,0,36,0,164,0,146,0,106,0,136,0,100,0,120,0,91,0,253,0,0,0,247,0,46,0,60,0,0,0,0,0,153,0,78,0,0,0,82,0,193,0,174,0,0,0,244,0,154,0,85,0,157,0,137,0,181,0,75,0,203,0,184,0,199,0,25,0,195,0,75,0,163,0,243,0,144,0,0,0,203,0,153,0,237,0,129,0);
signal scenario_full  : scenario_type := (220,31,214,31,51,31,200,31,46,31,210,31,201,31,236,31,9,31,47,31,124,31,124,30,41,31,21,31,206,31,52,31,52,30,73,31,73,30,73,29,213,31,8,31,124,31,124,30,124,29,124,28,12,31,12,30,108,31,108,30,132,31,82,31,87,31,87,30,57,31,187,31,154,31,56,31,80,31,111,31,180,31,180,30,168,31,147,31,112,31,249,31,116,31,116,30,255,31,248,31,248,30,187,31,132,31,138,31,93,31,24,31,96,31,96,30,93,31,82,31,6,31,195,31,230,31,230,30,41,31,41,30,41,29,166,31,153,31,153,31,153,30,253,31,253,30,227,31,198,31,198,30,198,29,6,31,221,31,155,31,206,31,216,31,163,31,122,31,124,31,79,31,19,31,206,31,206,30,167,31,175,31,234,31,239,31,239,30,194,31,194,30,221,31,221,30,221,29,128,31,23,31,141,31,141,30,254,31,215,31,135,31,93,31,215,31,215,30,21,31,166,31,166,30,134,31,9,31,174,31,204,31,73,31,94,31,245,31,150,31,150,30,119,31,207,31,30,31,204,31,50,31,206,31,206,30,206,29,84,31,197,31,189,31,167,31,51,31,226,31,170,31,187,31,222,31,222,30,222,29,198,31,28,31,85,31,246,31,89,31,90,31,212,31,45,31,11,31,239,31,86,31,61,31,61,30,197,31,115,31,115,30,94,31,179,31,169,31,244,31,57,31,57,30,28,31,49,31,49,30,93,31,145,31,10,31,120,31,214,31,9,31,217,31,134,31,97,31,61,31,20,31,100,31,118,31,213,31,218,31,117,31,58,31,2,31,191,31,247,31,34,31,81,31,86,31,96,31,234,31,42,31,174,31,23,31,140,31,213,31,176,31,204,31,6,31,97,31,16,31,9,31,163,31,83,31,199,31,61,31,39,31,39,30,145,31,161,31,14,31,1,31,95,31,95,30,214,31,229,31,164,31,234,31,16,31,164,31,48,31,80,31,80,30,98,31,123,31,75,31,75,30,32,31,79,31,101,31,4,31,7,31,189,31,1,31,33,31,135,31,219,31,178,31,226,31,172,31,172,30,67,31,244,31,247,31,190,31,9,31,9,30,110,31,48,31,48,30,160,31,95,31,95,30,95,29,59,31,69,31,240,31,155,31,81,31,151,31,151,30,151,29,232,31,154,31,139,31,139,30,139,29,103,31,103,30,78,31,128,31,78,31,66,31,130,31,55,31,37,31,70,31,219,31,17,31,238,31,216,31,124,31,133,31,214,31,167,31,167,30,210,31,16,31,63,31,248,31,220,31,220,30,82,31,82,30,82,29,40,31,81,31,197,31,197,30,144,31,36,31,69,31,232,31,102,31,229,31,229,30,229,29,32,31,251,31,234,31,94,31,96,31,204,31,205,31,154,31,218,31,250,31,32,31,230,31,230,30,250,31,43,31,43,30,187,31,187,30,243,31,211,31,169,31,22,31,177,31,186,31,186,30,52,31,29,31,29,30,142,31,1,31,1,30,48,31,49,31,118,31,248,31,248,30,118,31,118,30,203,31,149,31,86,31,252,31,97,31,218,31,177,31,149,31,69,31,69,30,98,31,115,31,201,31,18,31,156,31,28,31,179,31,130,31,201,31,73,31,130,31,206,31,21,31,142,31,174,31,50,31,148,31,89,31,214,31,76,31,76,30,76,29,147,31,181,31,181,30,151,31,104,31,150,31,138,31,59,31,103,31,134,31,134,30,212,31,5,31,61,31,21,31,162,31,130,31,237,31,237,30,222,31,24,31,56,31,231,31,115,31,115,31,115,30,250,31,250,30,9,31,247,31,75,31,43,31,43,30,23,31,66,31,247,31,145,31,196,31,203,31,14,31,210,31,90,31,64,31,149,31,69,31,230,31,230,30,230,29,236,31,112,31,112,31,122,31,196,31,204,31,58,31,58,30,102,31,40,31,75,31,168,31,35,31,52,31,43,31,43,30,251,31,251,30,153,31,153,30,153,29,49,31,19,31,158,31,100,31,100,30,26,31,116,31,116,30,74,31,222,31,207,31,14,31,175,31,93,31,131,31,164,31,93,31,93,30,93,29,198,31,166,31,83,31,89,31,76,31,76,30,76,29,9,31,9,30,62,31,62,30,213,31,234,31,37,31,155,31,128,31,249,31,249,30,178,31,178,30,7,31,7,30,176,31,176,30,176,29,176,31,93,31,115,31,126,31,197,31,50,31,50,30,193,31,114,31,146,31,19,31,119,31,245,31,24,31,117,31,93,31,93,30,92,31,157,31,157,30,157,29,185,31,121,31,96,31,202,31,34,31,204,31,204,30,95,31,95,30,133,31,207,31,56,31,122,31,154,31,223,31,117,31,171,31,171,30,171,29,171,28,171,27,39,31,205,31,206,31,78,31,172,31,28,31,213,31,144,31,144,30,16,31,130,31,12,31,12,30,87,31,26,31,168,31,223,31,212,31,24,31,218,31,218,30,218,29,218,28,229,31,215,31,244,31,44,31,56,31,82,31,195,31,195,30,212,31,222,31,222,30,134,31,113,31,17,31,121,31,12,31,12,30,50,31,50,30,142,31,169,31,240,31,131,31,217,31,41,31,163,31,60,31,155,31,202,31,33,31,33,30,33,29,138,31,88,31,88,30,74,31,74,30,138,31,173,31,72,31,239,31,33,31,213,31,97,31,79,31,63,31,41,31,41,30,204,31,196,31,190,31,190,30,115,31,191,31,31,31,31,30,213,31,178,31,80,31,163,31,171,31,213,31,122,31,197,31,139,31,178,31,42,31,112,31,112,30,26,31,190,31,190,30,190,29,216,31,156,31,156,30,106,31,159,31,99,31,151,31,84,31,84,30,53,31,88,31,126,31,77,31,59,31,110,31,110,30,82,31,82,30,82,29,80,31,115,31,228,31,209,31,209,30,118,31,118,30,15,31,127,31,111,31,206,31,118,31,254,31,116,31,61,31,61,30,162,31,112,31,95,31,94,31,94,30,20,31,20,30,98,31,98,30,42,31,215,31,101,31,159,31,74,31,74,30,89,31,143,31,174,31,131,31,240,31,240,30,14,31,14,30,176,31,191,31,211,31,147,31,201,31,145,31,63,31,235,31,121,31,92,31,197,31,191,31,176,31,63,31,63,30,16,31,139,31,145,31,101,31,101,30,247,31,184,31,8,31,54,31,128,31,128,30,128,29,210,31,196,31,149,31,241,31,54,31,227,31,227,30,195,31,7,31,161,31,19,31,48,31,184,31,184,30,184,29,253,31,168,31,14,31,89,31,27,31,160,31,159,31,34,31,209,31,102,31,155,31,190,31,168,31,108,31,108,30,37,31,180,31,180,30,83,31,80,31,227,31,224,31,36,31,164,31,146,31,106,31,136,31,100,31,120,31,91,31,253,31,253,30,247,31,46,31,60,31,60,30,60,29,153,31,78,31,78,30,82,31,193,31,174,31,174,30,244,31,154,31,85,31,157,31,137,31,181,31,75,31,203,31,184,31,199,31,25,31,195,31,75,31,163,31,243,31,144,31,144,30,203,31,153,31,237,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
