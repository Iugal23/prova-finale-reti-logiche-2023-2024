-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_617 is
end project_tb_617;

architecture project_tb_arch_617 of project_tb_617 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 571;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (82,0,78,0,17,0,48,0,74,0,209,0,44,0,220,0,0,0,9,0,10,0,0,0,148,0,157,0,142,0,119,0,109,0,0,0,193,0,22,0,104,0,99,0,164,0,217,0,114,0,106,0,156,0,130,0,197,0,0,0,165,0,125,0,32,0,140,0,133,0,52,0,211,0,182,0,198,0,0,0,0,0,0,0,0,0,180,0,0,0,90,0,179,0,0,0,51,0,222,0,57,0,252,0,0,0,129,0,48,0,162,0,98,0,195,0,187,0,0,0,56,0,5,0,188,0,156,0,251,0,145,0,3,0,139,0,0,0,23,0,99,0,0,0,25,0,203,0,146,0,200,0,2,0,0,0,11,0,65,0,140,0,35,0,210,0,54,0,128,0,89,0,226,0,0,0,28,0,114,0,83,0,120,0,156,0,24,0,0,0,34,0,187,0,69,0,29,0,112,0,99,0,142,0,22,0,187,0,234,0,147,0,64,0,0,0,229,0,69,0,211,0,246,0,0,0,222,0,39,0,251,0,230,0,177,0,44,0,95,0,44,0,48,0,251,0,138,0,0,0,90,0,89,0,162,0,0,0,0,0,87,0,33,0,0,0,242,0,39,0,58,0,39,0,102,0,0,0,65,0,0,0,135,0,0,0,21,0,239,0,110,0,244,0,96,0,183,0,77,0,112,0,87,0,97,0,194,0,252,0,187,0,221,0,0,0,173,0,128,0,0,0,91,0,244,0,0,0,248,0,0,0,208,0,85,0,80,0,190,0,214,0,0,0,243,0,90,0,0,0,0,0,0,0,121,0,156,0,30,0,0,0,201,0,246,0,150,0,0,0,59,0,253,0,0,0,97,0,236,0,0,0,0,0,0,0,0,0,118,0,74,0,208,0,150,0,78,0,219,0,116,0,0,0,57,0,139,0,134,0,0,0,174,0,47,0,210,0,0,0,182,0,0,0,211,0,0,0,0,0,133,0,0,0,0,0,88,0,114,0,59,0,115,0,204,0,25,0,182,0,0,0,125,0,162,0,108,0,246,0,16,0,224,0,106,0,224,0,143,0,78,0,85,0,31,0,105,0,1,0,0,0,156,0,160,0,56,0,0,0,252,0,113,0,87,0,160,0,5,0,0,0,0,0,139,0,160,0,13,0,166,0,23,0,240,0,237,0,0,0,41,0,31,0,161,0,0,0,235,0,234,0,199,0,73,0,140,0,2,0,60,0,0,0,157,0,0,0,83,0,62,0,151,0,83,0,114,0,68,0,0,0,172,0,202,0,0,0,158,0,60,0,106,0,102,0,188,0,59,0,221,0,0,0,50,0,0,0,169,0,60,0,118,0,82,0,42,0,0,0,166,0,47,0,245,0,136,0,155,0,168,0,102,0,131,0,158,0,79,0,207,0,180,0,50,0,0,0,251,0,156,0,215,0,138,0,97,0,0,0,168,0,234,0,40,0,199,0,71,0,72,0,0,0,0,0,0,0,0,0,0,0,118,0,237,0,155,0,31,0,0,0,51,0,119,0,100,0,232,0,35,0,0,0,211,0,0,0,0,0,21,0,154,0,0,0,204,0,158,0,0,0,10,0,0,0,111,0,229,0,87,0,0,0,41,0,87,0,0,0,228,0,113,0,143,0,103,0,197,0,102,0,219,0,169,0,0,0,251,0,142,0,163,0,213,0,136,0,20,0,123,0,156,0,54,0,149,0,0,0,0,0,205,0,116,0,216,0,36,0,184,0,65,0,224,0,194,0,23,0,109,0,96,0,255,0,232,0,209,0,230,0,80,0,107,0,0,0,190,0,216,0,44,0,167,0,72,0,149,0,9,0,215,0,0,0,240,0,136,0,95,0,43,0,128,0,0,0,232,0,0,0,120,0,90,0,58,0,172,0,9,0,114,0,89,0,131,0,0,0,88,0,0,0,0,0,232,0,0,0,220,0,63,0,0,0,42,0,113,0,126,0,204,0,192,0,194,0,247,0,79,0,226,0,181,0,168,0,0,0,146,0,0,0,0,0,244,0,238,0,168,0,160,0,0,0,91,0,44,0,0,0,240,0,89,0,0,0,17,0,33,0,0,0,0,0,143,0,224,0,210,0,95,0,47,0,112,0,187,0,0,0,229,0,53,0,27,0,0,0,4,0,3,0,177,0,106,0,135,0,241,0,58,0,40,0,211,0,25,0,120,0,54,0,142,0,66,0,229,0,16,0,0,0,46,0,0,0,0,0,213,0,169,0,59,0,113,0,218,0,0,0,44,0,169,0,147,0,132,0,83,0,0,0,126,0,0,0,250,0,160,0,147,0,0,0,176,0,215,0,142,0,216,0,92,0,209,0,110,0,53,0,102,0,166,0,158,0,16,0,56,0,62,0,215,0,11,0,0,0,240,0,130,0,138,0,64,0,73,0,196,0,0,0,0,0,150,0,113,0,85,0,248,0,158,0,0,0,72,0,126,0,113,0,125,0,0,0,188,0,203,0,250,0,0,0,0,0,162,0,0,0,142,0,160,0,221,0,63,0,88,0,7,0,4,0,0,0,115,0,0,0,210,0,20,0,68,0,182,0,48,0);
signal scenario_full  : scenario_type := (82,31,78,31,17,31,48,31,74,31,209,31,44,31,220,31,220,30,9,31,10,31,10,30,148,31,157,31,142,31,119,31,109,31,109,30,193,31,22,31,104,31,99,31,164,31,217,31,114,31,106,31,156,31,130,31,197,31,197,30,165,31,125,31,32,31,140,31,133,31,52,31,211,31,182,31,198,31,198,30,198,29,198,28,198,27,180,31,180,30,90,31,179,31,179,30,51,31,222,31,57,31,252,31,252,30,129,31,48,31,162,31,98,31,195,31,187,31,187,30,56,31,5,31,188,31,156,31,251,31,145,31,3,31,139,31,139,30,23,31,99,31,99,30,25,31,203,31,146,31,200,31,2,31,2,30,11,31,65,31,140,31,35,31,210,31,54,31,128,31,89,31,226,31,226,30,28,31,114,31,83,31,120,31,156,31,24,31,24,30,34,31,187,31,69,31,29,31,112,31,99,31,142,31,22,31,187,31,234,31,147,31,64,31,64,30,229,31,69,31,211,31,246,31,246,30,222,31,39,31,251,31,230,31,177,31,44,31,95,31,44,31,48,31,251,31,138,31,138,30,90,31,89,31,162,31,162,30,162,29,87,31,33,31,33,30,242,31,39,31,58,31,39,31,102,31,102,30,65,31,65,30,135,31,135,30,21,31,239,31,110,31,244,31,96,31,183,31,77,31,112,31,87,31,97,31,194,31,252,31,187,31,221,31,221,30,173,31,128,31,128,30,91,31,244,31,244,30,248,31,248,30,208,31,85,31,80,31,190,31,214,31,214,30,243,31,90,31,90,30,90,29,90,28,121,31,156,31,30,31,30,30,201,31,246,31,150,31,150,30,59,31,253,31,253,30,97,31,236,31,236,30,236,29,236,28,236,27,118,31,74,31,208,31,150,31,78,31,219,31,116,31,116,30,57,31,139,31,134,31,134,30,174,31,47,31,210,31,210,30,182,31,182,30,211,31,211,30,211,29,133,31,133,30,133,29,88,31,114,31,59,31,115,31,204,31,25,31,182,31,182,30,125,31,162,31,108,31,246,31,16,31,224,31,106,31,224,31,143,31,78,31,85,31,31,31,105,31,1,31,1,30,156,31,160,31,56,31,56,30,252,31,113,31,87,31,160,31,5,31,5,30,5,29,139,31,160,31,13,31,166,31,23,31,240,31,237,31,237,30,41,31,31,31,161,31,161,30,235,31,234,31,199,31,73,31,140,31,2,31,60,31,60,30,157,31,157,30,83,31,62,31,151,31,83,31,114,31,68,31,68,30,172,31,202,31,202,30,158,31,60,31,106,31,102,31,188,31,59,31,221,31,221,30,50,31,50,30,169,31,60,31,118,31,82,31,42,31,42,30,166,31,47,31,245,31,136,31,155,31,168,31,102,31,131,31,158,31,79,31,207,31,180,31,50,31,50,30,251,31,156,31,215,31,138,31,97,31,97,30,168,31,234,31,40,31,199,31,71,31,72,31,72,30,72,29,72,28,72,27,72,26,118,31,237,31,155,31,31,31,31,30,51,31,119,31,100,31,232,31,35,31,35,30,211,31,211,30,211,29,21,31,154,31,154,30,204,31,158,31,158,30,10,31,10,30,111,31,229,31,87,31,87,30,41,31,87,31,87,30,228,31,113,31,143,31,103,31,197,31,102,31,219,31,169,31,169,30,251,31,142,31,163,31,213,31,136,31,20,31,123,31,156,31,54,31,149,31,149,30,149,29,205,31,116,31,216,31,36,31,184,31,65,31,224,31,194,31,23,31,109,31,96,31,255,31,232,31,209,31,230,31,80,31,107,31,107,30,190,31,216,31,44,31,167,31,72,31,149,31,9,31,215,31,215,30,240,31,136,31,95,31,43,31,128,31,128,30,232,31,232,30,120,31,90,31,58,31,172,31,9,31,114,31,89,31,131,31,131,30,88,31,88,30,88,29,232,31,232,30,220,31,63,31,63,30,42,31,113,31,126,31,204,31,192,31,194,31,247,31,79,31,226,31,181,31,168,31,168,30,146,31,146,30,146,29,244,31,238,31,168,31,160,31,160,30,91,31,44,31,44,30,240,31,89,31,89,30,17,31,33,31,33,30,33,29,143,31,224,31,210,31,95,31,47,31,112,31,187,31,187,30,229,31,53,31,27,31,27,30,4,31,3,31,177,31,106,31,135,31,241,31,58,31,40,31,211,31,25,31,120,31,54,31,142,31,66,31,229,31,16,31,16,30,46,31,46,30,46,29,213,31,169,31,59,31,113,31,218,31,218,30,44,31,169,31,147,31,132,31,83,31,83,30,126,31,126,30,250,31,160,31,147,31,147,30,176,31,215,31,142,31,216,31,92,31,209,31,110,31,53,31,102,31,166,31,158,31,16,31,56,31,62,31,215,31,11,31,11,30,240,31,130,31,138,31,64,31,73,31,196,31,196,30,196,29,150,31,113,31,85,31,248,31,158,31,158,30,72,31,126,31,113,31,125,31,125,30,188,31,203,31,250,31,250,30,250,29,162,31,162,30,142,31,160,31,221,31,63,31,88,31,7,31,4,31,4,30,115,31,115,30,210,31,20,31,68,31,182,31,48,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
