-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 795;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (216,0,0,0,105,0,89,0,135,0,43,0,0,0,127,0,171,0,67,0,28,0,198,0,252,0,0,0,131,0,67,0,0,0,0,0,243,0,227,0,103,0,217,0,11,0,204,0,0,0,240,0,190,0,0,0,6,0,43,0,188,0,250,0,33,0,0,0,31,0,44,0,156,0,217,0,2,0,251,0,169,0,98,0,0,0,41,0,132,0,173,0,24,0,101,0,156,0,18,0,236,0,37,0,225,0,128,0,218,0,238,0,29,0,112,0,152,0,123,0,71,0,217,0,56,0,78,0,174,0,0,0,167,0,153,0,234,0,0,0,195,0,241,0,89,0,0,0,0,0,112,0,35,0,133,0,172,0,85,0,252,0,213,0,91,0,96,0,14,0,0,0,175,0,20,0,190,0,60,0,205,0,129,0,0,0,223,0,38,0,234,0,0,0,0,0,150,0,53,0,151,0,104,0,242,0,175,0,26,0,0,0,0,0,0,0,58,0,32,0,63,0,91,0,0,0,219,0,48,0,71,0,166,0,0,0,130,0,75,0,0,0,86,0,22,0,0,0,0,0,47,0,134,0,0,0,237,0,205,0,69,0,96,0,63,0,35,0,11,0,83,0,205,0,0,0,0,0,172,0,0,0,161,0,29,0,115,0,55,0,0,0,102,0,31,0,116,0,0,0,0,0,218,0,47,0,11,0,111,0,164,0,0,0,198,0,108,0,164,0,43,0,179,0,66,0,215,0,0,0,181,0,255,0,60,0,165,0,79,0,65,0,202,0,0,0,35,0,0,0,0,0,109,0,7,0,115,0,70,0,123,0,98,0,86,0,96,0,239,0,233,0,229,0,0,0,129,0,144,0,244,0,0,0,166,0,7,0,29,0,66,0,135,0,128,0,6,0,0,0,62,0,241,0,0,0,0,0,120,0,95,0,156,0,240,0,169,0,14,0,48,0,58,0,27,0,61,0,29,0,242,0,151,0,85,0,163,0,0,0,0,0,55,0,46,0,168,0,0,0,75,0,86,0,230,0,185,0,36,0,57,0,233,0,51,0,130,0,111,0,230,0,43,0,100,0,0,0,10,0,137,0,17,0,0,0,140,0,145,0,51,0,127,0,241,0,89,0,36,0,0,0,36,0,197,0,110,0,0,0,99,0,21,0,252,0,130,0,130,0,202,0,49,0,0,0,31,0,19,0,187,0,141,0,242,0,123,0,0,0,182,0,0,0,0,0,147,0,210,0,210,0,229,0,4,0,114,0,121,0,0,0,207,0,67,0,219,0,0,0,0,0,0,0,23,0,0,0,178,0,33,0,87,0,131,0,245,0,85,0,154,0,49,0,219,0,245,0,0,0,0,0,140,0,167,0,209,0,160,0,91,0,98,0,220,0,148,0,0,0,95,0,14,0,34,0,0,0,28,0,0,0,98,0,0,0,244,0,125,0,0,0,91,0,228,0,162,0,0,0,78,0,136,0,229,0,57,0,175,0,48,0,179,0,0,0,22,0,0,0,65,0,173,0,136,0,225,0,98,0,137,0,144,0,83,0,134,0,222,0,133,0,19,0,245,0,93,0,43,0,72,0,5,0,0,0,194,0,102,0,77,0,239,0,84,0,16,0,166,0,69,0,43,0,172,0,5,0,90,0,138,0,0,0,0,0,0,0,51,0,58,0,19,0,172,0,132,0,77,0,211,0,140,0,202,0,208,0,191,0,192,0,210,0,56,0,22,0,154,0,254,0,14,0,240,0,0,0,240,0,71,0,198,0,205,0,0,0,0,0,69,0,199,0,23,0,0,0,237,0,0,0,231,0,79,0,31,0,245,0,39,0,83,0,72,0,250,0,0,0,0,0,243,0,225,0,69,0,91,0,29,0,0,0,200,0,168,0,67,0,221,0,202,0,0,0,136,0,0,0,0,0,240,0,42,0,106,0,118,0,21,0,148,0,4,0,234,0,233,0,240,0,222,0,0,0,168,0,139,0,168,0,27,0,42,0,178,0,0,0,242,0,105,0,130,0,60,0,92,0,186,0,173,0,206,0,204,0,95,0,19,0,134,0,0,0,194,0,173,0,194,0,100,0,212,0,239,0,195,0,106,0,83,0,125,0,133,0,0,0,0,0,25,0,0,0,225,0,0,0,42,0,0,0,0,0,29,0,8,0,201,0,36,0,250,0,205,0,34,0,198,0,67,0,248,0,93,0,187,0,166,0,255,0,230,0,78,0,5,0,0,0,186,0,80,0,0,0,0,0,0,0,180,0,138,0,62,0,123,0,49,0,163,0,192,0,0,0,206,0,18,0,0,0,247,0,183,0,76,0,0,0,254,0,37,0,119,0,111,0,19,0,231,0,73,0,0,0,252,0,162,0,198,0,0,0,78,0,224,0,37,0,114,0,18,0,137,0,211,0,171,0,116,0,0,0,0,0,77,0,249,0,0,0,223,0,221,0,109,0,23,0,0,0,183,0,246,0,146,0,208,0,144,0,1,0,0,0,192,0,175,0,12,0,0,0,193,0,0,0,179,0,36,0,0,0,0,0,221,0,243,0,47,0,207,0,0,0,152,0,184,0,0,0,207,0,108,0,121,0,6,0,125,0,27,0,41,0,1,0,109,0,78,0,0,0,61,0,227,0,194,0,242,0,170,0,1,0,50,0,0,0,0,0,33,0,109,0,7,0,231,0,106,0,20,0,45,0,92,0,39,0,81,0,89,0,0,0,0,0,224,0,205,0,92,0,30,0,80,0,155,0,85,0,249,0,154,0,68,0,0,0,96,0,201,0,143,0,0,0,177,0,151,0,0,0,100,0,148,0,199,0,147,0,11,0,119,0,33,0,54,0,180,0,245,0,120,0,39,0,0,0,129,0,16,0,33,0,117,0,218,0,215,0,0,0,0,0,242,0,163,0,241,0,56,0,192,0,170,0,75,0,105,0,71,0,78,0,180,0,232,0,238,0,83,0,44,0,239,0,169,0,103,0,0,0,32,0,220,0,192,0,242,0,0,0,0,0,199,0,93,0,77,0,61,0,139,0,0,0,0,0,0,0,127,0,56,0,0,0,168,0,248,0,0,0,173,0,179,0,223,0,0,0,249,0,28,0,0,0,0,0,103,0,225,0,231,0,0,0,150,0,162,0,171,0,39,0,19,0,23,0,7,0,144,0,0,0,184,0,196,0,189,0,68,0,166,0,0,0,173,0,211,0,164,0,77,0,245,0,230,0,134,0,6,0,223,0,0,0,50,0,78,0,12,0,242,0,211,0,231,0,91,0,181,0,206,0,11,0,15,0,24,0,0,0,0,0,234,0,163,0,166,0,19,0,8,0,150,0,0,0,26,0,165,0,95,0,0,0,169,0,0,0,79,0,149,0,43,0,153,0,183,0,186,0,139,0,254,0,32,0,234,0,126,0,238,0,69,0,240,0,77,0,204,0,178,0,0,0,60,0,118,0,0,0,0,0,55,0,136,0,123,0,219,0,0,0,75,0,239,0,49,0,134,0,209,0,232,0,63,0,0,0,0,0,116,0,21,0,77,0,19,0,200,0,0,0,0,0,151,0,122,0,67,0,100,0,159,0);
signal scenario_full  : scenario_type := (216,31,216,30,105,31,89,31,135,31,43,31,43,30,127,31,171,31,67,31,28,31,198,31,252,31,252,30,131,31,67,31,67,30,67,29,243,31,227,31,103,31,217,31,11,31,204,31,204,30,240,31,190,31,190,30,6,31,43,31,188,31,250,31,33,31,33,30,31,31,44,31,156,31,217,31,2,31,251,31,169,31,98,31,98,30,41,31,132,31,173,31,24,31,101,31,156,31,18,31,236,31,37,31,225,31,128,31,218,31,238,31,29,31,112,31,152,31,123,31,71,31,217,31,56,31,78,31,174,31,174,30,167,31,153,31,234,31,234,30,195,31,241,31,89,31,89,30,89,29,112,31,35,31,133,31,172,31,85,31,252,31,213,31,91,31,96,31,14,31,14,30,175,31,20,31,190,31,60,31,205,31,129,31,129,30,223,31,38,31,234,31,234,30,234,29,150,31,53,31,151,31,104,31,242,31,175,31,26,31,26,30,26,29,26,28,58,31,32,31,63,31,91,31,91,30,219,31,48,31,71,31,166,31,166,30,130,31,75,31,75,30,86,31,22,31,22,30,22,29,47,31,134,31,134,30,237,31,205,31,69,31,96,31,63,31,35,31,11,31,83,31,205,31,205,30,205,29,172,31,172,30,161,31,29,31,115,31,55,31,55,30,102,31,31,31,116,31,116,30,116,29,218,31,47,31,11,31,111,31,164,31,164,30,198,31,108,31,164,31,43,31,179,31,66,31,215,31,215,30,181,31,255,31,60,31,165,31,79,31,65,31,202,31,202,30,35,31,35,30,35,29,109,31,7,31,115,31,70,31,123,31,98,31,86,31,96,31,239,31,233,31,229,31,229,30,129,31,144,31,244,31,244,30,166,31,7,31,29,31,66,31,135,31,128,31,6,31,6,30,62,31,241,31,241,30,241,29,120,31,95,31,156,31,240,31,169,31,14,31,48,31,58,31,27,31,61,31,29,31,242,31,151,31,85,31,163,31,163,30,163,29,55,31,46,31,168,31,168,30,75,31,86,31,230,31,185,31,36,31,57,31,233,31,51,31,130,31,111,31,230,31,43,31,100,31,100,30,10,31,137,31,17,31,17,30,140,31,145,31,51,31,127,31,241,31,89,31,36,31,36,30,36,31,197,31,110,31,110,30,99,31,21,31,252,31,130,31,130,31,202,31,49,31,49,30,31,31,19,31,187,31,141,31,242,31,123,31,123,30,182,31,182,30,182,29,147,31,210,31,210,31,229,31,4,31,114,31,121,31,121,30,207,31,67,31,219,31,219,30,219,29,219,28,23,31,23,30,178,31,33,31,87,31,131,31,245,31,85,31,154,31,49,31,219,31,245,31,245,30,245,29,140,31,167,31,209,31,160,31,91,31,98,31,220,31,148,31,148,30,95,31,14,31,34,31,34,30,28,31,28,30,98,31,98,30,244,31,125,31,125,30,91,31,228,31,162,31,162,30,78,31,136,31,229,31,57,31,175,31,48,31,179,31,179,30,22,31,22,30,65,31,173,31,136,31,225,31,98,31,137,31,144,31,83,31,134,31,222,31,133,31,19,31,245,31,93,31,43,31,72,31,5,31,5,30,194,31,102,31,77,31,239,31,84,31,16,31,166,31,69,31,43,31,172,31,5,31,90,31,138,31,138,30,138,29,138,28,51,31,58,31,19,31,172,31,132,31,77,31,211,31,140,31,202,31,208,31,191,31,192,31,210,31,56,31,22,31,154,31,254,31,14,31,240,31,240,30,240,31,71,31,198,31,205,31,205,30,205,29,69,31,199,31,23,31,23,30,237,31,237,30,231,31,79,31,31,31,245,31,39,31,83,31,72,31,250,31,250,30,250,29,243,31,225,31,69,31,91,31,29,31,29,30,200,31,168,31,67,31,221,31,202,31,202,30,136,31,136,30,136,29,240,31,42,31,106,31,118,31,21,31,148,31,4,31,234,31,233,31,240,31,222,31,222,30,168,31,139,31,168,31,27,31,42,31,178,31,178,30,242,31,105,31,130,31,60,31,92,31,186,31,173,31,206,31,204,31,95,31,19,31,134,31,134,30,194,31,173,31,194,31,100,31,212,31,239,31,195,31,106,31,83,31,125,31,133,31,133,30,133,29,25,31,25,30,225,31,225,30,42,31,42,30,42,29,29,31,8,31,201,31,36,31,250,31,205,31,34,31,198,31,67,31,248,31,93,31,187,31,166,31,255,31,230,31,78,31,5,31,5,30,186,31,80,31,80,30,80,29,80,28,180,31,138,31,62,31,123,31,49,31,163,31,192,31,192,30,206,31,18,31,18,30,247,31,183,31,76,31,76,30,254,31,37,31,119,31,111,31,19,31,231,31,73,31,73,30,252,31,162,31,198,31,198,30,78,31,224,31,37,31,114,31,18,31,137,31,211,31,171,31,116,31,116,30,116,29,77,31,249,31,249,30,223,31,221,31,109,31,23,31,23,30,183,31,246,31,146,31,208,31,144,31,1,31,1,30,192,31,175,31,12,31,12,30,193,31,193,30,179,31,36,31,36,30,36,29,221,31,243,31,47,31,207,31,207,30,152,31,184,31,184,30,207,31,108,31,121,31,6,31,125,31,27,31,41,31,1,31,109,31,78,31,78,30,61,31,227,31,194,31,242,31,170,31,1,31,50,31,50,30,50,29,33,31,109,31,7,31,231,31,106,31,20,31,45,31,92,31,39,31,81,31,89,31,89,30,89,29,224,31,205,31,92,31,30,31,80,31,155,31,85,31,249,31,154,31,68,31,68,30,96,31,201,31,143,31,143,30,177,31,151,31,151,30,100,31,148,31,199,31,147,31,11,31,119,31,33,31,54,31,180,31,245,31,120,31,39,31,39,30,129,31,16,31,33,31,117,31,218,31,215,31,215,30,215,29,242,31,163,31,241,31,56,31,192,31,170,31,75,31,105,31,71,31,78,31,180,31,232,31,238,31,83,31,44,31,239,31,169,31,103,31,103,30,32,31,220,31,192,31,242,31,242,30,242,29,199,31,93,31,77,31,61,31,139,31,139,30,139,29,139,28,127,31,56,31,56,30,168,31,248,31,248,30,173,31,179,31,223,31,223,30,249,31,28,31,28,30,28,29,103,31,225,31,231,31,231,30,150,31,162,31,171,31,39,31,19,31,23,31,7,31,144,31,144,30,184,31,196,31,189,31,68,31,166,31,166,30,173,31,211,31,164,31,77,31,245,31,230,31,134,31,6,31,223,31,223,30,50,31,78,31,12,31,242,31,211,31,231,31,91,31,181,31,206,31,11,31,15,31,24,31,24,30,24,29,234,31,163,31,166,31,19,31,8,31,150,31,150,30,26,31,165,31,95,31,95,30,169,31,169,30,79,31,149,31,43,31,153,31,183,31,186,31,139,31,254,31,32,31,234,31,126,31,238,31,69,31,240,31,77,31,204,31,178,31,178,30,60,31,118,31,118,30,118,29,55,31,136,31,123,31,219,31,219,30,75,31,239,31,49,31,134,31,209,31,232,31,63,31,63,30,63,29,116,31,21,31,77,31,19,31,200,31,200,30,200,29,151,31,122,31,67,31,100,31,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
