-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 754;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (72,0,255,0,0,0,148,0,0,0,204,0,118,0,222,0,174,0,212,0,14,0,95,0,43,0,0,0,33,0,226,0,143,0,114,0,22,0,115,0,0,0,139,0,78,0,227,0,10,0,145,0,164,0,93,0,0,0,23,0,0,0,58,0,0,0,39,0,48,0,174,0,217,0,109,0,0,0,191,0,52,0,68,0,171,0,217,0,0,0,111,0,54,0,0,0,161,0,222,0,52,0,0,0,0,0,241,0,85,0,7,0,120,0,36,0,123,0,11,0,175,0,0,0,218,0,0,0,0,0,201,0,20,0,216,0,21,0,137,0,54,0,0,0,53,0,136,0,2,0,223,0,239,0,190,0,199,0,252,0,28,0,0,0,138,0,23,0,237,0,76,0,202,0,0,0,28,0,72,0,83,0,196,0,73,0,87,0,0,0,217,0,0,0,158,0,0,0,0,0,0,0,185,0,137,0,243,0,115,0,64,0,194,0,176,0,59,0,30,0,138,0,108,0,0,0,121,0,200,0,249,0,0,0,0,0,191,0,197,0,118,0,249,0,117,0,10,0,6,0,128,0,36,0,0,0,94,0,72,0,122,0,112,0,241,0,0,0,93,0,224,0,101,0,0,0,0,0,225,0,33,0,4,0,51,0,121,0,0,0,0,0,0,0,110,0,0,0,120,0,132,0,222,0,61,0,136,0,220,0,0,0,244,0,4,0,0,0,69,0,0,0,0,0,85,0,175,0,60,0,239,0,153,0,50,0,82,0,94,0,145,0,210,0,0,0,120,0,229,0,221,0,138,0,156,0,31,0,12,0,221,0,57,0,0,0,201,0,59,0,54,0,200,0,0,0,175,0,213,0,202,0,1,0,252,0,252,0,69,0,178,0,5,0,0,0,105,0,87,0,123,0,211,0,67,0,81,0,24,0,209,0,11,0,233,0,0,0,150,0,151,0,0,0,161,0,39,0,0,0,38,0,81,0,229,0,122,0,141,0,14,0,146,0,26,0,21,0,196,0,139,0,96,0,0,0,0,0,0,0,107,0,84,0,169,0,0,0,36,0,103,0,84,0,3,0,2,0,25,0,3,0,39,0,150,0,84,0,0,0,213,0,5,0,208,0,174,0,65,0,190,0,34,0,196,0,53,0,93,0,130,0,0,0,190,0,58,0,211,0,70,0,118,0,129,0,185,0,239,0,247,0,0,0,17,0,203,0,19,0,0,0,155,0,166,0,194,0,0,0,87,0,69,0,145,0,55,0,3,0,114,0,120,0,59,0,255,0,55,0,181,0,104,0,128,0,0,0,88,0,15,0,45,0,154,0,160,0,34,0,0,0,189,0,30,0,54,0,156,0,159,0,21,0,0,0,126,0,44,0,193,0,136,0,0,0,62,0,0,0,100,0,69,0,53,0,33,0,42,0,239,0,180,0,205,0,79,0,96,0,0,0,163,0,5,0,213,0,207,0,74,0,0,0,154,0,109,0,0,0,0,0,128,0,61,0,0,0,0,0,137,0,45,0,93,0,0,0,85,0,10,0,133,0,100,0,0,0,228,0,211,0,92,0,0,0,86,0,0,0,0,0,95,0,59,0,22,0,0,0,143,0,24,0,147,0,118,0,0,0,0,0,160,0,220,0,103,0,211,0,25,0,201,0,239,0,159,0,0,0,157,0,221,0,0,0,62,0,0,0,0,0,5,0,163,0,165,0,35,0,100,0,63,0,0,0,34,0,58,0,33,0,43,0,155,0,0,0,44,0,137,0,213,0,26,0,140,0,119,0,0,0,34,0,227,0,153,0,3,0,131,0,113,0,38,0,144,0,138,0,196,0,128,0,197,0,0,0,161,0,131,0,5,0,0,0,169,0,0,0,35,0,0,0,52,0,162,0,193,0,179,0,17,0,14,0,137,0,0,0,142,0,234,0,48,0,216,0,188,0,206,0,33,0,0,0,132,0,196,0,171,0,230,0,86,0,34,0,177,0,10,0,0,0,0,0,66,0,49,0,195,0,61,0,198,0,68,0,123,0,125,0,115,0,187,0,0,0,172,0,122,0,124,0,0,0,190,0,200,0,0,0,147,0,0,0,246,0,93,0,0,0,0,0,73,0,58,0,56,0,0,0,14,0,137,0,0,0,188,0,56,0,20,0,88,0,181,0,90,0,145,0,254,0,0,0,0,0,8,0,0,0,9,0,114,0,202,0,75,0,0,0,0,0,72,0,12,0,171,0,219,0,0,0,203,0,126,0,0,0,0,0,33,0,235,0,109,0,69,0,232,0,159,0,173,0,116,0,197,0,156,0,0,0,0,0,241,0,192,0,83,0,0,0,10,0,129,0,85,0,0,0,175,0,183,0,137,0,3,0,86,0,47,0,0,0,78,0,172,0,14,0,34,0,0,0,11,0,126,0,25,0,216,0,12,0,237,0,226,0,159,0,87,0,10,0,0,0,50,0,109,0,223,0,111,0,44,0,0,0,96,0,15,0,63,0,254,0,0,0,239,0,222,0,163,0,52,0,199,0,95,0,76,0,223,0,50,0,44,0,122,0,40,0,0,0,150,0,209,0,239,0,156,0,122,0,74,0,149,0,255,0,8,0,0,0,24,0,0,0,47,0,170,0,0,0,1,0,45,0,0,0,0,0,70,0,0,0,70,0,0,0,171,0,70,0,163,0,0,0,211,0,157,0,113,0,147,0,1,0,32,0,36,0,184,0,241,0,37,0,159,0,26,0,0,0,222,0,95,0,82,0,0,0,220,0,165,0,227,0,0,0,0,0,143,0,0,0,206,0,0,0,2,0,57,0,107,0,82,0,189,0,0,0,0,0,59,0,230,0,224,0,167,0,0,0,254,0,123,0,37,0,232,0,206,0,52,0,97,0,214,0,18,0,156,0,79,0,72,0,237,0,0,0,242,0,209,0,115,0,199,0,0,0,77,0,233,0,241,0,92,0,127,0,101,0,233,0,23,0,253,0,221,0,3,0,151,0,45,0,188,0,166,0,0,0,2,0,67,0,81,0,0,0,244,0,73,0,22,0,22,0,220,0,0,0,0,0,129,0,92,0,91,0,90,0,13,0,26,0,129,0,0,0,133,0,19,0,22,0,194,0,253,0,0,0,166,0,2,0,0,0,0,0,0,0,0,0,254,0,35,0,0,0,22,0,139,0,57,0,180,0,165,0,20,0,187,0,125,0,200,0,130,0,81,0,0,0,1,0,29,0,143,0,57,0,161,0,128,0,0,0,141,0,175,0,240,0,100,0,0,0,176,0,12,0,182,0,254,0,6,0,178,0,0,0,52,0,224,0,0,0,136,0,76,0,0,0,63,0,191,0,76,0,105,0,10,0,107,0,0,0,128,0,66,0,45,0,244,0,59,0,0,0,179,0,49,0);
signal scenario_full  : scenario_type := (72,31,255,31,255,30,148,31,148,30,204,31,118,31,222,31,174,31,212,31,14,31,95,31,43,31,43,30,33,31,226,31,143,31,114,31,22,31,115,31,115,30,139,31,78,31,227,31,10,31,145,31,164,31,93,31,93,30,23,31,23,30,58,31,58,30,39,31,48,31,174,31,217,31,109,31,109,30,191,31,52,31,68,31,171,31,217,31,217,30,111,31,54,31,54,30,161,31,222,31,52,31,52,30,52,29,241,31,85,31,7,31,120,31,36,31,123,31,11,31,175,31,175,30,218,31,218,30,218,29,201,31,20,31,216,31,21,31,137,31,54,31,54,30,53,31,136,31,2,31,223,31,239,31,190,31,199,31,252,31,28,31,28,30,138,31,23,31,237,31,76,31,202,31,202,30,28,31,72,31,83,31,196,31,73,31,87,31,87,30,217,31,217,30,158,31,158,30,158,29,158,28,185,31,137,31,243,31,115,31,64,31,194,31,176,31,59,31,30,31,138,31,108,31,108,30,121,31,200,31,249,31,249,30,249,29,191,31,197,31,118,31,249,31,117,31,10,31,6,31,128,31,36,31,36,30,94,31,72,31,122,31,112,31,241,31,241,30,93,31,224,31,101,31,101,30,101,29,225,31,33,31,4,31,51,31,121,31,121,30,121,29,121,28,110,31,110,30,120,31,132,31,222,31,61,31,136,31,220,31,220,30,244,31,4,31,4,30,69,31,69,30,69,29,85,31,175,31,60,31,239,31,153,31,50,31,82,31,94,31,145,31,210,31,210,30,120,31,229,31,221,31,138,31,156,31,31,31,12,31,221,31,57,31,57,30,201,31,59,31,54,31,200,31,200,30,175,31,213,31,202,31,1,31,252,31,252,31,69,31,178,31,5,31,5,30,105,31,87,31,123,31,211,31,67,31,81,31,24,31,209,31,11,31,233,31,233,30,150,31,151,31,151,30,161,31,39,31,39,30,38,31,81,31,229,31,122,31,141,31,14,31,146,31,26,31,21,31,196,31,139,31,96,31,96,30,96,29,96,28,107,31,84,31,169,31,169,30,36,31,103,31,84,31,3,31,2,31,25,31,3,31,39,31,150,31,84,31,84,30,213,31,5,31,208,31,174,31,65,31,190,31,34,31,196,31,53,31,93,31,130,31,130,30,190,31,58,31,211,31,70,31,118,31,129,31,185,31,239,31,247,31,247,30,17,31,203,31,19,31,19,30,155,31,166,31,194,31,194,30,87,31,69,31,145,31,55,31,3,31,114,31,120,31,59,31,255,31,55,31,181,31,104,31,128,31,128,30,88,31,15,31,45,31,154,31,160,31,34,31,34,30,189,31,30,31,54,31,156,31,159,31,21,31,21,30,126,31,44,31,193,31,136,31,136,30,62,31,62,30,100,31,69,31,53,31,33,31,42,31,239,31,180,31,205,31,79,31,96,31,96,30,163,31,5,31,213,31,207,31,74,31,74,30,154,31,109,31,109,30,109,29,128,31,61,31,61,30,61,29,137,31,45,31,93,31,93,30,85,31,10,31,133,31,100,31,100,30,228,31,211,31,92,31,92,30,86,31,86,30,86,29,95,31,59,31,22,31,22,30,143,31,24,31,147,31,118,31,118,30,118,29,160,31,220,31,103,31,211,31,25,31,201,31,239,31,159,31,159,30,157,31,221,31,221,30,62,31,62,30,62,29,5,31,163,31,165,31,35,31,100,31,63,31,63,30,34,31,58,31,33,31,43,31,155,31,155,30,44,31,137,31,213,31,26,31,140,31,119,31,119,30,34,31,227,31,153,31,3,31,131,31,113,31,38,31,144,31,138,31,196,31,128,31,197,31,197,30,161,31,131,31,5,31,5,30,169,31,169,30,35,31,35,30,52,31,162,31,193,31,179,31,17,31,14,31,137,31,137,30,142,31,234,31,48,31,216,31,188,31,206,31,33,31,33,30,132,31,196,31,171,31,230,31,86,31,34,31,177,31,10,31,10,30,10,29,66,31,49,31,195,31,61,31,198,31,68,31,123,31,125,31,115,31,187,31,187,30,172,31,122,31,124,31,124,30,190,31,200,31,200,30,147,31,147,30,246,31,93,31,93,30,93,29,73,31,58,31,56,31,56,30,14,31,137,31,137,30,188,31,56,31,20,31,88,31,181,31,90,31,145,31,254,31,254,30,254,29,8,31,8,30,9,31,114,31,202,31,75,31,75,30,75,29,72,31,12,31,171,31,219,31,219,30,203,31,126,31,126,30,126,29,33,31,235,31,109,31,69,31,232,31,159,31,173,31,116,31,197,31,156,31,156,30,156,29,241,31,192,31,83,31,83,30,10,31,129,31,85,31,85,30,175,31,183,31,137,31,3,31,86,31,47,31,47,30,78,31,172,31,14,31,34,31,34,30,11,31,126,31,25,31,216,31,12,31,237,31,226,31,159,31,87,31,10,31,10,30,50,31,109,31,223,31,111,31,44,31,44,30,96,31,15,31,63,31,254,31,254,30,239,31,222,31,163,31,52,31,199,31,95,31,76,31,223,31,50,31,44,31,122,31,40,31,40,30,150,31,209,31,239,31,156,31,122,31,74,31,149,31,255,31,8,31,8,30,24,31,24,30,47,31,170,31,170,30,1,31,45,31,45,30,45,29,70,31,70,30,70,31,70,30,171,31,70,31,163,31,163,30,211,31,157,31,113,31,147,31,1,31,32,31,36,31,184,31,241,31,37,31,159,31,26,31,26,30,222,31,95,31,82,31,82,30,220,31,165,31,227,31,227,30,227,29,143,31,143,30,206,31,206,30,2,31,57,31,107,31,82,31,189,31,189,30,189,29,59,31,230,31,224,31,167,31,167,30,254,31,123,31,37,31,232,31,206,31,52,31,97,31,214,31,18,31,156,31,79,31,72,31,237,31,237,30,242,31,209,31,115,31,199,31,199,30,77,31,233,31,241,31,92,31,127,31,101,31,233,31,23,31,253,31,221,31,3,31,151,31,45,31,188,31,166,31,166,30,2,31,67,31,81,31,81,30,244,31,73,31,22,31,22,31,220,31,220,30,220,29,129,31,92,31,91,31,90,31,13,31,26,31,129,31,129,30,133,31,19,31,22,31,194,31,253,31,253,30,166,31,2,31,2,30,2,29,2,28,2,27,254,31,35,31,35,30,22,31,139,31,57,31,180,31,165,31,20,31,187,31,125,31,200,31,130,31,81,31,81,30,1,31,29,31,143,31,57,31,161,31,128,31,128,30,141,31,175,31,240,31,100,31,100,30,176,31,12,31,182,31,254,31,6,31,178,31,178,30,52,31,224,31,224,30,136,31,76,31,76,30,63,31,191,31,76,31,105,31,10,31,107,31,107,30,128,31,66,31,45,31,244,31,59,31,59,30,179,31,49,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
