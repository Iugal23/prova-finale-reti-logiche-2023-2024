-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 473;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,157,0,155,0,49,0,208,0,0,0,0,0,0,0,0,0,0,0,0,0,227,0,248,0,4,0,222,0,83,0,161,0,254,0,0,0,188,0,207,0,181,0,137,0,52,0,59,0,27,0,255,0,30,0,0,0,0,0,162,0,0,0,10,0,32,0,43,0,0,0,183,0,20,0,152,0,0,0,0,0,34,0,203,0,45,0,179,0,101,0,196,0,193,0,33,0,230,0,7,0,183,0,175,0,0,0,37,0,209,0,116,0,0,0,15,0,21,0,106,0,0,0,83,0,86,0,0,0,136,0,237,0,128,0,39,0,105,0,109,0,74,0,181,0,82,0,0,0,0,0,15,0,54,0,210,0,0,0,174,0,0,0,68,0,226,0,181,0,0,0,0,0,66,0,59,0,0,0,4,0,68,0,0,0,0,0,67,0,225,0,99,0,247,0,245,0,95,0,0,0,0,0,158,0,0,0,135,0,239,0,252,0,232,0,26,0,173,0,130,0,44,0,237,0,159,0,38,0,0,0,234,0,181,0,95,0,114,0,0,0,216,0,191,0,139,0,95,0,243,0,73,0,0,0,77,0,52,0,0,0,176,0,161,0,0,0,19,0,102,0,176,0,0,0,212,0,56,0,7,0,195,0,214,0,88,0,218,0,0,0,62,0,126,0,166,0,83,0,179,0,89,0,21,0,217,0,79,0,3,0,199,0,74,0,225,0,100,0,86,0,0,0,164,0,82,0,0,0,72,0,136,0,191,0,202,0,177,0,0,0,139,0,0,0,122,0,216,0,35,0,151,0,222,0,214,0,40,0,0,0,181,0,0,0,186,0,59,0,0,0,162,0,76,0,175,0,222,0,0,0,86,0,68,0,0,0,85,0,233,0,0,0,26,0,229,0,230,0,245,0,225,0,198,0,16,0,0,0,0,0,102,0,199,0,0,0,28,0,144,0,200,0,174,0,215,0,136,0,217,0,182,0,0,0,207,0,112,0,0,0,0,0,93,0,104,0,225,0,125,0,154,0,163,0,249,0,27,0,33,0,56,0,0,0,0,0,207,0,0,0,8,0,14,0,0,0,64,0,204,0,106,0,0,0,240,0,72,0,137,0,78,0,253,0,0,0,65,0,189,0,188,0,0,0,177,0,183,0,54,0,0,0,0,0,197,0,70,0,161,0,193,0,0,0,0,0,45,0,0,0,0,0,0,0,217,0,0,0,227,0,87,0,0,0,145,0,178,0,101,0,0,0,61,0,0,0,195,0,13,0,112,0,106,0,55,0,0,0,159,0,175,0,0,0,226,0,215,0,73,0,28,0,0,0,12,0,165,0,0,0,246,0,0,0,0,0,7,0,18,0,0,0,99,0,71,0,56,0,194,0,129,0,84,0,0,0,0,0,122,0,130,0,142,0,0,0,90,0,91,0,251,0,0,0,181,0,31,0,0,0,205,0,149,0,187,0,122,0,49,0,81,0,88,0,197,0,45,0,0,0,225,0,0,0,0,0,80,0,0,0,167,0,0,0,137,0,151,0,58,0,81,0,119,0,238,0,34,0,236,0,18,0,0,0,237,0,0,0,111,0,0,0,11,0,255,0,0,0,161,0,0,0,18,0,134,0,168,0,213,0,0,0,55,0,155,0,0,0,51,0,27,0,212,0,211,0,157,0,133,0,8,0,238,0,255,0,0,0,76,0,247,0,227,0,61,0,0,0,186,0,216,0,30,0,163,0,182,0,69,0,147,0,0,0,0,0,209,0,0,0,138,0,155,0,69,0,0,0,101,0,199,0,43,0,83,0,162,0,207,0,28,0,0,0,172,0,185,0,88,0,0,0,104,0,0,0,89,0,237,0,111,0,149,0,138,0,4,0,242,0,94,0,254,0,4,0,253,0,147,0,124,0,61,0,241,0,54,0,85,0,187,0,39,0,193,0,203,0,0,0,149,0,201,0,232,0,0,0,16,0,0,0,35,0,176,0,236,0,0,0,0,0,240,0,61,0,171,0,242,0,217,0,152,0,27,0,112,0,239,0,179,0,33,0,105,0,78,0,168,0,223,0,194,0,0,0,77,0,0,0,81,0,208,0,152,0,49,0,211,0,131,0,66,0,62,0,49,0,63,0,6,0,106,0);
signal scenario_full  : scenario_type := (250,31,157,31,155,31,49,31,208,31,208,30,208,29,208,28,208,27,208,26,208,25,227,31,248,31,4,31,222,31,83,31,161,31,254,31,254,30,188,31,207,31,181,31,137,31,52,31,59,31,27,31,255,31,30,31,30,30,30,29,162,31,162,30,10,31,32,31,43,31,43,30,183,31,20,31,152,31,152,30,152,29,34,31,203,31,45,31,179,31,101,31,196,31,193,31,33,31,230,31,7,31,183,31,175,31,175,30,37,31,209,31,116,31,116,30,15,31,21,31,106,31,106,30,83,31,86,31,86,30,136,31,237,31,128,31,39,31,105,31,109,31,74,31,181,31,82,31,82,30,82,29,15,31,54,31,210,31,210,30,174,31,174,30,68,31,226,31,181,31,181,30,181,29,66,31,59,31,59,30,4,31,68,31,68,30,68,29,67,31,225,31,99,31,247,31,245,31,95,31,95,30,95,29,158,31,158,30,135,31,239,31,252,31,232,31,26,31,173,31,130,31,44,31,237,31,159,31,38,31,38,30,234,31,181,31,95,31,114,31,114,30,216,31,191,31,139,31,95,31,243,31,73,31,73,30,77,31,52,31,52,30,176,31,161,31,161,30,19,31,102,31,176,31,176,30,212,31,56,31,7,31,195,31,214,31,88,31,218,31,218,30,62,31,126,31,166,31,83,31,179,31,89,31,21,31,217,31,79,31,3,31,199,31,74,31,225,31,100,31,86,31,86,30,164,31,82,31,82,30,72,31,136,31,191,31,202,31,177,31,177,30,139,31,139,30,122,31,216,31,35,31,151,31,222,31,214,31,40,31,40,30,181,31,181,30,186,31,59,31,59,30,162,31,76,31,175,31,222,31,222,30,86,31,68,31,68,30,85,31,233,31,233,30,26,31,229,31,230,31,245,31,225,31,198,31,16,31,16,30,16,29,102,31,199,31,199,30,28,31,144,31,200,31,174,31,215,31,136,31,217,31,182,31,182,30,207,31,112,31,112,30,112,29,93,31,104,31,225,31,125,31,154,31,163,31,249,31,27,31,33,31,56,31,56,30,56,29,207,31,207,30,8,31,14,31,14,30,64,31,204,31,106,31,106,30,240,31,72,31,137,31,78,31,253,31,253,30,65,31,189,31,188,31,188,30,177,31,183,31,54,31,54,30,54,29,197,31,70,31,161,31,193,31,193,30,193,29,45,31,45,30,45,29,45,28,217,31,217,30,227,31,87,31,87,30,145,31,178,31,101,31,101,30,61,31,61,30,195,31,13,31,112,31,106,31,55,31,55,30,159,31,175,31,175,30,226,31,215,31,73,31,28,31,28,30,12,31,165,31,165,30,246,31,246,30,246,29,7,31,18,31,18,30,99,31,71,31,56,31,194,31,129,31,84,31,84,30,84,29,122,31,130,31,142,31,142,30,90,31,91,31,251,31,251,30,181,31,31,31,31,30,205,31,149,31,187,31,122,31,49,31,81,31,88,31,197,31,45,31,45,30,225,31,225,30,225,29,80,31,80,30,167,31,167,30,137,31,151,31,58,31,81,31,119,31,238,31,34,31,236,31,18,31,18,30,237,31,237,30,111,31,111,30,11,31,255,31,255,30,161,31,161,30,18,31,134,31,168,31,213,31,213,30,55,31,155,31,155,30,51,31,27,31,212,31,211,31,157,31,133,31,8,31,238,31,255,31,255,30,76,31,247,31,227,31,61,31,61,30,186,31,216,31,30,31,163,31,182,31,69,31,147,31,147,30,147,29,209,31,209,30,138,31,155,31,69,31,69,30,101,31,199,31,43,31,83,31,162,31,207,31,28,31,28,30,172,31,185,31,88,31,88,30,104,31,104,30,89,31,237,31,111,31,149,31,138,31,4,31,242,31,94,31,254,31,4,31,253,31,147,31,124,31,61,31,241,31,54,31,85,31,187,31,39,31,193,31,203,31,203,30,149,31,201,31,232,31,232,30,16,31,16,30,35,31,176,31,236,31,236,30,236,29,240,31,61,31,171,31,242,31,217,31,152,31,27,31,112,31,239,31,179,31,33,31,105,31,78,31,168,31,223,31,194,31,194,30,77,31,77,30,81,31,208,31,152,31,49,31,211,31,131,31,66,31,62,31,49,31,63,31,6,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
