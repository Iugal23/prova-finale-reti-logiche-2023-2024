-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 254;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (124,0,78,0,0,0,0,0,135,0,0,0,0,0,104,0,2,0,29,0,132,0,0,0,102,0,0,0,110,0,170,0,136,0,109,0,0,0,0,0,240,0,79,0,139,0,22,0,0,0,214,0,192,0,191,0,228,0,0,0,21,0,30,0,193,0,173,0,0,0,95,0,0,0,199,0,191,0,0,0,129,0,141,0,0,0,89,0,0,0,72,0,96,0,140,0,30,0,59,0,0,0,19,0,233,0,126,0,0,0,159,0,0,0,0,0,27,0,29,0,173,0,188,0,107,0,29,0,0,0,0,0,25,0,220,0,97,0,175,0,0,0,0,0,70,0,74,0,252,0,85,0,0,0,249,0,2,0,55,0,211,0,0,0,166,0,29,0,0,0,92,0,0,0,76,0,146,0,0,0,0,0,114,0,149,0,0,0,117,0,41,0,77,0,148,0,236,0,144,0,44,0,172,0,161,0,148,0,199,0,218,0,72,0,0,0,99,0,207,0,75,0,146,0,116,0,0,0,206,0,178,0,20,0,98,0,0,0,0,0,0,0,0,0,97,0,0,0,140,0,0,0,82,0,0,0,231,0,166,0,147,0,88,0,59,0,0,0,126,0,187,0,3,0,0,0,102,0,24,0,88,0,31,0,211,0,0,0,119,0,201,0,214,0,70,0,60,0,21,0,0,0,102,0,27,0,52,0,24,0,222,0,21,0,147,0,137,0,199,0,251,0,0,0,126,0,72,0,130,0,11,0,20,0,28,0,0,0,37,0,141,0,73,0,43,0,199,0,65,0,219,0,245,0,0,0,205,0,45,0,0,0,54,0,75,0,160,0,235,0,216,0,216,0,138,0,37,0,0,0,0,0,0,0,239,0,69,0,251,0,190,0,61,0,0,0,226,0,106,0,167,0,1,0,0,0,0,0,128,0,0,0,108,0,0,0,246,0,0,0,188,0,75,0,90,0,8,0,240,0,127,0,247,0,243,0,8,0,218,0,147,0,120,0,168,0,190,0,0,0,0,0,200,0,130,0,187,0,159,0,162,0,0,0,183,0,224,0,254,0,136,0,83,0,40,0,118,0,125,0,205,0,232,0,18,0,109,0,156,0,66,0,65,0,238,0,4,0,0,0,0,0,0,0,97,0,75,0);
signal scenario_full  : scenario_type := (124,31,78,31,78,30,78,29,135,31,135,30,135,29,104,31,2,31,29,31,132,31,132,30,102,31,102,30,110,31,170,31,136,31,109,31,109,30,109,29,240,31,79,31,139,31,22,31,22,30,214,31,192,31,191,31,228,31,228,30,21,31,30,31,193,31,173,31,173,30,95,31,95,30,199,31,191,31,191,30,129,31,141,31,141,30,89,31,89,30,72,31,96,31,140,31,30,31,59,31,59,30,19,31,233,31,126,31,126,30,159,31,159,30,159,29,27,31,29,31,173,31,188,31,107,31,29,31,29,30,29,29,25,31,220,31,97,31,175,31,175,30,175,29,70,31,74,31,252,31,85,31,85,30,249,31,2,31,55,31,211,31,211,30,166,31,29,31,29,30,92,31,92,30,76,31,146,31,146,30,146,29,114,31,149,31,149,30,117,31,41,31,77,31,148,31,236,31,144,31,44,31,172,31,161,31,148,31,199,31,218,31,72,31,72,30,99,31,207,31,75,31,146,31,116,31,116,30,206,31,178,31,20,31,98,31,98,30,98,29,98,28,98,27,97,31,97,30,140,31,140,30,82,31,82,30,231,31,166,31,147,31,88,31,59,31,59,30,126,31,187,31,3,31,3,30,102,31,24,31,88,31,31,31,211,31,211,30,119,31,201,31,214,31,70,31,60,31,21,31,21,30,102,31,27,31,52,31,24,31,222,31,21,31,147,31,137,31,199,31,251,31,251,30,126,31,72,31,130,31,11,31,20,31,28,31,28,30,37,31,141,31,73,31,43,31,199,31,65,31,219,31,245,31,245,30,205,31,45,31,45,30,54,31,75,31,160,31,235,31,216,31,216,31,138,31,37,31,37,30,37,29,37,28,239,31,69,31,251,31,190,31,61,31,61,30,226,31,106,31,167,31,1,31,1,30,1,29,128,31,128,30,108,31,108,30,246,31,246,30,188,31,75,31,90,31,8,31,240,31,127,31,247,31,243,31,8,31,218,31,147,31,120,31,168,31,190,31,190,30,190,29,200,31,130,31,187,31,159,31,162,31,162,30,183,31,224,31,254,31,136,31,83,31,40,31,118,31,125,31,205,31,232,31,18,31,109,31,156,31,66,31,65,31,238,31,4,31,4,30,4,29,4,28,97,31,75,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
