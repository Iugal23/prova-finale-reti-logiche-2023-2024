-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_124 is
end project_tb_124;

architecture project_tb_arch_124 of project_tb_124 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 691;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,33,0,167,0,29,0,105,0,226,0,0,0,0,0,64,0,0,0,0,0,56,0,224,0,215,0,138,0,209,0,93,0,134,0,63,0,33,0,58,0,0,0,189,0,115,0,190,0,121,0,100,0,129,0,156,0,135,0,8,0,190,0,251,0,19,0,0,0,223,0,193,0,0,0,164,0,8,0,183,0,252,0,0,0,239,0,54,0,129,0,154,0,34,0,134,0,45,0,9,0,232,0,142,0,236,0,220,0,251,0,252,0,0,0,113,0,40,0,0,0,182,0,139,0,0,0,176,0,61,0,0,0,162,0,135,0,209,0,230,0,114,0,0,0,2,0,0,0,243,0,42,0,0,0,21,0,32,0,137,0,11,0,90,0,210,0,146,0,0,0,115,0,247,0,61,0,44,0,48,0,38,0,238,0,249,0,6,0,0,0,134,0,187,0,119,0,18,0,205,0,85,0,78,0,166,0,203,0,71,0,192,0,114,0,25,0,0,0,161,0,139,0,19,0,255,0,0,0,60,0,22,0,0,0,136,0,117,0,76,0,201,0,95,0,223,0,37,0,90,0,87,0,0,0,35,0,65,0,116,0,195,0,76,0,5,0,183,0,25,0,0,0,31,0,5,0,39,0,0,0,14,0,0,0,175,0,135,0,174,0,5,0,42,0,116,0,6,0,0,0,9,0,243,0,144,0,134,0,82,0,83,0,73,0,0,0,94,0,13,0,60,0,128,0,209,0,141,0,0,0,0,0,160,0,253,0,123,0,108,0,95,0,164,0,0,0,63,0,0,0,7,0,43,0,244,0,79,0,152,0,0,0,0,0,0,0,64,0,179,0,193,0,247,0,6,0,176,0,0,0,29,0,0,0,0,0,88,0,79,0,78,0,60,0,0,0,0,0,0,0,244,0,182,0,123,0,52,0,0,0,0,0,100,0,83,0,113,0,94,0,7,0,33,0,74,0,0,0,132,0,94,0,242,0,107,0,152,0,22,0,106,0,36,0,157,0,127,0,195,0,60,0,0,0,0,0,134,0,141,0,114,0,63,0,9,0,86,0,0,0,96,0,73,0,205,0,206,0,69,0,0,0,209,0,246,0,153,0,0,0,200,0,238,0,9,0,56,0,249,0,151,0,168,0,0,0,41,0,15,0,223,0,162,0,98,0,119,0,148,0,0,0,158,0,0,0,136,0,0,0,161,0,39,0,22,0,150,0,56,0,215,0,0,0,213,0,0,0,96,0,0,0,219,0,86,0,191,0,75,0,55,0,39,0,233,0,161,0,0,0,7,0,114,0,0,0,63,0,249,0,76,0,44,0,15,0,140,0,168,0,113,0,103,0,213,0,0,0,145,0,53,0,0,0,53,0,70,0,167,0,0,0,143,0,13,0,138,0,19,0,52,0,50,0,0,0,50,0,105,0,132,0,249,0,0,0,155,0,221,0,0,0,49,0,195,0,197,0,51,0,38,0,93,0,0,0,180,0,253,0,45,0,0,0,77,0,217,0,0,0,141,0,43,0,0,0,127,0,232,0,141,0,0,0,202,0,202,0,0,0,205,0,14,0,163,0,186,0,249,0,0,0,82,0,95,0,0,0,241,0,0,0,0,0,158,0,131,0,22,0,148,0,47,0,38,0,16,0,147,0,106,0,210,0,99,0,204,0,159,0,124,0,148,0,181,0,158,0,0,0,0,0,178,0,170,0,56,0,9,0,164,0,55,0,121,0,150,0,0,0,112,0,0,0,231,0,82,0,0,0,33,0,129,0,201,0,45,0,250,0,253,0,0,0,221,0,199,0,39,0,61,0,0,0,174,0,0,0,106,0,48,0,0,0,228,0,0,0,198,0,202,0,165,0,0,0,155,0,196,0,0,0,126,0,65,0,143,0,102,0,73,0,0,0,49,0,0,0,240,0,16,0,94,0,83,0,196,0,141,0,128,0,139,0,8,0,223,0,161,0,138,0,133,0,255,0,128,0,61,0,92,0,93,0,149,0,118,0,0,0,52,0,102,0,241,0,110,0,211,0,0,0,252,0,131,0,253,0,228,0,219,0,164,0,50,0,189,0,165,0,186,0,144,0,0,0,171,0,237,0,12,0,1,0,203,0,83,0,229,0,115,0,0,0,90,0,120,0,208,0,154,0,35,0,84,0,224,0,219,0,82,0,205,0,15,0,0,0,172,0,230,0,193,0,0,0,203,0,178,0,179,0,159,0,148,0,241,0,0,0,74,0,40,0,207,0,50,0,238,0,130,0,118,0,60,0,203,0,0,0,73,0,24,0,88,0,178,0,0,0,0,0,230,0,244,0,158,0,249,0,229,0,222,0,250,0,240,0,72,0,69,0,0,0,112,0,170,0,0,0,181,0,0,0,110,0,23,0,0,0,53,0,0,0,0,0,69,0,33,0,0,0,252,0,0,0,0,0,0,0,224,0,214,0,40,0,0,0,166,0,147,0,109,0,174,0,62,0,48,0,40,0,232,0,0,0,50,0,173,0,167,0,167,0,97,0,245,0,107,0,108,0,243,0,14,0,21,0,76,0,132,0,0,0,0,0,159,0,215,0,0,0,235,0,199,0,0,0,91,0,217,0,27,0,115,0,130,0,211,0,176,0,16,0,55,0,122,0,99,0,33,0,107,0,70,0,5,0,29,0,252,0,28,0,122,0,32,0,68,0,0,0,114,0,0,0,186,0,184,0,34,0,102,0,0,0,2,0,186,0,114,0,103,0,55,0,147,0,145,0,5,0,19,0,23,0,41,0,216,0,241,0,178,0,103,0,0,0,0,0,179,0,242,0,38,0,9,0,179,0,0,0,174,0,0,0,66,0,66,0,194,0,97,0,1,0,0,0,0,0,0,0,65,0,82,0,0,0,13,0,76,0,232,0,189,0,157,0,76,0,233,0,249,0,153,0,238,0,81,0,123,0,7,0,209,0,47,0,204,0,238,0,170,0,0,0,13,0,233,0,252,0,197,0,116,0,190,0,94,0,223,0,109,0,37,0,229,0,55,0,116,0,241,0,1,0,119,0,123,0,170,0,25,0,11,0,78,0,179,0,218,0,109,0,208,0,150,0,221,0,137,0,132,0,243,0,0,0,8,0);
signal scenario_full  : scenario_type := (136,31,33,31,167,31,29,31,105,31,226,31,226,30,226,29,64,31,64,30,64,29,56,31,224,31,215,31,138,31,209,31,93,31,134,31,63,31,33,31,58,31,58,30,189,31,115,31,190,31,121,31,100,31,129,31,156,31,135,31,8,31,190,31,251,31,19,31,19,30,223,31,193,31,193,30,164,31,8,31,183,31,252,31,252,30,239,31,54,31,129,31,154,31,34,31,134,31,45,31,9,31,232,31,142,31,236,31,220,31,251,31,252,31,252,30,113,31,40,31,40,30,182,31,139,31,139,30,176,31,61,31,61,30,162,31,135,31,209,31,230,31,114,31,114,30,2,31,2,30,243,31,42,31,42,30,21,31,32,31,137,31,11,31,90,31,210,31,146,31,146,30,115,31,247,31,61,31,44,31,48,31,38,31,238,31,249,31,6,31,6,30,134,31,187,31,119,31,18,31,205,31,85,31,78,31,166,31,203,31,71,31,192,31,114,31,25,31,25,30,161,31,139,31,19,31,255,31,255,30,60,31,22,31,22,30,136,31,117,31,76,31,201,31,95,31,223,31,37,31,90,31,87,31,87,30,35,31,65,31,116,31,195,31,76,31,5,31,183,31,25,31,25,30,31,31,5,31,39,31,39,30,14,31,14,30,175,31,135,31,174,31,5,31,42,31,116,31,6,31,6,30,9,31,243,31,144,31,134,31,82,31,83,31,73,31,73,30,94,31,13,31,60,31,128,31,209,31,141,31,141,30,141,29,160,31,253,31,123,31,108,31,95,31,164,31,164,30,63,31,63,30,7,31,43,31,244,31,79,31,152,31,152,30,152,29,152,28,64,31,179,31,193,31,247,31,6,31,176,31,176,30,29,31,29,30,29,29,88,31,79,31,78,31,60,31,60,30,60,29,60,28,244,31,182,31,123,31,52,31,52,30,52,29,100,31,83,31,113,31,94,31,7,31,33,31,74,31,74,30,132,31,94,31,242,31,107,31,152,31,22,31,106,31,36,31,157,31,127,31,195,31,60,31,60,30,60,29,134,31,141,31,114,31,63,31,9,31,86,31,86,30,96,31,73,31,205,31,206,31,69,31,69,30,209,31,246,31,153,31,153,30,200,31,238,31,9,31,56,31,249,31,151,31,168,31,168,30,41,31,15,31,223,31,162,31,98,31,119,31,148,31,148,30,158,31,158,30,136,31,136,30,161,31,39,31,22,31,150,31,56,31,215,31,215,30,213,31,213,30,96,31,96,30,219,31,86,31,191,31,75,31,55,31,39,31,233,31,161,31,161,30,7,31,114,31,114,30,63,31,249,31,76,31,44,31,15,31,140,31,168,31,113,31,103,31,213,31,213,30,145,31,53,31,53,30,53,31,70,31,167,31,167,30,143,31,13,31,138,31,19,31,52,31,50,31,50,30,50,31,105,31,132,31,249,31,249,30,155,31,221,31,221,30,49,31,195,31,197,31,51,31,38,31,93,31,93,30,180,31,253,31,45,31,45,30,77,31,217,31,217,30,141,31,43,31,43,30,127,31,232,31,141,31,141,30,202,31,202,31,202,30,205,31,14,31,163,31,186,31,249,31,249,30,82,31,95,31,95,30,241,31,241,30,241,29,158,31,131,31,22,31,148,31,47,31,38,31,16,31,147,31,106,31,210,31,99,31,204,31,159,31,124,31,148,31,181,31,158,31,158,30,158,29,178,31,170,31,56,31,9,31,164,31,55,31,121,31,150,31,150,30,112,31,112,30,231,31,82,31,82,30,33,31,129,31,201,31,45,31,250,31,253,31,253,30,221,31,199,31,39,31,61,31,61,30,174,31,174,30,106,31,48,31,48,30,228,31,228,30,198,31,202,31,165,31,165,30,155,31,196,31,196,30,126,31,65,31,143,31,102,31,73,31,73,30,49,31,49,30,240,31,16,31,94,31,83,31,196,31,141,31,128,31,139,31,8,31,223,31,161,31,138,31,133,31,255,31,128,31,61,31,92,31,93,31,149,31,118,31,118,30,52,31,102,31,241,31,110,31,211,31,211,30,252,31,131,31,253,31,228,31,219,31,164,31,50,31,189,31,165,31,186,31,144,31,144,30,171,31,237,31,12,31,1,31,203,31,83,31,229,31,115,31,115,30,90,31,120,31,208,31,154,31,35,31,84,31,224,31,219,31,82,31,205,31,15,31,15,30,172,31,230,31,193,31,193,30,203,31,178,31,179,31,159,31,148,31,241,31,241,30,74,31,40,31,207,31,50,31,238,31,130,31,118,31,60,31,203,31,203,30,73,31,24,31,88,31,178,31,178,30,178,29,230,31,244,31,158,31,249,31,229,31,222,31,250,31,240,31,72,31,69,31,69,30,112,31,170,31,170,30,181,31,181,30,110,31,23,31,23,30,53,31,53,30,53,29,69,31,33,31,33,30,252,31,252,30,252,29,252,28,224,31,214,31,40,31,40,30,166,31,147,31,109,31,174,31,62,31,48,31,40,31,232,31,232,30,50,31,173,31,167,31,167,31,97,31,245,31,107,31,108,31,243,31,14,31,21,31,76,31,132,31,132,30,132,29,159,31,215,31,215,30,235,31,199,31,199,30,91,31,217,31,27,31,115,31,130,31,211,31,176,31,16,31,55,31,122,31,99,31,33,31,107,31,70,31,5,31,29,31,252,31,28,31,122,31,32,31,68,31,68,30,114,31,114,30,186,31,184,31,34,31,102,31,102,30,2,31,186,31,114,31,103,31,55,31,147,31,145,31,5,31,19,31,23,31,41,31,216,31,241,31,178,31,103,31,103,30,103,29,179,31,242,31,38,31,9,31,179,31,179,30,174,31,174,30,66,31,66,31,194,31,97,31,1,31,1,30,1,29,1,28,65,31,82,31,82,30,13,31,76,31,232,31,189,31,157,31,76,31,233,31,249,31,153,31,238,31,81,31,123,31,7,31,209,31,47,31,204,31,238,31,170,31,170,30,13,31,233,31,252,31,197,31,116,31,190,31,94,31,223,31,109,31,37,31,229,31,55,31,116,31,241,31,1,31,119,31,123,31,170,31,25,31,11,31,78,31,179,31,218,31,109,31,208,31,150,31,221,31,137,31,132,31,243,31,243,30,8,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
