-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 919;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (10,0,173,0,148,0,209,0,253,0,213,0,99,0,34,0,38,0,148,0,217,0,150,0,107,0,121,0,226,0,170,0,110,0,88,0,219,0,56,0,0,0,0,0,153,0,166,0,224,0,0,0,0,0,215,0,0,0,213,0,103,0,0,0,70,0,115,0,143,0,0,0,160,0,232,0,0,0,81,0,114,0,0,0,227,0,0,0,236,0,41,0,42,0,135,0,10,0,8,0,205,0,76,0,209,0,203,0,252,0,218,0,0,0,0,0,0,0,25,0,0,0,7,0,82,0,191,0,0,0,38,0,0,0,0,0,0,0,167,0,244,0,0,0,247,0,88,0,220,0,216,0,47,0,0,0,0,0,122,0,155,0,252,0,151,0,53,0,255,0,172,0,173,0,0,0,190,0,26,0,9,0,110,0,0,0,218,0,218,0,67,0,147,0,238,0,159,0,224,0,0,0,146,0,0,0,220,0,203,0,163,0,0,0,239,0,6,0,47,0,113,0,67,0,156,0,0,0,246,0,251,0,30,0,0,0,253,0,167,0,128,0,0,0,252,0,20,0,0,0,0,0,191,0,122,0,0,0,36,0,0,0,169,0,166,0,251,0,179,0,0,0,164,0,4,0,58,0,21,0,191,0,87,0,110,0,170,0,23,0,0,0,137,0,167,0,0,0,153,0,205,0,41,0,157,0,191,0,13,0,0,0,170,0,0,0,229,0,0,0,204,0,36,0,5,0,182,0,0,0,242,0,80,0,245,0,38,0,0,0,41,0,94,0,111,0,26,0,0,0,0,0,0,0,0,0,161,0,175,0,98,0,226,0,0,0,239,0,0,0,0,0,174,0,189,0,8,0,6,0,0,0,193,0,55,0,206,0,202,0,35,0,140,0,204,0,21,0,93,0,251,0,0,0,119,0,0,0,197,0,0,0,186,0,157,0,53,0,0,0,169,0,0,0,48,0,6,0,0,0,7,0,168,0,0,0,0,0,172,0,192,0,32,0,0,0,0,0,166,0,49,0,185,0,126,0,165,0,13,0,211,0,205,0,190,0,48,0,0,0,0,0,210,0,224,0,0,0,233,0,163,0,2,0,76,0,214,0,72,0,251,0,209,0,125,0,15,0,0,0,0,0,205,0,32,0,235,0,30,0,110,0,191,0,71,0,83,0,253,0,17,0,0,0,212,0,232,0,199,0,218,0,131,0,254,0,0,0,86,0,251,0,177,0,12,0,118,0,50,0,41,0,0,0,0,0,215,0,153,0,0,0,129,0,0,0,88,0,74,0,0,0,0,0,86,0,58,0,249,0,245,0,52,0,0,0,93,0,0,0,130,0,0,0,60,0,0,0,65,0,224,0,194,0,22,0,79,0,0,0,191,0,0,0,125,0,0,0,218,0,167,0,104,0,197,0,88,0,18,0,0,0,12,0,225,0,209,0,122,0,42,0,110,0,156,0,130,0,75,0,85,0,26,0,207,0,47,0,59,0,0,0,53,0,248,0,58,0,0,0,153,0,0,0,0,0,18,0,132,0,0,0,113,0,99,0,228,0,236,0,220,0,117,0,151,0,0,0,49,0,40,0,0,0,0,0,0,0,0,0,79,0,182,0,186,0,0,0,152,0,254,0,109,0,158,0,153,0,0,0,222,0,88,0,137,0,50,0,179,0,46,0,76,0,226,0,57,0,146,0,0,0,97,0,0,0,215,0,0,0,29,0,237,0,0,0,0,0,47,0,59,0,79,0,82,0,209,0,0,0,0,0,95,0,0,0,147,0,0,0,118,0,0,0,0,0,102,0,224,0,168,0,23,0,238,0,4,0,242,0,128,0,18,0,205,0,85,0,0,0,136,0,0,0,115,0,215,0,42,0,16,0,165,0,130,0,113,0,75,0,112,0,198,0,0,0,0,0,84,0,47,0,0,0,0,0,1,0,198,0,181,0,0,0,0,0,66,0,107,0,40,0,218,0,235,0,0,0,117,0,120,0,0,0,171,0,161,0,102,0,250,0,0,0,65,0,239,0,11,0,6,0,0,0,72,0,57,0,103,0,244,0,76,0,90,0,186,0,14,0,118,0,234,0,133,0,201,0,54,0,172,0,0,0,153,0,0,0,134,0,0,0,102,0,171,0,0,0,139,0,96,0,240,0,0,0,159,0,154,0,142,0,196,0,37,0,45,0,105,0,53,0,31,0,0,0,39,0,42,0,119,0,246,0,249,0,2,0,245,0,134,0,184,0,240,0,243,0,0,0,146,0,158,0,73,0,37,0,0,0,241,0,0,0,55,0,0,0,233,0,245,0,188,0,0,0,199,0,0,0,133,0,197,0,0,0,0,0,0,0,210,0,166,0,199,0,0,0,46,0,46,0,21,0,222,0,196,0,0,0,24,0,81,0,5,0,94,0,155,0,104,0,97,0,26,0,125,0,0,0,77,0,207,0,0,0,155,0,57,0,126,0,188,0,131,0,254,0,133,0,177,0,0,0,110,0,193,0,106,0,227,0,0,0,0,0,84,0,12,0,130,0,164,0,96,0,39,0,140,0,55,0,210,0,115,0,177,0,41,0,0,0,104,0,87,0,0,0,78,0,59,0,163,0,68,0,43,0,0,0,81,0,92,0,239,0,39,0,0,0,44,0,41,0,34,0,71,0,18,0,60,0,42,0,38,0,159,0,37,0,185,0,239,0,31,0,218,0,0,0,0,0,163,0,110,0,0,0,0,0,117,0,0,0,33,0,214,0,92,0,248,0,37,0,0,0,244,0,35,0,0,0,53,0,0,0,72,0,0,0,69,0,0,0,179,0,20,0,0,0,15,0,125,0,74,0,125,0,0,0,0,0,0,0,0,0,24,0,100,0,0,0,7,0,0,0,182,0,68,0,118,0,0,0,81,0,0,0,157,0,235,0,155,0,123,0,34,0,231,0,54,0,221,0,233,0,26,0,0,0,51,0,147,0,130,0,154,0,204,0,99,0,100,0,78,0,131,0,153,0,0,0,251,0,44,0,0,0,153,0,167,0,0,0,113,0,0,0,127,0,47,0,67,0,61,0,47,0,0,0,143,0,86,0,111,0,191,0,196,0,125,0,170,0,254,0,156,0,238,0,0,0,237,0,0,0,0,0,102,0,95,0,203,0,0,0,128,0,254,0,136,0,0,0,115,0,83,0,55,0,110,0,144,0,228,0,147,0,51,0,110,0,88,0,0,0,200,0,18,0,72,0,187,0,197,0,0,0,241,0,191,0,102,0,32,0,0,0,51,0,213,0,0,0,103,0,138,0,234,0,63,0,121,0,12,0,159,0,0,0,247,0,34,0,0,0,174,0,155,0,17,0,0,0,0,0,160,0,93,0,0,0,59,0,0,0,19,0,60,0,24,0,0,0,55,0,83,0,1,0,0,0,18,0,173,0,54,0,211,0,0,0,101,0,255,0,26,0,145,0,66,0,186,0,0,0,0,0,74,0,68,0,92,0,76,0,110,0,129,0,129,0,155,0,134,0,115,0,160,0,73,0,245,0,0,0,86,0,214,0,0,0,0,0,241,0,56,0,0,0,112,0,32,0,147,0,224,0,0,0,172,0,0,0,51,0,236,0,112,0,0,0,243,0,132,0,236,0,0,0,76,0,249,0,178,0,0,0,161,0,67,0,214,0,250,0,12,0,176,0,111,0,0,0,181,0,173,0,0,0,185,0,155,0,62,0,89,0,189,0,169,0,156,0,84,0,139,0,238,0,0,0,0,0,181,0,180,0,45,0,133,0,0,0,133,0,234,0,234,0,0,0,212,0,0,0,242,0,229,0,81,0,0,0,96,0,82,0,108,0,185,0,33,0,77,0,4,0,58,0,191,0,19,0,71,0,216,0,0,0,98,0,0,0,147,0,132,0,252,0,248,0,137,0,108,0,0,0,56,0,5,0,23,0,0,0,19,0,0,0,168,0,103,0,115,0,25,0,0,0,118,0,247,0,245,0,28,0,42,0,193,0,54,0,43,0,35,0,69,0,0,0,0,0,0,0,0,0,0,0,63,0,0,0,0,0,10,0,214,0,66,0,206,0,9,0,0,0,0,0,245,0,74,0,170,0,75,0,143,0,0,0,94,0,142,0,0,0,0,0,228,0,0,0,128,0,0,0);
signal scenario_full  : scenario_type := (10,31,173,31,148,31,209,31,253,31,213,31,99,31,34,31,38,31,148,31,217,31,150,31,107,31,121,31,226,31,170,31,110,31,88,31,219,31,56,31,56,30,56,29,153,31,166,31,224,31,224,30,224,29,215,31,215,30,213,31,103,31,103,30,70,31,115,31,143,31,143,30,160,31,232,31,232,30,81,31,114,31,114,30,227,31,227,30,236,31,41,31,42,31,135,31,10,31,8,31,205,31,76,31,209,31,203,31,252,31,218,31,218,30,218,29,218,28,25,31,25,30,7,31,82,31,191,31,191,30,38,31,38,30,38,29,38,28,167,31,244,31,244,30,247,31,88,31,220,31,216,31,47,31,47,30,47,29,122,31,155,31,252,31,151,31,53,31,255,31,172,31,173,31,173,30,190,31,26,31,9,31,110,31,110,30,218,31,218,31,67,31,147,31,238,31,159,31,224,31,224,30,146,31,146,30,220,31,203,31,163,31,163,30,239,31,6,31,47,31,113,31,67,31,156,31,156,30,246,31,251,31,30,31,30,30,253,31,167,31,128,31,128,30,252,31,20,31,20,30,20,29,191,31,122,31,122,30,36,31,36,30,169,31,166,31,251,31,179,31,179,30,164,31,4,31,58,31,21,31,191,31,87,31,110,31,170,31,23,31,23,30,137,31,167,31,167,30,153,31,205,31,41,31,157,31,191,31,13,31,13,30,170,31,170,30,229,31,229,30,204,31,36,31,5,31,182,31,182,30,242,31,80,31,245,31,38,31,38,30,41,31,94,31,111,31,26,31,26,30,26,29,26,28,26,27,161,31,175,31,98,31,226,31,226,30,239,31,239,30,239,29,174,31,189,31,8,31,6,31,6,30,193,31,55,31,206,31,202,31,35,31,140,31,204,31,21,31,93,31,251,31,251,30,119,31,119,30,197,31,197,30,186,31,157,31,53,31,53,30,169,31,169,30,48,31,6,31,6,30,7,31,168,31,168,30,168,29,172,31,192,31,32,31,32,30,32,29,166,31,49,31,185,31,126,31,165,31,13,31,211,31,205,31,190,31,48,31,48,30,48,29,210,31,224,31,224,30,233,31,163,31,2,31,76,31,214,31,72,31,251,31,209,31,125,31,15,31,15,30,15,29,205,31,32,31,235,31,30,31,110,31,191,31,71,31,83,31,253,31,17,31,17,30,212,31,232,31,199,31,218,31,131,31,254,31,254,30,86,31,251,31,177,31,12,31,118,31,50,31,41,31,41,30,41,29,215,31,153,31,153,30,129,31,129,30,88,31,74,31,74,30,74,29,86,31,58,31,249,31,245,31,52,31,52,30,93,31,93,30,130,31,130,30,60,31,60,30,65,31,224,31,194,31,22,31,79,31,79,30,191,31,191,30,125,31,125,30,218,31,167,31,104,31,197,31,88,31,18,31,18,30,12,31,225,31,209,31,122,31,42,31,110,31,156,31,130,31,75,31,85,31,26,31,207,31,47,31,59,31,59,30,53,31,248,31,58,31,58,30,153,31,153,30,153,29,18,31,132,31,132,30,113,31,99,31,228,31,236,31,220,31,117,31,151,31,151,30,49,31,40,31,40,30,40,29,40,28,40,27,79,31,182,31,186,31,186,30,152,31,254,31,109,31,158,31,153,31,153,30,222,31,88,31,137,31,50,31,179,31,46,31,76,31,226,31,57,31,146,31,146,30,97,31,97,30,215,31,215,30,29,31,237,31,237,30,237,29,47,31,59,31,79,31,82,31,209,31,209,30,209,29,95,31,95,30,147,31,147,30,118,31,118,30,118,29,102,31,224,31,168,31,23,31,238,31,4,31,242,31,128,31,18,31,205,31,85,31,85,30,136,31,136,30,115,31,215,31,42,31,16,31,165,31,130,31,113,31,75,31,112,31,198,31,198,30,198,29,84,31,47,31,47,30,47,29,1,31,198,31,181,31,181,30,181,29,66,31,107,31,40,31,218,31,235,31,235,30,117,31,120,31,120,30,171,31,161,31,102,31,250,31,250,30,65,31,239,31,11,31,6,31,6,30,72,31,57,31,103,31,244,31,76,31,90,31,186,31,14,31,118,31,234,31,133,31,201,31,54,31,172,31,172,30,153,31,153,30,134,31,134,30,102,31,171,31,171,30,139,31,96,31,240,31,240,30,159,31,154,31,142,31,196,31,37,31,45,31,105,31,53,31,31,31,31,30,39,31,42,31,119,31,246,31,249,31,2,31,245,31,134,31,184,31,240,31,243,31,243,30,146,31,158,31,73,31,37,31,37,30,241,31,241,30,55,31,55,30,233,31,245,31,188,31,188,30,199,31,199,30,133,31,197,31,197,30,197,29,197,28,210,31,166,31,199,31,199,30,46,31,46,31,21,31,222,31,196,31,196,30,24,31,81,31,5,31,94,31,155,31,104,31,97,31,26,31,125,31,125,30,77,31,207,31,207,30,155,31,57,31,126,31,188,31,131,31,254,31,133,31,177,31,177,30,110,31,193,31,106,31,227,31,227,30,227,29,84,31,12,31,130,31,164,31,96,31,39,31,140,31,55,31,210,31,115,31,177,31,41,31,41,30,104,31,87,31,87,30,78,31,59,31,163,31,68,31,43,31,43,30,81,31,92,31,239,31,39,31,39,30,44,31,41,31,34,31,71,31,18,31,60,31,42,31,38,31,159,31,37,31,185,31,239,31,31,31,218,31,218,30,218,29,163,31,110,31,110,30,110,29,117,31,117,30,33,31,214,31,92,31,248,31,37,31,37,30,244,31,35,31,35,30,53,31,53,30,72,31,72,30,69,31,69,30,179,31,20,31,20,30,15,31,125,31,74,31,125,31,125,30,125,29,125,28,125,27,24,31,100,31,100,30,7,31,7,30,182,31,68,31,118,31,118,30,81,31,81,30,157,31,235,31,155,31,123,31,34,31,231,31,54,31,221,31,233,31,26,31,26,30,51,31,147,31,130,31,154,31,204,31,99,31,100,31,78,31,131,31,153,31,153,30,251,31,44,31,44,30,153,31,167,31,167,30,113,31,113,30,127,31,47,31,67,31,61,31,47,31,47,30,143,31,86,31,111,31,191,31,196,31,125,31,170,31,254,31,156,31,238,31,238,30,237,31,237,30,237,29,102,31,95,31,203,31,203,30,128,31,254,31,136,31,136,30,115,31,83,31,55,31,110,31,144,31,228,31,147,31,51,31,110,31,88,31,88,30,200,31,18,31,72,31,187,31,197,31,197,30,241,31,191,31,102,31,32,31,32,30,51,31,213,31,213,30,103,31,138,31,234,31,63,31,121,31,12,31,159,31,159,30,247,31,34,31,34,30,174,31,155,31,17,31,17,30,17,29,160,31,93,31,93,30,59,31,59,30,19,31,60,31,24,31,24,30,55,31,83,31,1,31,1,30,18,31,173,31,54,31,211,31,211,30,101,31,255,31,26,31,145,31,66,31,186,31,186,30,186,29,74,31,68,31,92,31,76,31,110,31,129,31,129,31,155,31,134,31,115,31,160,31,73,31,245,31,245,30,86,31,214,31,214,30,214,29,241,31,56,31,56,30,112,31,32,31,147,31,224,31,224,30,172,31,172,30,51,31,236,31,112,31,112,30,243,31,132,31,236,31,236,30,76,31,249,31,178,31,178,30,161,31,67,31,214,31,250,31,12,31,176,31,111,31,111,30,181,31,173,31,173,30,185,31,155,31,62,31,89,31,189,31,169,31,156,31,84,31,139,31,238,31,238,30,238,29,181,31,180,31,45,31,133,31,133,30,133,31,234,31,234,31,234,30,212,31,212,30,242,31,229,31,81,31,81,30,96,31,82,31,108,31,185,31,33,31,77,31,4,31,58,31,191,31,19,31,71,31,216,31,216,30,98,31,98,30,147,31,132,31,252,31,248,31,137,31,108,31,108,30,56,31,5,31,23,31,23,30,19,31,19,30,168,31,103,31,115,31,25,31,25,30,118,31,247,31,245,31,28,31,42,31,193,31,54,31,43,31,35,31,69,31,69,30,69,29,69,28,69,27,69,26,63,31,63,30,63,29,10,31,214,31,66,31,206,31,9,31,9,30,9,29,245,31,74,31,170,31,75,31,143,31,143,30,94,31,142,31,142,30,142,29,228,31,228,30,128,31,128,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
