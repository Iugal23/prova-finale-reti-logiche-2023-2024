-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_4 is
end project_tb_4;

architecture project_tb_arch_4 of project_tb_4 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 678;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,101,0,66,0,76,0,249,0,122,0,1,0,232,0,93,0,0,0,153,0,93,0,27,0,158,0,0,0,24,0,207,0,0,0,108,0,110,0,135,0,155,0,0,0,54,0,0,0,159,0,241,0,213,0,172,0,52,0,92,0,218,0,169,0,36,0,60,0,43,0,125,0,0,0,0,0,186,0,81,0,109,0,110,0,159,0,203,0,0,0,158,0,247,0,61,0,16,0,65,0,223,0,159,0,213,0,83,0,19,0,138,0,0,0,0,0,0,0,0,0,208,0,87,0,9,0,16,0,184,0,132,0,0,0,185,0,55,0,225,0,137,0,0,0,180,0,215,0,1,0,55,0,0,0,224,0,0,0,255,0,178,0,208,0,0,0,231,0,0,0,161,0,7,0,243,0,0,0,53,0,209,0,208,0,111,0,0,0,58,0,0,0,62,0,155,0,227,0,110,0,6,0,0,0,90,0,114,0,44,0,51,0,0,0,170,0,199,0,0,0,0,0,208,0,0,0,140,0,242,0,15,0,0,0,44,0,17,0,233,0,235,0,216,0,177,0,10,0,0,0,88,0,172,0,84,0,0,0,0,0,110,0,232,0,199,0,109,0,4,0,150,0,68,0,18,0,0,0,0,0,69,0,41,0,233,0,190,0,8,0,150,0,0,0,0,0,46,0,46,0,0,0,0,0,0,0,212,0,132,0,157,0,11,0,128,0,89,0,15,0,89,0,37,0,0,0,67,0,175,0,202,0,182,0,189,0,36,0,126,0,255,0,115,0,224,0,76,0,125,0,152,0,219,0,202,0,0,0,41,0,142,0,158,0,49,0,137,0,131,0,171,0,157,0,27,0,0,0,178,0,112,0,172,0,68,0,212,0,98,0,80,0,0,0,6,0,0,0,211,0,171,0,111,0,52,0,124,0,122,0,17,0,65,0,109,0,225,0,83,0,140,0,167,0,0,0,0,0,60,0,237,0,62,0,0,0,0,0,140,0,159,0,94,0,88,0,64,0,53,0,138,0,0,0,239,0,194,0,25,0,212,0,147,0,245,0,5,0,230,0,64,0,224,0,205,0,83,0,77,0,67,0,190,0,68,0,0,0,0,0,54,0,29,0,77,0,35,0,43,0,171,0,1,0,25,0,197,0,171,0,11,0,0,0,0,0,171,0,0,0,157,0,104,0,171,0,0,0,44,0,30,0,99,0,133,0,0,0,64,0,211,0,0,0,0,0,22,0,91,0,81,0,31,0,226,0,144,0,137,0,143,0,236,0,6,0,177,0,145,0,159,0,234,0,57,0,173,0,251,0,246,0,108,0,227,0,118,0,10,0,0,0,126,0,85,0,0,0,235,0,115,0,112,0,0,0,185,0,0,0,169,0,142,0,0,0,0,0,12,0,40,0,0,0,106,0,0,0,187,0,189,0,163,0,0,0,226,0,150,0,0,0,26,0,18,0,21,0,167,0,109,0,192,0,111,0,0,0,179,0,195,0,0,0,186,0,33,0,126,0,0,0,8,0,86,0,103,0,0,0,0,0,227,0,106,0,72,0,96,0,218,0,197,0,0,0,131,0,0,0,0,0,198,0,0,0,22,0,237,0,199,0,114,0,153,0,0,0,112,0,48,0,39,0,254,0,204,0,103,0,10,0,0,0,234,0,71,0,0,0,76,0,0,0,130,0,169,0,209,0,238,0,0,0,103,0,226,0,255,0,85,0,0,0,157,0,0,0,0,0,63,0,0,0,46,0,29,0,44,0,29,0,26,0,189,0,0,0,6,0,0,0,26,0,185,0,215,0,122,0,228,0,0,0,190,0,208,0,175,0,191,0,58,0,1,0,242,0,236,0,21,0,11,0,132,0,199,0,18,0,0,0,209,0,191,0,201,0,77,0,33,0,22,0,253,0,224,0,40,0,81,0,0,0,60,0,0,0,243,0,254,0,130,0,64,0,155,0,184,0,0,0,100,0,35,0,219,0,25,0,0,0,154,0,230,0,52,0,55,0,0,0,137,0,54,0,182,0,124,0,240,0,6,0,134,0,0,0,0,0,169,0,190,0,213,0,45,0,91,0,219,0,13,0,225,0,0,0,7,0,149,0,173,0,108,0,0,0,180,0,246,0,127,0,119,0,0,0,173,0,0,0,76,0,0,0,229,0,52,0,185,0,193,0,121,0,154,0,0,0,116,0,173,0,0,0,73,0,201,0,205,0,121,0,198,0,86,0,94,0,160,0,0,0,25,0,0,0,239,0,107,0,107,0,7,0,44,0,107,0,200,0,0,0,148,0,105,0,128,0,113,0,225,0,44,0,252,0,0,0,41,0,0,0,0,0,97,0,91,0,60,0,96,0,225,0,40,0,176,0,29,0,0,0,55,0,225,0,112,0,0,0,15,0,38,0,138,0,49,0,5,0,0,0,130,0,17,0,204,0,64,0,45,0,26,0,194,0,123,0,32,0,42,0,64,0,178,0,247,0,0,0,251,0,17,0,209,0,66,0,149,0,248,0,158,0,0,0,186,0,220,0,0,0,0,0,153,0,225,0,0,0,39,0,27,0,126,0,201,0,127,0,183,0,0,0,62,0,0,0,0,0,160,0,57,0,0,0,0,0,106,0,0,0,0,0,20,0,156,0,107,0,0,0,32,0,160,0,43,0,239,0,48,0,49,0,80,0,0,0,81,0,31,0,0,0,163,0,57,0,20,0,42,0,186,0,56,0,0,0,251,0,130,0,22,0,39,0,0,0,0,0,213,0,253,0,83,0,178,0,208,0,72,0,168,0,173,0,196,0,0,0,177,0,190,0,8,0,242,0,100,0,131,0,184,0,0,0,45,0,173,0,47,0,207,0,93,0,82,0,198,0,0,0,40,0,0,0,0,0,0,0,43,0,128,0,34,0,148,0,139,0,34,0,10,0,0,0,253,0,205,0,217,0,131,0,138,0,0,0,74,0,25,0,183,0,43,0,23,0,124,0,0,0,164,0,79,0,227,0,132,0,206,0,214,0,0,0,157,0,10,0,198,0,161,0,194,0,101,0,117,0,93,0);
signal scenario_full  : scenario_type := (0,0,101,31,66,31,76,31,249,31,122,31,1,31,232,31,93,31,93,30,153,31,93,31,27,31,158,31,158,30,24,31,207,31,207,30,108,31,110,31,135,31,155,31,155,30,54,31,54,30,159,31,241,31,213,31,172,31,52,31,92,31,218,31,169,31,36,31,60,31,43,31,125,31,125,30,125,29,186,31,81,31,109,31,110,31,159,31,203,31,203,30,158,31,247,31,61,31,16,31,65,31,223,31,159,31,213,31,83,31,19,31,138,31,138,30,138,29,138,28,138,27,208,31,87,31,9,31,16,31,184,31,132,31,132,30,185,31,55,31,225,31,137,31,137,30,180,31,215,31,1,31,55,31,55,30,224,31,224,30,255,31,178,31,208,31,208,30,231,31,231,30,161,31,7,31,243,31,243,30,53,31,209,31,208,31,111,31,111,30,58,31,58,30,62,31,155,31,227,31,110,31,6,31,6,30,90,31,114,31,44,31,51,31,51,30,170,31,199,31,199,30,199,29,208,31,208,30,140,31,242,31,15,31,15,30,44,31,17,31,233,31,235,31,216,31,177,31,10,31,10,30,88,31,172,31,84,31,84,30,84,29,110,31,232,31,199,31,109,31,4,31,150,31,68,31,18,31,18,30,18,29,69,31,41,31,233,31,190,31,8,31,150,31,150,30,150,29,46,31,46,31,46,30,46,29,46,28,212,31,132,31,157,31,11,31,128,31,89,31,15,31,89,31,37,31,37,30,67,31,175,31,202,31,182,31,189,31,36,31,126,31,255,31,115,31,224,31,76,31,125,31,152,31,219,31,202,31,202,30,41,31,142,31,158,31,49,31,137,31,131,31,171,31,157,31,27,31,27,30,178,31,112,31,172,31,68,31,212,31,98,31,80,31,80,30,6,31,6,30,211,31,171,31,111,31,52,31,124,31,122,31,17,31,65,31,109,31,225,31,83,31,140,31,167,31,167,30,167,29,60,31,237,31,62,31,62,30,62,29,140,31,159,31,94,31,88,31,64,31,53,31,138,31,138,30,239,31,194,31,25,31,212,31,147,31,245,31,5,31,230,31,64,31,224,31,205,31,83,31,77,31,67,31,190,31,68,31,68,30,68,29,54,31,29,31,77,31,35,31,43,31,171,31,1,31,25,31,197,31,171,31,11,31,11,30,11,29,171,31,171,30,157,31,104,31,171,31,171,30,44,31,30,31,99,31,133,31,133,30,64,31,211,31,211,30,211,29,22,31,91,31,81,31,31,31,226,31,144,31,137,31,143,31,236,31,6,31,177,31,145,31,159,31,234,31,57,31,173,31,251,31,246,31,108,31,227,31,118,31,10,31,10,30,126,31,85,31,85,30,235,31,115,31,112,31,112,30,185,31,185,30,169,31,142,31,142,30,142,29,12,31,40,31,40,30,106,31,106,30,187,31,189,31,163,31,163,30,226,31,150,31,150,30,26,31,18,31,21,31,167,31,109,31,192,31,111,31,111,30,179,31,195,31,195,30,186,31,33,31,126,31,126,30,8,31,86,31,103,31,103,30,103,29,227,31,106,31,72,31,96,31,218,31,197,31,197,30,131,31,131,30,131,29,198,31,198,30,22,31,237,31,199,31,114,31,153,31,153,30,112,31,48,31,39,31,254,31,204,31,103,31,10,31,10,30,234,31,71,31,71,30,76,31,76,30,130,31,169,31,209,31,238,31,238,30,103,31,226,31,255,31,85,31,85,30,157,31,157,30,157,29,63,31,63,30,46,31,29,31,44,31,29,31,26,31,189,31,189,30,6,31,6,30,26,31,185,31,215,31,122,31,228,31,228,30,190,31,208,31,175,31,191,31,58,31,1,31,242,31,236,31,21,31,11,31,132,31,199,31,18,31,18,30,209,31,191,31,201,31,77,31,33,31,22,31,253,31,224,31,40,31,81,31,81,30,60,31,60,30,243,31,254,31,130,31,64,31,155,31,184,31,184,30,100,31,35,31,219,31,25,31,25,30,154,31,230,31,52,31,55,31,55,30,137,31,54,31,182,31,124,31,240,31,6,31,134,31,134,30,134,29,169,31,190,31,213,31,45,31,91,31,219,31,13,31,225,31,225,30,7,31,149,31,173,31,108,31,108,30,180,31,246,31,127,31,119,31,119,30,173,31,173,30,76,31,76,30,229,31,52,31,185,31,193,31,121,31,154,31,154,30,116,31,173,31,173,30,73,31,201,31,205,31,121,31,198,31,86,31,94,31,160,31,160,30,25,31,25,30,239,31,107,31,107,31,7,31,44,31,107,31,200,31,200,30,148,31,105,31,128,31,113,31,225,31,44,31,252,31,252,30,41,31,41,30,41,29,97,31,91,31,60,31,96,31,225,31,40,31,176,31,29,31,29,30,55,31,225,31,112,31,112,30,15,31,38,31,138,31,49,31,5,31,5,30,130,31,17,31,204,31,64,31,45,31,26,31,194,31,123,31,32,31,42,31,64,31,178,31,247,31,247,30,251,31,17,31,209,31,66,31,149,31,248,31,158,31,158,30,186,31,220,31,220,30,220,29,153,31,225,31,225,30,39,31,27,31,126,31,201,31,127,31,183,31,183,30,62,31,62,30,62,29,160,31,57,31,57,30,57,29,106,31,106,30,106,29,20,31,156,31,107,31,107,30,32,31,160,31,43,31,239,31,48,31,49,31,80,31,80,30,81,31,31,31,31,30,163,31,57,31,20,31,42,31,186,31,56,31,56,30,251,31,130,31,22,31,39,31,39,30,39,29,213,31,253,31,83,31,178,31,208,31,72,31,168,31,173,31,196,31,196,30,177,31,190,31,8,31,242,31,100,31,131,31,184,31,184,30,45,31,173,31,47,31,207,31,93,31,82,31,198,31,198,30,40,31,40,30,40,29,40,28,43,31,128,31,34,31,148,31,139,31,34,31,10,31,10,30,253,31,205,31,217,31,131,31,138,31,138,30,74,31,25,31,183,31,43,31,23,31,124,31,124,30,164,31,79,31,227,31,132,31,206,31,214,31,214,30,157,31,10,31,198,31,161,31,194,31,101,31,117,31,93,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
