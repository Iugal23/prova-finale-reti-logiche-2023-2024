-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_91 is
end project_tb_91;

architecture project_tb_arch_91 of project_tb_91 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 786;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (37,0,216,0,0,0,232,0,84,0,0,0,196,0,227,0,30,0,0,0,248,0,253,0,0,0,71,0,202,0,143,0,89,0,3,0,125,0,186,0,48,0,0,0,245,0,229,0,210,0,210,0,185,0,197,0,186,0,68,0,95,0,16,0,41,0,207,0,254,0,64,0,249,0,0,0,182,0,180,0,166,0,51,0,35,0,250,0,0,0,61,0,1,0,120,0,173,0,145,0,0,0,239,0,37,0,180,0,77,0,141,0,16,0,118,0,121,0,93,0,165,0,51,0,98,0,0,0,233,0,113,0,171,0,29,0,87,0,190,0,79,0,15,0,5,0,0,0,242,0,79,0,5,0,245,0,33,0,141,0,61,0,253,0,187,0,178,0,71,0,227,0,127,0,0,0,121,0,149,0,132,0,0,0,211,0,254,0,221,0,234,0,11,0,147,0,78,0,0,0,79,0,154,0,48,0,84,0,73,0,182,0,186,0,0,0,67,0,0,0,0,0,255,0,198,0,229,0,56,0,241,0,69,0,0,0,0,0,93,0,207,0,117,0,83,0,226,0,160,0,138,0,215,0,40,0,79,0,83,0,87,0,84,0,0,0,223,0,0,0,0,0,36,0,206,0,142,0,178,0,222,0,142,0,98,0,159,0,103,0,126,0,152,0,254,0,47,0,100,0,131,0,0,0,238,0,175,0,238,0,84,0,121,0,132,0,114,0,183,0,231,0,244,0,93,0,237,0,199,0,130,0,31,0,52,0,0,0,250,0,191,0,17,0,156,0,0,0,252,0,233,0,0,0,42,0,154,0,37,0,93,0,0,0,69,0,0,0,62,0,0,0,141,0,83,0,46,0,197,0,215,0,127,0,252,0,67,0,208,0,0,0,112,0,144,0,37,0,106,0,150,0,224,0,169,0,0,0,99,0,0,0,235,0,0,0,81,0,223,0,0,0,0,0,175,0,59,0,69,0,146,0,219,0,175,0,160,0,191,0,176,0,0,0,161,0,83,0,0,0,77,0,231,0,0,0,112,0,161,0,145,0,33,0,53,0,30,0,92,0,188,0,181,0,153,0,0,0,0,0,240,0,103,0,0,0,114,0,107,0,244,0,61,0,21,0,17,0,56,0,255,0,122,0,55,0,179,0,0,0,0,0,249,0,251,0,197,0,19,0,162,0,0,0,23,0,108,0,225,0,65,0,0,0,68,0,230,0,101,0,245,0,35,0,0,0,0,0,0,0,240,0,146,0,33,0,175,0,0,0,45,0,0,0,47,0,81,0,76,0,121,0,219,0,83,0,0,0,83,0,0,0,244,0,231,0,0,0,0,0,206,0,19,0,0,0,141,0,111,0,93,0,11,0,181,0,225,0,0,0,121,0,247,0,0,0,220,0,170,0,166,0,80,0,244,0,0,0,73,0,175,0,165,0,193,0,163,0,167,0,77,0,207,0,0,0,0,0,24,0,167,0,182,0,251,0,53,0,54,0,173,0,2,0,61,0,167,0,156,0,0,0,0,0,137,0,134,0,15,0,100,0,0,0,211,0,87,0,215,0,50,0,245,0,219,0,0,0,159,0,234,0,138,0,77,0,216,0,28,0,40,0,44,0,255,0,220,0,202,0,132,0,220,0,172,0,111,0,108,0,0,0,87,0,124,0,235,0,111,0,0,0,91,0,38,0,33,0,74,0,0,0,178,0,10,0,0,0,182,0,12,0,49,0,46,0,34,0,238,0,44,0,246,0,6,0,159,0,55,0,0,0,215,0,60,0,116,0,181,0,68,0,24,0,150,0,0,0,0,0,179,0,14,0,0,0,0,0,171,0,214,0,122,0,253,0,4,0,138,0,0,0,0,0,77,0,0,0,56,0,31,0,128,0,190,0,206,0,153,0,133,0,78,0,6,0,138,0,240,0,110,0,0,0,0,0,0,0,0,0,114,0,0,0,7,0,0,0,229,0,0,0,6,0,0,0,26,0,0,0,110,0,0,0,38,0,0,0,0,0,35,0,0,0,145,0,238,0,164,0,129,0,59,0,108,0,199,0,147,0,16,0,54,0,147,0,85,0,84,0,89,0,67,0,205,0,196,0,116,0,46,0,0,0,31,0,0,0,245,0,55,0,42,0,12,0,0,0,245,0,149,0,113,0,123,0,236,0,107,0,89,0,197,0,0,0,172,0,175,0,0,0,168,0,0,0,0,0,36,0,25,0,127,0,0,0,235,0,212,0,251,0,19,0,195,0,90,0,13,0,0,0,132,0,41,0,0,0,0,0,126,0,179,0,68,0,34,0,233,0,232,0,0,0,242,0,228,0,0,0,21,0,105,0,74,0,0,0,150,0,80,0,154,0,0,0,146,0,130,0,52,0,41,0,63,0,86,0,115,0,186,0,229,0,82,0,143,0,171,0,105,0,22,0,0,0,73,0,49,0,197,0,114,0,0,0,91,0,119,0,138,0,110,0,0,0,96,0,91,0,151,0,3,0,181,0,250,0,126,0,0,0,207,0,116,0,69,0,135,0,127,0,0,0,3,0,9,0,4,0,0,0,166,0,5,0,237,0,174,0,60,0,0,0,81,0,0,0,248,0,205,0,250,0,148,0,93,0,0,0,231,0,35,0,160,0,26,0,136,0,0,0,86,0,193,0,0,0,227,0,0,0,208,0,62,0,162,0,131,0,253,0,230,0,0,0,115,0,143,0,222,0,28,0,0,0,12,0,254,0,178,0,0,0,8,0,196,0,128,0,116,0,14,0,248,0,241,0,8,0,190,0,68,0,0,0,228,0,0,0,0,0,233,0,135,0,0,0,160,0,7,0,0,0,3,0,0,0,0,0,0,0,0,0,11,0,155,0,116,0,111,0,244,0,147,0,0,0,93,0,141,0,198,0,0,0,55,0,0,0,180,0,107,0,231,0,155,0,20,0,7,0,40,0,0,0,120,0,0,0,16,0,64,0,0,0,15,0,0,0,41,0,6,0,87,0,0,0,125,0,25,0,210,0,79,0,180,0,37,0,209,0,177,0,240,0,131,0,0,0,144,0,218,0,0,0,0,0,33,0,222,0,105,0,175,0,0,0,208,0,0,0,98,0,108,0,103,0,218,0,40,0,105,0,137,0,142,0,195,0,231,0,112,0,212,0,200,0,221,0,157,0,225,0,66,0,206,0,181,0,7,0,17,0,198,0,33,0,130,0,242,0,231,0,179,0,182,0,213,0,137,0,240,0,27,0,0,0,247,0,0,0,152,0,0,0,152,0,184,0,204,0,17,0,152,0,249,0,69,0,18,0,219,0,213,0,60,0,80,0,122,0,63,0,194,0,220,0,7,0,244,0,156,0,199,0,84,0,101,0,92,0,0,0,123,0,10,0,140,0,26,0,23,0,8,0,217,0,132,0,147,0,0,0,17,0,212,0,0,0,32,0,100,0,160,0,174,0,63,0,116,0,41,0,93,0,239,0,197,0,11,0,141,0,158,0,25,0,110,0,95,0,184,0,115,0,152,0,248,0,44,0,36,0,205,0,0,0,115,0,223,0);
signal scenario_full  : scenario_type := (37,31,216,31,216,30,232,31,84,31,84,30,196,31,227,31,30,31,30,30,248,31,253,31,253,30,71,31,202,31,143,31,89,31,3,31,125,31,186,31,48,31,48,30,245,31,229,31,210,31,210,31,185,31,197,31,186,31,68,31,95,31,16,31,41,31,207,31,254,31,64,31,249,31,249,30,182,31,180,31,166,31,51,31,35,31,250,31,250,30,61,31,1,31,120,31,173,31,145,31,145,30,239,31,37,31,180,31,77,31,141,31,16,31,118,31,121,31,93,31,165,31,51,31,98,31,98,30,233,31,113,31,171,31,29,31,87,31,190,31,79,31,15,31,5,31,5,30,242,31,79,31,5,31,245,31,33,31,141,31,61,31,253,31,187,31,178,31,71,31,227,31,127,31,127,30,121,31,149,31,132,31,132,30,211,31,254,31,221,31,234,31,11,31,147,31,78,31,78,30,79,31,154,31,48,31,84,31,73,31,182,31,186,31,186,30,67,31,67,30,67,29,255,31,198,31,229,31,56,31,241,31,69,31,69,30,69,29,93,31,207,31,117,31,83,31,226,31,160,31,138,31,215,31,40,31,79,31,83,31,87,31,84,31,84,30,223,31,223,30,223,29,36,31,206,31,142,31,178,31,222,31,142,31,98,31,159,31,103,31,126,31,152,31,254,31,47,31,100,31,131,31,131,30,238,31,175,31,238,31,84,31,121,31,132,31,114,31,183,31,231,31,244,31,93,31,237,31,199,31,130,31,31,31,52,31,52,30,250,31,191,31,17,31,156,31,156,30,252,31,233,31,233,30,42,31,154,31,37,31,93,31,93,30,69,31,69,30,62,31,62,30,141,31,83,31,46,31,197,31,215,31,127,31,252,31,67,31,208,31,208,30,112,31,144,31,37,31,106,31,150,31,224,31,169,31,169,30,99,31,99,30,235,31,235,30,81,31,223,31,223,30,223,29,175,31,59,31,69,31,146,31,219,31,175,31,160,31,191,31,176,31,176,30,161,31,83,31,83,30,77,31,231,31,231,30,112,31,161,31,145,31,33,31,53,31,30,31,92,31,188,31,181,31,153,31,153,30,153,29,240,31,103,31,103,30,114,31,107,31,244,31,61,31,21,31,17,31,56,31,255,31,122,31,55,31,179,31,179,30,179,29,249,31,251,31,197,31,19,31,162,31,162,30,23,31,108,31,225,31,65,31,65,30,68,31,230,31,101,31,245,31,35,31,35,30,35,29,35,28,240,31,146,31,33,31,175,31,175,30,45,31,45,30,47,31,81,31,76,31,121,31,219,31,83,31,83,30,83,31,83,30,244,31,231,31,231,30,231,29,206,31,19,31,19,30,141,31,111,31,93,31,11,31,181,31,225,31,225,30,121,31,247,31,247,30,220,31,170,31,166,31,80,31,244,31,244,30,73,31,175,31,165,31,193,31,163,31,167,31,77,31,207,31,207,30,207,29,24,31,167,31,182,31,251,31,53,31,54,31,173,31,2,31,61,31,167,31,156,31,156,30,156,29,137,31,134,31,15,31,100,31,100,30,211,31,87,31,215,31,50,31,245,31,219,31,219,30,159,31,234,31,138,31,77,31,216,31,28,31,40,31,44,31,255,31,220,31,202,31,132,31,220,31,172,31,111,31,108,31,108,30,87,31,124,31,235,31,111,31,111,30,91,31,38,31,33,31,74,31,74,30,178,31,10,31,10,30,182,31,12,31,49,31,46,31,34,31,238,31,44,31,246,31,6,31,159,31,55,31,55,30,215,31,60,31,116,31,181,31,68,31,24,31,150,31,150,30,150,29,179,31,14,31,14,30,14,29,171,31,214,31,122,31,253,31,4,31,138,31,138,30,138,29,77,31,77,30,56,31,31,31,128,31,190,31,206,31,153,31,133,31,78,31,6,31,138,31,240,31,110,31,110,30,110,29,110,28,110,27,114,31,114,30,7,31,7,30,229,31,229,30,6,31,6,30,26,31,26,30,110,31,110,30,38,31,38,30,38,29,35,31,35,30,145,31,238,31,164,31,129,31,59,31,108,31,199,31,147,31,16,31,54,31,147,31,85,31,84,31,89,31,67,31,205,31,196,31,116,31,46,31,46,30,31,31,31,30,245,31,55,31,42,31,12,31,12,30,245,31,149,31,113,31,123,31,236,31,107,31,89,31,197,31,197,30,172,31,175,31,175,30,168,31,168,30,168,29,36,31,25,31,127,31,127,30,235,31,212,31,251,31,19,31,195,31,90,31,13,31,13,30,132,31,41,31,41,30,41,29,126,31,179,31,68,31,34,31,233,31,232,31,232,30,242,31,228,31,228,30,21,31,105,31,74,31,74,30,150,31,80,31,154,31,154,30,146,31,130,31,52,31,41,31,63,31,86,31,115,31,186,31,229,31,82,31,143,31,171,31,105,31,22,31,22,30,73,31,49,31,197,31,114,31,114,30,91,31,119,31,138,31,110,31,110,30,96,31,91,31,151,31,3,31,181,31,250,31,126,31,126,30,207,31,116,31,69,31,135,31,127,31,127,30,3,31,9,31,4,31,4,30,166,31,5,31,237,31,174,31,60,31,60,30,81,31,81,30,248,31,205,31,250,31,148,31,93,31,93,30,231,31,35,31,160,31,26,31,136,31,136,30,86,31,193,31,193,30,227,31,227,30,208,31,62,31,162,31,131,31,253,31,230,31,230,30,115,31,143,31,222,31,28,31,28,30,12,31,254,31,178,31,178,30,8,31,196,31,128,31,116,31,14,31,248,31,241,31,8,31,190,31,68,31,68,30,228,31,228,30,228,29,233,31,135,31,135,30,160,31,7,31,7,30,3,31,3,30,3,29,3,28,3,27,11,31,155,31,116,31,111,31,244,31,147,31,147,30,93,31,141,31,198,31,198,30,55,31,55,30,180,31,107,31,231,31,155,31,20,31,7,31,40,31,40,30,120,31,120,30,16,31,64,31,64,30,15,31,15,30,41,31,6,31,87,31,87,30,125,31,25,31,210,31,79,31,180,31,37,31,209,31,177,31,240,31,131,31,131,30,144,31,218,31,218,30,218,29,33,31,222,31,105,31,175,31,175,30,208,31,208,30,98,31,108,31,103,31,218,31,40,31,105,31,137,31,142,31,195,31,231,31,112,31,212,31,200,31,221,31,157,31,225,31,66,31,206,31,181,31,7,31,17,31,198,31,33,31,130,31,242,31,231,31,179,31,182,31,213,31,137,31,240,31,27,31,27,30,247,31,247,30,152,31,152,30,152,31,184,31,204,31,17,31,152,31,249,31,69,31,18,31,219,31,213,31,60,31,80,31,122,31,63,31,194,31,220,31,7,31,244,31,156,31,199,31,84,31,101,31,92,31,92,30,123,31,10,31,140,31,26,31,23,31,8,31,217,31,132,31,147,31,147,30,17,31,212,31,212,30,32,31,100,31,160,31,174,31,63,31,116,31,41,31,93,31,239,31,197,31,11,31,141,31,158,31,25,31,110,31,95,31,184,31,115,31,152,31,248,31,44,31,36,31,205,31,205,30,115,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
