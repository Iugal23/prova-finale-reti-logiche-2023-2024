-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 893;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,38,0,53,0,223,0,169,0,163,0,8,0,167,0,76,0,0,0,188,0,30,0,45,0,123,0,13,0,134,0,23,0,60,0,0,0,233,0,115,0,158,0,23,0,142,0,91,0,0,0,18,0,9,0,0,0,239,0,106,0,0,0,171,0,191,0,0,0,203,0,85,0,142,0,0,0,95,0,197,0,72,0,50,0,235,0,0,0,20,0,159,0,99,0,19,0,56,0,67,0,246,0,86,0,122,0,91,0,226,0,125,0,113,0,22,0,14,0,0,0,0,0,255,0,88,0,52,0,177,0,98,0,134,0,194,0,52,0,42,0,135,0,228,0,0,0,34,0,34,0,92,0,195,0,0,0,136,0,206,0,92,0,115,0,170,0,82,0,141,0,62,0,221,0,0,0,122,0,12,0,148,0,60,0,32,0,12,0,71,0,79,0,42,0,245,0,153,0,206,0,0,0,4,0,0,0,125,0,41,0,0,0,109,0,113,0,153,0,0,0,114,0,154,0,209,0,0,0,4,0,0,0,209,0,85,0,210,0,156,0,157,0,249,0,50,0,54,0,71,0,84,0,225,0,238,0,0,0,216,0,0,0,126,0,122,0,0,0,0,0,41,0,96,0,201,0,0,0,149,0,32,0,124,0,161,0,8,0,75,0,158,0,58,0,0,0,11,0,47,0,25,0,223,0,138,0,143,0,208,0,0,0,141,0,237,0,0,0,201,0,223,0,0,0,160,0,35,0,0,0,99,0,0,0,125,0,177,0,170,0,0,0,205,0,43,0,1,0,0,0,207,0,223,0,88,0,157,0,165,0,0,0,0,0,226,0,168,0,184,0,106,0,0,0,0,0,69,0,65,0,76,0,182,0,137,0,47,0,0,0,81,0,166,0,222,0,172,0,14,0,132,0,28,0,223,0,166,0,172,0,0,0,87,0,23,0,0,0,255,0,170,0,54,0,206,0,167,0,41,0,0,0,28,0,87,0,70,0,127,0,182,0,24,0,0,0,204,0,147,0,16,0,39,0,0,0,161,0,1,0,251,0,122,0,0,0,52,0,171,0,130,0,28,0,88,0,167,0,2,0,195,0,241,0,97,0,195,0,204,0,0,0,203,0,23,0,4,0,89,0,42,0,202,0,63,0,153,0,144,0,216,0,27,0,238,0,171,0,73,0,168,0,180,0,238,0,225,0,43,0,127,0,173,0,214,0,57,0,123,0,198,0,213,0,0,0,245,0,167,0,39,0,235,0,32,0,20,0,0,0,0,0,93,0,221,0,168,0,227,0,106,0,0,0,20,0,13,0,140,0,199,0,141,0,238,0,68,0,0,0,18,0,184,0,224,0,186,0,141,0,2,0,24,0,241,0,0,0,202,0,0,0,178,0,103,0,133,0,212,0,175,0,186,0,0,0,45,0,127,0,153,0,212,0,0,0,93,0,102,0,68,0,0,0,0,0,203,0,0,0,193,0,77,0,167,0,0,0,44,0,0,0,15,0,129,0,51,0,0,0,9,0,0,0,232,0,0,0,117,0,227,0,252,0,216,0,255,0,115,0,180,0,105,0,56,0,0,0,43,0,0,0,52,0,152,0,192,0,0,0,131,0,27,0,247,0,0,0,0,0,76,0,170,0,36,0,46,0,78,0,0,0,96,0,233,0,221,0,6,0,0,0,29,0,95,0,88,0,130,0,63,0,28,0,109,0,239,0,215,0,148,0,0,0,47,0,34,0,163,0,100,0,93,0,49,0,201,0,212,0,146,0,111,0,0,0,216,0,0,0,16,0,174,0,0,0,0,0,219,0,184,0,35,0,91,0,251,0,88,0,231,0,0,0,186,0,37,0,82,0,58,0,129,0,228,0,89,0,100,0,196,0,158,0,59,0,92,0,49,0,0,0,239,0,247,0,132,0,168,0,63,0,129,0,0,0,24,0,20,0,39,0,0,0,125,0,0,0,0,0,213,0,89,0,95,0,0,0,176,0,0,0,212,0,0,0,201,0,168,0,51,0,141,0,139,0,176,0,0,0,0,0,19,0,0,0,0,0,0,0,0,0,81,0,121,0,61,0,146,0,0,0,95,0,90,0,219,0,72,0,50,0,110,0,242,0,223,0,27,0,0,0,0,0,123,0,125,0,53,0,90,0,157,0,206,0,230,0,146,0,38,0,243,0,174,0,31,0,0,0,232,0,50,0,208,0,133,0,57,0,75,0,0,0,0,0,17,0,221,0,83,0,67,0,24,0,165,0,135,0,64,0,0,0,163,0,0,0,202,0,44,0,151,0,165,0,209,0,58,0,58,0,2,0,169,0,0,0,0,0,0,0,235,0,203,0,87,0,88,0,107,0,159,0,108,0,76,0,76,0,236,0,218,0,147,0,213,0,170,0,43,0,75,0,218,0,152,0,123,0,0,0,90,0,46,0,142,0,133,0,57,0,66,0,0,0,111,0,251,0,108,0,73,0,0,0,0,0,228,0,222,0,198,0,0,0,35,0,31,0,181,0,107,0,8,0,215,0,0,0,110,0,180,0,168,0,183,0,142,0,1,0,0,0,137,0,50,0,104,0,123,0,131,0,182,0,145,0,69,0,157,0,0,0,132,0,161,0,196,0,119,0,0,0,120,0,95,0,0,0,52,0,89,0,0,0,0,0,254,0,200,0,48,0,188,0,93,0,108,0,0,0,231,0,0,0,88,0,223,0,159,0,208,0,70,0,160,0,229,0,219,0,98,0,153,0,0,0,184,0,175,0,251,0,15,0,3,0,157,0,213,0,252,0,229,0,222,0,218,0,0,0,157,0,0,0,115,0,210,0,176,0,0,0,247,0,0,0,59,0,131,0,73,0,77,0,29,0,207,0,0,0,22,0,181,0,135,0,251,0,19,0,183,0,8,0,222,0,153,0,198,0,231,0,0,0,12,0,177,0,0,0,101,0,3,0,146,0,0,0,248,0,27,0,0,0,187,0,63,0,0,0,206,0,33,0,151,0,234,0,235,0,181,0,181,0,186,0,0,0,0,0,0,0,95,0,98,0,209,0,153,0,0,0,2,0,231,0,58,0,50,0,148,0,0,0,226,0,230,0,149,0,220,0,245,0,167,0,177,0,0,0,232,0,171,0,0,0,33,0,219,0,239,0,196,0,158,0,213,0,234,0,117,0,0,0,39,0,169,0,58,0,0,0,84,0,216,0,110,0,92,0,63,0,222,0,100,0,0,0,0,0,4,0,155,0,210,0,197,0,214,0,157,0,82,0,1,0,102,0,0,0,148,0,89,0,0,0,120,0,206,0,109,0,40,0,124,0,0,0,65,0,0,0,84,0,8,0,111,0,0,0,0,0,125,0,0,0,222,0,65,0,192,0,182,0,212,0,0,0,41,0,81,0,73,0,224,0,82,0,65,0,0,0,137,0,0,0,169,0,136,0,216,0,254,0,7,0,21,0,160,0,46,0,16,0,154,0,230,0,200,0,83,0,0,0,0,0,170,0,0,0,14,0,0,0,151,0,133,0,140,0,93,0,196,0,181,0,23,0,16,0,10,0,0,0,216,0,210,0,68,0,177,0,113,0,76,0,216,0,0,0,110,0,60,0,137,0,0,0,163,0,0,0,0,0,158,0,119,0,53,0,0,0,110,0,112,0,153,0,0,0,65,0,71,0,244,0,52,0,178,0,26,0,0,0,32,0,160,0,209,0,32,0,29,0,114,0,182,0,185,0,33,0,120,0,0,0,77,0,126,0,112,0,0,0,204,0,226,0,223,0,134,0,0,0,15,0,145,0,0,0,11,0,90,0,0,0,103,0,0,0,105,0,44,0,24,0,0,0,0,0,237,0,69,0,238,0,49,0,68,0,206,0,0,0,35,0,255,0,158,0,92,0,249,0,72,0,0,0,66,0,206,0,236,0,54,0,47,0,155,0,10,0,24,0,14,0,254,0,0,0,170,0,20,0,246,0,57,0,116,0,0,0,0,0,3,0,59,0,73,0,222,0,0,0,40,0,57,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,38,31,53,31,223,31,169,31,163,31,8,31,167,31,76,31,76,30,188,31,30,31,45,31,123,31,13,31,134,31,23,31,60,31,60,30,233,31,115,31,158,31,23,31,142,31,91,31,91,30,18,31,9,31,9,30,239,31,106,31,106,30,171,31,191,31,191,30,203,31,85,31,142,31,142,30,95,31,197,31,72,31,50,31,235,31,235,30,20,31,159,31,99,31,19,31,56,31,67,31,246,31,86,31,122,31,91,31,226,31,125,31,113,31,22,31,14,31,14,30,14,29,255,31,88,31,52,31,177,31,98,31,134,31,194,31,52,31,42,31,135,31,228,31,228,30,34,31,34,31,92,31,195,31,195,30,136,31,206,31,92,31,115,31,170,31,82,31,141,31,62,31,221,31,221,30,122,31,12,31,148,31,60,31,32,31,12,31,71,31,79,31,42,31,245,31,153,31,206,31,206,30,4,31,4,30,125,31,41,31,41,30,109,31,113,31,153,31,153,30,114,31,154,31,209,31,209,30,4,31,4,30,209,31,85,31,210,31,156,31,157,31,249,31,50,31,54,31,71,31,84,31,225,31,238,31,238,30,216,31,216,30,126,31,122,31,122,30,122,29,41,31,96,31,201,31,201,30,149,31,32,31,124,31,161,31,8,31,75,31,158,31,58,31,58,30,11,31,47,31,25,31,223,31,138,31,143,31,208,31,208,30,141,31,237,31,237,30,201,31,223,31,223,30,160,31,35,31,35,30,99,31,99,30,125,31,177,31,170,31,170,30,205,31,43,31,1,31,1,30,207,31,223,31,88,31,157,31,165,31,165,30,165,29,226,31,168,31,184,31,106,31,106,30,106,29,69,31,65,31,76,31,182,31,137,31,47,31,47,30,81,31,166,31,222,31,172,31,14,31,132,31,28,31,223,31,166,31,172,31,172,30,87,31,23,31,23,30,255,31,170,31,54,31,206,31,167,31,41,31,41,30,28,31,87,31,70,31,127,31,182,31,24,31,24,30,204,31,147,31,16,31,39,31,39,30,161,31,1,31,251,31,122,31,122,30,52,31,171,31,130,31,28,31,88,31,167,31,2,31,195,31,241,31,97,31,195,31,204,31,204,30,203,31,23,31,4,31,89,31,42,31,202,31,63,31,153,31,144,31,216,31,27,31,238,31,171,31,73,31,168,31,180,31,238,31,225,31,43,31,127,31,173,31,214,31,57,31,123,31,198,31,213,31,213,30,245,31,167,31,39,31,235,31,32,31,20,31,20,30,20,29,93,31,221,31,168,31,227,31,106,31,106,30,20,31,13,31,140,31,199,31,141,31,238,31,68,31,68,30,18,31,184,31,224,31,186,31,141,31,2,31,24,31,241,31,241,30,202,31,202,30,178,31,103,31,133,31,212,31,175,31,186,31,186,30,45,31,127,31,153,31,212,31,212,30,93,31,102,31,68,31,68,30,68,29,203,31,203,30,193,31,77,31,167,31,167,30,44,31,44,30,15,31,129,31,51,31,51,30,9,31,9,30,232,31,232,30,117,31,227,31,252,31,216,31,255,31,115,31,180,31,105,31,56,31,56,30,43,31,43,30,52,31,152,31,192,31,192,30,131,31,27,31,247,31,247,30,247,29,76,31,170,31,36,31,46,31,78,31,78,30,96,31,233,31,221,31,6,31,6,30,29,31,95,31,88,31,130,31,63,31,28,31,109,31,239,31,215,31,148,31,148,30,47,31,34,31,163,31,100,31,93,31,49,31,201,31,212,31,146,31,111,31,111,30,216,31,216,30,16,31,174,31,174,30,174,29,219,31,184,31,35,31,91,31,251,31,88,31,231,31,231,30,186,31,37,31,82,31,58,31,129,31,228,31,89,31,100,31,196,31,158,31,59,31,92,31,49,31,49,30,239,31,247,31,132,31,168,31,63,31,129,31,129,30,24,31,20,31,39,31,39,30,125,31,125,30,125,29,213,31,89,31,95,31,95,30,176,31,176,30,212,31,212,30,201,31,168,31,51,31,141,31,139,31,176,31,176,30,176,29,19,31,19,30,19,29,19,28,19,27,81,31,121,31,61,31,146,31,146,30,95,31,90,31,219,31,72,31,50,31,110,31,242,31,223,31,27,31,27,30,27,29,123,31,125,31,53,31,90,31,157,31,206,31,230,31,146,31,38,31,243,31,174,31,31,31,31,30,232,31,50,31,208,31,133,31,57,31,75,31,75,30,75,29,17,31,221,31,83,31,67,31,24,31,165,31,135,31,64,31,64,30,163,31,163,30,202,31,44,31,151,31,165,31,209,31,58,31,58,31,2,31,169,31,169,30,169,29,169,28,235,31,203,31,87,31,88,31,107,31,159,31,108,31,76,31,76,31,236,31,218,31,147,31,213,31,170,31,43,31,75,31,218,31,152,31,123,31,123,30,90,31,46,31,142,31,133,31,57,31,66,31,66,30,111,31,251,31,108,31,73,31,73,30,73,29,228,31,222,31,198,31,198,30,35,31,31,31,181,31,107,31,8,31,215,31,215,30,110,31,180,31,168,31,183,31,142,31,1,31,1,30,137,31,50,31,104,31,123,31,131,31,182,31,145,31,69,31,157,31,157,30,132,31,161,31,196,31,119,31,119,30,120,31,95,31,95,30,52,31,89,31,89,30,89,29,254,31,200,31,48,31,188,31,93,31,108,31,108,30,231,31,231,30,88,31,223,31,159,31,208,31,70,31,160,31,229,31,219,31,98,31,153,31,153,30,184,31,175,31,251,31,15,31,3,31,157,31,213,31,252,31,229,31,222,31,218,31,218,30,157,31,157,30,115,31,210,31,176,31,176,30,247,31,247,30,59,31,131,31,73,31,77,31,29,31,207,31,207,30,22,31,181,31,135,31,251,31,19,31,183,31,8,31,222,31,153,31,198,31,231,31,231,30,12,31,177,31,177,30,101,31,3,31,146,31,146,30,248,31,27,31,27,30,187,31,63,31,63,30,206,31,33,31,151,31,234,31,235,31,181,31,181,31,186,31,186,30,186,29,186,28,95,31,98,31,209,31,153,31,153,30,2,31,231,31,58,31,50,31,148,31,148,30,226,31,230,31,149,31,220,31,245,31,167,31,177,31,177,30,232,31,171,31,171,30,33,31,219,31,239,31,196,31,158,31,213,31,234,31,117,31,117,30,39,31,169,31,58,31,58,30,84,31,216,31,110,31,92,31,63,31,222,31,100,31,100,30,100,29,4,31,155,31,210,31,197,31,214,31,157,31,82,31,1,31,102,31,102,30,148,31,89,31,89,30,120,31,206,31,109,31,40,31,124,31,124,30,65,31,65,30,84,31,8,31,111,31,111,30,111,29,125,31,125,30,222,31,65,31,192,31,182,31,212,31,212,30,41,31,81,31,73,31,224,31,82,31,65,31,65,30,137,31,137,30,169,31,136,31,216,31,254,31,7,31,21,31,160,31,46,31,16,31,154,31,230,31,200,31,83,31,83,30,83,29,170,31,170,30,14,31,14,30,151,31,133,31,140,31,93,31,196,31,181,31,23,31,16,31,10,31,10,30,216,31,210,31,68,31,177,31,113,31,76,31,216,31,216,30,110,31,60,31,137,31,137,30,163,31,163,30,163,29,158,31,119,31,53,31,53,30,110,31,112,31,153,31,153,30,65,31,71,31,244,31,52,31,178,31,26,31,26,30,32,31,160,31,209,31,32,31,29,31,114,31,182,31,185,31,33,31,120,31,120,30,77,31,126,31,112,31,112,30,204,31,226,31,223,31,134,31,134,30,15,31,145,31,145,30,11,31,90,31,90,30,103,31,103,30,105,31,44,31,24,31,24,30,24,29,237,31,69,31,238,31,49,31,68,31,206,31,206,30,35,31,255,31,158,31,92,31,249,31,72,31,72,30,66,31,206,31,236,31,54,31,47,31,155,31,10,31,24,31,14,31,254,31,254,30,170,31,20,31,246,31,57,31,116,31,116,30,116,29,3,31,59,31,73,31,222,31,222,30,40,31,57,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
