-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (199,0,40,0,251,0,180,0,216,0,90,0,36,0,123,0,215,0,237,0,0,0,110,0,225,0,115,0,0,0,17,0,5,0,161,0,178,0,104,0,0,0,195,0,0,0,77,0,112,0,75,0,101,0,54,0,0,0,224,0,0,0,140,0,199,0,0,0,0,0,149,0,184,0,155,0,174,0,127,0,0,0,226,0,74,0,0,0,209,0,68,0,94,0,17,0,94,0,155,0,41,0,115,0,99,0,109,0,0,0,56,0,236,0,0,0,31,0,255,0,17,0,0,0,229,0,14,0,56,0,249,0,237,0,110,0,38,0,195,0,238,0,218,0,0,0,8,0,61,0,73,0,184,0,4,0,0,0,76,0,55,0,72,0,245,0,88,0,50,0,0,0,0,0,6,0,220,0,150,0,136,0,192,0,251,0,0,0,0,0,0,0,0,0,89,0,0,0,140,0,129,0,223,0,246,0,0,0,124,0,133,0,0,0,163,0,115,0,90,0,245,0,233,0,95,0,202,0,63,0,23,0,177,0,171,0,0,0,170,0,3,0,37,0,144,0,23,0,77,0,56,0,56,0,0,0,155,0,161,0,44,0,194,0,89,0,0,0,143,0,221,0,42,0,170,0,246,0,76,0,231,0,205,0,124,0,126,0,117,0,178,0,127,0,144,0,106,0,146,0,114,0,105,0,0,0,143,0,30,0,109,0,121,0,0,0,207,0,97,0,159,0,45,0,136,0,187,0,38,0,216,0,49,0,21,0,113,0,35,0,28,0,58,0,0,0,0,0,10,0,157,0,248,0,146,0,78,0,120,0,54,0,0,0,0,0,169,0,182,0,160,0,185,0,58,0,88,0,143,0,3,0,255,0,78,0,38,0,17,0,0,0,176,0,0,0,132,0,75,0,0,0,27,0,55,0,237,0,192,0,67,0,0,0,53,0,67,0,116,0,114,0,217,0,183,0,148,0,0,0,37,0,58,0,202,0,34,0,163,0,16,0,246,0,0,0,14,0,0,0,0,0,0,0,252,0,78,0,43,0,247,0,0,0,0,0,189,0,255,0,169,0,114,0,245,0,89,0,0,0,117,0,0,0,160,0,187,0,4,0,88,0,239,0,149,0,148,0,226,0,116,0,63,0,25,0,22,0,199,0,6,0,209,0,248,0,0,0,219,0,43,0,198,0,31,0,0,0,252,0,0,0,184,0,241,0,182,0,27,0,136,0,0,0,236,0,169,0,84,0,217,0,0,0,178,0,99,0,0,0,189,0,0,0,208,0,105,0,182,0,142,0,0,0,106,0,0,0,137,0,194,0,0,0,241,0,67,0,128,0,123,0,115,0,29,0,219,0,225,0,215,0,0,0,248,0,82,0,0,0,61,0,84,0,96,0,49,0,29,0,82,0,240,0,224,0,137,0,78,0,216,0,50,0,255,0,46,0,0,0,107,0,75,0,0,0,157,0,133,0,0,0,10,0,202,0,107,0,99,0,123,0,18,0,103,0,55,0,79,0,29,0,223,0,197,0,234,0,210,0,0,0,100,0,117,0,20,0,59,0,3,0,116,0,165,0,129,0,138,0,244,0,0,0,66,0,72,0,246,0,56,0,208,0,0,0,75,0,8,0,39,0,20,0,178,0,160,0,182,0,247,0,228,0,131,0,247,0,94,0,249,0,73,0,99,0,225,0,0,0,217,0,111,0,182,0,34,0,30,0,245,0,185,0,11,0,19,0,18,0,190,0,79,0,23,0,0,0,5,0,150,0,0,0,160,0,0,0,0,0,20,0,198,0,111,0,0,0,208,0,159,0,161,0,240,0,0,0,0,0,41,0,0,0,0,0,132,0,14,0,182,0,235,0,84,0,80,0,243,0,68,0,76,0,0,0,0,0,0,0,47,0,43,0,189,0,105,0,153,0,172,0,0,0,11,0,165,0,151,0,211,0,0,0,97,0,198,0,162,0,26,0,22,0,61,0,7,0,37,0,1,0,179,0,0,0,0,0,94,0,153,0,158,0,0,0,241,0,0,0,0,0,129,0,0,0,0,0,192,0,217,0,0,0,119,0,133,0,15,0,137,0,18,0,11,0,207,0,188,0,70,0,10,0,0,0,24,0,15,0,2,0,178,0,175,0,86,0,17,0,197,0,70,0,143,0,179,0,232,0,113,0,192,0,0,0,121,0,0,0,251,0,186,0,36,0,209,0,32,0,26,0,87,0,182,0,202,0,248,0,49,0,0,0,113,0,78,0,130,0,96,0,74,0,0,0,104,0,13,0,0,0,0,0,5,0,12,0,0,0,247,0,197,0,208,0,118,0,253,0,101,0,0,0,175,0,131,0,199,0,148,0,12,0,139,0,0,0,84,0,209,0,194,0,0,0,96,0,0,0,185,0,0,0,161,0,98,0,46,0,217,0,195,0,164,0,0,0,58,0,0,0,0,0,161,0,241,0,0,0,225,0,88,0,221,0,189,0,133,0,210,0,0,0,231,0,120,0,0,0,0,0,104,0,103,0,194,0,43,0,17,0,152,0,22,0,149,0,45,0,58,0,85,0,129,0,6,0,0,0,0,0,21,0,25,0,247,0,69,0,44,0,161,0,238,0,206,0,100,0,13,0,194,0,53,0,8,0,70,0,0,0,0,0,104,0,41,0,155,0,44,0,53,0,93,0,78,0,252,0,200,0,204,0,15,0,94,0,24,0,87,0,3,0,45,0,74,0,94,0,96,0,74,0,90,0,0,0,187,0,208,0,204,0,0,0,106,0,217,0,0,0,232,0,111,0,163,0,251,0,112,0,244,0,149,0,18,0,185,0,24,0,196,0,210,0,0,0,194,0,213,0,133,0,135,0,0,0,0,0,0,0,12,0,0,0,68,0,246,0,50,0,230,0,203,0,115,0,124,0,98,0,0,0,46,0,74,0,0,0,87,0,0,0,69,0,0,0,250,0,169,0,252,0,0,0,97,0,220,0,0,0,0,0,0,0,14,0,66,0,58,0,123,0,190,0,111,0,15,0,10,0,79,0,142,0,203,0,137,0,132,0,126,0,93,0,30,0,129,0,0,0,107,0,166,0,100,0,28,0,215,0,152,0,181,0,212,0,91,0,29,0,76,0,14,0,139,0,103,0,44,0,0,0,138,0,50,0,148,0,0,0,28,0,73,0,131,0,246,0,13,0,0,0,64,0,80,0,0,0,168,0,88,0,77,0,159,0,120,0,16,0,166,0,171,0,196,0,30,0,90,0,89,0,89,0,254,0,0,0,230,0,143,0,2,0,36,0,0,0,0,0,0,0,0,0,0,0,220,0,130,0,149,0,133,0,125,0,0,0,0,0,67,0,186,0,217,0,219,0,152,0,183,0,14,0,9,0,106,0,63,0,182,0,78,0,0,0,0,0,0,0,97,0,194,0,11,0,2,0,105,0,115,0,96,0,254,0,115,0,132,0,140,0,13,0,96,0,48,0,54,0,21,0,226,0,253,0,1,0,232,0,53,0,92,0,47,0,20,0,74,0,245,0,0,0,54,0,247,0,0,0,108,0,254,0,89,0,0,0,237,0,98,0,96,0,42,0,228,0,0,0,65,0,239,0,192,0,0,0,141,0,158,0,28,0,19,0,0,0,0,0,0,0,151,0,26,0,148,0,194,0,97,0,97,0,32,0,173,0,30,0,0,0,17,0,162,0,213,0,66,0,0,0,105,0,0,0,131,0,0,0,85,0,31,0,99,0,1,0,169,0,214,0,233,0,182,0,0,0,172,0,0,0,234,0,254,0,132,0,49,0,225,0,216,0,147,0,27,0,0,0,172,0,120,0,54,0,33,0,0,0,215,0,32,0,235,0,179,0,216,0,205,0,24,0,74,0,55,0,212,0,21,0,208,0,141,0,173,0,93,0,0,0,162,0,40,0,245,0,133,0,188,0,191,0,22,0,173,0,236,0,80,0,20,0,82,0,0,0,0,0,225,0,156,0,0,0,56,0,68,0,0,0,0,0,116,0,74,0,42,0,0,0,124,0,0,0,79,0,47,0,241,0,238,0,146,0,119,0,189,0,0,0,78,0,205,0,65,0,142,0,73,0,11,0,211,0,16,0,0,0,0,0,175,0,236,0,0,0,0,0,71,0,0,0,118,0,68,0,123,0,117,0,234,0,0,0,91,0,255,0,169,0,105,0,162,0,251,0,65,0,15,0,153,0,0,0,165,0,0,0,211,0,75,0,136,0,0,0,0,0,0,0,91,0,196,0,93,0,55,0,236,0,89,0,79,0,0,0,54,0,189,0,8,0,156,0,11,0,59,0,71,0,16,0,49,0,145,0,77,0,224,0,187,0,152,0,250,0,134,0,39,0,153,0,177,0,49,0,253,0,0,0,212,0,138,0,43,0);
signal scenario_full  : scenario_type := (199,31,40,31,251,31,180,31,216,31,90,31,36,31,123,31,215,31,237,31,237,30,110,31,225,31,115,31,115,30,17,31,5,31,161,31,178,31,104,31,104,30,195,31,195,30,77,31,112,31,75,31,101,31,54,31,54,30,224,31,224,30,140,31,199,31,199,30,199,29,149,31,184,31,155,31,174,31,127,31,127,30,226,31,74,31,74,30,209,31,68,31,94,31,17,31,94,31,155,31,41,31,115,31,99,31,109,31,109,30,56,31,236,31,236,30,31,31,255,31,17,31,17,30,229,31,14,31,56,31,249,31,237,31,110,31,38,31,195,31,238,31,218,31,218,30,8,31,61,31,73,31,184,31,4,31,4,30,76,31,55,31,72,31,245,31,88,31,50,31,50,30,50,29,6,31,220,31,150,31,136,31,192,31,251,31,251,30,251,29,251,28,251,27,89,31,89,30,140,31,129,31,223,31,246,31,246,30,124,31,133,31,133,30,163,31,115,31,90,31,245,31,233,31,95,31,202,31,63,31,23,31,177,31,171,31,171,30,170,31,3,31,37,31,144,31,23,31,77,31,56,31,56,31,56,30,155,31,161,31,44,31,194,31,89,31,89,30,143,31,221,31,42,31,170,31,246,31,76,31,231,31,205,31,124,31,126,31,117,31,178,31,127,31,144,31,106,31,146,31,114,31,105,31,105,30,143,31,30,31,109,31,121,31,121,30,207,31,97,31,159,31,45,31,136,31,187,31,38,31,216,31,49,31,21,31,113,31,35,31,28,31,58,31,58,30,58,29,10,31,157,31,248,31,146,31,78,31,120,31,54,31,54,30,54,29,169,31,182,31,160,31,185,31,58,31,88,31,143,31,3,31,255,31,78,31,38,31,17,31,17,30,176,31,176,30,132,31,75,31,75,30,27,31,55,31,237,31,192,31,67,31,67,30,53,31,67,31,116,31,114,31,217,31,183,31,148,31,148,30,37,31,58,31,202,31,34,31,163,31,16,31,246,31,246,30,14,31,14,30,14,29,14,28,252,31,78,31,43,31,247,31,247,30,247,29,189,31,255,31,169,31,114,31,245,31,89,31,89,30,117,31,117,30,160,31,187,31,4,31,88,31,239,31,149,31,148,31,226,31,116,31,63,31,25,31,22,31,199,31,6,31,209,31,248,31,248,30,219,31,43,31,198,31,31,31,31,30,252,31,252,30,184,31,241,31,182,31,27,31,136,31,136,30,236,31,169,31,84,31,217,31,217,30,178,31,99,31,99,30,189,31,189,30,208,31,105,31,182,31,142,31,142,30,106,31,106,30,137,31,194,31,194,30,241,31,67,31,128,31,123,31,115,31,29,31,219,31,225,31,215,31,215,30,248,31,82,31,82,30,61,31,84,31,96,31,49,31,29,31,82,31,240,31,224,31,137,31,78,31,216,31,50,31,255,31,46,31,46,30,107,31,75,31,75,30,157,31,133,31,133,30,10,31,202,31,107,31,99,31,123,31,18,31,103,31,55,31,79,31,29,31,223,31,197,31,234,31,210,31,210,30,100,31,117,31,20,31,59,31,3,31,116,31,165,31,129,31,138,31,244,31,244,30,66,31,72,31,246,31,56,31,208,31,208,30,75,31,8,31,39,31,20,31,178,31,160,31,182,31,247,31,228,31,131,31,247,31,94,31,249,31,73,31,99,31,225,31,225,30,217,31,111,31,182,31,34,31,30,31,245,31,185,31,11,31,19,31,18,31,190,31,79,31,23,31,23,30,5,31,150,31,150,30,160,31,160,30,160,29,20,31,198,31,111,31,111,30,208,31,159,31,161,31,240,31,240,30,240,29,41,31,41,30,41,29,132,31,14,31,182,31,235,31,84,31,80,31,243,31,68,31,76,31,76,30,76,29,76,28,47,31,43,31,189,31,105,31,153,31,172,31,172,30,11,31,165,31,151,31,211,31,211,30,97,31,198,31,162,31,26,31,22,31,61,31,7,31,37,31,1,31,179,31,179,30,179,29,94,31,153,31,158,31,158,30,241,31,241,30,241,29,129,31,129,30,129,29,192,31,217,31,217,30,119,31,133,31,15,31,137,31,18,31,11,31,207,31,188,31,70,31,10,31,10,30,24,31,15,31,2,31,178,31,175,31,86,31,17,31,197,31,70,31,143,31,179,31,232,31,113,31,192,31,192,30,121,31,121,30,251,31,186,31,36,31,209,31,32,31,26,31,87,31,182,31,202,31,248,31,49,31,49,30,113,31,78,31,130,31,96,31,74,31,74,30,104,31,13,31,13,30,13,29,5,31,12,31,12,30,247,31,197,31,208,31,118,31,253,31,101,31,101,30,175,31,131,31,199,31,148,31,12,31,139,31,139,30,84,31,209,31,194,31,194,30,96,31,96,30,185,31,185,30,161,31,98,31,46,31,217,31,195,31,164,31,164,30,58,31,58,30,58,29,161,31,241,31,241,30,225,31,88,31,221,31,189,31,133,31,210,31,210,30,231,31,120,31,120,30,120,29,104,31,103,31,194,31,43,31,17,31,152,31,22,31,149,31,45,31,58,31,85,31,129,31,6,31,6,30,6,29,21,31,25,31,247,31,69,31,44,31,161,31,238,31,206,31,100,31,13,31,194,31,53,31,8,31,70,31,70,30,70,29,104,31,41,31,155,31,44,31,53,31,93,31,78,31,252,31,200,31,204,31,15,31,94,31,24,31,87,31,3,31,45,31,74,31,94,31,96,31,74,31,90,31,90,30,187,31,208,31,204,31,204,30,106,31,217,31,217,30,232,31,111,31,163,31,251,31,112,31,244,31,149,31,18,31,185,31,24,31,196,31,210,31,210,30,194,31,213,31,133,31,135,31,135,30,135,29,135,28,12,31,12,30,68,31,246,31,50,31,230,31,203,31,115,31,124,31,98,31,98,30,46,31,74,31,74,30,87,31,87,30,69,31,69,30,250,31,169,31,252,31,252,30,97,31,220,31,220,30,220,29,220,28,14,31,66,31,58,31,123,31,190,31,111,31,15,31,10,31,79,31,142,31,203,31,137,31,132,31,126,31,93,31,30,31,129,31,129,30,107,31,166,31,100,31,28,31,215,31,152,31,181,31,212,31,91,31,29,31,76,31,14,31,139,31,103,31,44,31,44,30,138,31,50,31,148,31,148,30,28,31,73,31,131,31,246,31,13,31,13,30,64,31,80,31,80,30,168,31,88,31,77,31,159,31,120,31,16,31,166,31,171,31,196,31,30,31,90,31,89,31,89,31,254,31,254,30,230,31,143,31,2,31,36,31,36,30,36,29,36,28,36,27,36,26,220,31,130,31,149,31,133,31,125,31,125,30,125,29,67,31,186,31,217,31,219,31,152,31,183,31,14,31,9,31,106,31,63,31,182,31,78,31,78,30,78,29,78,28,97,31,194,31,11,31,2,31,105,31,115,31,96,31,254,31,115,31,132,31,140,31,13,31,96,31,48,31,54,31,21,31,226,31,253,31,1,31,232,31,53,31,92,31,47,31,20,31,74,31,245,31,245,30,54,31,247,31,247,30,108,31,254,31,89,31,89,30,237,31,98,31,96,31,42,31,228,31,228,30,65,31,239,31,192,31,192,30,141,31,158,31,28,31,19,31,19,30,19,29,19,28,151,31,26,31,148,31,194,31,97,31,97,31,32,31,173,31,30,31,30,30,17,31,162,31,213,31,66,31,66,30,105,31,105,30,131,31,131,30,85,31,31,31,99,31,1,31,169,31,214,31,233,31,182,31,182,30,172,31,172,30,234,31,254,31,132,31,49,31,225,31,216,31,147,31,27,31,27,30,172,31,120,31,54,31,33,31,33,30,215,31,32,31,235,31,179,31,216,31,205,31,24,31,74,31,55,31,212,31,21,31,208,31,141,31,173,31,93,31,93,30,162,31,40,31,245,31,133,31,188,31,191,31,22,31,173,31,236,31,80,31,20,31,82,31,82,30,82,29,225,31,156,31,156,30,56,31,68,31,68,30,68,29,116,31,74,31,42,31,42,30,124,31,124,30,79,31,47,31,241,31,238,31,146,31,119,31,189,31,189,30,78,31,205,31,65,31,142,31,73,31,11,31,211,31,16,31,16,30,16,29,175,31,236,31,236,30,236,29,71,31,71,30,118,31,68,31,123,31,117,31,234,31,234,30,91,31,255,31,169,31,105,31,162,31,251,31,65,31,15,31,153,31,153,30,165,31,165,30,211,31,75,31,136,31,136,30,136,29,136,28,91,31,196,31,93,31,55,31,236,31,89,31,79,31,79,30,54,31,189,31,8,31,156,31,11,31,59,31,71,31,16,31,49,31,145,31,77,31,224,31,187,31,152,31,250,31,134,31,39,31,153,31,177,31,49,31,253,31,253,30,212,31,138,31,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
