-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 693;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (115,0,0,0,58,0,230,0,26,0,123,0,25,0,192,0,71,0,198,0,230,0,135,0,0,0,0,0,183,0,192,0,0,0,169,0,39,0,0,0,242,0,223,0,0,0,122,0,155,0,111,0,240,0,0,0,51,0,121,0,248,0,198,0,0,0,125,0,138,0,94,0,51,0,223,0,0,0,0,0,16,0,0,0,119,0,0,0,0,0,93,0,152,0,230,0,107,0,99,0,65,0,191,0,10,0,161,0,43,0,113,0,195,0,212,0,0,0,0,0,0,0,195,0,21,0,118,0,118,0,203,0,0,0,139,0,212,0,174,0,14,0,241,0,56,0,110,0,65,0,0,0,0,0,80,0,147,0,66,0,20,0,51,0,135,0,183,0,0,0,217,0,100,0,175,0,73,0,133,0,0,0,187,0,0,0,93,0,28,0,0,0,87,0,112,0,181,0,242,0,231,0,254,0,31,0,240,0,0,0,221,0,0,0,0,0,115,0,78,0,104,0,112,0,10,0,93,0,225,0,183,0,102,0,0,0,0,0,89,0,225,0,0,0,0,0,134,0,110,0,85,0,0,0,192,0,34,0,65,0,165,0,190,0,0,0,0,0,0,0,161,0,0,0,137,0,174,0,73,0,0,0,0,0,220,0,75,0,105,0,0,0,246,0,84,0,169,0,113,0,152,0,111,0,0,0,153,0,35,0,48,0,220,0,115,0,234,0,204,0,4,0,29,0,167,0,47,0,0,0,195,0,28,0,123,0,114,0,233,0,0,0,172,0,218,0,216,0,0,0,0,0,12,0,222,0,0,0,0,0,34,0,250,0,50,0,100,0,80,0,40,0,215,0,0,0,49,0,164,0,253,0,130,0,183,0,148,0,78,0,50,0,213,0,92,0,19,0,12,0,0,0,135,0,220,0,32,0,191,0,221,0,189,0,187,0,233,0,164,0,101,0,70,0,0,0,0,0,59,0,74,0,121,0,124,0,253,0,0,0,0,0,107,0,111,0,146,0,229,0,58,0,57,0,185,0,90,0,0,0,143,0,0,0,196,0,0,0,45,0,0,0,0,0,43,0,50,0,0,0,166,0,127,0,160,0,0,0,207,0,239,0,45,0,183,0,148,0,108,0,53,0,131,0,0,0,165,0,10,0,28,0,23,0,143,0,127,0,134,0,0,0,14,0,155,0,46,0,181,0,21,0,0,0,47,0,187,0,0,0,172,0,236,0,81,0,53,0,0,0,86,0,41,0,0,0,0,0,67,0,16,0,3,0,0,0,30,0,50,0,123,0,0,0,250,0,8,0,45,0,0,0,160,0,42,0,29,0,0,0,55,0,44,0,0,0,15,0,54,0,108,0,194,0,0,0,229,0,26,0,0,0,215,0,220,0,179,0,78,0,173,0,138,0,241,0,236,0,153,0,168,0,66,0,204,0,176,0,70,0,199,0,254,0,241,0,175,0,155,0,0,0,0,0,0,0,37,0,218,0,120,0,115,0,235,0,168,0,8,0,0,0,149,0,0,0,247,0,183,0,93,0,88,0,165,0,228,0,214,0,221,0,150,0,122,0,21,0,186,0,55,0,255,0,209,0,25,0,194,0,0,0,29,0,55,0,145,0,116,0,120,0,52,0,102,0,0,0,28,0,215,0,196,0,0,0,0,0,1,0,168,0,0,0,215,0,107,0,76,0,185,0,200,0,149,0,0,0,132,0,0,0,175,0,90,0,0,0,212,0,0,0,0,0,89,0,122,0,144,0,68,0,0,0,163,0,129,0,225,0,0,0,0,0,61,0,122,0,0,0,3,0,143,0,82,0,13,0,12,0,225,0,39,0,152,0,0,0,79,0,254,0,10,0,185,0,0,0,46,0,75,0,0,0,0,0,0,0,132,0,0,0,118,0,0,0,160,0,193,0,0,0,0,0,0,0,88,0,42,0,0,0,33,0,0,0,149,0,0,0,123,0,77,0,54,0,0,0,124,0,43,0,0,0,230,0,132,0,200,0,182,0,129,0,0,0,112,0,243,0,0,0,0,0,216,0,0,0,130,0,60,0,136,0,198,0,179,0,150,0,193,0,87,0,12,0,158,0,96,0,77,0,0,0,0,0,232,0,197,0,173,0,0,0,6,0,78,0,238,0,174,0,0,0,170,0,227,0,127,0,172,0,20,0,0,0,212,0,66,0,117,0,48,0,219,0,216,0,158,0,26,0,0,0,29,0,94,0,169,0,32,0,137,0,40,0,0,0,0,0,13,0,251,0,245,0,254,0,0,0,88,0,0,0,75,0,136,0,0,0,0,0,25,0,213,0,7,0,137,0,252,0,32,0,95,0,4,0,175,0,142,0,153,0,0,0,58,0,0,0,0,0,153,0,0,0,6,0,87,0,142,0,1,0,66,0,114,0,0,0,0,0,239,0,85,0,74,0,0,0,222,0,0,0,177,0,14,0,214,0,0,0,0,0,139,0,138,0,169,0,177,0,203,0,156,0,172,0,145,0,100,0,253,0,0,0,150,0,24,0,176,0,16,0,95,0,5,0,116,0,128,0,115,0,227,0,0,0,0,0,8,0,136,0,29,0,0,0,0,0,0,0,60,0,0,0,102,0,0,0,149,0,52,0,249,0,83,0,213,0,232,0,133,0,58,0,75,0,0,0,111,0,0,0,209,0,242,0,217,0,136,0,253,0,120,0,130,0,0,0,100,0,166,0,121,0,118,0,60,0,189,0,2,0,63,0,97,0,0,0,22,0,77,0,239,0,30,0,132,0,137,0,23,0,106,0,195,0,0,0,154,0,233,0,127,0,240,0,208,0,0,0,212,0,184,0,0,0,174,0,58,0,63,0,126,0,165,0,53,0,123,0,118,0,0,0,0,0,0,0,144,0,0,0,157,0,3,0,142,0,214,0,163,0,154,0,214,0,0,0,105,0,121,0,147,0,218,0,0,0,108,0,0,0,102,0,234,0,71,0,41,0,0,0,36,0,60,0,158,0,191,0,221,0,202,0,171,0,194,0,189,0,0,0,188,0,111,0,135,0,0,0,20,0,41,0,234,0,220,0,6,0,90,0,96,0,163,0,21,0,89,0,0,0,139,0,0,0,195,0,77,0,101,0,40,0);
signal scenario_full  : scenario_type := (115,31,115,30,58,31,230,31,26,31,123,31,25,31,192,31,71,31,198,31,230,31,135,31,135,30,135,29,183,31,192,31,192,30,169,31,39,31,39,30,242,31,223,31,223,30,122,31,155,31,111,31,240,31,240,30,51,31,121,31,248,31,198,31,198,30,125,31,138,31,94,31,51,31,223,31,223,30,223,29,16,31,16,30,119,31,119,30,119,29,93,31,152,31,230,31,107,31,99,31,65,31,191,31,10,31,161,31,43,31,113,31,195,31,212,31,212,30,212,29,212,28,195,31,21,31,118,31,118,31,203,31,203,30,139,31,212,31,174,31,14,31,241,31,56,31,110,31,65,31,65,30,65,29,80,31,147,31,66,31,20,31,51,31,135,31,183,31,183,30,217,31,100,31,175,31,73,31,133,31,133,30,187,31,187,30,93,31,28,31,28,30,87,31,112,31,181,31,242,31,231,31,254,31,31,31,240,31,240,30,221,31,221,30,221,29,115,31,78,31,104,31,112,31,10,31,93,31,225,31,183,31,102,31,102,30,102,29,89,31,225,31,225,30,225,29,134,31,110,31,85,31,85,30,192,31,34,31,65,31,165,31,190,31,190,30,190,29,190,28,161,31,161,30,137,31,174,31,73,31,73,30,73,29,220,31,75,31,105,31,105,30,246,31,84,31,169,31,113,31,152,31,111,31,111,30,153,31,35,31,48,31,220,31,115,31,234,31,204,31,4,31,29,31,167,31,47,31,47,30,195,31,28,31,123,31,114,31,233,31,233,30,172,31,218,31,216,31,216,30,216,29,12,31,222,31,222,30,222,29,34,31,250,31,50,31,100,31,80,31,40,31,215,31,215,30,49,31,164,31,253,31,130,31,183,31,148,31,78,31,50,31,213,31,92,31,19,31,12,31,12,30,135,31,220,31,32,31,191,31,221,31,189,31,187,31,233,31,164,31,101,31,70,31,70,30,70,29,59,31,74,31,121,31,124,31,253,31,253,30,253,29,107,31,111,31,146,31,229,31,58,31,57,31,185,31,90,31,90,30,143,31,143,30,196,31,196,30,45,31,45,30,45,29,43,31,50,31,50,30,166,31,127,31,160,31,160,30,207,31,239,31,45,31,183,31,148,31,108,31,53,31,131,31,131,30,165,31,10,31,28,31,23,31,143,31,127,31,134,31,134,30,14,31,155,31,46,31,181,31,21,31,21,30,47,31,187,31,187,30,172,31,236,31,81,31,53,31,53,30,86,31,41,31,41,30,41,29,67,31,16,31,3,31,3,30,30,31,50,31,123,31,123,30,250,31,8,31,45,31,45,30,160,31,42,31,29,31,29,30,55,31,44,31,44,30,15,31,54,31,108,31,194,31,194,30,229,31,26,31,26,30,215,31,220,31,179,31,78,31,173,31,138,31,241,31,236,31,153,31,168,31,66,31,204,31,176,31,70,31,199,31,254,31,241,31,175,31,155,31,155,30,155,29,155,28,37,31,218,31,120,31,115,31,235,31,168,31,8,31,8,30,149,31,149,30,247,31,183,31,93,31,88,31,165,31,228,31,214,31,221,31,150,31,122,31,21,31,186,31,55,31,255,31,209,31,25,31,194,31,194,30,29,31,55,31,145,31,116,31,120,31,52,31,102,31,102,30,28,31,215,31,196,31,196,30,196,29,1,31,168,31,168,30,215,31,107,31,76,31,185,31,200,31,149,31,149,30,132,31,132,30,175,31,90,31,90,30,212,31,212,30,212,29,89,31,122,31,144,31,68,31,68,30,163,31,129,31,225,31,225,30,225,29,61,31,122,31,122,30,3,31,143,31,82,31,13,31,12,31,225,31,39,31,152,31,152,30,79,31,254,31,10,31,185,31,185,30,46,31,75,31,75,30,75,29,75,28,132,31,132,30,118,31,118,30,160,31,193,31,193,30,193,29,193,28,88,31,42,31,42,30,33,31,33,30,149,31,149,30,123,31,77,31,54,31,54,30,124,31,43,31,43,30,230,31,132,31,200,31,182,31,129,31,129,30,112,31,243,31,243,30,243,29,216,31,216,30,130,31,60,31,136,31,198,31,179,31,150,31,193,31,87,31,12,31,158,31,96,31,77,31,77,30,77,29,232,31,197,31,173,31,173,30,6,31,78,31,238,31,174,31,174,30,170,31,227,31,127,31,172,31,20,31,20,30,212,31,66,31,117,31,48,31,219,31,216,31,158,31,26,31,26,30,29,31,94,31,169,31,32,31,137,31,40,31,40,30,40,29,13,31,251,31,245,31,254,31,254,30,88,31,88,30,75,31,136,31,136,30,136,29,25,31,213,31,7,31,137,31,252,31,32,31,95,31,4,31,175,31,142,31,153,31,153,30,58,31,58,30,58,29,153,31,153,30,6,31,87,31,142,31,1,31,66,31,114,31,114,30,114,29,239,31,85,31,74,31,74,30,222,31,222,30,177,31,14,31,214,31,214,30,214,29,139,31,138,31,169,31,177,31,203,31,156,31,172,31,145,31,100,31,253,31,253,30,150,31,24,31,176,31,16,31,95,31,5,31,116,31,128,31,115,31,227,31,227,30,227,29,8,31,136,31,29,31,29,30,29,29,29,28,60,31,60,30,102,31,102,30,149,31,52,31,249,31,83,31,213,31,232,31,133,31,58,31,75,31,75,30,111,31,111,30,209,31,242,31,217,31,136,31,253,31,120,31,130,31,130,30,100,31,166,31,121,31,118,31,60,31,189,31,2,31,63,31,97,31,97,30,22,31,77,31,239,31,30,31,132,31,137,31,23,31,106,31,195,31,195,30,154,31,233,31,127,31,240,31,208,31,208,30,212,31,184,31,184,30,174,31,58,31,63,31,126,31,165,31,53,31,123,31,118,31,118,30,118,29,118,28,144,31,144,30,157,31,3,31,142,31,214,31,163,31,154,31,214,31,214,30,105,31,121,31,147,31,218,31,218,30,108,31,108,30,102,31,234,31,71,31,41,31,41,30,36,31,60,31,158,31,191,31,221,31,202,31,171,31,194,31,189,31,189,30,188,31,111,31,135,31,135,30,20,31,41,31,234,31,220,31,6,31,90,31,96,31,163,31,21,31,89,31,89,30,139,31,139,30,195,31,77,31,101,31,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
