-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 836;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,168,0,9,0,56,0,214,0,255,0,237,0,204,0,190,0,170,0,235,0,0,0,115,0,96,0,53,0,252,0,74,0,45,0,160,0,12,0,208,0,237,0,178,0,212,0,0,0,220,0,123,0,35,0,0,0,83,0,243,0,250,0,158,0,135,0,145,0,183,0,68,0,178,0,92,0,85,0,0,0,240,0,89,0,8,0,189,0,102,0,0,0,0,0,161,0,56,0,220,0,172,0,0,0,0,0,226,0,206,0,0,0,27,0,13,0,69,0,101,0,39,0,0,0,215,0,29,0,0,0,80,0,64,0,50,0,0,0,116,0,11,0,121,0,63,0,81,0,246,0,139,0,226,0,228,0,0,0,0,0,191,0,213,0,0,0,0,0,53,0,24,0,197,0,19,0,145,0,249,0,247,0,246,0,186,0,140,0,201,0,21,0,141,0,6,0,59,0,223,0,185,0,42,0,216,0,0,0,194,0,86,0,38,0,77,0,183,0,34,0,223,0,105,0,82,0,163,0,0,0,2,0,205,0,232,0,61,0,30,0,19,0,125,0,171,0,13,0,202,0,0,0,148,0,187,0,56,0,252,0,0,0,173,0,142,0,169,0,182,0,126,0,66,0,105,0,252,0,191,0,238,0,41,0,178,0,0,0,220,0,0,0,167,0,0,0,63,0,0,0,0,0,40,0,32,0,147,0,115,0,7,0,62,0,161,0,156,0,0,0,145,0,0,0,219,0,0,0,201,0,187,0,187,0,169,0,0,0,197,0,163,0,0,0,12,0,0,0,0,0,54,0,86,0,242,0,116,0,45,0,38,0,42,0,94,0,0,0,158,0,27,0,59,0,201,0,0,0,155,0,23,0,60,0,203,0,10,0,86,0,75,0,185,0,87,0,239,0,79,0,123,0,198,0,161,0,117,0,147,0,0,0,0,0,252,0,0,0,198,0,72,0,0,0,82,0,139,0,16,0,51,0,11,0,254,0,164,0,205,0,142,0,0,0,21,0,0,0,180,0,203,0,0,0,131,0,203,0,80,0,0,0,196,0,11,0,189,0,23,0,120,0,231,0,119,0,195,0,59,0,0,0,158,0,15,0,0,0,240,0,0,0,140,0,161,0,149,0,0,0,178,0,0,0,0,0,0,0,179,0,236,0,18,0,0,0,55,0,133,0,251,0,215,0,54,0,189,0,6,0,0,0,101,0,130,0,0,0,0,0,75,0,50,0,58,0,59,0,14,0,0,0,62,0,224,0,206,0,192,0,207,0,239,0,0,0,41,0,0,0,0,0,117,0,103,0,54,0,112,0,190,0,107,0,98,0,0,0,140,0,42,0,255,0,0,0,180,0,64,0,126,0,15,0,0,0,200,0,0,0,19,0,5,0,133,0,64,0,255,0,1,0,46,0,51,0,95,0,231,0,132,0,92,0,18,0,0,0,0,0,149,0,14,0,158,0,252,0,129,0,221,0,0,0,146,0,25,0,0,0,98,0,0,0,37,0,37,0,63,0,91,0,160,0,0,0,200,0,17,0,244,0,68,0,120,0,0,0,112,0,126,0,210,0,178,0,5,0,96,0,0,0,0,0,112,0,112,0,186,0,229,0,0,0,23,0,1,0,21,0,27,0,180,0,181,0,23,0,95,0,205,0,242,0,0,0,132,0,189,0,69,0,210,0,54,0,40,0,14,0,31,0,54,0,108,0,13,0,0,0,67,0,138,0,135,0,232,0,198,0,77,0,235,0,0,0,54,0,232,0,0,0,189,0,247,0,89,0,16,0,32,0,14,0,242,0,0,0,119,0,140,0,186,0,153,0,94,0,183,0,147,0,54,0,92,0,105,0,183,0,0,0,212,0,111,0,0,0,0,0,66,0,62,0,131,0,231,0,121,0,50,0,0,0,242,0,177,0,3,0,206,0,223,0,246,0,224,0,0,0,241,0,147,0,236,0,123,0,39,0,0,0,76,0,114,0,242,0,21,0,162,0,171,0,40,0,113,0,53,0,222,0,47,0,40,0,17,0,121,0,238,0,94,0,36,0,134,0,54,0,86,0,106,0,0,0,68,0,0,0,119,0,250,0,47,0,215,0,0,0,227,0,139,0,156,0,92,0,0,0,72,0,172,0,202,0,0,0,104,0,116,0,0,0,143,0,60,0,0,0,0,0,0,0,169,0,133,0,225,0,14,0,2,0,32,0,0,0,186,0,206,0,0,0,12,0,0,0,223,0,168,0,231,0,85,0,56,0,116,0,105,0,54,0,0,0,190,0,97,0,168,0,37,0,215,0,144,0,200,0,251,0,0,0,82,0,232,0,249,0,38,0,32,0,0,0,0,0,144,0,81,0,223,0,0,0,165,0,115,0,176,0,87,0,0,0,65,0,67,0,53,0,193,0,12,0,175,0,23,0,205,0,101,0,50,0,0,0,188,0,236,0,189,0,103,0,0,0,0,0,199,0,200,0,177,0,133,0,200,0,61,0,154,0,158,0,0,0,102,0,242,0,57,0,0,0,119,0,98,0,2,0,232,0,0,0,57,0,51,0,84,0,130,0,192,0,0,0,212,0,175,0,0,0,1,0,98,0,50,0,243,0,156,0,223,0,125,0,180,0,190,0,36,0,76,0,0,0,14,0,252,0,174,0,65,0,101,0,61,0,87,0,231,0,165,0,0,0,105,0,10,0,0,0,252,0,0,0,137,0,55,0,135,0,0,0,219,0,0,0,233,0,144,0,182,0,6,0,0,0,246,0,48,0,41,0,71,0,0,0,0,0,57,0,27,0,241,0,19,0,0,0,36,0,216,0,214,0,132,0,197,0,0,0,95,0,212,0,146,0,232,0,212,0,163,0,231,0,91,0,2,0,207,0,164,0,0,0,0,0,0,0,29,0,144,0,32,0,237,0,95,0,0,0,131,0,88,0,203,0,207,0,229,0,171,0,207,0,168,0,0,0,14,0,153,0,190,0,189,0,204,0,13,0,98,0,62,0,49,0,0,0,131,0,235,0,195,0,120,0,102,0,171,0,0,0,66,0,48,0,234,0,39,0,13,0,163,0,96,0,202,0,202,0,21,0,153,0,0,0,16,0,13,0,181,0,0,0,0,0,173,0,23,0,34,0,142,0,143,0,53,0,0,0,157,0,44,0,225,0,241,0,102,0,108,0,68,0,0,0,1,0,0,0,205,0,0,0,0,0,3,0,138,0,19,0,165,0,45,0,162,0,100,0,230,0,51,0,77,0,110,0,0,0,0,0,163,0,87,0,68,0,224,0,0,0,196,0,13,0,94,0,194,0,29,0,43,0,170,0,0,0,233,0,132,0,203,0,97,0,58,0,231,0,53,0,245,0,120,0,0,0,0,0,172,0,73,0,67,0,95,0,153,0,224,0,186,0,111,0,81,0,0,0,203,0,20,0,189,0,169,0,187,0,139,0,138,0,35,0,70,0,218,0,0,0,0,0,110,0,167,0,189,0,160,0,22,0,29,0,89,0,65,0,190,0,44,0,0,0,0,0,146,0,230,0,0,0,41,0,0,0,242,0,149,0,201,0,218,0,63,0,0,0,47,0,228,0,206,0,118,0,0,0,0,0,39,0,151,0,18,0,5,0,224,0,252,0,184,0,140,0,0,0,160,0,69,0,108,0,0,0,194,0,216,0,76,0,47,0,0,0,74,0,104,0,131,0,121,0,198,0,0,0,0,0,83,0,60,0,219,0,22,0,0,0,181,0,168,0,49,0,30,0,0,0,65,0,102,0);
signal scenario_full  : scenario_type := (250,31,168,31,9,31,56,31,214,31,255,31,237,31,204,31,190,31,170,31,235,31,235,30,115,31,96,31,53,31,252,31,74,31,45,31,160,31,12,31,208,31,237,31,178,31,212,31,212,30,220,31,123,31,35,31,35,30,83,31,243,31,250,31,158,31,135,31,145,31,183,31,68,31,178,31,92,31,85,31,85,30,240,31,89,31,8,31,189,31,102,31,102,30,102,29,161,31,56,31,220,31,172,31,172,30,172,29,226,31,206,31,206,30,27,31,13,31,69,31,101,31,39,31,39,30,215,31,29,31,29,30,80,31,64,31,50,31,50,30,116,31,11,31,121,31,63,31,81,31,246,31,139,31,226,31,228,31,228,30,228,29,191,31,213,31,213,30,213,29,53,31,24,31,197,31,19,31,145,31,249,31,247,31,246,31,186,31,140,31,201,31,21,31,141,31,6,31,59,31,223,31,185,31,42,31,216,31,216,30,194,31,86,31,38,31,77,31,183,31,34,31,223,31,105,31,82,31,163,31,163,30,2,31,205,31,232,31,61,31,30,31,19,31,125,31,171,31,13,31,202,31,202,30,148,31,187,31,56,31,252,31,252,30,173,31,142,31,169,31,182,31,126,31,66,31,105,31,252,31,191,31,238,31,41,31,178,31,178,30,220,31,220,30,167,31,167,30,63,31,63,30,63,29,40,31,32,31,147,31,115,31,7,31,62,31,161,31,156,31,156,30,145,31,145,30,219,31,219,30,201,31,187,31,187,31,169,31,169,30,197,31,163,31,163,30,12,31,12,30,12,29,54,31,86,31,242,31,116,31,45,31,38,31,42,31,94,31,94,30,158,31,27,31,59,31,201,31,201,30,155,31,23,31,60,31,203,31,10,31,86,31,75,31,185,31,87,31,239,31,79,31,123,31,198,31,161,31,117,31,147,31,147,30,147,29,252,31,252,30,198,31,72,31,72,30,82,31,139,31,16,31,51,31,11,31,254,31,164,31,205,31,142,31,142,30,21,31,21,30,180,31,203,31,203,30,131,31,203,31,80,31,80,30,196,31,11,31,189,31,23,31,120,31,231,31,119,31,195,31,59,31,59,30,158,31,15,31,15,30,240,31,240,30,140,31,161,31,149,31,149,30,178,31,178,30,178,29,178,28,179,31,236,31,18,31,18,30,55,31,133,31,251,31,215,31,54,31,189,31,6,31,6,30,101,31,130,31,130,30,130,29,75,31,50,31,58,31,59,31,14,31,14,30,62,31,224,31,206,31,192,31,207,31,239,31,239,30,41,31,41,30,41,29,117,31,103,31,54,31,112,31,190,31,107,31,98,31,98,30,140,31,42,31,255,31,255,30,180,31,64,31,126,31,15,31,15,30,200,31,200,30,19,31,5,31,133,31,64,31,255,31,1,31,46,31,51,31,95,31,231,31,132,31,92,31,18,31,18,30,18,29,149,31,14,31,158,31,252,31,129,31,221,31,221,30,146,31,25,31,25,30,98,31,98,30,37,31,37,31,63,31,91,31,160,31,160,30,200,31,17,31,244,31,68,31,120,31,120,30,112,31,126,31,210,31,178,31,5,31,96,31,96,30,96,29,112,31,112,31,186,31,229,31,229,30,23,31,1,31,21,31,27,31,180,31,181,31,23,31,95,31,205,31,242,31,242,30,132,31,189,31,69,31,210,31,54,31,40,31,14,31,31,31,54,31,108,31,13,31,13,30,67,31,138,31,135,31,232,31,198,31,77,31,235,31,235,30,54,31,232,31,232,30,189,31,247,31,89,31,16,31,32,31,14,31,242,31,242,30,119,31,140,31,186,31,153,31,94,31,183,31,147,31,54,31,92,31,105,31,183,31,183,30,212,31,111,31,111,30,111,29,66,31,62,31,131,31,231,31,121,31,50,31,50,30,242,31,177,31,3,31,206,31,223,31,246,31,224,31,224,30,241,31,147,31,236,31,123,31,39,31,39,30,76,31,114,31,242,31,21,31,162,31,171,31,40,31,113,31,53,31,222,31,47,31,40,31,17,31,121,31,238,31,94,31,36,31,134,31,54,31,86,31,106,31,106,30,68,31,68,30,119,31,250,31,47,31,215,31,215,30,227,31,139,31,156,31,92,31,92,30,72,31,172,31,202,31,202,30,104,31,116,31,116,30,143,31,60,31,60,30,60,29,60,28,169,31,133,31,225,31,14,31,2,31,32,31,32,30,186,31,206,31,206,30,12,31,12,30,223,31,168,31,231,31,85,31,56,31,116,31,105,31,54,31,54,30,190,31,97,31,168,31,37,31,215,31,144,31,200,31,251,31,251,30,82,31,232,31,249,31,38,31,32,31,32,30,32,29,144,31,81,31,223,31,223,30,165,31,115,31,176,31,87,31,87,30,65,31,67,31,53,31,193,31,12,31,175,31,23,31,205,31,101,31,50,31,50,30,188,31,236,31,189,31,103,31,103,30,103,29,199,31,200,31,177,31,133,31,200,31,61,31,154,31,158,31,158,30,102,31,242,31,57,31,57,30,119,31,98,31,2,31,232,31,232,30,57,31,51,31,84,31,130,31,192,31,192,30,212,31,175,31,175,30,1,31,98,31,50,31,243,31,156,31,223,31,125,31,180,31,190,31,36,31,76,31,76,30,14,31,252,31,174,31,65,31,101,31,61,31,87,31,231,31,165,31,165,30,105,31,10,31,10,30,252,31,252,30,137,31,55,31,135,31,135,30,219,31,219,30,233,31,144,31,182,31,6,31,6,30,246,31,48,31,41,31,71,31,71,30,71,29,57,31,27,31,241,31,19,31,19,30,36,31,216,31,214,31,132,31,197,31,197,30,95,31,212,31,146,31,232,31,212,31,163,31,231,31,91,31,2,31,207,31,164,31,164,30,164,29,164,28,29,31,144,31,32,31,237,31,95,31,95,30,131,31,88,31,203,31,207,31,229,31,171,31,207,31,168,31,168,30,14,31,153,31,190,31,189,31,204,31,13,31,98,31,62,31,49,31,49,30,131,31,235,31,195,31,120,31,102,31,171,31,171,30,66,31,48,31,234,31,39,31,13,31,163,31,96,31,202,31,202,31,21,31,153,31,153,30,16,31,13,31,181,31,181,30,181,29,173,31,23,31,34,31,142,31,143,31,53,31,53,30,157,31,44,31,225,31,241,31,102,31,108,31,68,31,68,30,1,31,1,30,205,31,205,30,205,29,3,31,138,31,19,31,165,31,45,31,162,31,100,31,230,31,51,31,77,31,110,31,110,30,110,29,163,31,87,31,68,31,224,31,224,30,196,31,13,31,94,31,194,31,29,31,43,31,170,31,170,30,233,31,132,31,203,31,97,31,58,31,231,31,53,31,245,31,120,31,120,30,120,29,172,31,73,31,67,31,95,31,153,31,224,31,186,31,111,31,81,31,81,30,203,31,20,31,189,31,169,31,187,31,139,31,138,31,35,31,70,31,218,31,218,30,218,29,110,31,167,31,189,31,160,31,22,31,29,31,89,31,65,31,190,31,44,31,44,30,44,29,146,31,230,31,230,30,41,31,41,30,242,31,149,31,201,31,218,31,63,31,63,30,47,31,228,31,206,31,118,31,118,30,118,29,39,31,151,31,18,31,5,31,224,31,252,31,184,31,140,31,140,30,160,31,69,31,108,31,108,30,194,31,216,31,76,31,47,31,47,30,74,31,104,31,131,31,121,31,198,31,198,30,198,29,83,31,60,31,219,31,22,31,22,30,181,31,168,31,49,31,30,31,30,30,65,31,102,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
