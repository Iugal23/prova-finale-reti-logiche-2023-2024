-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_358 is
end project_tb_358;

architecture project_tb_arch_358 of project_tb_358 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 238;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (204,0,212,0,245,0,0,0,0,0,0,0,145,0,59,0,185,0,2,0,97,0,208,0,0,0,174,0,110,0,215,0,91,0,253,0,0,0,0,0,0,0,0,0,142,0,111,0,135,0,204,0,88,0,39,0,45,0,0,0,216,0,253,0,86,0,15,0,14,0,17,0,23,0,0,0,144,0,38,0,0,0,178,0,93,0,168,0,208,0,36,0,76,0,176,0,255,0,253,0,54,0,156,0,186,0,137,0,46,0,0,0,88,0,0,0,231,0,174,0,121,0,0,0,27,0,94,0,0,0,234,0,36,0,254,0,66,0,17,0,201,0,0,0,20,0,166,0,114,0,105,0,0,0,0,0,141,0,192,0,146,0,69,0,7,0,140,0,180,0,107,0,243,0,56,0,64,0,0,0,209,0,34,0,0,0,60,0,0,0,0,0,56,0,0,0,118,0,254,0,224,0,0,0,182,0,103,0,231,0,139,0,121,0,0,0,0,0,53,0,58,0,113,0,118,0,242,0,63,0,222,0,39,0,232,0,189,0,202,0,27,0,205,0,68,0,1,0,0,0,198,0,0,0,0,0,148,0,0,0,235,0,0,0,32,0,0,0,249,0,242,0,212,0,125,0,0,0,201,0,145,0,0,0,205,0,191,0,8,0,83,0,48,0,61,0,0,0,134,0,254,0,224,0,131,0,0,0,203,0,145,0,229,0,76,0,245,0,6,0,252,0,88,0,224,0,0,0,126,0,75,0,128,0,226,0,237,0,0,0,223,0,62,0,60,0,0,0,93,0,75,0,29,0,127,0,97,0,232,0,54,0,0,0,148,0,132,0,87,0,103,0,137,0,229,0,207,0,100,0,178,0,143,0,73,0,253,0,79,0,181,0,241,0,106,0,168,0,224,0,199,0,3,0,114,0,175,0,63,0,141,0,107,0,0,0,0,0,30,0,158,0,0,0,124,0,212,0,162,0,224,0,236,0,157,0,0,0,43,0,228,0,224,0,45,0,190,0,0,0,0,0,27,0,0,0,126,0,36,0,202,0,40,0,78,0,250,0,0,0,0,0,120,0,0,0);
signal scenario_full  : scenario_type := (204,31,212,31,245,31,245,30,245,29,245,28,145,31,59,31,185,31,2,31,97,31,208,31,208,30,174,31,110,31,215,31,91,31,253,31,253,30,253,29,253,28,253,27,142,31,111,31,135,31,204,31,88,31,39,31,45,31,45,30,216,31,253,31,86,31,15,31,14,31,17,31,23,31,23,30,144,31,38,31,38,30,178,31,93,31,168,31,208,31,36,31,76,31,176,31,255,31,253,31,54,31,156,31,186,31,137,31,46,31,46,30,88,31,88,30,231,31,174,31,121,31,121,30,27,31,94,31,94,30,234,31,36,31,254,31,66,31,17,31,201,31,201,30,20,31,166,31,114,31,105,31,105,30,105,29,141,31,192,31,146,31,69,31,7,31,140,31,180,31,107,31,243,31,56,31,64,31,64,30,209,31,34,31,34,30,60,31,60,30,60,29,56,31,56,30,118,31,254,31,224,31,224,30,182,31,103,31,231,31,139,31,121,31,121,30,121,29,53,31,58,31,113,31,118,31,242,31,63,31,222,31,39,31,232,31,189,31,202,31,27,31,205,31,68,31,1,31,1,30,198,31,198,30,198,29,148,31,148,30,235,31,235,30,32,31,32,30,249,31,242,31,212,31,125,31,125,30,201,31,145,31,145,30,205,31,191,31,8,31,83,31,48,31,61,31,61,30,134,31,254,31,224,31,131,31,131,30,203,31,145,31,229,31,76,31,245,31,6,31,252,31,88,31,224,31,224,30,126,31,75,31,128,31,226,31,237,31,237,30,223,31,62,31,60,31,60,30,93,31,75,31,29,31,127,31,97,31,232,31,54,31,54,30,148,31,132,31,87,31,103,31,137,31,229,31,207,31,100,31,178,31,143,31,73,31,253,31,79,31,181,31,241,31,106,31,168,31,224,31,199,31,3,31,114,31,175,31,63,31,141,31,107,31,107,30,107,29,30,31,158,31,158,30,124,31,212,31,162,31,224,31,236,31,157,31,157,30,43,31,228,31,224,31,45,31,190,31,190,30,190,29,27,31,27,30,126,31,36,31,202,31,40,31,78,31,250,31,250,30,250,29,120,31,120,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
