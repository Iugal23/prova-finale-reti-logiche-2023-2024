-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_778 is
end project_tb_778;

architecture project_tb_arch_778 of project_tb_778 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 604;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,190,0,0,0,33,0,194,0,142,0,103,0,26,0,3,0,0,0,0,0,39,0,61,0,0,0,48,0,100,0,190,0,227,0,136,0,6,0,141,0,190,0,157,0,0,0,140,0,129,0,32,0,70,0,125,0,26,0,9,0,0,0,68,0,129,0,235,0,154,0,178,0,216,0,215,0,0,0,75,0,134,0,10,0,239,0,214,0,0,0,151,0,242,0,155,0,179,0,214,0,147,0,113,0,123,0,0,0,4,0,141,0,165,0,106,0,135,0,26,0,156,0,20,0,0,0,17,0,203,0,229,0,233,0,0,0,190,0,0,0,0,0,201,0,20,0,110,0,207,0,133,0,220,0,14,0,160,0,49,0,3,0,226,0,214,0,51,0,116,0,77,0,178,0,0,0,7,0,0,0,49,0,7,0,44,0,124,0,37,0,142,0,177,0,0,0,118,0,226,0,220,0,84,0,200,0,180,0,104,0,184,0,0,0,231,0,0,0,59,0,200,0,185,0,133,0,0,0,244,0,122,0,53,0,36,0,24,0,94,0,0,0,0,0,0,0,200,0,139,0,232,0,75,0,155,0,246,0,79,0,54,0,189,0,13,0,125,0,125,0,27,0,154,0,48,0,0,0,122,0,125,0,245,0,24,0,0,0,19,0,21,0,96,0,0,0,189,0,232,0,8,0,0,0,123,0,0,0,164,0,237,0,224,0,158,0,216,0,0,0,66,0,182,0,248,0,0,0,49,0,28,0,0,0,113,0,28,0,234,0,46,0,208,0,0,0,111,0,215,0,147,0,118,0,83,0,124,0,108,0,107,0,0,0,121,0,1,0,161,0,107,0,177,0,0,0,240,0,175,0,6,0,86,0,0,0,176,0,0,0,61,0,0,0,75,0,0,0,62,0,0,0,69,0,235,0,172,0,140,0,159,0,37,0,190,0,127,0,249,0,206,0,63,0,28,0,201,0,36,0,232,0,45,0,227,0,217,0,0,0,53,0,0,0,240,0,231,0,0,0,91,0,163,0,0,0,36,0,15,0,154,0,11,0,126,0,199,0,186,0,0,0,19,0,0,0,212,0,111,0,157,0,0,0,0,0,0,0,131,0,10,0,227,0,136,0,176,0,117,0,118,0,255,0,46,0,45,0,0,0,223,0,215,0,0,0,79,0,113,0,0,0,53,0,6,0,74,0,52,0,60,0,125,0,0,0,0,0,76,0,127,0,154,0,0,0,80,0,120,0,31,0,90,0,252,0,248,0,0,0,78,0,7,0,7,0,239,0,237,0,226,0,194,0,183,0,178,0,134,0,171,0,189,0,0,0,189,0,0,0,191,0,94,0,177,0,216,0,245,0,113,0,102,0,239,0,0,0,219,0,0,0,7,0,37,0,0,0,24,0,119,0,0,0,45,0,240,0,251,0,0,0,66,0,151,0,176,0,0,0,0,0,0,0,187,0,108,0,213,0,0,0,0,0,179,0,15,0,206,0,5,0,38,0,171,0,15,0,0,0,1,0,0,0,95,0,122,0,243,0,153,0,3,0,162,0,0,0,215,0,129,0,184,0,181,0,64,0,95,0,71,0,231,0,60,0,0,0,0,0,106,0,0,0,0,0,0,0,0,0,128,0,0,0,118,0,150,0,207,0,0,0,220,0,27,0,55,0,188,0,56,0,91,0,146,0,48,0,0,0,112,0,56,0,109,0,56,0,51,0,71,0,0,0,91,0,94,0,109,0,244,0,67,0,183,0,201,0,224,0,0,0,158,0,36,0,196,0,111,0,127,0,0,0,52,0,0,0,178,0,106,0,215,0,231,0,0,0,155,0,0,0,4,0,182,0,234,0,103,0,175,0,0,0,120,0,201,0,0,0,32,0,200,0,44,0,120,0,0,0,59,0,61,0,160,0,0,0,26,0,0,0,78,0,249,0,0,0,2,0,65,0,0,0,209,0,0,0,118,0,38,0,0,0,0,0,172,0,222,0,60,0,176,0,29,0,0,0,244,0,112,0,167,0,140,0,225,0,112,0,172,0,154,0,232,0,0,0,123,0,61,0,4,0,174,0,204,0,0,0,2,0,0,0,130,0,54,0,198,0,31,0,89,0,191,0,17,0,235,0,202,0,198,0,0,0,183,0,8,0,137,0,91,0,112,0,0,0,194,0,0,0,154,0,166,0,198,0,92,0,186,0,144,0,0,0,0,0,87,0,119,0,75,0,54,0,0,0,95,0,0,0,69,0,0,0,162,0,0,0,56,0,0,0,201,0,0,0,160,0,164,0,0,0,0,0,237,0,172,0,0,0,123,0,0,0,186,0,81,0,226,0,85,0,49,0,181,0,171,0,0,0,0,0,96,0,0,0,0,0,214,0,0,0,78,0,0,0,68,0,0,0,236,0,142,0,0,0,160,0,41,0,134,0,248,0,17,0,11,0,25,0,225,0,70,0,54,0,73,0,53,0,34,0,184,0,119,0,0,0,153,0,107,0,0,0,40,0,183,0,227,0,39,0,40,0,247,0,46,0,19,0,31,0,186,0,51,0,157,0,248,0,52,0,134,0,35,0,0,0,2,0,86,0,252,0,0,0,244,0,171,0,46,0,0,0,10,0,220,0,153,0,80,0,0,0,139,0,183,0,209,0,0,0,180,0,145,0,211,0,219,0,125,0,7,0,0,0,0,0,142,0,190,0,0,0,218,0,0,0,38,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,190,31,190,30,33,31,194,31,142,31,103,31,26,31,3,31,3,30,3,29,39,31,61,31,61,30,48,31,100,31,190,31,227,31,136,31,6,31,141,31,190,31,157,31,157,30,140,31,129,31,32,31,70,31,125,31,26,31,9,31,9,30,68,31,129,31,235,31,154,31,178,31,216,31,215,31,215,30,75,31,134,31,10,31,239,31,214,31,214,30,151,31,242,31,155,31,179,31,214,31,147,31,113,31,123,31,123,30,4,31,141,31,165,31,106,31,135,31,26,31,156,31,20,31,20,30,17,31,203,31,229,31,233,31,233,30,190,31,190,30,190,29,201,31,20,31,110,31,207,31,133,31,220,31,14,31,160,31,49,31,3,31,226,31,214,31,51,31,116,31,77,31,178,31,178,30,7,31,7,30,49,31,7,31,44,31,124,31,37,31,142,31,177,31,177,30,118,31,226,31,220,31,84,31,200,31,180,31,104,31,184,31,184,30,231,31,231,30,59,31,200,31,185,31,133,31,133,30,244,31,122,31,53,31,36,31,24,31,94,31,94,30,94,29,94,28,200,31,139,31,232,31,75,31,155,31,246,31,79,31,54,31,189,31,13,31,125,31,125,31,27,31,154,31,48,31,48,30,122,31,125,31,245,31,24,31,24,30,19,31,21,31,96,31,96,30,189,31,232,31,8,31,8,30,123,31,123,30,164,31,237,31,224,31,158,31,216,31,216,30,66,31,182,31,248,31,248,30,49,31,28,31,28,30,113,31,28,31,234,31,46,31,208,31,208,30,111,31,215,31,147,31,118,31,83,31,124,31,108,31,107,31,107,30,121,31,1,31,161,31,107,31,177,31,177,30,240,31,175,31,6,31,86,31,86,30,176,31,176,30,61,31,61,30,75,31,75,30,62,31,62,30,69,31,235,31,172,31,140,31,159,31,37,31,190,31,127,31,249,31,206,31,63,31,28,31,201,31,36,31,232,31,45,31,227,31,217,31,217,30,53,31,53,30,240,31,231,31,231,30,91,31,163,31,163,30,36,31,15,31,154,31,11,31,126,31,199,31,186,31,186,30,19,31,19,30,212,31,111,31,157,31,157,30,157,29,157,28,131,31,10,31,227,31,136,31,176,31,117,31,118,31,255,31,46,31,45,31,45,30,223,31,215,31,215,30,79,31,113,31,113,30,53,31,6,31,74,31,52,31,60,31,125,31,125,30,125,29,76,31,127,31,154,31,154,30,80,31,120,31,31,31,90,31,252,31,248,31,248,30,78,31,7,31,7,31,239,31,237,31,226,31,194,31,183,31,178,31,134,31,171,31,189,31,189,30,189,31,189,30,191,31,94,31,177,31,216,31,245,31,113,31,102,31,239,31,239,30,219,31,219,30,7,31,37,31,37,30,24,31,119,31,119,30,45,31,240,31,251,31,251,30,66,31,151,31,176,31,176,30,176,29,176,28,187,31,108,31,213,31,213,30,213,29,179,31,15,31,206,31,5,31,38,31,171,31,15,31,15,30,1,31,1,30,95,31,122,31,243,31,153,31,3,31,162,31,162,30,215,31,129,31,184,31,181,31,64,31,95,31,71,31,231,31,60,31,60,30,60,29,106,31,106,30,106,29,106,28,106,27,128,31,128,30,118,31,150,31,207,31,207,30,220,31,27,31,55,31,188,31,56,31,91,31,146,31,48,31,48,30,112,31,56,31,109,31,56,31,51,31,71,31,71,30,91,31,94,31,109,31,244,31,67,31,183,31,201,31,224,31,224,30,158,31,36,31,196,31,111,31,127,31,127,30,52,31,52,30,178,31,106,31,215,31,231,31,231,30,155,31,155,30,4,31,182,31,234,31,103,31,175,31,175,30,120,31,201,31,201,30,32,31,200,31,44,31,120,31,120,30,59,31,61,31,160,31,160,30,26,31,26,30,78,31,249,31,249,30,2,31,65,31,65,30,209,31,209,30,118,31,38,31,38,30,38,29,172,31,222,31,60,31,176,31,29,31,29,30,244,31,112,31,167,31,140,31,225,31,112,31,172,31,154,31,232,31,232,30,123,31,61,31,4,31,174,31,204,31,204,30,2,31,2,30,130,31,54,31,198,31,31,31,89,31,191,31,17,31,235,31,202,31,198,31,198,30,183,31,8,31,137,31,91,31,112,31,112,30,194,31,194,30,154,31,166,31,198,31,92,31,186,31,144,31,144,30,144,29,87,31,119,31,75,31,54,31,54,30,95,31,95,30,69,31,69,30,162,31,162,30,56,31,56,30,201,31,201,30,160,31,164,31,164,30,164,29,237,31,172,31,172,30,123,31,123,30,186,31,81,31,226,31,85,31,49,31,181,31,171,31,171,30,171,29,96,31,96,30,96,29,214,31,214,30,78,31,78,30,68,31,68,30,236,31,142,31,142,30,160,31,41,31,134,31,248,31,17,31,11,31,25,31,225,31,70,31,54,31,73,31,53,31,34,31,184,31,119,31,119,30,153,31,107,31,107,30,40,31,183,31,227,31,39,31,40,31,247,31,46,31,19,31,31,31,186,31,51,31,157,31,248,31,52,31,134,31,35,31,35,30,2,31,86,31,252,31,252,30,244,31,171,31,46,31,46,30,10,31,220,31,153,31,80,31,80,30,139,31,183,31,209,31,209,30,180,31,145,31,211,31,219,31,125,31,7,31,7,30,7,29,142,31,190,31,190,30,218,31,218,30,38,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
