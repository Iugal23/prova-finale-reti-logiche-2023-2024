-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 648;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (144,0,153,0,81,0,222,0,0,0,19,0,21,0,55,0,0,0,21,0,247,0,112,0,35,0,248,0,227,0,204,0,43,0,172,0,135,0,50,0,196,0,247,0,201,0,116,0,166,0,222,0,109,0,4,0,165,0,89,0,222,0,99,0,2,0,0,0,205,0,223,0,178,0,86,0,238,0,201,0,0,0,164,0,5,0,34,0,229,0,169,0,219,0,206,0,52,0,27,0,232,0,0,0,163,0,44,0,112,0,220,0,0,0,6,0,201,0,253,0,0,0,14,0,65,0,204,0,77,0,0,0,84,0,0,0,229,0,221,0,0,0,0,0,164,0,43,0,0,0,238,0,191,0,122,0,10,0,225,0,0,0,134,0,129,0,148,0,0,0,74,0,61,0,102,0,136,0,97,0,40,0,0,0,194,0,216,0,51,0,4,0,156,0,89,0,47,0,34,0,0,0,232,0,0,0,79,0,226,0,38,0,234,0,233,0,230,0,0,0,16,0,0,0,4,0,0,0,153,0,210,0,206,0,164,0,233,0,208,0,184,0,222,0,0,0,156,0,41,0,34,0,10,0,181,0,222,0,12,0,47,0,122,0,97,0,225,0,214,0,44,0,249,0,78,0,235,0,230,0,238,0,0,0,84,0,35,0,192,0,82,0,44,0,100,0,213,0,77,0,96,0,130,0,183,0,248,0,233,0,249,0,43,0,0,0,110,0,125,0,188,0,40,0,63,0,175,0,0,0,3,0,41,0,230,0,186,0,254,0,253,0,0,0,92,0,232,0,211,0,87,0,185,0,0,0,92,0,37,0,151,0,96,0,0,0,205,0,5,0,221,0,131,0,0,0,74,0,0,0,39,0,0,0,39,0,141,0,110,0,78,0,197,0,0,0,0,0,168,0,45,0,39,0,239,0,101,0,217,0,128,0,168,0,177,0,165,0,250,0,132,0,37,0,0,0,0,0,0,0,24,0,0,0,17,0,236,0,133,0,65,0,250,0,9,0,0,0,213,0,0,0,86,0,0,0,45,0,0,0,0,0,55,0,214,0,242,0,175,0,114,0,162,0,73,0,0,0,87,0,163,0,0,0,87,0,69,0,12,0,96,0,199,0,87,0,0,0,143,0,0,0,0,0,244,0,18,0,244,0,242,0,0,0,0,0,199,0,239,0,116,0,0,0,42,0,0,0,52,0,0,0,63,0,53,0,78,0,0,0,80,0,137,0,40,0,25,0,0,0,48,0,103,0,191,0,102,0,1,0,0,0,91,0,140,0,98,0,93,0,149,0,223,0,136,0,0,0,0,0,131,0,0,0,61,0,3,0,177,0,250,0,0,0,72,0,139,0,190,0,250,0,0,0,0,0,221,0,0,0,113,0,55,0,106,0,33,0,211,0,0,0,96,0,83,0,0,0,4,0,177,0,10,0,206,0,16,0,0,0,186,0,92,0,89,0,126,0,197,0,185,0,80,0,43,0,65,0,45,0,0,0,31,0,135,0,0,0,13,0,0,0,249,0,11,0,0,0,143,0,3,0,234,0,96,0,0,0,246,0,45,0,114,0,28,0,201,0,151,0,230,0,0,0,69,0,204,0,0,0,178,0,19,0,88,0,154,0,20,0,66,0,248,0,156,0,149,0,198,0,0,0,207,0,51,0,22,0,236,0,231,0,47,0,18,0,30,0,243,0,247,0,218,0,104,0,110,0,227,0,213,0,0,0,217,0,77,0,242,0,0,0,76,0,197,0,0,0,124,0,0,0,79,0,114,0,0,0,124,0,210,0,72,0,181,0,53,0,0,0,72,0,0,0,168,0,171,0,213,0,138,0,40,0,79,0,241,0,44,0,5,0,108,0,0,0,113,0,0,0,226,0,87,0,125,0,65,0,64,0,6,0,122,0,243,0,186,0,52,0,23,0,0,0,0,0,0,0,173,0,201,0,57,0,232,0,88,0,94,0,142,0,204,0,85,0,121,0,166,0,54,0,132,0,0,0,146,0,178,0,156,0,0,0,0,0,159,0,58,0,119,0,0,0,0,0,35,0,153,0,102,0,110,0,51,0,154,0,0,0,152,0,155,0,0,0,208,0,191,0,74,0,86,0,6,0,0,0,82,0,202,0,209,0,0,0,59,0,189,0,0,0,0,0,113,0,134,0,57,0,136,0,125,0,218,0,223,0,81,0,0,0,87,0,43,0,192,0,149,0,51,0,0,0,0,0,197,0,169,0,187,0,240,0,0,0,46,0,182,0,1,0,29,0,79,0,55,0,73,0,0,0,150,0,2,0,17,0,85,0,0,0,72,0,152,0,131,0,20,0,0,0,0,0,245,0,153,0,185,0,12,0,242,0,173,0,240,0,111,0,172,0,105,0,201,0,182,0,40,0,137,0,112,0,52,0,71,0,197,0,97,0,130,0,243,0,201,0,0,0,9,0,146,0,195,0,29,0,84,0,205,0,5,0,173,0,117,0,113,0,78,0,0,0,163,0,0,0,24,0,189,0,99,0,7,0,91,0,0,0,92,0,149,0,150,0,117,0,112,0,193,0,96,0,236,0,248,0,229,0,176,0,128,0,51,0,158,0,0,0,254,0,169,0,5,0,221,0,16,0,165,0,184,0,113,0,168,0,195,0,206,0,0,0,0,0,206,0,0,0,55,0,16,0,87,0,146,0,0,0,0,0,81,0,0,0,217,0,93,0,79,0,206,0,16,0,235,0,223,0,0,0,88,0,0,0,245,0,73,0,98,0,39,0,0,0,0,0,249,0,85,0,218,0,3,0,29,0,215,0,146,0,56,0,189,0,137,0,125,0,203,0,130,0,38,0,166,0,222,0,190,0,35,0,40,0,8,0,31,0,27,0,228,0,29,0,0,0,0,0,0,0,253,0,182,0,0,0,0,0,0,0,96,0,148,0);
signal scenario_full  : scenario_type := (144,31,153,31,81,31,222,31,222,30,19,31,21,31,55,31,55,30,21,31,247,31,112,31,35,31,248,31,227,31,204,31,43,31,172,31,135,31,50,31,196,31,247,31,201,31,116,31,166,31,222,31,109,31,4,31,165,31,89,31,222,31,99,31,2,31,2,30,205,31,223,31,178,31,86,31,238,31,201,31,201,30,164,31,5,31,34,31,229,31,169,31,219,31,206,31,52,31,27,31,232,31,232,30,163,31,44,31,112,31,220,31,220,30,6,31,201,31,253,31,253,30,14,31,65,31,204,31,77,31,77,30,84,31,84,30,229,31,221,31,221,30,221,29,164,31,43,31,43,30,238,31,191,31,122,31,10,31,225,31,225,30,134,31,129,31,148,31,148,30,74,31,61,31,102,31,136,31,97,31,40,31,40,30,194,31,216,31,51,31,4,31,156,31,89,31,47,31,34,31,34,30,232,31,232,30,79,31,226,31,38,31,234,31,233,31,230,31,230,30,16,31,16,30,4,31,4,30,153,31,210,31,206,31,164,31,233,31,208,31,184,31,222,31,222,30,156,31,41,31,34,31,10,31,181,31,222,31,12,31,47,31,122,31,97,31,225,31,214,31,44,31,249,31,78,31,235,31,230,31,238,31,238,30,84,31,35,31,192,31,82,31,44,31,100,31,213,31,77,31,96,31,130,31,183,31,248,31,233,31,249,31,43,31,43,30,110,31,125,31,188,31,40,31,63,31,175,31,175,30,3,31,41,31,230,31,186,31,254,31,253,31,253,30,92,31,232,31,211,31,87,31,185,31,185,30,92,31,37,31,151,31,96,31,96,30,205,31,5,31,221,31,131,31,131,30,74,31,74,30,39,31,39,30,39,31,141,31,110,31,78,31,197,31,197,30,197,29,168,31,45,31,39,31,239,31,101,31,217,31,128,31,168,31,177,31,165,31,250,31,132,31,37,31,37,30,37,29,37,28,24,31,24,30,17,31,236,31,133,31,65,31,250,31,9,31,9,30,213,31,213,30,86,31,86,30,45,31,45,30,45,29,55,31,214,31,242,31,175,31,114,31,162,31,73,31,73,30,87,31,163,31,163,30,87,31,69,31,12,31,96,31,199,31,87,31,87,30,143,31,143,30,143,29,244,31,18,31,244,31,242,31,242,30,242,29,199,31,239,31,116,31,116,30,42,31,42,30,52,31,52,30,63,31,53,31,78,31,78,30,80,31,137,31,40,31,25,31,25,30,48,31,103,31,191,31,102,31,1,31,1,30,91,31,140,31,98,31,93,31,149,31,223,31,136,31,136,30,136,29,131,31,131,30,61,31,3,31,177,31,250,31,250,30,72,31,139,31,190,31,250,31,250,30,250,29,221,31,221,30,113,31,55,31,106,31,33,31,211,31,211,30,96,31,83,31,83,30,4,31,177,31,10,31,206,31,16,31,16,30,186,31,92,31,89,31,126,31,197,31,185,31,80,31,43,31,65,31,45,31,45,30,31,31,135,31,135,30,13,31,13,30,249,31,11,31,11,30,143,31,3,31,234,31,96,31,96,30,246,31,45,31,114,31,28,31,201,31,151,31,230,31,230,30,69,31,204,31,204,30,178,31,19,31,88,31,154,31,20,31,66,31,248,31,156,31,149,31,198,31,198,30,207,31,51,31,22,31,236,31,231,31,47,31,18,31,30,31,243,31,247,31,218,31,104,31,110,31,227,31,213,31,213,30,217,31,77,31,242,31,242,30,76,31,197,31,197,30,124,31,124,30,79,31,114,31,114,30,124,31,210,31,72,31,181,31,53,31,53,30,72,31,72,30,168,31,171,31,213,31,138,31,40,31,79,31,241,31,44,31,5,31,108,31,108,30,113,31,113,30,226,31,87,31,125,31,65,31,64,31,6,31,122,31,243,31,186,31,52,31,23,31,23,30,23,29,23,28,173,31,201,31,57,31,232,31,88,31,94,31,142,31,204,31,85,31,121,31,166,31,54,31,132,31,132,30,146,31,178,31,156,31,156,30,156,29,159,31,58,31,119,31,119,30,119,29,35,31,153,31,102,31,110,31,51,31,154,31,154,30,152,31,155,31,155,30,208,31,191,31,74,31,86,31,6,31,6,30,82,31,202,31,209,31,209,30,59,31,189,31,189,30,189,29,113,31,134,31,57,31,136,31,125,31,218,31,223,31,81,31,81,30,87,31,43,31,192,31,149,31,51,31,51,30,51,29,197,31,169,31,187,31,240,31,240,30,46,31,182,31,1,31,29,31,79,31,55,31,73,31,73,30,150,31,2,31,17,31,85,31,85,30,72,31,152,31,131,31,20,31,20,30,20,29,245,31,153,31,185,31,12,31,242,31,173,31,240,31,111,31,172,31,105,31,201,31,182,31,40,31,137,31,112,31,52,31,71,31,197,31,97,31,130,31,243,31,201,31,201,30,9,31,146,31,195,31,29,31,84,31,205,31,5,31,173,31,117,31,113,31,78,31,78,30,163,31,163,30,24,31,189,31,99,31,7,31,91,31,91,30,92,31,149,31,150,31,117,31,112,31,193,31,96,31,236,31,248,31,229,31,176,31,128,31,51,31,158,31,158,30,254,31,169,31,5,31,221,31,16,31,165,31,184,31,113,31,168,31,195,31,206,31,206,30,206,29,206,31,206,30,55,31,16,31,87,31,146,31,146,30,146,29,81,31,81,30,217,31,93,31,79,31,206,31,16,31,235,31,223,31,223,30,88,31,88,30,245,31,73,31,98,31,39,31,39,30,39,29,249,31,85,31,218,31,3,31,29,31,215,31,146,31,56,31,189,31,137,31,125,31,203,31,130,31,38,31,166,31,222,31,190,31,35,31,40,31,8,31,31,31,27,31,228,31,29,31,29,30,29,29,29,28,253,31,182,31,182,30,182,29,182,28,96,31,148,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
