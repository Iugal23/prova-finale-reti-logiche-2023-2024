-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 659;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,0,0,201,0,103,0,0,0,0,0,34,0,143,0,18,0,0,0,88,0,157,0,0,0,164,0,89,0,251,0,15,0,0,0,81,0,153,0,0,0,0,0,208,0,118,0,0,0,132,0,163,0,80,0,0,0,0,0,32,0,60,0,159,0,219,0,66,0,0,0,216,0,238,0,135,0,247,0,34,0,13,0,191,0,135,0,2,0,191,0,1,0,211,0,65,0,232,0,217,0,214,0,112,0,77,0,5,0,49,0,23,0,0,0,107,0,237,0,134,0,0,0,150,0,133,0,121,0,158,0,227,0,132,0,163,0,113,0,245,0,8,0,204,0,99,0,245,0,41,0,37,0,55,0,52,0,118,0,12,0,195,0,137,0,132,0,0,0,144,0,207,0,84,0,13,0,134,0,199,0,187,0,32,0,0,0,0,0,62,0,103,0,40,0,237,0,221,0,199,0,0,0,33,0,27,0,249,0,8,0,162,0,30,0,107,0,149,0,37,0,145,0,163,0,127,0,235,0,4,0,113,0,0,0,207,0,0,0,10,0,238,0,0,0,167,0,119,0,57,0,187,0,75,0,169,0,72,0,17,0,105,0,0,0,203,0,131,0,0,0,205,0,6,0,237,0,249,0,81,0,232,0,67,0,0,0,0,0,158,0,76,0,0,0,39,0,170,0,0,0,0,0,74,0,72,0,26,0,251,0,33,0,114,0,67,0,99,0,76,0,96,0,203,0,151,0,47,0,128,0,205,0,114,0,253,0,0,0,172,0,170,0,0,0,0,0,0,0,241,0,212,0,110,0,194,0,34,0,149,0,140,0,194,0,0,0,112,0,84,0,82,0,2,0,90,0,0,0,253,0,182,0,0,0,38,0,105,0,51,0,0,0,233,0,71,0,28,0,19,0,241,0,35,0,230,0,144,0,46,0,202,0,78,0,254,0,183,0,56,0,6,0,0,0,179,0,0,0,3,0,116,0,176,0,117,0,38,0,13,0,71,0,19,0,127,0,0,0,0,0,160,0,139,0,241,0,130,0,203,0,225,0,94,0,0,0,0,0,41,0,0,0,34,0,0,0,247,0,10,0,208,0,204,0,0,0,87,0,0,0,63,0,223,0,5,0,139,0,77,0,251,0,132,0,104,0,251,0,212,0,105,0,0,0,24,0,149,0,232,0,104,0,121,0,91,0,0,0,69,0,251,0,198,0,0,0,157,0,0,0,178,0,190,0,210,0,132,0,137,0,0,0,254,0,105,0,102,0,105,0,189,0,153,0,168,0,244,0,144,0,236,0,140,0,234,0,184,0,0,0,0,0,76,0,162,0,12,0,138,0,153,0,197,0,82,0,0,0,1,0,0,0,28,0,0,0,0,0,180,0,139,0,55,0,0,0,155,0,109,0,0,0,45,0,0,0,150,0,231,0,196,0,241,0,17,0,10,0,77,0,223,0,131,0,0,0,227,0,25,0,18,0,0,0,8,0,128,0,90,0,58,0,29,0,27,0,73,0,120,0,86,0,34,0,186,0,100,0,0,0,239,0,61,0,24,0,205,0,174,0,147,0,240,0,143,0,85,0,18,0,0,0,77,0,50,0,0,0,182,0,0,0,16,0,55,0,50,0,62,0,93,0,0,0,0,0,91,0,0,0,122,0,59,0,145,0,70,0,181,0,239,0,173,0,245,0,0,0,11,0,0,0,30,0,165,0,116,0,177,0,188,0,45,0,71,0,0,0,0,0,181,0,15,0,19,0,110,0,0,0,0,0,169,0,154,0,127,0,0,0,231,0,75,0,97,0,118,0,206,0,98,0,140,0,61,0,100,0,141,0,217,0,160,0,24,0,217,0,97,0,30,0,234,0,190,0,0,0,54,0,0,0,0,0,212,0,242,0,207,0,108,0,113,0,47,0,13,0,65,0,190,0,78,0,238,0,67,0,164,0,126,0,206,0,85,0,169,0,83,0,0,0,247,0,108,0,0,0,239,0,192,0,0,0,0,0,248,0,0,0,129,0,42,0,0,0,159,0,147,0,206,0,77,0,97,0,71,0,68,0,0,0,112,0,36,0,24,0,108,0,155,0,242,0,245,0,233,0,193,0,2,0,80,0,243,0,70,0,0,0,199,0,176,0,163,0,140,0,68,0,112,0,56,0,203,0,0,0,0,0,100,0,237,0,0,0,0,0,9,0,0,0,135,0,45,0,119,0,0,0,170,0,11,0,235,0,244,0,240,0,153,0,136,0,200,0,224,0,125,0,0,0,114,0,0,0,108,0,14,0,0,0,100,0,186,0,85,0,182,0,218,0,145,0,3,0,142,0,0,0,81,0,56,0,183,0,197,0,201,0,96,0,37,0,10,0,125,0,33,0,28,0,251,0,106,0,137,0,155,0,66,0,0,0,55,0,83,0,233,0,248,0,0,0,46,0,72,0,0,0,41,0,70,0,22,0,14,0,34,0,43,0,15,0,201,0,20,0,7,0,75,0,206,0,23,0,0,0,0,0,84,0,106,0,0,0,245,0,194,0,0,0,0,0,222,0,90,0,0,0,66,0,0,0,174,0,142,0,244,0,186,0,174,0,75,0,72,0,73,0,15,0,167,0,238,0,134,0,251,0,242,0,49,0,195,0,44,0,51,0,0,0,18,0,198,0,73,0,135,0,94,0,39,0,184,0,0,0,0,0,198,0,0,0,217,0,0,0,241,0,220,0,71,0,179,0,143,0,120,0,201,0,34,0,38,0,0,0,105,0,167,0,253,0,73,0,37,0,147,0,51,0,32,0,190,0,252,0,1,0,0,0,0,0,124,0,238,0,88,0,55,0,36,0,12,0,49,0,0,0,73,0,90,0,149,0,29,0,129,0,0,0,32,0,210,0,96,0,0,0,0,0,0,0,0,0,62,0,220,0,1,0,0,0,0,0,36,0,164,0,45,0,211,0,235,0,63,0,0,0,51,0,187,0,96,0);
signal scenario_full  : scenario_type := (35,31,35,30,201,31,103,31,103,30,103,29,34,31,143,31,18,31,18,30,88,31,157,31,157,30,164,31,89,31,251,31,15,31,15,30,81,31,153,31,153,30,153,29,208,31,118,31,118,30,132,31,163,31,80,31,80,30,80,29,32,31,60,31,159,31,219,31,66,31,66,30,216,31,238,31,135,31,247,31,34,31,13,31,191,31,135,31,2,31,191,31,1,31,211,31,65,31,232,31,217,31,214,31,112,31,77,31,5,31,49,31,23,31,23,30,107,31,237,31,134,31,134,30,150,31,133,31,121,31,158,31,227,31,132,31,163,31,113,31,245,31,8,31,204,31,99,31,245,31,41,31,37,31,55,31,52,31,118,31,12,31,195,31,137,31,132,31,132,30,144,31,207,31,84,31,13,31,134,31,199,31,187,31,32,31,32,30,32,29,62,31,103,31,40,31,237,31,221,31,199,31,199,30,33,31,27,31,249,31,8,31,162,31,30,31,107,31,149,31,37,31,145,31,163,31,127,31,235,31,4,31,113,31,113,30,207,31,207,30,10,31,238,31,238,30,167,31,119,31,57,31,187,31,75,31,169,31,72,31,17,31,105,31,105,30,203,31,131,31,131,30,205,31,6,31,237,31,249,31,81,31,232,31,67,31,67,30,67,29,158,31,76,31,76,30,39,31,170,31,170,30,170,29,74,31,72,31,26,31,251,31,33,31,114,31,67,31,99,31,76,31,96,31,203,31,151,31,47,31,128,31,205,31,114,31,253,31,253,30,172,31,170,31,170,30,170,29,170,28,241,31,212,31,110,31,194,31,34,31,149,31,140,31,194,31,194,30,112,31,84,31,82,31,2,31,90,31,90,30,253,31,182,31,182,30,38,31,105,31,51,31,51,30,233,31,71,31,28,31,19,31,241,31,35,31,230,31,144,31,46,31,202,31,78,31,254,31,183,31,56,31,6,31,6,30,179,31,179,30,3,31,116,31,176,31,117,31,38,31,13,31,71,31,19,31,127,31,127,30,127,29,160,31,139,31,241,31,130,31,203,31,225,31,94,31,94,30,94,29,41,31,41,30,34,31,34,30,247,31,10,31,208,31,204,31,204,30,87,31,87,30,63,31,223,31,5,31,139,31,77,31,251,31,132,31,104,31,251,31,212,31,105,31,105,30,24,31,149,31,232,31,104,31,121,31,91,31,91,30,69,31,251,31,198,31,198,30,157,31,157,30,178,31,190,31,210,31,132,31,137,31,137,30,254,31,105,31,102,31,105,31,189,31,153,31,168,31,244,31,144,31,236,31,140,31,234,31,184,31,184,30,184,29,76,31,162,31,12,31,138,31,153,31,197,31,82,31,82,30,1,31,1,30,28,31,28,30,28,29,180,31,139,31,55,31,55,30,155,31,109,31,109,30,45,31,45,30,150,31,231,31,196,31,241,31,17,31,10,31,77,31,223,31,131,31,131,30,227,31,25,31,18,31,18,30,8,31,128,31,90,31,58,31,29,31,27,31,73,31,120,31,86,31,34,31,186,31,100,31,100,30,239,31,61,31,24,31,205,31,174,31,147,31,240,31,143,31,85,31,18,31,18,30,77,31,50,31,50,30,182,31,182,30,16,31,55,31,50,31,62,31,93,31,93,30,93,29,91,31,91,30,122,31,59,31,145,31,70,31,181,31,239,31,173,31,245,31,245,30,11,31,11,30,30,31,165,31,116,31,177,31,188,31,45,31,71,31,71,30,71,29,181,31,15,31,19,31,110,31,110,30,110,29,169,31,154,31,127,31,127,30,231,31,75,31,97,31,118,31,206,31,98,31,140,31,61,31,100,31,141,31,217,31,160,31,24,31,217,31,97,31,30,31,234,31,190,31,190,30,54,31,54,30,54,29,212,31,242,31,207,31,108,31,113,31,47,31,13,31,65,31,190,31,78,31,238,31,67,31,164,31,126,31,206,31,85,31,169,31,83,31,83,30,247,31,108,31,108,30,239,31,192,31,192,30,192,29,248,31,248,30,129,31,42,31,42,30,159,31,147,31,206,31,77,31,97,31,71,31,68,31,68,30,112,31,36,31,24,31,108,31,155,31,242,31,245,31,233,31,193,31,2,31,80,31,243,31,70,31,70,30,199,31,176,31,163,31,140,31,68,31,112,31,56,31,203,31,203,30,203,29,100,31,237,31,237,30,237,29,9,31,9,30,135,31,45,31,119,31,119,30,170,31,11,31,235,31,244,31,240,31,153,31,136,31,200,31,224,31,125,31,125,30,114,31,114,30,108,31,14,31,14,30,100,31,186,31,85,31,182,31,218,31,145,31,3,31,142,31,142,30,81,31,56,31,183,31,197,31,201,31,96,31,37,31,10,31,125,31,33,31,28,31,251,31,106,31,137,31,155,31,66,31,66,30,55,31,83,31,233,31,248,31,248,30,46,31,72,31,72,30,41,31,70,31,22,31,14,31,34,31,43,31,15,31,201,31,20,31,7,31,75,31,206,31,23,31,23,30,23,29,84,31,106,31,106,30,245,31,194,31,194,30,194,29,222,31,90,31,90,30,66,31,66,30,174,31,142,31,244,31,186,31,174,31,75,31,72,31,73,31,15,31,167,31,238,31,134,31,251,31,242,31,49,31,195,31,44,31,51,31,51,30,18,31,198,31,73,31,135,31,94,31,39,31,184,31,184,30,184,29,198,31,198,30,217,31,217,30,241,31,220,31,71,31,179,31,143,31,120,31,201,31,34,31,38,31,38,30,105,31,167,31,253,31,73,31,37,31,147,31,51,31,32,31,190,31,252,31,1,31,1,30,1,29,124,31,238,31,88,31,55,31,36,31,12,31,49,31,49,30,73,31,90,31,149,31,29,31,129,31,129,30,32,31,210,31,96,31,96,30,96,29,96,28,96,27,62,31,220,31,1,31,1,30,1,29,36,31,164,31,45,31,211,31,235,31,63,31,63,30,51,31,187,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
