-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 812;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (184,0,89,0,206,0,0,0,162,0,106,0,23,0,82,0,22,0,201,0,60,0,0,0,207,0,13,0,192,0,166,0,142,0,227,0,108,0,94,0,52,0,112,0,98,0,245,0,168,0,182,0,119,0,0,0,245,0,98,0,229,0,76,0,0,0,249,0,22,0,27,0,130,0,169,0,253,0,91,0,0,0,39,0,143,0,192,0,103,0,87,0,246,0,206,0,21,0,24,0,222,0,56,0,125,0,186,0,0,0,0,0,149,0,0,0,0,0,134,0,0,0,197,0,217,0,125,0,149,0,9,0,9,0,0,0,192,0,123,0,2,0,87,0,130,0,39,0,64,0,5,0,105,0,0,0,0,0,112,0,111,0,36,0,0,0,70,0,82,0,0,0,148,0,69,0,231,0,223,0,143,0,0,0,244,0,0,0,72,0,153,0,18,0,136,0,25,0,157,0,96,0,0,0,142,0,62,0,179,0,72,0,33,0,205,0,0,0,106,0,30,0,122,0,217,0,0,0,0,0,0,0,135,0,249,0,0,0,195,0,102,0,0,0,51,0,158,0,103,0,174,0,0,0,0,0,0,0,230,0,104,0,0,0,0,0,0,0,179,0,226,0,156,0,0,0,26,0,190,0,113,0,47,0,0,0,220,0,37,0,154,0,238,0,180,0,78,0,0,0,192,0,0,0,147,0,68,0,174,0,73,0,0,0,166,0,10,0,114,0,184,0,120,0,232,0,80,0,210,0,71,0,0,0,0,0,224,0,233,0,167,0,205,0,82,0,110,0,255,0,64,0,197,0,38,0,0,0,167,0,54,0,224,0,233,0,67,0,3,0,138,0,0,0,93,0,121,0,108,0,140,0,0,0,123,0,0,0,222,0,101,0,197,0,0,0,241,0,3,0,0,0,67,0,59,0,62,0,104,0,204,0,0,0,4,0,163,0,145,0,96,0,112,0,151,0,102,0,139,0,219,0,211,0,185,0,110,0,9,0,26,0,19,0,205,0,223,0,173,0,93,0,166,0,255,0,0,0,151,0,129,0,220,0,0,0,28,0,145,0,106,0,201,0,252,0,236,0,213,0,0,0,123,0,15,0,247,0,10,0,227,0,0,0,0,0,199,0,247,0,151,0,242,0,141,0,73,0,230,0,48,0,201,0,65,0,66,0,201,0,25,0,126,0,34,0,20,0,88,0,0,0,38,0,0,0,0,0,0,0,0,0,0,0,0,0,153,0,0,0,202,0,152,0,198,0,51,0,137,0,240,0,237,0,57,0,47,0,6,0,52,0,0,0,0,0,173,0,220,0,231,0,15,0,116,0,94,0,52,0,20,0,73,0,0,0,0,0,0,0,69,0,182,0,150,0,219,0,98,0,228,0,108,0,192,0,0,0,52,0,127,0,22,0,59,0,52,0,0,0,0,0,255,0,0,0,219,0,250,0,138,0,155,0,174,0,157,0,8,0,41,0,60,0,117,0,47,0,112,0,58,0,227,0,91,0,122,0,185,0,0,0,199,0,172,0,214,0,133,0,3,0,196,0,188,0,250,0,61,0,215,0,135,0,235,0,0,0,170,0,37,0,11,0,239,0,0,0,83,0,188,0,64,0,216,0,190,0,42,0,230,0,55,0,0,0,0,0,162,0,237,0,253,0,219,0,239,0,169,0,96,0,163,0,223,0,116,0,0,0,248,0,220,0,79,0,0,0,0,0,118,0,65,0,227,0,0,0,250,0,227,0,60,0,0,0,119,0,0,0,199,0,40,0,1,0,92,0,53,0,172,0,0,0,155,0,0,0,244,0,216,0,120,0,33,0,190,0,210,0,10,0,158,0,103,0,17,0,249,0,46,0,1,0,245,0,0,0,0,0,22,0,216,0,17,0,81,0,9,0,0,0,183,0,13,0,178,0,117,0,73,0,0,0,243,0,0,0,205,0,101,0,94,0,245,0,0,0,45,0,232,0,0,0,0,0,246,0,0,0,215,0,194,0,160,0,211,0,173,0,178,0,151,0,69,0,0,0,0,0,110,0,86,0,0,0,131,0,41,0,254,0,209,0,125,0,42,0,50,0,130,0,0,0,0,0,77,0,227,0,83,0,0,0,0,0,187,0,255,0,130,0,0,0,126,0,0,0,3,0,112,0,0,0,0,0,112,0,179,0,0,0,50,0,139,0,22,0,161,0,9,0,96,0,227,0,0,0,174,0,220,0,208,0,61,0,106,0,22,0,0,0,171,0,150,0,0,0,0,0,0,0,205,0,26,0,0,0,131,0,54,0,86,0,80,0,13,0,205,0,22,0,238,0,0,0,1,0,249,0,104,0,226,0,87,0,179,0,0,0,0,0,0,0,159,0,0,0,17,0,0,0,0,0,0,0,51,0,93,0,42,0,55,0,13,0,21,0,36,0,0,0,0,0,0,0,150,0,5,0,192,0,201,0,177,0,145,0,1,0,19,0,126,0,201,0,36,0,6,0,58,0,194,0,223,0,15,0,0,0,143,0,76,0,228,0,0,0,70,0,91,0,250,0,200,0,142,0,195,0,56,0,193,0,230,0,74,0,94,0,166,0,125,0,145,0,60,0,153,0,204,0,239,0,15,0,0,0,62,0,209,0,213,0,0,0,193,0,54,0,192,0,186,0,97,0,122,0,181,0,41,0,239,0,78,0,143,0,123,0,236,0,0,0,206,0,142,0,56,0,97,0,102,0,236,0,244,0,12,0,18,0,220,0,47,0,152,0,0,0,21,0,19,0,232,0,161,0,0,0,121,0,230,0,0,0,18,0,244,0,0,0,24,0,240,0,127,0,0,0,206,0,232,0,20,0,41,0,76,0,67,0,116,0,153,0,177,0,0,0,0,0,247,0,206,0,32,0,245,0,0,0,50,0,213,0,71,0,126,0,51,0,172,0,231,0,117,0,166,0,86,0,208,0,175,0,50,0,140,0,223,0,244,0,163,0,40,0,126,0,157,0,29,0,187,0,94,0,0,0,90,0,0,0,0,0,191,0,0,0,90,0,112,0,42,0,160,0,10,0,246,0,97,0,39,0,0,0,133,0,97,0,0,0,0,0,0,0,238,0,255,0,165,0,0,0,157,0,235,0,247,0,110,0,0,0,0,0,165,0,148,0,0,0,19,0,32,0,204,0,129,0,214,0,155,0,0,0,169,0,167,0,0,0,44,0,234,0,199,0,0,0,210,0,0,0,214,0,186,0,30,0,46,0,174,0,81,0,211,0,211,0,255,0,0,0,100,0,100,0,211,0,232,0,19,0,201,0,0,0,63,0,32,0,21,0,100,0,149,0,59,0,221,0,143,0,121,0,66,0,206,0,0,0,135,0,247,0,247,0,149,0,56,0,123,0,125,0,0,0,171,0,7,0,52,0,68,0,56,0,79,0,183,0,200,0,98,0,173,0,193,0,230,0,3,0,36,0,30,0,150,0,149,0,190,0,183,0,199,0,171,0,158,0,85,0,20,0,199,0,0,0,21,0,0,0,205,0,129,0,127,0,67,0,0,0,153,0,5,0,0,0,0,0,218,0,36,0,185,0,233,0,131,0,0,0,72,0,0,0,156,0,126,0,172,0,131,0,239,0,227,0,12,0,0,0,240,0,111,0,212,0,3,0,131,0,48,0,252,0,70,0,0,0);
signal scenario_full  : scenario_type := (184,31,89,31,206,31,206,30,162,31,106,31,23,31,82,31,22,31,201,31,60,31,60,30,207,31,13,31,192,31,166,31,142,31,227,31,108,31,94,31,52,31,112,31,98,31,245,31,168,31,182,31,119,31,119,30,245,31,98,31,229,31,76,31,76,30,249,31,22,31,27,31,130,31,169,31,253,31,91,31,91,30,39,31,143,31,192,31,103,31,87,31,246,31,206,31,21,31,24,31,222,31,56,31,125,31,186,31,186,30,186,29,149,31,149,30,149,29,134,31,134,30,197,31,217,31,125,31,149,31,9,31,9,31,9,30,192,31,123,31,2,31,87,31,130,31,39,31,64,31,5,31,105,31,105,30,105,29,112,31,111,31,36,31,36,30,70,31,82,31,82,30,148,31,69,31,231,31,223,31,143,31,143,30,244,31,244,30,72,31,153,31,18,31,136,31,25,31,157,31,96,31,96,30,142,31,62,31,179,31,72,31,33,31,205,31,205,30,106,31,30,31,122,31,217,31,217,30,217,29,217,28,135,31,249,31,249,30,195,31,102,31,102,30,51,31,158,31,103,31,174,31,174,30,174,29,174,28,230,31,104,31,104,30,104,29,104,28,179,31,226,31,156,31,156,30,26,31,190,31,113,31,47,31,47,30,220,31,37,31,154,31,238,31,180,31,78,31,78,30,192,31,192,30,147,31,68,31,174,31,73,31,73,30,166,31,10,31,114,31,184,31,120,31,232,31,80,31,210,31,71,31,71,30,71,29,224,31,233,31,167,31,205,31,82,31,110,31,255,31,64,31,197,31,38,31,38,30,167,31,54,31,224,31,233,31,67,31,3,31,138,31,138,30,93,31,121,31,108,31,140,31,140,30,123,31,123,30,222,31,101,31,197,31,197,30,241,31,3,31,3,30,67,31,59,31,62,31,104,31,204,31,204,30,4,31,163,31,145,31,96,31,112,31,151,31,102,31,139,31,219,31,211,31,185,31,110,31,9,31,26,31,19,31,205,31,223,31,173,31,93,31,166,31,255,31,255,30,151,31,129,31,220,31,220,30,28,31,145,31,106,31,201,31,252,31,236,31,213,31,213,30,123,31,15,31,247,31,10,31,227,31,227,30,227,29,199,31,247,31,151,31,242,31,141,31,73,31,230,31,48,31,201,31,65,31,66,31,201,31,25,31,126,31,34,31,20,31,88,31,88,30,38,31,38,30,38,29,38,28,38,27,38,26,38,25,153,31,153,30,202,31,152,31,198,31,51,31,137,31,240,31,237,31,57,31,47,31,6,31,52,31,52,30,52,29,173,31,220,31,231,31,15,31,116,31,94,31,52,31,20,31,73,31,73,30,73,29,73,28,69,31,182,31,150,31,219,31,98,31,228,31,108,31,192,31,192,30,52,31,127,31,22,31,59,31,52,31,52,30,52,29,255,31,255,30,219,31,250,31,138,31,155,31,174,31,157,31,8,31,41,31,60,31,117,31,47,31,112,31,58,31,227,31,91,31,122,31,185,31,185,30,199,31,172,31,214,31,133,31,3,31,196,31,188,31,250,31,61,31,215,31,135,31,235,31,235,30,170,31,37,31,11,31,239,31,239,30,83,31,188,31,64,31,216,31,190,31,42,31,230,31,55,31,55,30,55,29,162,31,237,31,253,31,219,31,239,31,169,31,96,31,163,31,223,31,116,31,116,30,248,31,220,31,79,31,79,30,79,29,118,31,65,31,227,31,227,30,250,31,227,31,60,31,60,30,119,31,119,30,199,31,40,31,1,31,92,31,53,31,172,31,172,30,155,31,155,30,244,31,216,31,120,31,33,31,190,31,210,31,10,31,158,31,103,31,17,31,249,31,46,31,1,31,245,31,245,30,245,29,22,31,216,31,17,31,81,31,9,31,9,30,183,31,13,31,178,31,117,31,73,31,73,30,243,31,243,30,205,31,101,31,94,31,245,31,245,30,45,31,232,31,232,30,232,29,246,31,246,30,215,31,194,31,160,31,211,31,173,31,178,31,151,31,69,31,69,30,69,29,110,31,86,31,86,30,131,31,41,31,254,31,209,31,125,31,42,31,50,31,130,31,130,30,130,29,77,31,227,31,83,31,83,30,83,29,187,31,255,31,130,31,130,30,126,31,126,30,3,31,112,31,112,30,112,29,112,31,179,31,179,30,50,31,139,31,22,31,161,31,9,31,96,31,227,31,227,30,174,31,220,31,208,31,61,31,106,31,22,31,22,30,171,31,150,31,150,30,150,29,150,28,205,31,26,31,26,30,131,31,54,31,86,31,80,31,13,31,205,31,22,31,238,31,238,30,1,31,249,31,104,31,226,31,87,31,179,31,179,30,179,29,179,28,159,31,159,30,17,31,17,30,17,29,17,28,51,31,93,31,42,31,55,31,13,31,21,31,36,31,36,30,36,29,36,28,150,31,5,31,192,31,201,31,177,31,145,31,1,31,19,31,126,31,201,31,36,31,6,31,58,31,194,31,223,31,15,31,15,30,143,31,76,31,228,31,228,30,70,31,91,31,250,31,200,31,142,31,195,31,56,31,193,31,230,31,74,31,94,31,166,31,125,31,145,31,60,31,153,31,204,31,239,31,15,31,15,30,62,31,209,31,213,31,213,30,193,31,54,31,192,31,186,31,97,31,122,31,181,31,41,31,239,31,78,31,143,31,123,31,236,31,236,30,206,31,142,31,56,31,97,31,102,31,236,31,244,31,12,31,18,31,220,31,47,31,152,31,152,30,21,31,19,31,232,31,161,31,161,30,121,31,230,31,230,30,18,31,244,31,244,30,24,31,240,31,127,31,127,30,206,31,232,31,20,31,41,31,76,31,67,31,116,31,153,31,177,31,177,30,177,29,247,31,206,31,32,31,245,31,245,30,50,31,213,31,71,31,126,31,51,31,172,31,231,31,117,31,166,31,86,31,208,31,175,31,50,31,140,31,223,31,244,31,163,31,40,31,126,31,157,31,29,31,187,31,94,31,94,30,90,31,90,30,90,29,191,31,191,30,90,31,112,31,42,31,160,31,10,31,246,31,97,31,39,31,39,30,133,31,97,31,97,30,97,29,97,28,238,31,255,31,165,31,165,30,157,31,235,31,247,31,110,31,110,30,110,29,165,31,148,31,148,30,19,31,32,31,204,31,129,31,214,31,155,31,155,30,169,31,167,31,167,30,44,31,234,31,199,31,199,30,210,31,210,30,214,31,186,31,30,31,46,31,174,31,81,31,211,31,211,31,255,31,255,30,100,31,100,31,211,31,232,31,19,31,201,31,201,30,63,31,32,31,21,31,100,31,149,31,59,31,221,31,143,31,121,31,66,31,206,31,206,30,135,31,247,31,247,31,149,31,56,31,123,31,125,31,125,30,171,31,7,31,52,31,68,31,56,31,79,31,183,31,200,31,98,31,173,31,193,31,230,31,3,31,36,31,30,31,150,31,149,31,190,31,183,31,199,31,171,31,158,31,85,31,20,31,199,31,199,30,21,31,21,30,205,31,129,31,127,31,67,31,67,30,153,31,5,31,5,30,5,29,218,31,36,31,185,31,233,31,131,31,131,30,72,31,72,30,156,31,126,31,172,31,131,31,239,31,227,31,12,31,12,30,240,31,111,31,212,31,3,31,131,31,48,31,252,31,70,31,70,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
