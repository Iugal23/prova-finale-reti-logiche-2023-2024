-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_312 is
end project_tb_312;

architecture project_tb_arch_312 of project_tb_312 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 451;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (203,0,0,0,108,0,22,0,117,0,28,0,234,0,53,0,238,0,90,0,0,0,36,0,106,0,88,0,33,0,110,0,65,0,110,0,0,0,228,0,104,0,212,0,0,0,73,0,96,0,67,0,192,0,146,0,61,0,66,0,0,0,0,0,161,0,0,0,61,0,92,0,105,0,0,0,71,0,217,0,0,0,13,0,197,0,37,0,0,0,135,0,168,0,41,0,144,0,151,0,81,0,28,0,122,0,156,0,33,0,7,0,227,0,128,0,53,0,0,0,0,0,240,0,9,0,246,0,197,0,248,0,0,0,234,0,59,0,122,0,181,0,0,0,166,0,0,0,39,0,0,0,0,0,92,0,119,0,0,0,72,0,129,0,203,0,181,0,137,0,174,0,222,0,209,0,196,0,160,0,0,0,0,0,81,0,125,0,210,0,67,0,181,0,0,0,134,0,200,0,54,0,206,0,52,0,0,0,246,0,236,0,214,0,217,0,226,0,3,0,230,0,0,0,134,0,0,0,197,0,0,0,151,0,22,0,193,0,0,0,114,0,65,0,103,0,82,0,0,0,193,0,65,0,123,0,94,0,206,0,40,0,109,0,86,0,167,0,199,0,186,0,144,0,69,0,160,0,98,0,255,0,0,0,93,0,54,0,9,0,88,0,0,0,146,0,85,0,0,0,0,0,55,0,0,0,14,0,124,0,111,0,220,0,187,0,202,0,229,0,20,0,230,0,94,0,194,0,111,0,105,0,54,0,35,0,72,0,54,0,178,0,70,0,184,0,0,0,203,0,114,0,14,0,0,0,159,0,172,0,223,0,194,0,71,0,23,0,0,0,255,0,122,0,0,0,143,0,241,0,45,0,65,0,41,0,37,0,0,0,0,0,137,0,105,0,0,0,248,0,0,0,208,0,118,0,172,0,43,0,177,0,162,0,101,0,161,0,58,0,57,0,107,0,227,0,144,0,138,0,221,0,0,0,34,0,179,0,50,0,34,0,104,0,0,0,0,0,140,0,177,0,123,0,0,0,9,0,122,0,4,0,198,0,47,0,19,0,131,0,189,0,25,0,0,0,255,0,168,0,219,0,0,0,217,0,0,0,78,0,118,0,110,0,137,0,168,0,238,0,164,0,130,0,0,0,81,0,98,0,244,0,242,0,128,0,96,0,0,0,0,0,28,0,0,0,0,0,147,0,212,0,160,0,113,0,92,0,0,0,69,0,160,0,0,0,0,0,63,0,174,0,92,0,253,0,236,0,155,0,0,0,178,0,213,0,88,0,231,0,209,0,166,0,31,0,0,0,94,0,30,0,95,0,94,0,109,0,129,0,163,0,171,0,227,0,34,0,134,0,36,0,240,0,77,0,63,0,125,0,104,0,2,0,120,0,81,0,140,0,173,0,90,0,41,0,32,0,139,0,85,0,43,0,94,0,24,0,244,0,0,0,219,0,0,0,7,0,208,0,13,0,101,0,0,0,68,0,165,0,30,0,57,0,230,0,226,0,115,0,13,0,234,0,171,0,74,0,203,0,191,0,3,0,26,0,0,0,0,0,54,0,138,0,197,0,48,0,210,0,199,0,0,0,56,0,246,0,121,0,185,0,177,0,137,0,25,0,157,0,172,0,0,0,240,0,56,0,0,0,50,0,147,0,0,0,184,0,29,0,0,0,8,0,10,0,204,0,27,0,2,0,35,0,0,0,60,0,71,0,213,0,194,0,167,0,48,0,0,0,0,0,148,0,86,0,245,0,6,0,146,0,0,0,82,0,167,0,241,0,197,0,48,0,131,0,221,0,96,0,77,0,182,0,127,0,254,0,91,0,0,0,116,0,70,0,127,0,7,0,41,0,239,0,123,0,0,0,124,0,227,0,94,0,192,0,18,0,15,0,37,0,44,0,45,0,147,0,0,0,76,0,234,0,0,0,0,0,7,0,142,0,0,0,0,0,3,0,21,0,70,0,99,0,0,0,247,0,218,0,206,0,0,0,166,0,210,0,0,0,131,0,162,0,221,0,156,0,91,0,0,0);
signal scenario_full  : scenario_type := (203,31,203,30,108,31,22,31,117,31,28,31,234,31,53,31,238,31,90,31,90,30,36,31,106,31,88,31,33,31,110,31,65,31,110,31,110,30,228,31,104,31,212,31,212,30,73,31,96,31,67,31,192,31,146,31,61,31,66,31,66,30,66,29,161,31,161,30,61,31,92,31,105,31,105,30,71,31,217,31,217,30,13,31,197,31,37,31,37,30,135,31,168,31,41,31,144,31,151,31,81,31,28,31,122,31,156,31,33,31,7,31,227,31,128,31,53,31,53,30,53,29,240,31,9,31,246,31,197,31,248,31,248,30,234,31,59,31,122,31,181,31,181,30,166,31,166,30,39,31,39,30,39,29,92,31,119,31,119,30,72,31,129,31,203,31,181,31,137,31,174,31,222,31,209,31,196,31,160,31,160,30,160,29,81,31,125,31,210,31,67,31,181,31,181,30,134,31,200,31,54,31,206,31,52,31,52,30,246,31,236,31,214,31,217,31,226,31,3,31,230,31,230,30,134,31,134,30,197,31,197,30,151,31,22,31,193,31,193,30,114,31,65,31,103,31,82,31,82,30,193,31,65,31,123,31,94,31,206,31,40,31,109,31,86,31,167,31,199,31,186,31,144,31,69,31,160,31,98,31,255,31,255,30,93,31,54,31,9,31,88,31,88,30,146,31,85,31,85,30,85,29,55,31,55,30,14,31,124,31,111,31,220,31,187,31,202,31,229,31,20,31,230,31,94,31,194,31,111,31,105,31,54,31,35,31,72,31,54,31,178,31,70,31,184,31,184,30,203,31,114,31,14,31,14,30,159,31,172,31,223,31,194,31,71,31,23,31,23,30,255,31,122,31,122,30,143,31,241,31,45,31,65,31,41,31,37,31,37,30,37,29,137,31,105,31,105,30,248,31,248,30,208,31,118,31,172,31,43,31,177,31,162,31,101,31,161,31,58,31,57,31,107,31,227,31,144,31,138,31,221,31,221,30,34,31,179,31,50,31,34,31,104,31,104,30,104,29,140,31,177,31,123,31,123,30,9,31,122,31,4,31,198,31,47,31,19,31,131,31,189,31,25,31,25,30,255,31,168,31,219,31,219,30,217,31,217,30,78,31,118,31,110,31,137,31,168,31,238,31,164,31,130,31,130,30,81,31,98,31,244,31,242,31,128,31,96,31,96,30,96,29,28,31,28,30,28,29,147,31,212,31,160,31,113,31,92,31,92,30,69,31,160,31,160,30,160,29,63,31,174,31,92,31,253,31,236,31,155,31,155,30,178,31,213,31,88,31,231,31,209,31,166,31,31,31,31,30,94,31,30,31,95,31,94,31,109,31,129,31,163,31,171,31,227,31,34,31,134,31,36,31,240,31,77,31,63,31,125,31,104,31,2,31,120,31,81,31,140,31,173,31,90,31,41,31,32,31,139,31,85,31,43,31,94,31,24,31,244,31,244,30,219,31,219,30,7,31,208,31,13,31,101,31,101,30,68,31,165,31,30,31,57,31,230,31,226,31,115,31,13,31,234,31,171,31,74,31,203,31,191,31,3,31,26,31,26,30,26,29,54,31,138,31,197,31,48,31,210,31,199,31,199,30,56,31,246,31,121,31,185,31,177,31,137,31,25,31,157,31,172,31,172,30,240,31,56,31,56,30,50,31,147,31,147,30,184,31,29,31,29,30,8,31,10,31,204,31,27,31,2,31,35,31,35,30,60,31,71,31,213,31,194,31,167,31,48,31,48,30,48,29,148,31,86,31,245,31,6,31,146,31,146,30,82,31,167,31,241,31,197,31,48,31,131,31,221,31,96,31,77,31,182,31,127,31,254,31,91,31,91,30,116,31,70,31,127,31,7,31,41,31,239,31,123,31,123,30,124,31,227,31,94,31,192,31,18,31,15,31,37,31,44,31,45,31,147,31,147,30,76,31,234,31,234,30,234,29,7,31,142,31,142,30,142,29,3,31,21,31,70,31,99,31,99,30,247,31,218,31,206,31,206,30,166,31,210,31,210,30,131,31,162,31,221,31,156,31,91,31,91,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
