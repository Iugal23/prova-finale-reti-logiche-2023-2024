-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_342 is
end project_tb_342;

architecture project_tb_arch_342 of project_tb_342 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 723;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (138,0,0,0,30,0,244,0,111,0,0,0,240,0,166,0,0,0,207,0,0,0,0,0,42,0,9,0,21,0,9,0,81,0,0,0,184,0,252,0,42,0,56,0,139,0,45,0,209,0,138,0,0,0,17,0,220,0,0,0,0,0,52,0,224,0,109,0,0,0,40,0,85,0,249,0,66,0,236,0,70,0,213,0,41,0,125,0,200,0,0,0,115,0,80,0,94,0,0,0,0,0,68,0,252,0,0,0,207,0,59,0,168,0,50,0,161,0,59,0,88,0,0,0,0,0,0,0,74,0,131,0,0,0,103,0,0,0,221,0,69,0,185,0,0,0,196,0,172,0,197,0,231,0,34,0,84,0,180,0,171,0,79,0,62,0,7,0,203,0,11,0,0,0,92,0,78,0,146,0,188,0,0,0,62,0,131,0,146,0,144,0,0,0,182,0,162,0,0,0,104,0,43,0,0,0,0,0,153,0,232,0,0,0,119,0,164,0,232,0,135,0,128,0,166,0,151,0,0,0,92,0,203,0,42,0,114,0,12,0,203,0,55,0,204,0,0,0,0,0,0,0,20,0,155,0,87,0,23,0,0,0,26,0,239,0,211,0,184,0,137,0,140,0,231,0,0,0,211,0,81,0,48,0,138,0,160,0,15,0,37,0,110,0,0,0,0,0,221,0,0,0,0,0,133,0,183,0,224,0,165,0,77,0,0,0,102,0,81,0,76,0,163,0,37,0,214,0,50,0,211,0,1,0,58,0,185,0,248,0,0,0,11,0,0,0,80,0,210,0,0,0,95,0,133,0,1,0,161,0,103,0,31,0,143,0,140,0,0,0,0,0,35,0,38,0,72,0,0,0,237,0,0,0,207,0,92,0,0,0,21,0,38,0,0,0,0,0,237,0,0,0,97,0,224,0,58,0,101,0,201,0,0,0,196,0,23,0,244,0,69,0,192,0,214,0,109,0,0,0,164,0,0,0,11,0,214,0,0,0,253,0,71,0,130,0,145,0,108,0,70,0,37,0,181,0,70,0,245,0,138,0,120,0,137,0,235,0,205,0,0,0,213,0,0,0,95,0,82,0,179,0,159,0,53,0,163,0,234,0,1,0,107,0,111,0,255,0,20,0,7,0,158,0,185,0,148,0,67,0,253,0,0,0,23,0,172,0,36,0,92,0,0,0,0,0,0,0,188,0,58,0,29,0,153,0,162,0,66,0,0,0,67,0,200,0,0,0,236,0,62,0,14,0,0,0,7,0,28,0,0,0,0,0,96,0,0,0,0,0,0,0,0,0,0,0,0,0,134,0,147,0,0,0,77,0,22,0,47,0,173,0,0,0,0,0,52,0,63,0,110,0,147,0,182,0,118,0,37,0,76,0,101,0,142,0,248,0,31,0,101,0,0,0,0,0,228,0,117,0,16,0,222,0,223,0,0,0,91,0,220,0,133,0,30,0,248,0,24,0,162,0,227,0,165,0,160,0,104,0,40,0,216,0,208,0,80,0,192,0,150,0,77,0,84,0,114,0,220,0,62,0,205,0,110,0,135,0,55,0,214,0,127,0,85,0,109,0,69,0,193,0,200,0,57,0,239,0,198,0,126,0,174,0,225,0,140,0,2,0,241,0,143,0,65,0,0,0,0,0,239,0,0,0,0,0,0,0,69,0,140,0,3,0,0,0,184,0,0,0,194,0,3,0,17,0,251,0,66,0,211,0,56,0,180,0,53,0,92,0,108,0,188,0,185,0,171,0,0,0,204,0,155,0,103,0,234,0,0,0,94,0,157,0,0,0,0,0,116,0,0,0,70,0,43,0,255,0,253,0,0,0,70,0,29,0,58,0,72,0,0,0,3,0,0,0,189,0,159,0,68,0,95,0,45,0,252,0,0,0,80,0,6,0,0,0,0,0,138,0,24,0,192,0,30,0,160,0,172,0,61,0,219,0,0,0,33,0,40,0,218,0,186,0,146,0,154,0,52,0,45,0,16,0,142,0,0,0,0,0,243,0,116,0,173,0,142,0,84,0,16,0,191,0,200,0,28,0,29,0,207,0,97,0,0,0,221,0,232,0,155,0,66,0,42,0,88,0,198,0,215,0,91,0,194,0,147,0,185,0,0,0,0,0,16,0,85,0,0,0,228,0,69,0,18,0,159,0,220,0,30,0,240,0,0,0,183,0,22,0,158,0,0,0,39,0,197,0,34,0,22,0,220,0,217,0,62,0,218,0,79,0,196,0,19,0,0,0,127,0,0,0,110,0,197,0,209,0,218,0,49,0,72,0,117,0,0,0,28,0,86,0,54,0,190,0,186,0,0,0,181,0,115,0,148,0,59,0,64,0,40,0,125,0,0,0,0,0,250,0,167,0,45,0,209,0,0,0,119,0,73,0,0,0,66,0,223,0,0,0,154,0,96,0,0,0,95,0,34,0,47,0,75,0,156,0,117,0,114,0,109,0,0,0,231,0,208,0,213,0,109,0,212,0,0,0,0,0,141,0,106,0,35,0,91,0,169,0,190,0,0,0,87,0,86,0,0,0,209,0,33,0,171,0,0,0,0,0,0,0,0,0,120,0,83,0,226,0,239,0,0,0,139,0,182,0,28,0,56,0,153,0,0,0,0,0,64,0,36,0,176,0,195,0,125,0,127,0,9,0,157,0,0,0,0,0,228,0,161,0,222,0,109,0,141,0,34,0,241,0,217,0,0,0,105,0,0,0,110,0,132,0,115,0,183,0,133,0,114,0,0,0,0,0,47,0,108,0,121,0,0,0,0,0,210,0,42,0,156,0,27,0,93,0,131,0,143,0,27,0,127,0,31,0,100,0,109,0,69,0,152,0,149,0,76,0,28,0,7,0,196,0,149,0,228,0,197,0,151,0,27,0,0,0,80,0,194,0,253,0,107,0,101,0,184,0,237,0,80,0,109,0,120,0,89,0,15,0,228,0,237,0,0,0,205,0,0,0,1,0,7,0,187,0,176,0,0,0,157,0,0,0,255,0,9,0,16,0,30,0,26,0,0,0,195,0,69,0,125,0,0,0,202,0,157,0,0,0,237,0,0,0,98,0,220,0,0,0,0,0,147,0,116,0,114,0,226,0,118,0,31,0,121,0,180,0,98,0,109,0,0,0,47,0,27,0,2,0,0,0,0,0,162,0,173,0,237,0,99,0,146,0,0,0,37,0,93,0,0,0,116,0,92,0,149,0,161,0,186,0,253,0,0,0,251,0,158,0,145,0,87,0,0,0,144,0);
signal scenario_full  : scenario_type := (138,31,138,30,30,31,244,31,111,31,111,30,240,31,166,31,166,30,207,31,207,30,207,29,42,31,9,31,21,31,9,31,81,31,81,30,184,31,252,31,42,31,56,31,139,31,45,31,209,31,138,31,138,30,17,31,220,31,220,30,220,29,52,31,224,31,109,31,109,30,40,31,85,31,249,31,66,31,236,31,70,31,213,31,41,31,125,31,200,31,200,30,115,31,80,31,94,31,94,30,94,29,68,31,252,31,252,30,207,31,59,31,168,31,50,31,161,31,59,31,88,31,88,30,88,29,88,28,74,31,131,31,131,30,103,31,103,30,221,31,69,31,185,31,185,30,196,31,172,31,197,31,231,31,34,31,84,31,180,31,171,31,79,31,62,31,7,31,203,31,11,31,11,30,92,31,78,31,146,31,188,31,188,30,62,31,131,31,146,31,144,31,144,30,182,31,162,31,162,30,104,31,43,31,43,30,43,29,153,31,232,31,232,30,119,31,164,31,232,31,135,31,128,31,166,31,151,31,151,30,92,31,203,31,42,31,114,31,12,31,203,31,55,31,204,31,204,30,204,29,204,28,20,31,155,31,87,31,23,31,23,30,26,31,239,31,211,31,184,31,137,31,140,31,231,31,231,30,211,31,81,31,48,31,138,31,160,31,15,31,37,31,110,31,110,30,110,29,221,31,221,30,221,29,133,31,183,31,224,31,165,31,77,31,77,30,102,31,81,31,76,31,163,31,37,31,214,31,50,31,211,31,1,31,58,31,185,31,248,31,248,30,11,31,11,30,80,31,210,31,210,30,95,31,133,31,1,31,161,31,103,31,31,31,143,31,140,31,140,30,140,29,35,31,38,31,72,31,72,30,237,31,237,30,207,31,92,31,92,30,21,31,38,31,38,30,38,29,237,31,237,30,97,31,224,31,58,31,101,31,201,31,201,30,196,31,23,31,244,31,69,31,192,31,214,31,109,31,109,30,164,31,164,30,11,31,214,31,214,30,253,31,71,31,130,31,145,31,108,31,70,31,37,31,181,31,70,31,245,31,138,31,120,31,137,31,235,31,205,31,205,30,213,31,213,30,95,31,82,31,179,31,159,31,53,31,163,31,234,31,1,31,107,31,111,31,255,31,20,31,7,31,158,31,185,31,148,31,67,31,253,31,253,30,23,31,172,31,36,31,92,31,92,30,92,29,92,28,188,31,58,31,29,31,153,31,162,31,66,31,66,30,67,31,200,31,200,30,236,31,62,31,14,31,14,30,7,31,28,31,28,30,28,29,96,31,96,30,96,29,96,28,96,27,96,26,96,25,134,31,147,31,147,30,77,31,22,31,47,31,173,31,173,30,173,29,52,31,63,31,110,31,147,31,182,31,118,31,37,31,76,31,101,31,142,31,248,31,31,31,101,31,101,30,101,29,228,31,117,31,16,31,222,31,223,31,223,30,91,31,220,31,133,31,30,31,248,31,24,31,162,31,227,31,165,31,160,31,104,31,40,31,216,31,208,31,80,31,192,31,150,31,77,31,84,31,114,31,220,31,62,31,205,31,110,31,135,31,55,31,214,31,127,31,85,31,109,31,69,31,193,31,200,31,57,31,239,31,198,31,126,31,174,31,225,31,140,31,2,31,241,31,143,31,65,31,65,30,65,29,239,31,239,30,239,29,239,28,69,31,140,31,3,31,3,30,184,31,184,30,194,31,3,31,17,31,251,31,66,31,211,31,56,31,180,31,53,31,92,31,108,31,188,31,185,31,171,31,171,30,204,31,155,31,103,31,234,31,234,30,94,31,157,31,157,30,157,29,116,31,116,30,70,31,43,31,255,31,253,31,253,30,70,31,29,31,58,31,72,31,72,30,3,31,3,30,189,31,159,31,68,31,95,31,45,31,252,31,252,30,80,31,6,31,6,30,6,29,138,31,24,31,192,31,30,31,160,31,172,31,61,31,219,31,219,30,33,31,40,31,218,31,186,31,146,31,154,31,52,31,45,31,16,31,142,31,142,30,142,29,243,31,116,31,173,31,142,31,84,31,16,31,191,31,200,31,28,31,29,31,207,31,97,31,97,30,221,31,232,31,155,31,66,31,42,31,88,31,198,31,215,31,91,31,194,31,147,31,185,31,185,30,185,29,16,31,85,31,85,30,228,31,69,31,18,31,159,31,220,31,30,31,240,31,240,30,183,31,22,31,158,31,158,30,39,31,197,31,34,31,22,31,220,31,217,31,62,31,218,31,79,31,196,31,19,31,19,30,127,31,127,30,110,31,197,31,209,31,218,31,49,31,72,31,117,31,117,30,28,31,86,31,54,31,190,31,186,31,186,30,181,31,115,31,148,31,59,31,64,31,40,31,125,31,125,30,125,29,250,31,167,31,45,31,209,31,209,30,119,31,73,31,73,30,66,31,223,31,223,30,154,31,96,31,96,30,95,31,34,31,47,31,75,31,156,31,117,31,114,31,109,31,109,30,231,31,208,31,213,31,109,31,212,31,212,30,212,29,141,31,106,31,35,31,91,31,169,31,190,31,190,30,87,31,86,31,86,30,209,31,33,31,171,31,171,30,171,29,171,28,171,27,120,31,83,31,226,31,239,31,239,30,139,31,182,31,28,31,56,31,153,31,153,30,153,29,64,31,36,31,176,31,195,31,125,31,127,31,9,31,157,31,157,30,157,29,228,31,161,31,222,31,109,31,141,31,34,31,241,31,217,31,217,30,105,31,105,30,110,31,132,31,115,31,183,31,133,31,114,31,114,30,114,29,47,31,108,31,121,31,121,30,121,29,210,31,42,31,156,31,27,31,93,31,131,31,143,31,27,31,127,31,31,31,100,31,109,31,69,31,152,31,149,31,76,31,28,31,7,31,196,31,149,31,228,31,197,31,151,31,27,31,27,30,80,31,194,31,253,31,107,31,101,31,184,31,237,31,80,31,109,31,120,31,89,31,15,31,228,31,237,31,237,30,205,31,205,30,1,31,7,31,187,31,176,31,176,30,157,31,157,30,255,31,9,31,16,31,30,31,26,31,26,30,195,31,69,31,125,31,125,30,202,31,157,31,157,30,237,31,237,30,98,31,220,31,220,30,220,29,147,31,116,31,114,31,226,31,118,31,31,31,121,31,180,31,98,31,109,31,109,30,47,31,27,31,2,31,2,30,2,29,162,31,173,31,237,31,99,31,146,31,146,30,37,31,93,31,93,30,116,31,92,31,149,31,161,31,186,31,253,31,253,30,251,31,158,31,145,31,87,31,87,30,144,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
