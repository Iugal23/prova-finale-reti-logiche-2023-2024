-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 909;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,210,0,132,0,124,0,0,0,69,0,83,0,24,0,129,0,197,0,0,0,206,0,121,0,33,0,50,0,0,0,0,0,23,0,204,0,28,0,194,0,146,0,247,0,0,0,0,0,182,0,25,0,163,0,9,0,239,0,0,0,230,0,31,0,144,0,166,0,233,0,13,0,0,0,70,0,31,0,157,0,171,0,106,0,255,0,81,0,72,0,153,0,199,0,85,0,0,0,204,0,35,0,6,0,33,0,21,0,0,0,7,0,30,0,246,0,219,0,179,0,181,0,170,0,75,0,152,0,96,0,95,0,0,0,0,0,66,0,31,0,79,0,172,0,121,0,46,0,36,0,172,0,147,0,245,0,163,0,204,0,2,0,79,0,0,0,234,0,68,0,76,0,154,0,0,0,140,0,113,0,120,0,244,0,0,0,150,0,93,0,206,0,49,0,126,0,240,0,37,0,71,0,22,0,231,0,0,0,0,0,239,0,115,0,190,0,246,0,223,0,159,0,55,0,74,0,98,0,80,0,137,0,46,0,0,0,0,0,0,0,67,0,0,0,167,0,217,0,0,0,186,0,162,0,59,0,77,0,74,0,35,0,122,0,41,0,107,0,0,0,0,0,220,0,0,0,76,0,0,0,4,0,0,0,80,0,238,0,219,0,62,0,123,0,62,0,0,0,94,0,0,0,80,0,95,0,0,0,0,0,105,0,247,0,148,0,109,0,172,0,193,0,149,0,168,0,104,0,136,0,98,0,179,0,57,0,119,0,252,0,2,0,33,0,174,0,240,0,0,0,39,0,0,0,4,0,147,0,70,0,27,0,158,0,156,0,109,0,166,0,234,0,0,0,243,0,184,0,188,0,109,0,0,0,89,0,0,0,0,0,0,0,68,0,30,0,0,0,0,0,120,0,250,0,35,0,182,0,0,0,69,0,79,0,0,0,81,0,164,0,0,0,105,0,242,0,15,0,223,0,206,0,117,0,105,0,191,0,0,0,0,0,0,0,163,0,144,0,181,0,131,0,236,0,233,0,132,0,170,0,187,0,0,0,49,0,167,0,67,0,136,0,227,0,121,0,144,0,44,0,43,0,30,0,0,0,30,0,0,0,40,0,147,0,145,0,0,0,20,0,133,0,18,0,59,0,169,0,53,0,142,0,196,0,50,0,229,0,0,0,136,0,82,0,148,0,203,0,140,0,58,0,236,0,237,0,221,0,189,0,63,0,160,0,32,0,197,0,216,0,215,0,243,0,1,0,0,0,237,0,190,0,233,0,0,0,102,0,0,0,83,0,1,0,40,0,49,0,35,0,0,0,54,0,92,0,210,0,184,0,29,0,216,0,0,0,187,0,111,0,0,0,65,0,16,0,0,0,147,0,0,0,209,0,144,0,0,0,23,0,64,0,231,0,44,0,21,0,0,0,34,0,127,0,0,0,100,0,249,0,0,0,153,0,36,0,6,0,171,0,0,0,41,0,240,0,81,0,236,0,0,0,8,0,27,0,49,0,174,0,39,0,207,0,67,0,0,0,69,0,57,0,227,0,0,0,103,0,0,0,45,0,220,0,16,0,147,0,123,0,237,0,80,0,212,0,0,0,80,0,204,0,220,0,239,0,11,0,0,0,51,0,3,0,0,0,0,0,93,0,181,0,213,0,161,0,108,0,93,0,174,0,169,0,0,0,0,0,135,0,0,0,253,0,251,0,89,0,0,0,62,0,9,0,116,0,0,0,0,0,37,0,67,0,98,0,181,0,74,0,136,0,242,0,206,0,253,0,123,0,0,0,70,0,0,0,0,0,68,0,163,0,69,0,0,0,147,0,0,0,0,0,55,0,145,0,107,0,130,0,47,0,161,0,55,0,0,0,0,0,33,0,173,0,44,0,215,0,0,0,195,0,1,0,199,0,31,0,127,0,107,0,192,0,153,0,200,0,194,0,0,0,237,0,221,0,0,0,146,0,10,0,38,0,234,0,174,0,111,0,242,0,94,0,245,0,0,0,227,0,0,0,67,0,0,0,229,0,29,0,169,0,114,0,7,0,159,0,225,0,226,0,0,0,141,0,21,0,0,0,134,0,47,0,101,0,97,0,0,0,182,0,100,0,158,0,80,0,183,0,158,0,162,0,14,0,8,0,0,0,0,0,7,0,155,0,0,0,181,0,199,0,146,0,100,0,0,0,183,0,66,0,112,0,47,0,228,0,0,0,0,0,167,0,0,0,62,0,0,0,100,0,0,0,6,0,116,0,5,0,0,0,110,0,104,0,0,0,185,0,128,0,86,0,0,0,73,0,236,0,246,0,164,0,232,0,150,0,163,0,0,0,201,0,0,0,84,0,112,0,105,0,0,0,0,0,20,0,168,0,112,0,32,0,0,0,111,0,0,0,168,0,174,0,134,0,0,0,81,0,0,0,131,0,105,0,0,0,0,0,146,0,0,0,135,0,30,0,139,0,201,0,193,0,233,0,0,0,216,0,39,0,119,0,227,0,0,0,102,0,121,0,84,0,229,0,235,0,44,0,97,0,98,0,131,0,248,0,185,0,13,0,152,0,0,0,35,0,64,0,50,0,238,0,77,0,107,0,6,0,124,0,225,0,206,0,75,0,241,0,237,0,236,0,185,0,78,0,12,0,206,0,62,0,129,0,45,0,61,0,0,0,202,0,194,0,146,0,109,0,19,0,182,0,193,0,124,0,41,0,170,0,173,0,199,0,64,0,232,0,55,0,0,0,107,0,0,0,113,0,66,0,124,0,6,0,208,0,113,0,252,0,238,0,171,0,13,0,123,0,95,0,150,0,218,0,252,0,164,0,175,0,161,0,122,0,253,0,0,0,179,0,78,0,226,0,0,0,255,0,94,0,94,0,0,0,0,0,0,0,0,0,148,0,127,0,0,0,144,0,194,0,0,0,2,0,197,0,197,0,110,0,89,0,0,0,0,0,130,0,96,0,21,0,22,0,0,0,28,0,212,0,67,0,0,0,38,0,90,0,11,0,241,0,0,0,0,0,174,0,4,0,54,0,186,0,15,0,1,0,0,0,113,0,163,0,118,0,81,0,170,0,0,0,137,0,214,0,2,0,155,0,117,0,192,0,189,0,38,0,14,0,130,0,144,0,200,0,54,0,0,0,84,0,127,0,0,0,95,0,0,0,158,0,22,0,20,0,246,0,72,0,0,0,0,0,202,0,0,0,0,0,0,0,0,0,153,0,136,0,163,0,0,0,25,0,136,0,253,0,0,0,62,0,34,0,101,0,103,0,0,0,0,0,216,0,172,0,0,0,171,0,0,0,208,0,30,0,220,0,23,0,0,0,130,0,195,0,90,0,120,0,69,0,42,0,245,0,67,0,128,0,47,0,29,0,0,0,150,0,184,0,0,0,0,0,0,0,67,0,128,0,0,0,0,0,62,0,44,0,146,0,174,0,166,0,86,0,133,0,118,0,239,0,103,0,0,0,217,0,37,0,24,0,180,0,84,0,20,0,0,0,0,0,237,0,47,0,0,0,122,0,219,0,77,0,166,0,0,0,128,0,227,0,159,0,0,0,201,0,113,0,184,0,206,0,157,0,0,0,142,0,109,0,37,0,0,0,0,0,101,0,0,0,60,0,0,0,65,0,0,0,253,0,113,0,0,0,0,0,0,0,90,0,0,0,26,0,236,0,104,0,177,0,33,0,41,0,246,0,172,0,201,0,64,0,184,0,220,0,248,0,79,0,49,0,60,0,0,0,0,0,196,0,174,0,0,0,226,0,161,0,61,0,206,0,52,0,206,0,38,0,82,0,210,0,51,0,248,0,246,0,233,0,36,0,121,0,179,0,238,0,48,0,29,0,237,0,157,0,95,0,0,0,0,0,66,0,170,0,184,0,16,0,31,0,29,0,0,0,216,0,179,0,0,0,119,0,169,0,23,0,21,0,24,0,20,0,0,0,238,0,3,0,115,0,109,0,193,0,0,0,111,0,0,0,97,0,127,0,0,0,134,0,61,0,190,0,67,0,0,0,223,0,0,0,117,0,94,0,200,0,0,0,197,0,201,0,224,0,136,0,33,0,150,0,73,0,205,0,20,0,124,0);
signal scenario_full  : scenario_type := (0,0,0,0,210,31,132,31,124,31,124,30,69,31,83,31,24,31,129,31,197,31,197,30,206,31,121,31,33,31,50,31,50,30,50,29,23,31,204,31,28,31,194,31,146,31,247,31,247,30,247,29,182,31,25,31,163,31,9,31,239,31,239,30,230,31,31,31,144,31,166,31,233,31,13,31,13,30,70,31,31,31,157,31,171,31,106,31,255,31,81,31,72,31,153,31,199,31,85,31,85,30,204,31,35,31,6,31,33,31,21,31,21,30,7,31,30,31,246,31,219,31,179,31,181,31,170,31,75,31,152,31,96,31,95,31,95,30,95,29,66,31,31,31,79,31,172,31,121,31,46,31,36,31,172,31,147,31,245,31,163,31,204,31,2,31,79,31,79,30,234,31,68,31,76,31,154,31,154,30,140,31,113,31,120,31,244,31,244,30,150,31,93,31,206,31,49,31,126,31,240,31,37,31,71,31,22,31,231,31,231,30,231,29,239,31,115,31,190,31,246,31,223,31,159,31,55,31,74,31,98,31,80,31,137,31,46,31,46,30,46,29,46,28,67,31,67,30,167,31,217,31,217,30,186,31,162,31,59,31,77,31,74,31,35,31,122,31,41,31,107,31,107,30,107,29,220,31,220,30,76,31,76,30,4,31,4,30,80,31,238,31,219,31,62,31,123,31,62,31,62,30,94,31,94,30,80,31,95,31,95,30,95,29,105,31,247,31,148,31,109,31,172,31,193,31,149,31,168,31,104,31,136,31,98,31,179,31,57,31,119,31,252,31,2,31,33,31,174,31,240,31,240,30,39,31,39,30,4,31,147,31,70,31,27,31,158,31,156,31,109,31,166,31,234,31,234,30,243,31,184,31,188,31,109,31,109,30,89,31,89,30,89,29,89,28,68,31,30,31,30,30,30,29,120,31,250,31,35,31,182,31,182,30,69,31,79,31,79,30,81,31,164,31,164,30,105,31,242,31,15,31,223,31,206,31,117,31,105,31,191,31,191,30,191,29,191,28,163,31,144,31,181,31,131,31,236,31,233,31,132,31,170,31,187,31,187,30,49,31,167,31,67,31,136,31,227,31,121,31,144,31,44,31,43,31,30,31,30,30,30,31,30,30,40,31,147,31,145,31,145,30,20,31,133,31,18,31,59,31,169,31,53,31,142,31,196,31,50,31,229,31,229,30,136,31,82,31,148,31,203,31,140,31,58,31,236,31,237,31,221,31,189,31,63,31,160,31,32,31,197,31,216,31,215,31,243,31,1,31,1,30,237,31,190,31,233,31,233,30,102,31,102,30,83,31,1,31,40,31,49,31,35,31,35,30,54,31,92,31,210,31,184,31,29,31,216,31,216,30,187,31,111,31,111,30,65,31,16,31,16,30,147,31,147,30,209,31,144,31,144,30,23,31,64,31,231,31,44,31,21,31,21,30,34,31,127,31,127,30,100,31,249,31,249,30,153,31,36,31,6,31,171,31,171,30,41,31,240,31,81,31,236,31,236,30,8,31,27,31,49,31,174,31,39,31,207,31,67,31,67,30,69,31,57,31,227,31,227,30,103,31,103,30,45,31,220,31,16,31,147,31,123,31,237,31,80,31,212,31,212,30,80,31,204,31,220,31,239,31,11,31,11,30,51,31,3,31,3,30,3,29,93,31,181,31,213,31,161,31,108,31,93,31,174,31,169,31,169,30,169,29,135,31,135,30,253,31,251,31,89,31,89,30,62,31,9,31,116,31,116,30,116,29,37,31,67,31,98,31,181,31,74,31,136,31,242,31,206,31,253,31,123,31,123,30,70,31,70,30,70,29,68,31,163,31,69,31,69,30,147,31,147,30,147,29,55,31,145,31,107,31,130,31,47,31,161,31,55,31,55,30,55,29,33,31,173,31,44,31,215,31,215,30,195,31,1,31,199,31,31,31,127,31,107,31,192,31,153,31,200,31,194,31,194,30,237,31,221,31,221,30,146,31,10,31,38,31,234,31,174,31,111,31,242,31,94,31,245,31,245,30,227,31,227,30,67,31,67,30,229,31,29,31,169,31,114,31,7,31,159,31,225,31,226,31,226,30,141,31,21,31,21,30,134,31,47,31,101,31,97,31,97,30,182,31,100,31,158,31,80,31,183,31,158,31,162,31,14,31,8,31,8,30,8,29,7,31,155,31,155,30,181,31,199,31,146,31,100,31,100,30,183,31,66,31,112,31,47,31,228,31,228,30,228,29,167,31,167,30,62,31,62,30,100,31,100,30,6,31,116,31,5,31,5,30,110,31,104,31,104,30,185,31,128,31,86,31,86,30,73,31,236,31,246,31,164,31,232,31,150,31,163,31,163,30,201,31,201,30,84,31,112,31,105,31,105,30,105,29,20,31,168,31,112,31,32,31,32,30,111,31,111,30,168,31,174,31,134,31,134,30,81,31,81,30,131,31,105,31,105,30,105,29,146,31,146,30,135,31,30,31,139,31,201,31,193,31,233,31,233,30,216,31,39,31,119,31,227,31,227,30,102,31,121,31,84,31,229,31,235,31,44,31,97,31,98,31,131,31,248,31,185,31,13,31,152,31,152,30,35,31,64,31,50,31,238,31,77,31,107,31,6,31,124,31,225,31,206,31,75,31,241,31,237,31,236,31,185,31,78,31,12,31,206,31,62,31,129,31,45,31,61,31,61,30,202,31,194,31,146,31,109,31,19,31,182,31,193,31,124,31,41,31,170,31,173,31,199,31,64,31,232,31,55,31,55,30,107,31,107,30,113,31,66,31,124,31,6,31,208,31,113,31,252,31,238,31,171,31,13,31,123,31,95,31,150,31,218,31,252,31,164,31,175,31,161,31,122,31,253,31,253,30,179,31,78,31,226,31,226,30,255,31,94,31,94,31,94,30,94,29,94,28,94,27,148,31,127,31,127,30,144,31,194,31,194,30,2,31,197,31,197,31,110,31,89,31,89,30,89,29,130,31,96,31,21,31,22,31,22,30,28,31,212,31,67,31,67,30,38,31,90,31,11,31,241,31,241,30,241,29,174,31,4,31,54,31,186,31,15,31,1,31,1,30,113,31,163,31,118,31,81,31,170,31,170,30,137,31,214,31,2,31,155,31,117,31,192,31,189,31,38,31,14,31,130,31,144,31,200,31,54,31,54,30,84,31,127,31,127,30,95,31,95,30,158,31,22,31,20,31,246,31,72,31,72,30,72,29,202,31,202,30,202,29,202,28,202,27,153,31,136,31,163,31,163,30,25,31,136,31,253,31,253,30,62,31,34,31,101,31,103,31,103,30,103,29,216,31,172,31,172,30,171,31,171,30,208,31,30,31,220,31,23,31,23,30,130,31,195,31,90,31,120,31,69,31,42,31,245,31,67,31,128,31,47,31,29,31,29,30,150,31,184,31,184,30,184,29,184,28,67,31,128,31,128,30,128,29,62,31,44,31,146,31,174,31,166,31,86,31,133,31,118,31,239,31,103,31,103,30,217,31,37,31,24,31,180,31,84,31,20,31,20,30,20,29,237,31,47,31,47,30,122,31,219,31,77,31,166,31,166,30,128,31,227,31,159,31,159,30,201,31,113,31,184,31,206,31,157,31,157,30,142,31,109,31,37,31,37,30,37,29,101,31,101,30,60,31,60,30,65,31,65,30,253,31,113,31,113,30,113,29,113,28,90,31,90,30,26,31,236,31,104,31,177,31,33,31,41,31,246,31,172,31,201,31,64,31,184,31,220,31,248,31,79,31,49,31,60,31,60,30,60,29,196,31,174,31,174,30,226,31,161,31,61,31,206,31,52,31,206,31,38,31,82,31,210,31,51,31,248,31,246,31,233,31,36,31,121,31,179,31,238,31,48,31,29,31,237,31,157,31,95,31,95,30,95,29,66,31,170,31,184,31,16,31,31,31,29,31,29,30,216,31,179,31,179,30,119,31,169,31,23,31,21,31,24,31,20,31,20,30,238,31,3,31,115,31,109,31,193,31,193,30,111,31,111,30,97,31,127,31,127,30,134,31,61,31,190,31,67,31,67,30,223,31,223,30,117,31,94,31,200,31,200,30,197,31,201,31,224,31,136,31,33,31,150,31,73,31,205,31,20,31,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
