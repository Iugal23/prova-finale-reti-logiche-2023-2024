-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_3 is
end project_tb_3;

architecture project_tb_arch_3 of project_tb_3 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 808;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,40,0,242,0,149,0,150,0,186,0,6,0,138,0,0,0,36,0,248,0,135,0,35,0,177,0,105,0,178,0,181,0,177,0,152,0,0,0,248,0,238,0,100,0,164,0,53,0,211,0,17,0,185,0,0,0,119,0,4,0,0,0,117,0,84,0,0,0,218,0,83,0,222,0,240,0,0,0,161,0,0,0,112,0,194,0,126,0,91,0,62,0,14,0,86,0,115,0,33,0,123,0,0,0,214,0,251,0,12,0,241,0,26,0,133,0,0,0,147,0,51,0,205,0,62,0,11,0,3,0,0,0,135,0,151,0,85,0,81,0,188,0,108,0,0,0,117,0,242,0,129,0,74,0,211,0,208,0,8,0,47,0,135,0,174,0,105,0,103,0,201,0,68,0,234,0,145,0,92,0,16,0,24,0,0,0,166,0,65,0,22,0,138,0,96,0,111,0,64,0,21,0,23,0,222,0,199,0,0,0,139,0,165,0,78,0,148,0,6,0,118,0,219,0,29,0,0,0,124,0,242,0,205,0,0,0,56,0,194,0,203,0,0,0,83,0,26,0,53,0,217,0,12,0,0,0,158,0,174,0,227,0,50,0,125,0,241,0,139,0,198,0,208,0,36,0,0,0,7,0,90,0,131,0,0,0,99,0,216,0,0,0,251,0,181,0,120,0,73,0,245,0,21,0,75,0,79,0,174,0,14,0,166,0,251,0,31,0,235,0,0,0,69,0,0,0,0,0,0,0,0,0,155,0,0,0,189,0,233,0,11,0,191,0,243,0,91,0,0,0,0,0,0,0,98,0,77,0,13,0,184,0,17,0,0,0,74,0,0,0,0,0,40,0,110,0,8,0,200,0,60,0,177,0,115,0,83,0,0,0,10,0,179,0,3,0,82,0,119,0,223,0,143,0,177,0,255,0,4,0,55,0,0,0,39,0,81,0,22,0,151,0,0,0,62,0,0,0,0,0,108,0,99,0,115,0,116,0,2,0,73,0,29,0,233,0,253,0,85,0,139,0,0,0,86,0,102,0,122,0,39,0,0,0,50,0,128,0,4,0,246,0,154,0,231,0,231,0,116,0,31,0,221,0,31,0,178,0,186,0,0,0,56,0,9,0,21,0,41,0,143,0,56,0,97,0,127,0,0,0,194,0,145,0,226,0,61,0,91,0,110,0,127,0,37,0,0,0,129,0,118,0,0,0,164,0,127,0,70,0,177,0,26,0,0,0,208,0,135,0,146,0,103,0,24,0,62,0,188,0,239,0,77,0,75,0,185,0,214,0,0,0,0,0,181,0,60,0,0,0,247,0,79,0,175,0,164,0,198,0,107,0,92,0,75,0,35,0,136,0,73,0,155,0,0,0,84,0,0,0,0,0,120,0,113,0,196,0,89,0,27,0,52,0,83,0,240,0,132,0,0,0,0,0,0,0,101,0,178,0,0,0,180,0,124,0,0,0,143,0,195,0,0,0,79,0,88,0,150,0,144,0,125,0,168,0,243,0,88,0,111,0,50,0,180,0,12,0,15,0,14,0,0,0,77,0,0,0,107,0,145,0,199,0,188,0,237,0,54,0,176,0,0,0,0,0,69,0,216,0,186,0,65,0,165,0,0,0,14,0,0,0,162,0,188,0,38,0,198,0,121,0,112,0,39,0,176,0,164,0,88,0,95,0,213,0,10,0,168,0,53,0,0,0,107,0,190,0,221,0,91,0,166,0,126,0,229,0,147,0,105,0,139,0,0,0,49,0,249,0,194,0,195,0,199,0,34,0,34,0,36,0,178,0,232,0,0,0,176,0,182,0,0,0,0,0,144,0,201,0,7,0,0,0,141,0,131,0,16,0,251,0,255,0,0,0,36,0,241,0,17,0,113,0,0,0,214,0,184,0,199,0,50,0,188,0,234,0,224,0,0,0,15,0,0,0,148,0,0,0,0,0,0,0,209,0,58,0,200,0,108,0,142,0,222,0,34,0,56,0,182,0,72,0,211,0,0,0,19,0,181,0,94,0,71,0,144,0,98,0,0,0,95,0,0,0,104,0,210,0,218,0,92,0,52,0,216,0,199,0,10,0,229,0,121,0,42,0,0,0,14,0,47,0,141,0,207,0,0,0,120,0,145,0,232,0,28,0,0,0,52,0,217,0,34,0,225,0,134,0,210,0,0,0,98,0,93,0,140,0,40,0,31,0,110,0,236,0,65,0,216,0,16,0,0,0,135,0,223,0,0,0,150,0,52,0,79,0,0,0,177,0,146,0,0,0,200,0,217,0,213,0,0,0,13,0,0,0,0,0,193,0,0,0,159,0,13,0,0,0,114,0,147,0,231,0,255,0,144,0,0,0,70,0,188,0,103,0,152,0,0,0,0,0,213,0,237,0,137,0,160,0,125,0,75,0,0,0,28,0,197,0,216,0,22,0,33,0,196,0,254,0,31,0,0,0,144,0,49,0,108,0,168,0,201,0,38,0,137,0,149,0,0,0,73,0,13,0,0,0,19,0,159,0,12,0,0,0,79,0,111,0,0,0,38,0,206,0,0,0,90,0,130,0,234,0,0,0,189,0,0,0,0,0,81,0,109,0,113,0,143,0,0,0,10,0,162,0,98,0,247,0,42,0,205,0,222,0,114,0,47,0,242,0,0,0,148,0,82,0,248,0,176,0,254,0,12,0,104,0,149,0,43,0,0,0,231,0,13,0,0,0,200,0,177,0,1,0,174,0,59,0,186,0,19,0,66,0,158,0,89,0,21,0,83,0,122,0,13,0,61,0,0,0,0,0,0,0,38,0,139,0,112,0,104,0,0,0,0,0,63,0,130,0,32,0,170,0,84,0,61,0,247,0,61,0,96,0,62,0,101,0,0,0,0,0,0,0,159,0,38,0,119,0,23,0,216,0,0,0,217,0,28,0,149,0,0,0,0,0,121,0,103,0,0,0,147,0,107,0,0,0,0,0,67,0,0,0,46,0,78,0,0,0,232,0,211,0,69,0,199,0,110,0,7,0,250,0,191,0,0,0,138,0,22,0,124,0,8,0,240,0,149,0,187,0,242,0,227,0,124,0,192,0,207,0,12,0,213,0,166,0,190,0,130,0,23,0,213,0,159,0,0,0,141,0,128,0,168,0,126,0,0,0,190,0,179,0,251,0,93,0,0,0,120,0,247,0,80,0,84,0,0,0,182,0,194,0,207,0,189,0,213,0,154,0,17,0,231,0,135,0,0,0,88,0,80,0,205,0,102,0,25,0,82,0,37,0,132,0,8,0,182,0,203,0,139,0,0,0,145,0,247,0,227,0,37,0,108,0,186,0,67,0,50,0,0,0,64,0,101,0,24,0,0,0,221,0,16,0,167,0,0,0,95,0,55,0,130,0,95,0,181,0,0,0,0,0,172,0,50,0,148,0,127,0,93,0,103,0,230,0,0,0,251,0,0,0,148,0,28,0,0,0,39,0,0,0,191,0,106,0,69,0,30,0,15,0,41,0,56,0,152,0,173,0,144,0,14,0,182,0,43,0,212,0,37,0,63,0,30,0,0,0,49,0,224,0,226,0,230,0,218,0,196,0,29,0,132,0,50,0,113,0,88,0,214,0,123,0,25,0,206,0,105,0,150,0,41,0,24,0,205,0);
signal scenario_full  : scenario_type := (0,0,40,31,242,31,149,31,150,31,186,31,6,31,138,31,138,30,36,31,248,31,135,31,35,31,177,31,105,31,178,31,181,31,177,31,152,31,152,30,248,31,238,31,100,31,164,31,53,31,211,31,17,31,185,31,185,30,119,31,4,31,4,30,117,31,84,31,84,30,218,31,83,31,222,31,240,31,240,30,161,31,161,30,112,31,194,31,126,31,91,31,62,31,14,31,86,31,115,31,33,31,123,31,123,30,214,31,251,31,12,31,241,31,26,31,133,31,133,30,147,31,51,31,205,31,62,31,11,31,3,31,3,30,135,31,151,31,85,31,81,31,188,31,108,31,108,30,117,31,242,31,129,31,74,31,211,31,208,31,8,31,47,31,135,31,174,31,105,31,103,31,201,31,68,31,234,31,145,31,92,31,16,31,24,31,24,30,166,31,65,31,22,31,138,31,96,31,111,31,64,31,21,31,23,31,222,31,199,31,199,30,139,31,165,31,78,31,148,31,6,31,118,31,219,31,29,31,29,30,124,31,242,31,205,31,205,30,56,31,194,31,203,31,203,30,83,31,26,31,53,31,217,31,12,31,12,30,158,31,174,31,227,31,50,31,125,31,241,31,139,31,198,31,208,31,36,31,36,30,7,31,90,31,131,31,131,30,99,31,216,31,216,30,251,31,181,31,120,31,73,31,245,31,21,31,75,31,79,31,174,31,14,31,166,31,251,31,31,31,235,31,235,30,69,31,69,30,69,29,69,28,69,27,155,31,155,30,189,31,233,31,11,31,191,31,243,31,91,31,91,30,91,29,91,28,98,31,77,31,13,31,184,31,17,31,17,30,74,31,74,30,74,29,40,31,110,31,8,31,200,31,60,31,177,31,115,31,83,31,83,30,10,31,179,31,3,31,82,31,119,31,223,31,143,31,177,31,255,31,4,31,55,31,55,30,39,31,81,31,22,31,151,31,151,30,62,31,62,30,62,29,108,31,99,31,115,31,116,31,2,31,73,31,29,31,233,31,253,31,85,31,139,31,139,30,86,31,102,31,122,31,39,31,39,30,50,31,128,31,4,31,246,31,154,31,231,31,231,31,116,31,31,31,221,31,31,31,178,31,186,31,186,30,56,31,9,31,21,31,41,31,143,31,56,31,97,31,127,31,127,30,194,31,145,31,226,31,61,31,91,31,110,31,127,31,37,31,37,30,129,31,118,31,118,30,164,31,127,31,70,31,177,31,26,31,26,30,208,31,135,31,146,31,103,31,24,31,62,31,188,31,239,31,77,31,75,31,185,31,214,31,214,30,214,29,181,31,60,31,60,30,247,31,79,31,175,31,164,31,198,31,107,31,92,31,75,31,35,31,136,31,73,31,155,31,155,30,84,31,84,30,84,29,120,31,113,31,196,31,89,31,27,31,52,31,83,31,240,31,132,31,132,30,132,29,132,28,101,31,178,31,178,30,180,31,124,31,124,30,143,31,195,31,195,30,79,31,88,31,150,31,144,31,125,31,168,31,243,31,88,31,111,31,50,31,180,31,12,31,15,31,14,31,14,30,77,31,77,30,107,31,145,31,199,31,188,31,237,31,54,31,176,31,176,30,176,29,69,31,216,31,186,31,65,31,165,31,165,30,14,31,14,30,162,31,188,31,38,31,198,31,121,31,112,31,39,31,176,31,164,31,88,31,95,31,213,31,10,31,168,31,53,31,53,30,107,31,190,31,221,31,91,31,166,31,126,31,229,31,147,31,105,31,139,31,139,30,49,31,249,31,194,31,195,31,199,31,34,31,34,31,36,31,178,31,232,31,232,30,176,31,182,31,182,30,182,29,144,31,201,31,7,31,7,30,141,31,131,31,16,31,251,31,255,31,255,30,36,31,241,31,17,31,113,31,113,30,214,31,184,31,199,31,50,31,188,31,234,31,224,31,224,30,15,31,15,30,148,31,148,30,148,29,148,28,209,31,58,31,200,31,108,31,142,31,222,31,34,31,56,31,182,31,72,31,211,31,211,30,19,31,181,31,94,31,71,31,144,31,98,31,98,30,95,31,95,30,104,31,210,31,218,31,92,31,52,31,216,31,199,31,10,31,229,31,121,31,42,31,42,30,14,31,47,31,141,31,207,31,207,30,120,31,145,31,232,31,28,31,28,30,52,31,217,31,34,31,225,31,134,31,210,31,210,30,98,31,93,31,140,31,40,31,31,31,110,31,236,31,65,31,216,31,16,31,16,30,135,31,223,31,223,30,150,31,52,31,79,31,79,30,177,31,146,31,146,30,200,31,217,31,213,31,213,30,13,31,13,30,13,29,193,31,193,30,159,31,13,31,13,30,114,31,147,31,231,31,255,31,144,31,144,30,70,31,188,31,103,31,152,31,152,30,152,29,213,31,237,31,137,31,160,31,125,31,75,31,75,30,28,31,197,31,216,31,22,31,33,31,196,31,254,31,31,31,31,30,144,31,49,31,108,31,168,31,201,31,38,31,137,31,149,31,149,30,73,31,13,31,13,30,19,31,159,31,12,31,12,30,79,31,111,31,111,30,38,31,206,31,206,30,90,31,130,31,234,31,234,30,189,31,189,30,189,29,81,31,109,31,113,31,143,31,143,30,10,31,162,31,98,31,247,31,42,31,205,31,222,31,114,31,47,31,242,31,242,30,148,31,82,31,248,31,176,31,254,31,12,31,104,31,149,31,43,31,43,30,231,31,13,31,13,30,200,31,177,31,1,31,174,31,59,31,186,31,19,31,66,31,158,31,89,31,21,31,83,31,122,31,13,31,61,31,61,30,61,29,61,28,38,31,139,31,112,31,104,31,104,30,104,29,63,31,130,31,32,31,170,31,84,31,61,31,247,31,61,31,96,31,62,31,101,31,101,30,101,29,101,28,159,31,38,31,119,31,23,31,216,31,216,30,217,31,28,31,149,31,149,30,149,29,121,31,103,31,103,30,147,31,107,31,107,30,107,29,67,31,67,30,46,31,78,31,78,30,232,31,211,31,69,31,199,31,110,31,7,31,250,31,191,31,191,30,138,31,22,31,124,31,8,31,240,31,149,31,187,31,242,31,227,31,124,31,192,31,207,31,12,31,213,31,166,31,190,31,130,31,23,31,213,31,159,31,159,30,141,31,128,31,168,31,126,31,126,30,190,31,179,31,251,31,93,31,93,30,120,31,247,31,80,31,84,31,84,30,182,31,194,31,207,31,189,31,213,31,154,31,17,31,231,31,135,31,135,30,88,31,80,31,205,31,102,31,25,31,82,31,37,31,132,31,8,31,182,31,203,31,139,31,139,30,145,31,247,31,227,31,37,31,108,31,186,31,67,31,50,31,50,30,64,31,101,31,24,31,24,30,221,31,16,31,167,31,167,30,95,31,55,31,130,31,95,31,181,31,181,30,181,29,172,31,50,31,148,31,127,31,93,31,103,31,230,31,230,30,251,31,251,30,148,31,28,31,28,30,39,31,39,30,191,31,106,31,69,31,30,31,15,31,41,31,56,31,152,31,173,31,144,31,14,31,182,31,43,31,212,31,37,31,63,31,30,31,30,30,49,31,224,31,226,31,230,31,218,31,196,31,29,31,132,31,50,31,113,31,88,31,214,31,123,31,25,31,206,31,105,31,150,31,41,31,24,31,205,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
