-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_854 is
end project_tb_854;

architecture project_tb_arch_854 of project_tb_854 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 392;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (99,0,103,0,48,0,0,0,177,0,0,0,192,0,226,0,132,0,7,0,255,0,141,0,44,0,86,0,186,0,88,0,38,0,70,0,112,0,0,0,185,0,57,0,65,0,150,0,214,0,74,0,172,0,162,0,84,0,84,0,0,0,0,0,170,0,84,0,26,0,104,0,5,0,198,0,206,0,93,0,153,0,0,0,0,0,29,0,32,0,33,0,155,0,177,0,118,0,56,0,218,0,0,0,0,0,146,0,142,0,217,0,250,0,216,0,161,0,54,0,217,0,156,0,93,0,43,0,129,0,75,0,0,0,16,0,12,0,184,0,76,0,242,0,112,0,16,0,0,0,93,0,0,0,95,0,255,0,130,0,229,0,1,0,150,0,0,0,124,0,185,0,17,0,53,0,32,0,0,0,180,0,0,0,106,0,0,0,0,0,0,0,96,0,179,0,0,0,155,0,41,0,239,0,110,0,215,0,68,0,0,0,0,0,12,0,154,0,121,0,0,0,85,0,227,0,38,0,248,0,0,0,1,0,253,0,76,0,208,0,172,0,0,0,69,0,162,0,94,0,81,0,4,0,87,0,107,0,134,0,35,0,0,0,5,0,252,0,65,0,48,0,30,0,66,0,0,0,0,0,250,0,6,0,8,0,201,0,9,0,214,0,236,0,65,0,138,0,244,0,250,0,64,0,3,0,78,0,0,0,0,0,0,0,0,0,81,0,71,0,24,0,29,0,137,0,235,0,185,0,131,0,183,0,43,0,201,0,119,0,83,0,161,0,37,0,0,0,156,0,121,0,130,0,1,0,25,0,102,0,211,0,136,0,125,0,176,0,139,0,42,0,222,0,0,0,119,0,253,0,77,0,74,0,166,0,227,0,14,0,141,0,123,0,186,0,54,0,126,0,0,0,238,0,230,0,52,0,254,0,0,0,165,0,4,0,39,0,30,0,220,0,208,0,102,0,0,0,144,0,50,0,116,0,218,0,132,0,106,0,140,0,0,0,39,0,75,0,198,0,31,0,12,0,227,0,254,0,69,0,91,0,81,0,0,0,155,0,0,0,147,0,0,0,211,0,36,0,14,0,54,0,31,0,36,0,242,0,40,0,0,0,30,0,212,0,181,0,19,0,252,0,125,0,0,0,0,0,113,0,244,0,209,0,135,0,37,0,49,0,216,0,199,0,9,0,0,0,129,0,84,0,0,0,229,0,0,0,48,0,33,0,171,0,43,0,0,0,74,0,76,0,0,0,174,0,143,0,164,0,106,0,0,0,59,0,34,0,137,0,0,0,11,0,13,0,1,0,82,0,129,0,168,0,128,0,116,0,56,0,194,0,0,0,50,0,138,0,6,0,109,0,73,0,0,0,255,0,61,0,25,0,137,0,176,0,219,0,119,0,94,0,50,0,0,0,0,0,204,0,0,0,135,0,233,0,198,0,149,0,182,0,0,0,0,0,0,0,226,0,73,0,55,0,110,0,161,0,0,0,40,0,46,0,180,0,206,0,0,0,120,0,17,0,0,0,34,0,61,0,0,0,120,0,180,0,85,0,4,0,249,0,95,0,111,0,28,0,0,0,179,0,134,0,106,0,108,0,0,0,111,0,8,0,10,0,0,0,0,0,49,0,223,0,216,0,82,0,85,0,0,0,25,0,160,0,252,0,204,0,171,0,130,0,0,0,0,0,0,0,42,0,0,0,147,0,0,0,199,0,75,0,134,0,0,0,11,0,69,0,91,0,174,0,62,0,137,0,8,0,57,0,11,0);
signal scenario_full  : scenario_type := (99,31,103,31,48,31,48,30,177,31,177,30,192,31,226,31,132,31,7,31,255,31,141,31,44,31,86,31,186,31,88,31,38,31,70,31,112,31,112,30,185,31,57,31,65,31,150,31,214,31,74,31,172,31,162,31,84,31,84,31,84,30,84,29,170,31,84,31,26,31,104,31,5,31,198,31,206,31,93,31,153,31,153,30,153,29,29,31,32,31,33,31,155,31,177,31,118,31,56,31,218,31,218,30,218,29,146,31,142,31,217,31,250,31,216,31,161,31,54,31,217,31,156,31,93,31,43,31,129,31,75,31,75,30,16,31,12,31,184,31,76,31,242,31,112,31,16,31,16,30,93,31,93,30,95,31,255,31,130,31,229,31,1,31,150,31,150,30,124,31,185,31,17,31,53,31,32,31,32,30,180,31,180,30,106,31,106,30,106,29,106,28,96,31,179,31,179,30,155,31,41,31,239,31,110,31,215,31,68,31,68,30,68,29,12,31,154,31,121,31,121,30,85,31,227,31,38,31,248,31,248,30,1,31,253,31,76,31,208,31,172,31,172,30,69,31,162,31,94,31,81,31,4,31,87,31,107,31,134,31,35,31,35,30,5,31,252,31,65,31,48,31,30,31,66,31,66,30,66,29,250,31,6,31,8,31,201,31,9,31,214,31,236,31,65,31,138,31,244,31,250,31,64,31,3,31,78,31,78,30,78,29,78,28,78,27,81,31,71,31,24,31,29,31,137,31,235,31,185,31,131,31,183,31,43,31,201,31,119,31,83,31,161,31,37,31,37,30,156,31,121,31,130,31,1,31,25,31,102,31,211,31,136,31,125,31,176,31,139,31,42,31,222,31,222,30,119,31,253,31,77,31,74,31,166,31,227,31,14,31,141,31,123,31,186,31,54,31,126,31,126,30,238,31,230,31,52,31,254,31,254,30,165,31,4,31,39,31,30,31,220,31,208,31,102,31,102,30,144,31,50,31,116,31,218,31,132,31,106,31,140,31,140,30,39,31,75,31,198,31,31,31,12,31,227,31,254,31,69,31,91,31,81,31,81,30,155,31,155,30,147,31,147,30,211,31,36,31,14,31,54,31,31,31,36,31,242,31,40,31,40,30,30,31,212,31,181,31,19,31,252,31,125,31,125,30,125,29,113,31,244,31,209,31,135,31,37,31,49,31,216,31,199,31,9,31,9,30,129,31,84,31,84,30,229,31,229,30,48,31,33,31,171,31,43,31,43,30,74,31,76,31,76,30,174,31,143,31,164,31,106,31,106,30,59,31,34,31,137,31,137,30,11,31,13,31,1,31,82,31,129,31,168,31,128,31,116,31,56,31,194,31,194,30,50,31,138,31,6,31,109,31,73,31,73,30,255,31,61,31,25,31,137,31,176,31,219,31,119,31,94,31,50,31,50,30,50,29,204,31,204,30,135,31,233,31,198,31,149,31,182,31,182,30,182,29,182,28,226,31,73,31,55,31,110,31,161,31,161,30,40,31,46,31,180,31,206,31,206,30,120,31,17,31,17,30,34,31,61,31,61,30,120,31,180,31,85,31,4,31,249,31,95,31,111,31,28,31,28,30,179,31,134,31,106,31,108,31,108,30,111,31,8,31,10,31,10,30,10,29,49,31,223,31,216,31,82,31,85,31,85,30,25,31,160,31,252,31,204,31,171,31,130,31,130,30,130,29,130,28,42,31,42,30,147,31,147,30,199,31,75,31,134,31,134,30,11,31,69,31,91,31,174,31,62,31,137,31,8,31,57,31,11,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
