-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 781;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (22,0,64,0,0,0,107,0,0,0,137,0,0,0,29,0,159,0,32,0,164,0,216,0,241,0,90,0,62,0,121,0,233,0,149,0,0,0,204,0,95,0,187,0,8,0,172,0,147,0,0,0,40,0,113,0,1,0,254,0,56,0,0,0,125,0,60,0,34,0,37,0,106,0,0,0,163,0,208,0,10,0,99,0,91,0,60,0,48,0,251,0,19,0,21,0,243,0,64,0,124,0,172,0,243,0,52,0,0,0,241,0,218,0,20,0,76,0,93,0,190,0,78,0,0,0,214,0,54,0,58,0,0,0,189,0,229,0,197,0,13,0,124,0,201,0,48,0,204,0,123,0,105,0,176,0,0,0,0,0,0,0,64,0,219,0,144,0,198,0,87,0,0,0,13,0,152,0,0,0,121,0,0,0,0,0,0,0,0,0,155,0,77,0,204,0,130,0,252,0,107,0,80,0,230,0,211,0,80,0,116,0,0,0,47,0,122,0,123,0,173,0,0,0,196,0,118,0,127,0,210,0,0,0,105,0,136,0,0,0,142,0,14,0,98,0,190,0,73,0,71,0,154,0,205,0,0,0,254,0,231,0,50,0,7,0,149,0,157,0,6,0,102,0,53,0,0,0,0,0,237,0,34,0,0,0,0,0,38,0,199,0,49,0,0,0,229,0,196,0,213,0,89,0,220,0,54,0,168,0,0,0,152,0,25,0,186,0,0,0,127,0,25,0,223,0,20,0,6,0,238,0,154,0,3,0,195,0,37,0,243,0,198,0,174,0,198,0,232,0,0,0,22,0,113,0,128,0,200,0,180,0,0,0,0,0,69,0,227,0,230,0,19,0,174,0,0,0,0,0,166,0,194,0,210,0,79,0,58,0,97,0,135,0,92,0,250,0,0,0,28,0,77,0,223,0,0,0,146,0,182,0,224,0,0,0,144,0,55,0,106,0,40,0,0,0,91,0,81,0,52,0,75,0,171,0,71,0,206,0,162,0,97,0,131,0,184,0,177,0,50,0,131,0,0,0,178,0,119,0,15,0,192,0,0,0,46,0,131,0,0,0,0,0,46,0,90,0,57,0,159,0,226,0,39,0,95,0,0,0,211,0,226,0,167,0,99,0,226,0,19,0,67,0,14,0,34,0,107,0,0,0,226,0,0,0,106,0,20,0,0,0,152,0,248,0,179,0,118,0,84,0,0,0,198,0,229,0,149,0,94,0,138,0,76,0,0,0,247,0,175,0,127,0,27,0,0,0,176,0,0,0,152,0,0,0,142,0,212,0,141,0,230,0,101,0,0,0,0,0,225,0,104,0,141,0,20,0,47,0,252,0,92,0,225,0,38,0,242,0,60,0,199,0,125,0,121,0,92,0,140,0,248,0,0,0,221,0,119,0,47,0,154,0,23,0,11,0,254,0,169,0,116,0,0,0,0,0,151,0,123,0,0,0,0,0,35,0,159,0,173,0,163,0,241,0,0,0,0,0,229,0,61,0,216,0,169,0,165,0,117,0,0,0,129,0,0,0,203,0,35,0,0,0,0,0,197,0,103,0,0,0,139,0,67,0,4,0,164,0,201,0,48,0,62,0,43,0,57,0,0,0,180,0,0,0,0,0,185,0,197,0,136,0,113,0,229,0,3,0,190,0,63,0,203,0,213,0,0,0,246,0,32,0,164,0,0,0,214,0,0,0,167,0,46,0,0,0,4,0,226,0,183,0,0,0,76,0,144,0,33,0,72,0,23,0,13,0,0,0,168,0,0,0,209,0,0,0,182,0,87,0,215,0,101,0,0,0,228,0,5,0,192,0,0,0,16,0,95,0,65,0,0,0,60,0,136,0,4,0,138,0,205,0,218,0,181,0,131,0,64,0,41,0,219,0,150,0,0,0,253,0,213,0,59,0,181,0,162,0,135,0,64,0,0,0,251,0,28,0,66,0,0,0,153,0,201,0,0,0,205,0,29,0,110,0,192,0,166,0,106,0,0,0,159,0,0,0,4,0,152,0,219,0,0,0,217,0,1,0,0,0,250,0,29,0,48,0,122,0,126,0,94,0,8,0,103,0,117,0,12,0,133,0,69,0,33,0,0,0,122,0,44,0,253,0,196,0,190,0,138,0,14,0,154,0,149,0,125,0,208,0,133,0,0,0,0,0,41,0,209,0,22,0,0,0,84,0,194,0,144,0,73,0,185,0,25,0,79,0,93,0,112,0,196,0,200,0,223,0,0,0,109,0,247,0,53,0,80,0,124,0,0,0,114,0,228,0,19,0,39,0,119,0,81,0,238,0,155,0,61,0,13,0,66,0,91,0,225,0,99,0,177,0,0,0,213,0,0,0,0,0,103,0,0,0,30,0,148,0,0,0,231,0,0,0,176,0,150,0,66,0,0,0,251,0,0,0,172,0,98,0,145,0,14,0,0,0,151,0,66,0,58,0,0,0,175,0,65,0,211,0,18,0,36,0,63,0,150,0,109,0,112,0,244,0,0,0,233,0,9,0,28,0,185,0,62,0,0,0,102,0,65,0,0,0,24,0,132,0,218,0,0,0,1,0,0,0,0,0,162,0,0,0,79,0,230,0,209,0,231,0,38,0,0,0,0,0,4,0,200,0,0,0,0,0,0,0,132,0,72,0,219,0,50,0,6,0,232,0,127,0,121,0,125,0,156,0,36,0,0,0,112,0,206,0,58,0,0,0,100,0,132,0,5,0,114,0,0,0,100,0,202,0,30,0,209,0,140,0,93,0,0,0,166,0,52,0,62,0,92,0,109,0,121,0,212,0,80,0,103,0,39,0,30,0,96,0,0,0,0,0,0,0,0,0,20,0,246,0,3,0,103,0,142,0,240,0,85,0,179,0,54,0,74,0,188,0,42,0,83,0,135,0,20,0,237,0,27,0,196,0,83,0,199,0,101,0,0,0,253,0,0,0,0,0,18,0,65,0,228,0,191,0,251,0,6,0,68,0,27,0,0,0,0,0,0,0,106,0,85,0,167,0,22,0,133,0,155,0,62,0,0,0,61,0,114,0,180,0,0,0,231,0,249,0,0,0,95,0,0,0,80,0,31,0,71,0,3,0,62,0,79,0,72,0,139,0,201,0,0,0,189,0,147,0,176,0,247,0,188,0,0,0,0,0,0,0,14,0,134,0,148,0,0,0,165,0,176,0,87,0,64,0,151,0,162,0,0,0,42,0,0,0,110,0,253,0,140,0,40,0,164,0,66,0,98,0,99,0,165,0,138,0,0,0,236,0,0,0,200,0,68,0,207,0,49,0,116,0,171,0,222,0,75,0,156,0,68,0,98,0,25,0,89,0,210,0,182,0,71,0,234,0,197,0,0,0,67,0,85,0,248,0,41,0,153,0,220,0,86,0,136,0,85,0,19,0,26,0,224,0,0,0,170,0,120,0,0,0,253,0,51,0,176,0,120,0,0,0,0,0,107,0,44,0,124,0,111,0,0,0,185,0,158,0,211,0,150,0,154,0,204,0,73,0,0,0,206,0,44,0);
signal scenario_full  : scenario_type := (22,31,64,31,64,30,107,31,107,30,137,31,137,30,29,31,159,31,32,31,164,31,216,31,241,31,90,31,62,31,121,31,233,31,149,31,149,30,204,31,95,31,187,31,8,31,172,31,147,31,147,30,40,31,113,31,1,31,254,31,56,31,56,30,125,31,60,31,34,31,37,31,106,31,106,30,163,31,208,31,10,31,99,31,91,31,60,31,48,31,251,31,19,31,21,31,243,31,64,31,124,31,172,31,243,31,52,31,52,30,241,31,218,31,20,31,76,31,93,31,190,31,78,31,78,30,214,31,54,31,58,31,58,30,189,31,229,31,197,31,13,31,124,31,201,31,48,31,204,31,123,31,105,31,176,31,176,30,176,29,176,28,64,31,219,31,144,31,198,31,87,31,87,30,13,31,152,31,152,30,121,31,121,30,121,29,121,28,121,27,155,31,77,31,204,31,130,31,252,31,107,31,80,31,230,31,211,31,80,31,116,31,116,30,47,31,122,31,123,31,173,31,173,30,196,31,118,31,127,31,210,31,210,30,105,31,136,31,136,30,142,31,14,31,98,31,190,31,73,31,71,31,154,31,205,31,205,30,254,31,231,31,50,31,7,31,149,31,157,31,6,31,102,31,53,31,53,30,53,29,237,31,34,31,34,30,34,29,38,31,199,31,49,31,49,30,229,31,196,31,213,31,89,31,220,31,54,31,168,31,168,30,152,31,25,31,186,31,186,30,127,31,25,31,223,31,20,31,6,31,238,31,154,31,3,31,195,31,37,31,243,31,198,31,174,31,198,31,232,31,232,30,22,31,113,31,128,31,200,31,180,31,180,30,180,29,69,31,227,31,230,31,19,31,174,31,174,30,174,29,166,31,194,31,210,31,79,31,58,31,97,31,135,31,92,31,250,31,250,30,28,31,77,31,223,31,223,30,146,31,182,31,224,31,224,30,144,31,55,31,106,31,40,31,40,30,91,31,81,31,52,31,75,31,171,31,71,31,206,31,162,31,97,31,131,31,184,31,177,31,50,31,131,31,131,30,178,31,119,31,15,31,192,31,192,30,46,31,131,31,131,30,131,29,46,31,90,31,57,31,159,31,226,31,39,31,95,31,95,30,211,31,226,31,167,31,99,31,226,31,19,31,67,31,14,31,34,31,107,31,107,30,226,31,226,30,106,31,20,31,20,30,152,31,248,31,179,31,118,31,84,31,84,30,198,31,229,31,149,31,94,31,138,31,76,31,76,30,247,31,175,31,127,31,27,31,27,30,176,31,176,30,152,31,152,30,142,31,212,31,141,31,230,31,101,31,101,30,101,29,225,31,104,31,141,31,20,31,47,31,252,31,92,31,225,31,38,31,242,31,60,31,199,31,125,31,121,31,92,31,140,31,248,31,248,30,221,31,119,31,47,31,154,31,23,31,11,31,254,31,169,31,116,31,116,30,116,29,151,31,123,31,123,30,123,29,35,31,159,31,173,31,163,31,241,31,241,30,241,29,229,31,61,31,216,31,169,31,165,31,117,31,117,30,129,31,129,30,203,31,35,31,35,30,35,29,197,31,103,31,103,30,139,31,67,31,4,31,164,31,201,31,48,31,62,31,43,31,57,31,57,30,180,31,180,30,180,29,185,31,197,31,136,31,113,31,229,31,3,31,190,31,63,31,203,31,213,31,213,30,246,31,32,31,164,31,164,30,214,31,214,30,167,31,46,31,46,30,4,31,226,31,183,31,183,30,76,31,144,31,33,31,72,31,23,31,13,31,13,30,168,31,168,30,209,31,209,30,182,31,87,31,215,31,101,31,101,30,228,31,5,31,192,31,192,30,16,31,95,31,65,31,65,30,60,31,136,31,4,31,138,31,205,31,218,31,181,31,131,31,64,31,41,31,219,31,150,31,150,30,253,31,213,31,59,31,181,31,162,31,135,31,64,31,64,30,251,31,28,31,66,31,66,30,153,31,201,31,201,30,205,31,29,31,110,31,192,31,166,31,106,31,106,30,159,31,159,30,4,31,152,31,219,31,219,30,217,31,1,31,1,30,250,31,29,31,48,31,122,31,126,31,94,31,8,31,103,31,117,31,12,31,133,31,69,31,33,31,33,30,122,31,44,31,253,31,196,31,190,31,138,31,14,31,154,31,149,31,125,31,208,31,133,31,133,30,133,29,41,31,209,31,22,31,22,30,84,31,194,31,144,31,73,31,185,31,25,31,79,31,93,31,112,31,196,31,200,31,223,31,223,30,109,31,247,31,53,31,80,31,124,31,124,30,114,31,228,31,19,31,39,31,119,31,81,31,238,31,155,31,61,31,13,31,66,31,91,31,225,31,99,31,177,31,177,30,213,31,213,30,213,29,103,31,103,30,30,31,148,31,148,30,231,31,231,30,176,31,150,31,66,31,66,30,251,31,251,30,172,31,98,31,145,31,14,31,14,30,151,31,66,31,58,31,58,30,175,31,65,31,211,31,18,31,36,31,63,31,150,31,109,31,112,31,244,31,244,30,233,31,9,31,28,31,185,31,62,31,62,30,102,31,65,31,65,30,24,31,132,31,218,31,218,30,1,31,1,30,1,29,162,31,162,30,79,31,230,31,209,31,231,31,38,31,38,30,38,29,4,31,200,31,200,30,200,29,200,28,132,31,72,31,219,31,50,31,6,31,232,31,127,31,121,31,125,31,156,31,36,31,36,30,112,31,206,31,58,31,58,30,100,31,132,31,5,31,114,31,114,30,100,31,202,31,30,31,209,31,140,31,93,31,93,30,166,31,52,31,62,31,92,31,109,31,121,31,212,31,80,31,103,31,39,31,30,31,96,31,96,30,96,29,96,28,96,27,20,31,246,31,3,31,103,31,142,31,240,31,85,31,179,31,54,31,74,31,188,31,42,31,83,31,135,31,20,31,237,31,27,31,196,31,83,31,199,31,101,31,101,30,253,31,253,30,253,29,18,31,65,31,228,31,191,31,251,31,6,31,68,31,27,31,27,30,27,29,27,28,106,31,85,31,167,31,22,31,133,31,155,31,62,31,62,30,61,31,114,31,180,31,180,30,231,31,249,31,249,30,95,31,95,30,80,31,31,31,71,31,3,31,62,31,79,31,72,31,139,31,201,31,201,30,189,31,147,31,176,31,247,31,188,31,188,30,188,29,188,28,14,31,134,31,148,31,148,30,165,31,176,31,87,31,64,31,151,31,162,31,162,30,42,31,42,30,110,31,253,31,140,31,40,31,164,31,66,31,98,31,99,31,165,31,138,31,138,30,236,31,236,30,200,31,68,31,207,31,49,31,116,31,171,31,222,31,75,31,156,31,68,31,98,31,25,31,89,31,210,31,182,31,71,31,234,31,197,31,197,30,67,31,85,31,248,31,41,31,153,31,220,31,86,31,136,31,85,31,19,31,26,31,224,31,224,30,170,31,120,31,120,30,253,31,51,31,176,31,120,31,120,30,120,29,107,31,44,31,124,31,111,31,111,30,185,31,158,31,211,31,150,31,154,31,204,31,73,31,73,30,206,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
