-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 822;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (30,0,0,0,155,0,243,0,240,0,143,0,0,0,118,0,0,0,23,0,216,0,77,0,73,0,11,0,0,0,55,0,93,0,183,0,83,0,250,0,0,0,0,0,84,0,160,0,226,0,15,0,70,0,155,0,66,0,91,0,212,0,0,0,0,0,0,0,96,0,125,0,234,0,0,0,39,0,244,0,148,0,79,0,107,0,119,0,0,0,162,0,157,0,0,0,0,0,144,0,245,0,132,0,0,0,159,0,222,0,160,0,83,0,95,0,252,0,0,0,61,0,214,0,0,0,12,0,149,0,0,0,169,0,163,0,255,0,52,0,23,0,246,0,0,0,170,0,3,0,62,0,17,0,12,0,38,0,146,0,72,0,19,0,0,0,16,0,103,0,154,0,137,0,21,0,4,0,131,0,126,0,241,0,125,0,153,0,36,0,14,0,0,0,235,0,248,0,127,0,147,0,255,0,251,0,233,0,80,0,0,0,174,0,143,0,94,0,38,0,0,0,143,0,178,0,144,0,171,0,98,0,247,0,240,0,30,0,0,0,236,0,13,0,0,0,159,0,229,0,136,0,0,0,162,0,86,0,208,0,173,0,13,0,168,0,115,0,27,0,154,0,0,0,40,0,60,0,65,0,0,0,23,0,170,0,110,0,0,0,161,0,162,0,5,0,44,0,184,0,0,0,150,0,0,0,123,0,198,0,254,0,174,0,0,0,122,0,110,0,0,0,20,0,9,0,0,0,201,0,180,0,180,0,156,0,160,0,4,0,118,0,35,0,135,0,85,0,0,0,61,0,93,0,250,0,221,0,155,0,146,0,0,0,38,0,130,0,219,0,152,0,96,0,166,0,191,0,0,0,219,0,187,0,127,0,0,0,0,0,46,0,49,0,135,0,223,0,0,0,70,0,16,0,139,0,36,0,221,0,168,0,61,0,157,0,0,0,17,0,69,0,222,0,36,0,22,0,8,0,238,0,104,0,122,0,195,0,181,0,167,0,46,0,144,0,202,0,109,0,115,0,23,0,113,0,0,0,72,0,37,0,30,0,132,0,0,0,0,0,242,0,48,0,236,0,130,0,88,0,187,0,0,0,231,0,237,0,188,0,219,0,0,0,92,0,130,0,3,0,20,0,238,0,0,0,110,0,243,0,52,0,134,0,0,0,185,0,4,0,191,0,8,0,0,0,236,0,132,0,199,0,19,0,0,0,133,0,72,0,250,0,187,0,97,0,0,0,183,0,77,0,12,0,0,0,114,0,129,0,11,0,251,0,87,0,56,0,53,0,231,0,0,0,73,0,252,0,130,0,118,0,0,0,242,0,54,0,50,0,229,0,185,0,173,0,4,0,136,0,0,0,8,0,153,0,118,0,64,0,203,0,2,0,0,0,101,0,54,0,104,0,116,0,92,0,249,0,81,0,141,0,0,0,126,0,69,0,0,0,98,0,16,0,177,0,173,0,0,0,81,0,0,0,120,0,82,0,28,0,205,0,228,0,199,0,0,0,154,0,250,0,0,0,165,0,109,0,241,0,6,0,214,0,121,0,217,0,154,0,35,0,0,0,16,0,0,0,165,0,239,0,0,0,199,0,80,0,218,0,173,0,0,0,36,0,191,0,106,0,112,0,170,0,162,0,169,0,98,0,59,0,0,0,175,0,112,0,64,0,164,0,207,0,249,0,225,0,0,0,187,0,249,0,65,0,0,0,151,0,78,0,180,0,0,0,129,0,191,0,72,0,215,0,20,0,235,0,12,0,148,0,25,0,0,0,42,0,95,0,122,0,0,0,210,0,44,0,39,0,234,0,104,0,131,0,3,0,35,0,154,0,131,0,59,0,116,0,117,0,66,0,215,0,133,0,0,0,194,0,183,0,56,0,47,0,178,0,10,0,0,0,207,0,121,0,226,0,130,0,0,0,115,0,123,0,0,0,0,0,63,0,99,0,63,0,24,0,8,0,108,0,0,0,230,0,201,0,6,0,88,0,207,0,158,0,100,0,205,0,124,0,0,0,24,0,0,0,0,0,100,0,140,0,28,0,7,0,4,0,153,0,141,0,207,0,103,0,0,0,80,0,131,0,0,0,217,0,193,0,233,0,33,0,203,0,161,0,197,0,0,0,195,0,228,0,174,0,197,0,0,0,0,0,0,0,67,0,0,0,55,0,214,0,236,0,174,0,217,0,125,0,129,0,0,0,0,0,238,0,181,0,104,0,126,0,246,0,0,0,72,0,232,0,0,0,240,0,179,0,218,0,131,0,146,0,164,0,218,0,0,0,165,0,224,0,71,0,196,0,79,0,0,0,0,0,250,0,140,0,46,0,7,0,8,0,101,0,74,0,0,0,36,0,146,0,0,0,66,0,175,0,227,0,0,0,0,0,0,0,0,0,128,0,214,0,57,0,0,0,124,0,53,0,49,0,0,0,0,0,58,0,0,0,0,0,90,0,235,0,13,0,119,0,202,0,210,0,139,0,216,0,0,0,179,0,214,0,91,0,127,0,112,0,0,0,103,0,67,0,97,0,85,0,111,0,224,0,136,0,203,0,42,0,70,0,39,0,244,0,5,0,235,0,96,0,134,0,194,0,162,0,152,0,24,0,95,0,0,0,209,0,0,0,62,0,11,0,121,0,46,0,62,0,239,0,45,0,59,0,108,0,134,0,233,0,238,0,12,0,194,0,241,0,106,0,249,0,155,0,82,0,16,0,54,0,0,0,247,0,0,0,0,0,176,0,88,0,0,0,12,0,37,0,246,0,35,0,0,0,0,0,0,0,0,0,0,0,37,0,37,0,55,0,148,0,126,0,0,0,0,0,213,0,197,0,31,0,0,0,0,0,210,0,98,0,168,0,205,0,0,0,0,0,57,0,0,0,88,0,239,0,18,0,0,0,92,0,76,0,19,0,242,0,154,0,27,0,54,0,0,0,230,0,37,0,238,0,76,0,34,0,107,0,161,0,101,0,251,0,245,0,136,0,151,0,202,0,4,0,138,0,2,0,63,0,25,0,2,0,126,0,99,0,109,0,191,0,104,0,157,0,0,0,0,0,166,0,177,0,62,0,101,0,96,0,100,0,242,0,5,0,81,0,0,0,252,0,27,0,79,0,157,0,154,0,23,0,30,0,34,0,196,0,240,0,59,0,0,0,161,0,38,0,208,0,1,0,174,0,0,0,225,0,188,0,189,0,48,0,206,0,30,0,200,0,41,0,198,0,0,0,255,0,242,0,88,0,131,0,149,0,227,0,177,0,41,0,0,0,59,0,245,0,241,0,122,0,212,0,109,0,0,0,0,0,237,0,154,0,131,0,0,0,94,0,198,0,212,0,32,0,33,0,178,0,37,0,139,0,0,0,0,0,0,0,103,0,245,0,38,0,188,0,251,0,244,0,228,0,0,0,95,0,91,0,196,0,246,0,244,0,53,0,92,0,151,0,0,0,206,0,119,0,165,0,24,0,182,0,0,0,147,0,0,0,16,0,61,0,130,0,21,0,17,0,183,0,193,0,225,0,0,0,33,0,94,0,82,0,126,0,184,0,0,0,68,0,0,0,2,0,237,0,237,0,212,0,211,0,0,0,91,0,238,0,136,0,0,0,5,0,81,0,232,0,0,0,102,0,0,0,168,0,140,0,171,0,41,0,18,0,163,0,0,0,16,0,70,0,74,0,52,0,115,0,158,0,40,0,34,0,0,0);
signal scenario_full  : scenario_type := (30,31,30,30,155,31,243,31,240,31,143,31,143,30,118,31,118,30,23,31,216,31,77,31,73,31,11,31,11,30,55,31,93,31,183,31,83,31,250,31,250,30,250,29,84,31,160,31,226,31,15,31,70,31,155,31,66,31,91,31,212,31,212,30,212,29,212,28,96,31,125,31,234,31,234,30,39,31,244,31,148,31,79,31,107,31,119,31,119,30,162,31,157,31,157,30,157,29,144,31,245,31,132,31,132,30,159,31,222,31,160,31,83,31,95,31,252,31,252,30,61,31,214,31,214,30,12,31,149,31,149,30,169,31,163,31,255,31,52,31,23,31,246,31,246,30,170,31,3,31,62,31,17,31,12,31,38,31,146,31,72,31,19,31,19,30,16,31,103,31,154,31,137,31,21,31,4,31,131,31,126,31,241,31,125,31,153,31,36,31,14,31,14,30,235,31,248,31,127,31,147,31,255,31,251,31,233,31,80,31,80,30,174,31,143,31,94,31,38,31,38,30,143,31,178,31,144,31,171,31,98,31,247,31,240,31,30,31,30,30,236,31,13,31,13,30,159,31,229,31,136,31,136,30,162,31,86,31,208,31,173,31,13,31,168,31,115,31,27,31,154,31,154,30,40,31,60,31,65,31,65,30,23,31,170,31,110,31,110,30,161,31,162,31,5,31,44,31,184,31,184,30,150,31,150,30,123,31,198,31,254,31,174,31,174,30,122,31,110,31,110,30,20,31,9,31,9,30,201,31,180,31,180,31,156,31,160,31,4,31,118,31,35,31,135,31,85,31,85,30,61,31,93,31,250,31,221,31,155,31,146,31,146,30,38,31,130,31,219,31,152,31,96,31,166,31,191,31,191,30,219,31,187,31,127,31,127,30,127,29,46,31,49,31,135,31,223,31,223,30,70,31,16,31,139,31,36,31,221,31,168,31,61,31,157,31,157,30,17,31,69,31,222,31,36,31,22,31,8,31,238,31,104,31,122,31,195,31,181,31,167,31,46,31,144,31,202,31,109,31,115,31,23,31,113,31,113,30,72,31,37,31,30,31,132,31,132,30,132,29,242,31,48,31,236,31,130,31,88,31,187,31,187,30,231,31,237,31,188,31,219,31,219,30,92,31,130,31,3,31,20,31,238,31,238,30,110,31,243,31,52,31,134,31,134,30,185,31,4,31,191,31,8,31,8,30,236,31,132,31,199,31,19,31,19,30,133,31,72,31,250,31,187,31,97,31,97,30,183,31,77,31,12,31,12,30,114,31,129,31,11,31,251,31,87,31,56,31,53,31,231,31,231,30,73,31,252,31,130,31,118,31,118,30,242,31,54,31,50,31,229,31,185,31,173,31,4,31,136,31,136,30,8,31,153,31,118,31,64,31,203,31,2,31,2,30,101,31,54,31,104,31,116,31,92,31,249,31,81,31,141,31,141,30,126,31,69,31,69,30,98,31,16,31,177,31,173,31,173,30,81,31,81,30,120,31,82,31,28,31,205,31,228,31,199,31,199,30,154,31,250,31,250,30,165,31,109,31,241,31,6,31,214,31,121,31,217,31,154,31,35,31,35,30,16,31,16,30,165,31,239,31,239,30,199,31,80,31,218,31,173,31,173,30,36,31,191,31,106,31,112,31,170,31,162,31,169,31,98,31,59,31,59,30,175,31,112,31,64,31,164,31,207,31,249,31,225,31,225,30,187,31,249,31,65,31,65,30,151,31,78,31,180,31,180,30,129,31,191,31,72,31,215,31,20,31,235,31,12,31,148,31,25,31,25,30,42,31,95,31,122,31,122,30,210,31,44,31,39,31,234,31,104,31,131,31,3,31,35,31,154,31,131,31,59,31,116,31,117,31,66,31,215,31,133,31,133,30,194,31,183,31,56,31,47,31,178,31,10,31,10,30,207,31,121,31,226,31,130,31,130,30,115,31,123,31,123,30,123,29,63,31,99,31,63,31,24,31,8,31,108,31,108,30,230,31,201,31,6,31,88,31,207,31,158,31,100,31,205,31,124,31,124,30,24,31,24,30,24,29,100,31,140,31,28,31,7,31,4,31,153,31,141,31,207,31,103,31,103,30,80,31,131,31,131,30,217,31,193,31,233,31,33,31,203,31,161,31,197,31,197,30,195,31,228,31,174,31,197,31,197,30,197,29,197,28,67,31,67,30,55,31,214,31,236,31,174,31,217,31,125,31,129,31,129,30,129,29,238,31,181,31,104,31,126,31,246,31,246,30,72,31,232,31,232,30,240,31,179,31,218,31,131,31,146,31,164,31,218,31,218,30,165,31,224,31,71,31,196,31,79,31,79,30,79,29,250,31,140,31,46,31,7,31,8,31,101,31,74,31,74,30,36,31,146,31,146,30,66,31,175,31,227,31,227,30,227,29,227,28,227,27,128,31,214,31,57,31,57,30,124,31,53,31,49,31,49,30,49,29,58,31,58,30,58,29,90,31,235,31,13,31,119,31,202,31,210,31,139,31,216,31,216,30,179,31,214,31,91,31,127,31,112,31,112,30,103,31,67,31,97,31,85,31,111,31,224,31,136,31,203,31,42,31,70,31,39,31,244,31,5,31,235,31,96,31,134,31,194,31,162,31,152,31,24,31,95,31,95,30,209,31,209,30,62,31,11,31,121,31,46,31,62,31,239,31,45,31,59,31,108,31,134,31,233,31,238,31,12,31,194,31,241,31,106,31,249,31,155,31,82,31,16,31,54,31,54,30,247,31,247,30,247,29,176,31,88,31,88,30,12,31,37,31,246,31,35,31,35,30,35,29,35,28,35,27,35,26,37,31,37,31,55,31,148,31,126,31,126,30,126,29,213,31,197,31,31,31,31,30,31,29,210,31,98,31,168,31,205,31,205,30,205,29,57,31,57,30,88,31,239,31,18,31,18,30,92,31,76,31,19,31,242,31,154,31,27,31,54,31,54,30,230,31,37,31,238,31,76,31,34,31,107,31,161,31,101,31,251,31,245,31,136,31,151,31,202,31,4,31,138,31,2,31,63,31,25,31,2,31,126,31,99,31,109,31,191,31,104,31,157,31,157,30,157,29,166,31,177,31,62,31,101,31,96,31,100,31,242,31,5,31,81,31,81,30,252,31,27,31,79,31,157,31,154,31,23,31,30,31,34,31,196,31,240,31,59,31,59,30,161,31,38,31,208,31,1,31,174,31,174,30,225,31,188,31,189,31,48,31,206,31,30,31,200,31,41,31,198,31,198,30,255,31,242,31,88,31,131,31,149,31,227,31,177,31,41,31,41,30,59,31,245,31,241,31,122,31,212,31,109,31,109,30,109,29,237,31,154,31,131,31,131,30,94,31,198,31,212,31,32,31,33,31,178,31,37,31,139,31,139,30,139,29,139,28,103,31,245,31,38,31,188,31,251,31,244,31,228,31,228,30,95,31,91,31,196,31,246,31,244,31,53,31,92,31,151,31,151,30,206,31,119,31,165,31,24,31,182,31,182,30,147,31,147,30,16,31,61,31,130,31,21,31,17,31,183,31,193,31,225,31,225,30,33,31,94,31,82,31,126,31,184,31,184,30,68,31,68,30,2,31,237,31,237,31,212,31,211,31,211,30,91,31,238,31,136,31,136,30,5,31,81,31,232,31,232,30,102,31,102,30,168,31,140,31,171,31,41,31,18,31,163,31,163,30,16,31,70,31,74,31,52,31,115,31,158,31,40,31,34,31,34,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
