-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 348;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,36,0,192,0,207,0,225,0,223,0,0,0,72,0,226,0,191,0,118,0,82,0,86,0,185,0,115,0,166,0,0,0,162,0,188,0,0,0,59,0,124,0,0,0,0,0,145,0,125,0,0,0,0,0,0,0,119,0,93,0,29,0,69,0,26,0,174,0,9,0,56,0,240,0,0,0,99,0,195,0,222,0,76,0,0,0,0,0,83,0,88,0,219,0,0,0,0,0,232,0,20,0,254,0,89,0,0,0,181,0,91,0,136,0,170,0,73,0,0,0,95,0,3,0,107,0,197,0,248,0,117,0,0,0,0,0,74,0,6,0,91,0,0,0,0,0,0,0,77,0,11,0,244,0,111,0,218,0,10,0,216,0,47,0,33,0,44,0,0,0,233,0,0,0,0,0,29,0,200,0,237,0,134,0,226,0,186,0,84,0,56,0,12,0,13,0,219,0,87,0,212,0,77,0,126,0,83,0,151,0,0,0,101,0,180,0,205,0,234,0,194,0,228,0,91,0,42,0,246,0,128,0,0,0,81,0,141,0,223,0,139,0,217,0,171,0,153,0,237,0,41,0,205,0,61,0,216,0,146,0,112,0,34,0,150,0,14,0,108,0,27,0,221,0,173,0,63,0,189,0,82,0,13,0,205,0,175,0,234,0,0,0,197,0,152,0,10,0,0,0,5,0,181,0,44,0,217,0,43,0,208,0,120,0,47,0,223,0,23,0,209,0,190,0,76,0,240,0,147,0,231,0,197,0,146,0,210,0,148,0,46,0,0,0,217,0,154,0,22,0,0,0,226,0,48,0,107,0,165,0,60,0,48,0,163,0,246,0,2,0,58,0,0,0,18,0,86,0,182,0,0,0,60,0,0,0,201,0,35,0,15,0,177,0,0,0,0,0,70,0,126,0,0,0,122,0,215,0,19,0,25,0,204,0,196,0,82,0,0,0,0,0,0,0,0,0,8,0,144,0,203,0,93,0,112,0,11,0,0,0,211,0,233,0,216,0,76,0,62,0,15,0,32,0,12,0,245,0,194,0,0,0,151,0,74,0,66,0,137,0,0,0,0,0,167,0,180,0,114,0,57,0,133,0,227,0,62,0,0,0,0,0,0,0,166,0,145,0,142,0,0,0,237,0,123,0,146,0,132,0,104,0,162,0,18,0,60,0,43,0,198,0,211,0,205,0,182,0,0,0,39,0,0,0,176,0,217,0,23,0,14,0,207,0,18,0,48,0,14,0,43,0,24,0,89,0,223,0,139,0,150,0,194,0,72,0,185,0,117,0,252,0,0,0,57,0,237,0,7,0,147,0,58,0,0,0,191,0,0,0,23,0,123,0,0,0,3,0,210,0,113,0,145,0,164,0,103,0,0,0,0,0,76,0,202,0,182,0,0,0,0,0,193,0,155,0,63,0,206,0,90,0,149,0,87,0,202,0,80,0,0,0,0,0,104,0,162,0,195,0,111,0,131,0,0,0,40,0,67,0,200,0,133,0,49,0,77,0,15,0,18,0,16,0,201,0,155,0,52,0,0,0,23,0,0,0,112,0,203,0,243,0,104,0);
signal scenario_full  : scenario_type := (0,0,36,31,192,31,207,31,225,31,223,31,223,30,72,31,226,31,191,31,118,31,82,31,86,31,185,31,115,31,166,31,166,30,162,31,188,31,188,30,59,31,124,31,124,30,124,29,145,31,125,31,125,30,125,29,125,28,119,31,93,31,29,31,69,31,26,31,174,31,9,31,56,31,240,31,240,30,99,31,195,31,222,31,76,31,76,30,76,29,83,31,88,31,219,31,219,30,219,29,232,31,20,31,254,31,89,31,89,30,181,31,91,31,136,31,170,31,73,31,73,30,95,31,3,31,107,31,197,31,248,31,117,31,117,30,117,29,74,31,6,31,91,31,91,30,91,29,91,28,77,31,11,31,244,31,111,31,218,31,10,31,216,31,47,31,33,31,44,31,44,30,233,31,233,30,233,29,29,31,200,31,237,31,134,31,226,31,186,31,84,31,56,31,12,31,13,31,219,31,87,31,212,31,77,31,126,31,83,31,151,31,151,30,101,31,180,31,205,31,234,31,194,31,228,31,91,31,42,31,246,31,128,31,128,30,81,31,141,31,223,31,139,31,217,31,171,31,153,31,237,31,41,31,205,31,61,31,216,31,146,31,112,31,34,31,150,31,14,31,108,31,27,31,221,31,173,31,63,31,189,31,82,31,13,31,205,31,175,31,234,31,234,30,197,31,152,31,10,31,10,30,5,31,181,31,44,31,217,31,43,31,208,31,120,31,47,31,223,31,23,31,209,31,190,31,76,31,240,31,147,31,231,31,197,31,146,31,210,31,148,31,46,31,46,30,217,31,154,31,22,31,22,30,226,31,48,31,107,31,165,31,60,31,48,31,163,31,246,31,2,31,58,31,58,30,18,31,86,31,182,31,182,30,60,31,60,30,201,31,35,31,15,31,177,31,177,30,177,29,70,31,126,31,126,30,122,31,215,31,19,31,25,31,204,31,196,31,82,31,82,30,82,29,82,28,82,27,8,31,144,31,203,31,93,31,112,31,11,31,11,30,211,31,233,31,216,31,76,31,62,31,15,31,32,31,12,31,245,31,194,31,194,30,151,31,74,31,66,31,137,31,137,30,137,29,167,31,180,31,114,31,57,31,133,31,227,31,62,31,62,30,62,29,62,28,166,31,145,31,142,31,142,30,237,31,123,31,146,31,132,31,104,31,162,31,18,31,60,31,43,31,198,31,211,31,205,31,182,31,182,30,39,31,39,30,176,31,217,31,23,31,14,31,207,31,18,31,48,31,14,31,43,31,24,31,89,31,223,31,139,31,150,31,194,31,72,31,185,31,117,31,252,31,252,30,57,31,237,31,7,31,147,31,58,31,58,30,191,31,191,30,23,31,123,31,123,30,3,31,210,31,113,31,145,31,164,31,103,31,103,30,103,29,76,31,202,31,182,31,182,30,182,29,193,31,155,31,63,31,206,31,90,31,149,31,87,31,202,31,80,31,80,30,80,29,104,31,162,31,195,31,111,31,131,31,131,30,40,31,67,31,200,31,133,31,49,31,77,31,15,31,18,31,16,31,201,31,155,31,52,31,52,30,23,31,23,30,112,31,203,31,243,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
