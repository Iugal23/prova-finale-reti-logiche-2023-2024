-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 661;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,155,0,0,0,101,0,173,0,147,0,124,0,40,0,126,0,0,0,102,0,127,0,196,0,241,0,13,0,160,0,242,0,23,0,105,0,0,0,218,0,0,0,45,0,36,0,0,0,0,0,0,0,0,0,0,0,206,0,114,0,0,0,33,0,173,0,128,0,12,0,96,0,192,0,46,0,198,0,3,0,131,0,47,0,114,0,174,0,60,0,0,0,0,0,0,0,35,0,101,0,197,0,152,0,185,0,27,0,0,0,152,0,0,0,16,0,74,0,72,0,252,0,165,0,0,0,58,0,162,0,212,0,71,0,28,0,208,0,249,0,223,0,0,0,167,0,0,0,171,0,54,0,0,0,0,0,42,0,10,0,224,0,152,0,109,0,60,0,83,0,194,0,107,0,32,0,201,0,0,0,220,0,41,0,102,0,127,0,32,0,176,0,127,0,0,0,0,0,202,0,238,0,51,0,97,0,18,0,100,0,250,0,0,0,0,0,100,0,0,0,89,0,0,0,118,0,129,0,114,0,0,0,0,0,250,0,91,0,91,0,244,0,13,0,178,0,175,0,0,0,106,0,0,0,77,0,157,0,67,0,26,0,0,0,217,0,0,0,130,0,27,0,169,0,242,0,96,0,172,0,146,0,32,0,0,0,218,0,152,0,236,0,98,0,0,0,0,0,227,0,178,0,216,0,235,0,165,0,0,0,91,0,0,0,95,0,0,0,194,0,34,0,0,0,64,0,212,0,186,0,230,0,21,0,213,0,0,0,0,0,0,0,214,0,111,0,0,0,191,0,155,0,224,0,204,0,0,0,235,0,19,0,89,0,92,0,167,0,56,0,243,0,34,0,82,0,195,0,0,0,248,0,112,0,34,0,73,0,163,0,245,0,237,0,0,0,118,0,151,0,141,0,0,0,54,0,248,0,180,0,200,0,245,0,226,0,0,0,0,0,14,0,0,0,73,0,52,0,0,0,157,0,0,0,158,0,0,0,8,0,0,0,0,0,125,0,69,0,0,0,0,0,216,0,172,0,27,0,16,0,79,0,0,0,0,0,191,0,0,0,141,0,21,0,165,0,198,0,79,0,78,0,115,0,0,0,7,0,0,0,234,0,11,0,187,0,196,0,69,0,0,0,200,0,76,0,218,0,21,0,7,0,82,0,179,0,18,0,175,0,155,0,0,0,0,0,117,0,0,0,71,0,0,0,47,0,153,0,135,0,245,0,0,0,0,0,53,0,196,0,0,0,92,0,244,0,0,0,197,0,120,0,47,0,38,0,229,0,162,0,50,0,183,0,224,0,0,0,0,0,0,0,149,0,0,0,15,0,62,0,144,0,0,0,55,0,176,0,0,0,247,0,247,0,0,0,61,0,105,0,73,0,12,0,131,0,36,0,194,0,0,0,140,0,214,0,206,0,195,0,29,0,11,0,117,0,195,0,120,0,166,0,109,0,90,0,21,0,28,0,53,0,42,0,199,0,93,0,0,0,52,0,130,0,2,0,44,0,0,0,0,0,70,0,239,0,166,0,144,0,0,0,47,0,0,0,87,0,45,0,73,0,226,0,206,0,47,0,0,0,42,0,0,0,18,0,13,0,17,0,0,0,202,0,5,0,193,0,204,0,60,0,24,0,29,0,144,0,248,0,190,0,168,0,152,0,208,0,0,0,242,0,165,0,81,0,6,0,185,0,0,0,44,0,139,0,246,0,0,0,94,0,40,0,24,0,11,0,73,0,4,0,198,0,89,0,76,0,39,0,0,0,130,0,221,0,146,0,167,0,0,0,80,0,236,0,113,0,35,0,123,0,0,0,96,0,0,0,0,0,47,0,234,0,110,0,0,0,225,0,141,0,241,0,0,0,173,0,147,0,175,0,115,0,20,0,79,0,183,0,234,0,0,0,244,0,0,0,107,0,209,0,117,0,185,0,0,0,156,0,101,0,90,0,7,0,10,0,96,0,206,0,101,0,24,0,63,0,0,0,179,0,29,0,0,0,42,0,0,0,83,0,209,0,186,0,214,0,0,0,177,0,0,0,0,0,0,0,245,0,144,0,170,0,151,0,129,0,109,0,235,0,31,0,161,0,148,0,0,0,246,0,22,0,147,0,0,0,241,0,174,0,249,0,125,0,81,0,0,0,250,0,172,0,235,0,28,0,0,0,99,0,236,0,41,0,128,0,57,0,150,0,0,0,239,0,123,0,137,0,28,0,240,0,86,0,213,0,0,0,71,0,104,0,56,0,151,0,216,0,253,0,127,0,11,0,87,0,153,0,238,0,32,0,0,0,119,0,0,0,196,0,159,0,135,0,17,0,202,0,15,0,39,0,0,0,149,0,0,0,0,0,117,0,90,0,83,0,32,0,20,0,0,0,191,0,0,0,87,0,121,0,97,0,0,0,89,0,221,0,46,0,27,0,44,0,104,0,0,0,0,0,0,0,0,0,162,0,0,0,227,0,249,0,234,0,209,0,130,0,83,0,0,0,0,0,201,0,0,0,89,0,113,0,0,0,175,0,60,0,46,0,117,0,150,0,200,0,31,0,197,0,109,0,98,0,39,0,7,0,39,0,151,0,74,0,0,0,114,0,99,0,0,0,14,0,123,0,238,0,43,0,0,0,118,0,53,0,23,0,64,0,147,0,180,0,0,0,110,0,231,0,0,0,230,0,15,0,234,0,241,0,217,0,154,0,135,0,210,0,215,0,142,0,166,0,254,0,0,0,44,0,86,0,193,0,0,0,65,0,0,0,12,0,239,0,163,0,235,0,145,0,219,0,0,0,58,0,0,0,183,0,241,0,39,0,206,0,124,0,215,0,191,0,192,0,126,0,211,0,80,0,24,0,75,0,2,0,0,0,239,0,0,0,202,0,190,0,66,0,132,0,166,0,253,0,19,0,132,0,74,0,54,0,0,0,254,0,0,0,226,0,53,0,57,0,245,0,67,0,166,0,0,0,189,0,92,0,178,0);
signal scenario_full  : scenario_type := (0,0,155,31,155,30,101,31,173,31,147,31,124,31,40,31,126,31,126,30,102,31,127,31,196,31,241,31,13,31,160,31,242,31,23,31,105,31,105,30,218,31,218,30,45,31,36,31,36,30,36,29,36,28,36,27,36,26,206,31,114,31,114,30,33,31,173,31,128,31,12,31,96,31,192,31,46,31,198,31,3,31,131,31,47,31,114,31,174,31,60,31,60,30,60,29,60,28,35,31,101,31,197,31,152,31,185,31,27,31,27,30,152,31,152,30,16,31,74,31,72,31,252,31,165,31,165,30,58,31,162,31,212,31,71,31,28,31,208,31,249,31,223,31,223,30,167,31,167,30,171,31,54,31,54,30,54,29,42,31,10,31,224,31,152,31,109,31,60,31,83,31,194,31,107,31,32,31,201,31,201,30,220,31,41,31,102,31,127,31,32,31,176,31,127,31,127,30,127,29,202,31,238,31,51,31,97,31,18,31,100,31,250,31,250,30,250,29,100,31,100,30,89,31,89,30,118,31,129,31,114,31,114,30,114,29,250,31,91,31,91,31,244,31,13,31,178,31,175,31,175,30,106,31,106,30,77,31,157,31,67,31,26,31,26,30,217,31,217,30,130,31,27,31,169,31,242,31,96,31,172,31,146,31,32,31,32,30,218,31,152,31,236,31,98,31,98,30,98,29,227,31,178,31,216,31,235,31,165,31,165,30,91,31,91,30,95,31,95,30,194,31,34,31,34,30,64,31,212,31,186,31,230,31,21,31,213,31,213,30,213,29,213,28,214,31,111,31,111,30,191,31,155,31,224,31,204,31,204,30,235,31,19,31,89,31,92,31,167,31,56,31,243,31,34,31,82,31,195,31,195,30,248,31,112,31,34,31,73,31,163,31,245,31,237,31,237,30,118,31,151,31,141,31,141,30,54,31,248,31,180,31,200,31,245,31,226,31,226,30,226,29,14,31,14,30,73,31,52,31,52,30,157,31,157,30,158,31,158,30,8,31,8,30,8,29,125,31,69,31,69,30,69,29,216,31,172,31,27,31,16,31,79,31,79,30,79,29,191,31,191,30,141,31,21,31,165,31,198,31,79,31,78,31,115,31,115,30,7,31,7,30,234,31,11,31,187,31,196,31,69,31,69,30,200,31,76,31,218,31,21,31,7,31,82,31,179,31,18,31,175,31,155,31,155,30,155,29,117,31,117,30,71,31,71,30,47,31,153,31,135,31,245,31,245,30,245,29,53,31,196,31,196,30,92,31,244,31,244,30,197,31,120,31,47,31,38,31,229,31,162,31,50,31,183,31,224,31,224,30,224,29,224,28,149,31,149,30,15,31,62,31,144,31,144,30,55,31,176,31,176,30,247,31,247,31,247,30,61,31,105,31,73,31,12,31,131,31,36,31,194,31,194,30,140,31,214,31,206,31,195,31,29,31,11,31,117,31,195,31,120,31,166,31,109,31,90,31,21,31,28,31,53,31,42,31,199,31,93,31,93,30,52,31,130,31,2,31,44,31,44,30,44,29,70,31,239,31,166,31,144,31,144,30,47,31,47,30,87,31,45,31,73,31,226,31,206,31,47,31,47,30,42,31,42,30,18,31,13,31,17,31,17,30,202,31,5,31,193,31,204,31,60,31,24,31,29,31,144,31,248,31,190,31,168,31,152,31,208,31,208,30,242,31,165,31,81,31,6,31,185,31,185,30,44,31,139,31,246,31,246,30,94,31,40,31,24,31,11,31,73,31,4,31,198,31,89,31,76,31,39,31,39,30,130,31,221,31,146,31,167,31,167,30,80,31,236,31,113,31,35,31,123,31,123,30,96,31,96,30,96,29,47,31,234,31,110,31,110,30,225,31,141,31,241,31,241,30,173,31,147,31,175,31,115,31,20,31,79,31,183,31,234,31,234,30,244,31,244,30,107,31,209,31,117,31,185,31,185,30,156,31,101,31,90,31,7,31,10,31,96,31,206,31,101,31,24,31,63,31,63,30,179,31,29,31,29,30,42,31,42,30,83,31,209,31,186,31,214,31,214,30,177,31,177,30,177,29,177,28,245,31,144,31,170,31,151,31,129,31,109,31,235,31,31,31,161,31,148,31,148,30,246,31,22,31,147,31,147,30,241,31,174,31,249,31,125,31,81,31,81,30,250,31,172,31,235,31,28,31,28,30,99,31,236,31,41,31,128,31,57,31,150,31,150,30,239,31,123,31,137,31,28,31,240,31,86,31,213,31,213,30,71,31,104,31,56,31,151,31,216,31,253,31,127,31,11,31,87,31,153,31,238,31,32,31,32,30,119,31,119,30,196,31,159,31,135,31,17,31,202,31,15,31,39,31,39,30,149,31,149,30,149,29,117,31,90,31,83,31,32,31,20,31,20,30,191,31,191,30,87,31,121,31,97,31,97,30,89,31,221,31,46,31,27,31,44,31,104,31,104,30,104,29,104,28,104,27,162,31,162,30,227,31,249,31,234,31,209,31,130,31,83,31,83,30,83,29,201,31,201,30,89,31,113,31,113,30,175,31,60,31,46,31,117,31,150,31,200,31,31,31,197,31,109,31,98,31,39,31,7,31,39,31,151,31,74,31,74,30,114,31,99,31,99,30,14,31,123,31,238,31,43,31,43,30,118,31,53,31,23,31,64,31,147,31,180,31,180,30,110,31,231,31,231,30,230,31,15,31,234,31,241,31,217,31,154,31,135,31,210,31,215,31,142,31,166,31,254,31,254,30,44,31,86,31,193,31,193,30,65,31,65,30,12,31,239,31,163,31,235,31,145,31,219,31,219,30,58,31,58,30,183,31,241,31,39,31,206,31,124,31,215,31,191,31,192,31,126,31,211,31,80,31,24,31,75,31,2,31,2,30,239,31,239,30,202,31,190,31,66,31,132,31,166,31,253,31,19,31,132,31,74,31,54,31,54,30,254,31,254,30,226,31,53,31,57,31,245,31,67,31,166,31,166,30,189,31,92,31,178,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
