-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 779;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (228,0,223,0,115,0,111,0,81,0,95,0,152,0,0,0,115,0,0,0,65,0,0,0,255,0,0,0,195,0,0,0,0,0,196,0,0,0,79,0,0,0,212,0,219,0,222,0,0,0,204,0,26,0,0,0,53,0,186,0,54,0,202,0,182,0,0,0,0,0,225,0,223,0,192,0,0,0,232,0,13,0,184,0,95,0,228,0,198,0,214,0,162,0,23,0,165,0,178,0,230,0,31,0,100,0,62,0,94,0,173,0,226,0,146,0,97,0,109,0,140,0,0,0,28,0,208,0,15,0,148,0,211,0,145,0,83,0,43,0,0,0,80,0,148,0,127,0,237,0,91,0,113,0,0,0,128,0,134,0,0,0,144,0,0,0,71,0,234,0,123,0,0,0,159,0,240,0,0,0,189,0,0,0,250,0,160,0,242,0,215,0,148,0,120,0,63,0,69,0,0,0,60,0,195,0,0,0,87,0,165,0,114,0,206,0,140,0,219,0,121,0,115,0,0,0,244,0,0,0,78,0,0,0,81,0,8,0,0,0,0,0,0,0,202,0,252,0,0,0,0,0,90,0,0,0,1,0,0,0,67,0,121,0,94,0,191,0,133,0,0,0,0,0,137,0,90,0,44,0,29,0,208,0,224,0,158,0,140,0,173,0,152,0,175,0,42,0,59,0,83,0,199,0,181,0,0,0,244,0,184,0,178,0,136,0,164,0,0,0,226,0,0,0,140,0,0,0,138,0,160,0,207,0,136,0,38,0,157,0,211,0,0,0,153,0,3,0,225,0,213,0,0,0,180,0,0,0,212,0,230,0,17,0,26,0,233,0,158,0,238,0,0,0,50,0,163,0,72,0,138,0,184,0,0,0,0,0,107,0,148,0,0,0,121,0,85,0,202,0,0,0,0,0,177,0,0,0,53,0,107,0,155,0,0,0,70,0,173,0,185,0,168,0,86,0,141,0,78,0,244,0,112,0,129,0,182,0,178,0,205,0,0,0,230,0,104,0,0,0,34,0,120,0,243,0,222,0,26,0,143,0,150,0,0,0,46,0,203,0,155,0,194,0,1,0,100,0,12,0,0,0,0,0,228,0,33,0,220,0,55,0,209,0,85,0,131,0,241,0,0,0,0,0,52,0,147,0,171,0,0,0,52,0,252,0,70,0,178,0,126,0,36,0,26,0,64,0,0,0,0,0,157,0,230,0,0,0,28,0,0,0,203,0,147,0,0,0,0,0,116,0,147,0,198,0,0,0,231,0,119,0,154,0,81,0,0,0,135,0,0,0,134,0,0,0,89,0,92,0,45,0,90,0,105,0,147,0,48,0,0,0,81,0,92,0,0,0,113,0,12,0,225,0,155,0,0,0,100,0,132,0,113,0,58,0,107,0,80,0,0,0,35,0,162,0,180,0,208,0,146,0,151,0,160,0,129,0,0,0,29,0,52,0,0,0,185,0,216,0,146,0,225,0,58,0,212,0,44,0,250,0,83,0,211,0,184,0,45,0,0,0,8,0,160,0,146,0,17,0,73,0,0,0,0,0,15,0,7,0,59,0,21,0,0,0,0,0,236,0,16,0,33,0,240,0,137,0,181,0,71,0,142,0,134,0,0,0,8,0,64,0,195,0,150,0,26,0,137,0,0,0,140,0,124,0,92,0,159,0,54,0,196,0,98,0,76,0,162,0,69,0,175,0,21,0,220,0,136,0,61,0,163,0,119,0,65,0,230,0,168,0,244,0,12,0,140,0,245,0,88,0,188,0,5,0,33,0,126,0,191,0,26,0,1,0,169,0,58,0,13,0,6,0,100,0,19,0,0,0,197,0,0,0,20,0,0,0,29,0,89,0,165,0,26,0,45,0,53,0,73,0,0,0,22,0,124,0,222,0,244,0,196,0,230,0,236,0,0,0,199,0,63,0,162,0,0,0,249,0,251,0,165,0,78,0,210,0,241,0,0,0,28,0,254,0,223,0,245,0,149,0,120,0,147,0,209,0,0,0,0,0,10,0,247,0,222,0,237,0,67,0,32,0,204,0,90,0,0,0,104,0,102,0,246,0,135,0,168,0,151,0,186,0,0,0,112,0,12,0,19,0,203,0,143,0,64,0,28,0,120,0,232,0,131,0,228,0,250,0,0,0,0,0,0,0,156,0,225,0,18,0,0,0,0,0,194,0,232,0,0,0,62,0,59,0,87,0,99,0,209,0,12,0,220,0,0,0,239,0,0,0,99,0,216,0,0,0,201,0,145,0,66,0,141,0,69,0,205,0,17,0,89,0,185,0,220,0,180,0,0,0,48,0,84,0,112,0,151,0,239,0,57,0,130,0,227,0,90,0,15,0,0,0,206,0,0,0,3,0,34,0,126,0,32,0,0,0,91,0,170,0,0,0,15,0,123,0,191,0,129,0,180,0,168,0,205,0,0,0,82,0,0,0,211,0,63,0,235,0,114,0,104,0,5,0,157,0,26,0,6,0,0,0,112,0,246,0,62,0,0,0,0,0,18,0,14,0,246,0,52,0,100,0,0,0,77,0,144,0,78,0,0,0,173,0,39,0,5,0,27,0,81,0,106,0,202,0,90,0,215,0,245,0,0,0,191,0,0,0,0,0,157,0,0,0,226,0,216,0,171,0,146,0,196,0,17,0,135,0,216,0,206,0,0,0,0,0,142,0,56,0,223,0,108,0,188,0,0,0,0,0,237,0,104,0,0,0,217,0,83,0,0,0,71,0,102,0,0,0,195,0,219,0,0,0,0,0,97,0,213,0,157,0,195,0,39,0,215,0,9,0,3,0,224,0,0,0,103,0,148,0,0,0,120,0,180,0,0,0,66,0,78,0,0,0,128,0,22,0,186,0,254,0,238,0,115,0,0,0,197,0,49,0,43,0,171,0,130,0,65,0,0,0,252,0,31,0,72,0,234,0,0,0,0,0,155,0,164,0,177,0,0,0,31,0,141,0,110,0,225,0,149,0,0,0,175,0,231,0,151,0,0,0,33,0,26,0,159,0,138,0,184,0,0,0,0,0,0,0,247,0,0,0,209,0,249,0,17,0,166,0,0,0,66,0,0,0,121,0,0,0,254,0,192,0,0,0,207,0,14,0,0,0,164,0,200,0,201,0,204,0,199,0,152,0,0,0,197,0,21,0,0,0,150,0,164,0,223,0,195,0,189,0,223,0,169,0,50,0,104,0,0,0,81,0,151,0,217,0,240,0,201,0,55,0,232,0,0,0,87,0,70,0,116,0,137,0,222,0,232,0,203,0,224,0,12,0,70,0,85,0,118,0,170,0,155,0,0,0,3,0,36,0,0,0,187,0,168,0,122,0,0,0,162,0,190,0,240,0,48,0,0,0,39,0,31,0,0,0,17,0,86,0,120,0,69,0,0,0,64,0,0,0,69,0,239,0,85,0,41,0,76,0,175,0,216,0,100,0,234,0,86,0,0,0,155,0,238,0,249,0,49,0,141,0,3,0,154,0,221,0,14,0,242,0,0,0);
signal scenario_full  : scenario_type := (228,31,223,31,115,31,111,31,81,31,95,31,152,31,152,30,115,31,115,30,65,31,65,30,255,31,255,30,195,31,195,30,195,29,196,31,196,30,79,31,79,30,212,31,219,31,222,31,222,30,204,31,26,31,26,30,53,31,186,31,54,31,202,31,182,31,182,30,182,29,225,31,223,31,192,31,192,30,232,31,13,31,184,31,95,31,228,31,198,31,214,31,162,31,23,31,165,31,178,31,230,31,31,31,100,31,62,31,94,31,173,31,226,31,146,31,97,31,109,31,140,31,140,30,28,31,208,31,15,31,148,31,211,31,145,31,83,31,43,31,43,30,80,31,148,31,127,31,237,31,91,31,113,31,113,30,128,31,134,31,134,30,144,31,144,30,71,31,234,31,123,31,123,30,159,31,240,31,240,30,189,31,189,30,250,31,160,31,242,31,215,31,148,31,120,31,63,31,69,31,69,30,60,31,195,31,195,30,87,31,165,31,114,31,206,31,140,31,219,31,121,31,115,31,115,30,244,31,244,30,78,31,78,30,81,31,8,31,8,30,8,29,8,28,202,31,252,31,252,30,252,29,90,31,90,30,1,31,1,30,67,31,121,31,94,31,191,31,133,31,133,30,133,29,137,31,90,31,44,31,29,31,208,31,224,31,158,31,140,31,173,31,152,31,175,31,42,31,59,31,83,31,199,31,181,31,181,30,244,31,184,31,178,31,136,31,164,31,164,30,226,31,226,30,140,31,140,30,138,31,160,31,207,31,136,31,38,31,157,31,211,31,211,30,153,31,3,31,225,31,213,31,213,30,180,31,180,30,212,31,230,31,17,31,26,31,233,31,158,31,238,31,238,30,50,31,163,31,72,31,138,31,184,31,184,30,184,29,107,31,148,31,148,30,121,31,85,31,202,31,202,30,202,29,177,31,177,30,53,31,107,31,155,31,155,30,70,31,173,31,185,31,168,31,86,31,141,31,78,31,244,31,112,31,129,31,182,31,178,31,205,31,205,30,230,31,104,31,104,30,34,31,120,31,243,31,222,31,26,31,143,31,150,31,150,30,46,31,203,31,155,31,194,31,1,31,100,31,12,31,12,30,12,29,228,31,33,31,220,31,55,31,209,31,85,31,131,31,241,31,241,30,241,29,52,31,147,31,171,31,171,30,52,31,252,31,70,31,178,31,126,31,36,31,26,31,64,31,64,30,64,29,157,31,230,31,230,30,28,31,28,30,203,31,147,31,147,30,147,29,116,31,147,31,198,31,198,30,231,31,119,31,154,31,81,31,81,30,135,31,135,30,134,31,134,30,89,31,92,31,45,31,90,31,105,31,147,31,48,31,48,30,81,31,92,31,92,30,113,31,12,31,225,31,155,31,155,30,100,31,132,31,113,31,58,31,107,31,80,31,80,30,35,31,162,31,180,31,208,31,146,31,151,31,160,31,129,31,129,30,29,31,52,31,52,30,185,31,216,31,146,31,225,31,58,31,212,31,44,31,250,31,83,31,211,31,184,31,45,31,45,30,8,31,160,31,146,31,17,31,73,31,73,30,73,29,15,31,7,31,59,31,21,31,21,30,21,29,236,31,16,31,33,31,240,31,137,31,181,31,71,31,142,31,134,31,134,30,8,31,64,31,195,31,150,31,26,31,137,31,137,30,140,31,124,31,92,31,159,31,54,31,196,31,98,31,76,31,162,31,69,31,175,31,21,31,220,31,136,31,61,31,163,31,119,31,65,31,230,31,168,31,244,31,12,31,140,31,245,31,88,31,188,31,5,31,33,31,126,31,191,31,26,31,1,31,169,31,58,31,13,31,6,31,100,31,19,31,19,30,197,31,197,30,20,31,20,30,29,31,89,31,165,31,26,31,45,31,53,31,73,31,73,30,22,31,124,31,222,31,244,31,196,31,230,31,236,31,236,30,199,31,63,31,162,31,162,30,249,31,251,31,165,31,78,31,210,31,241,31,241,30,28,31,254,31,223,31,245,31,149,31,120,31,147,31,209,31,209,30,209,29,10,31,247,31,222,31,237,31,67,31,32,31,204,31,90,31,90,30,104,31,102,31,246,31,135,31,168,31,151,31,186,31,186,30,112,31,12,31,19,31,203,31,143,31,64,31,28,31,120,31,232,31,131,31,228,31,250,31,250,30,250,29,250,28,156,31,225,31,18,31,18,30,18,29,194,31,232,31,232,30,62,31,59,31,87,31,99,31,209,31,12,31,220,31,220,30,239,31,239,30,99,31,216,31,216,30,201,31,145,31,66,31,141,31,69,31,205,31,17,31,89,31,185,31,220,31,180,31,180,30,48,31,84,31,112,31,151,31,239,31,57,31,130,31,227,31,90,31,15,31,15,30,206,31,206,30,3,31,34,31,126,31,32,31,32,30,91,31,170,31,170,30,15,31,123,31,191,31,129,31,180,31,168,31,205,31,205,30,82,31,82,30,211,31,63,31,235,31,114,31,104,31,5,31,157,31,26,31,6,31,6,30,112,31,246,31,62,31,62,30,62,29,18,31,14,31,246,31,52,31,100,31,100,30,77,31,144,31,78,31,78,30,173,31,39,31,5,31,27,31,81,31,106,31,202,31,90,31,215,31,245,31,245,30,191,31,191,30,191,29,157,31,157,30,226,31,216,31,171,31,146,31,196,31,17,31,135,31,216,31,206,31,206,30,206,29,142,31,56,31,223,31,108,31,188,31,188,30,188,29,237,31,104,31,104,30,217,31,83,31,83,30,71,31,102,31,102,30,195,31,219,31,219,30,219,29,97,31,213,31,157,31,195,31,39,31,215,31,9,31,3,31,224,31,224,30,103,31,148,31,148,30,120,31,180,31,180,30,66,31,78,31,78,30,128,31,22,31,186,31,254,31,238,31,115,31,115,30,197,31,49,31,43,31,171,31,130,31,65,31,65,30,252,31,31,31,72,31,234,31,234,30,234,29,155,31,164,31,177,31,177,30,31,31,141,31,110,31,225,31,149,31,149,30,175,31,231,31,151,31,151,30,33,31,26,31,159,31,138,31,184,31,184,30,184,29,184,28,247,31,247,30,209,31,249,31,17,31,166,31,166,30,66,31,66,30,121,31,121,30,254,31,192,31,192,30,207,31,14,31,14,30,164,31,200,31,201,31,204,31,199,31,152,31,152,30,197,31,21,31,21,30,150,31,164,31,223,31,195,31,189,31,223,31,169,31,50,31,104,31,104,30,81,31,151,31,217,31,240,31,201,31,55,31,232,31,232,30,87,31,70,31,116,31,137,31,222,31,232,31,203,31,224,31,12,31,70,31,85,31,118,31,170,31,155,31,155,30,3,31,36,31,36,30,187,31,168,31,122,31,122,30,162,31,190,31,240,31,48,31,48,30,39,31,31,31,31,30,17,31,86,31,120,31,69,31,69,30,64,31,64,30,69,31,239,31,85,31,41,31,76,31,175,31,216,31,100,31,234,31,86,31,86,30,155,31,238,31,249,31,49,31,141,31,3,31,154,31,221,31,14,31,242,31,242,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
