-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 393;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,97,0,0,0,181,0,215,0,85,0,190,0,45,0,49,0,155,0,170,0,25,0,206,0,132,0,106,0,239,0,91,0,52,0,0,0,13,0,138,0,193,0,242,0,197,0,151,0,0,0,169,0,0,0,252,0,90,0,251,0,108,0,0,0,163,0,5,0,51,0,0,0,197,0,69,0,96,0,232,0,9,0,80,0,255,0,157,0,206,0,187,0,42,0,203,0,179,0,101,0,0,0,24,0,209,0,136,0,146,0,102,0,190,0,72,0,145,0,115,0,17,0,189,0,0,0,241,0,50,0,89,0,0,0,181,0,0,0,78,0,123,0,22,0,0,0,210,0,0,0,194,0,104,0,52,0,229,0,131,0,0,0,183,0,198,0,206,0,52,0,34,0,160,0,225,0,218,0,0,0,116,0,132,0,148,0,81,0,236,0,85,0,63,0,66,0,0,0,109,0,48,0,0,0,146,0,9,0,126,0,246,0,197,0,102,0,116,0,116,0,157,0,0,0,72,0,171,0,48,0,217,0,27,0,0,0,19,0,195,0,40,0,150,0,85,0,117,0,0,0,159,0,36,0,0,0,151,0,25,0,57,0,56,0,151,0,171,0,169,0,0,0,0,0,240,0,70,0,0,0,41,0,249,0,49,0,0,0,64,0,61,0,111,0,76,0,173,0,30,0,0,0,162,0,22,0,0,0,108,0,74,0,36,0,242,0,0,0,214,0,54,0,125,0,74,0,179,0,222,0,186,0,0,0,192,0,9,0,46,0,0,0,233,0,22,0,176,0,110,0,190,0,186,0,0,0,74,0,2,0,0,0,165,0,46,0,0,0,178,0,118,0,0,0,154,0,64,0,197,0,0,0,237,0,96,0,0,0,197,0,114,0,99,0,3,0,218,0,154,0,236,0,203,0,0,0,7,0,16,0,155,0,197,0,197,0,32,0,187,0,14,0,0,0,103,0,81,0,147,0,84,0,0,0,116,0,198,0,125,0,0,0,110,0,154,0,42,0,104,0,200,0,181,0,18,0,0,0,218,0,0,0,29,0,0,0,162,0,220,0,224,0,214,0,225,0,46,0,39,0,64,0,231,0,0,0,137,0,11,0,195,0,0,0,110,0,246,0,95,0,77,0,62,0,220,0,79,0,30,0,79,0,166,0,0,0,0,0,201,0,194,0,180,0,248,0,144,0,168,0,93,0,221,0,0,0,0,0,0,0,23,0,178,0,0,0,0,0,87,0,218,0,207,0,142,0,41,0,104,0,0,0,19,0,188,0,118,0,211,0,183,0,0,0,249,0,0,0,189,0,179,0,128,0,106,0,203,0,228,0,45,0,146,0,168,0,189,0,196,0,186,0,209,0,222,0,41,0,150,0,124,0,179,0,0,0,169,0,212,0,137,0,251,0,110,0,71,0,0,0,216,0,57,0,40,0,0,0,34,0,0,0,64,0,154,0,0,0,57,0,129,0,0,0,128,0,56,0,39,0,186,0,71,0,139,0,82,0,1,0,67,0,198,0,147,0,234,0,227,0,0,0,0,0,129,0,197,0,52,0,67,0,0,0,25,0,171,0,27,0,164,0,152,0,236,0,133,0,92,0,170,0,217,0,45,0,0,0,0,0,3,0,29,0,135,0,138,0,0,0,246,0,204,0,207,0,170,0,0,0,0,0,190,0,217,0,0,0,78,0,0,0,89,0,0,0,0,0,113,0,248,0,149,0,254,0,17,0,251,0,175,0,4,0,60,0,91,0,63,0,83,0,76,0);
signal scenario_full  : scenario_type := (0,0,97,31,97,30,181,31,215,31,85,31,190,31,45,31,49,31,155,31,170,31,25,31,206,31,132,31,106,31,239,31,91,31,52,31,52,30,13,31,138,31,193,31,242,31,197,31,151,31,151,30,169,31,169,30,252,31,90,31,251,31,108,31,108,30,163,31,5,31,51,31,51,30,197,31,69,31,96,31,232,31,9,31,80,31,255,31,157,31,206,31,187,31,42,31,203,31,179,31,101,31,101,30,24,31,209,31,136,31,146,31,102,31,190,31,72,31,145,31,115,31,17,31,189,31,189,30,241,31,50,31,89,31,89,30,181,31,181,30,78,31,123,31,22,31,22,30,210,31,210,30,194,31,104,31,52,31,229,31,131,31,131,30,183,31,198,31,206,31,52,31,34,31,160,31,225,31,218,31,218,30,116,31,132,31,148,31,81,31,236,31,85,31,63,31,66,31,66,30,109,31,48,31,48,30,146,31,9,31,126,31,246,31,197,31,102,31,116,31,116,31,157,31,157,30,72,31,171,31,48,31,217,31,27,31,27,30,19,31,195,31,40,31,150,31,85,31,117,31,117,30,159,31,36,31,36,30,151,31,25,31,57,31,56,31,151,31,171,31,169,31,169,30,169,29,240,31,70,31,70,30,41,31,249,31,49,31,49,30,64,31,61,31,111,31,76,31,173,31,30,31,30,30,162,31,22,31,22,30,108,31,74,31,36,31,242,31,242,30,214,31,54,31,125,31,74,31,179,31,222,31,186,31,186,30,192,31,9,31,46,31,46,30,233,31,22,31,176,31,110,31,190,31,186,31,186,30,74,31,2,31,2,30,165,31,46,31,46,30,178,31,118,31,118,30,154,31,64,31,197,31,197,30,237,31,96,31,96,30,197,31,114,31,99,31,3,31,218,31,154,31,236,31,203,31,203,30,7,31,16,31,155,31,197,31,197,31,32,31,187,31,14,31,14,30,103,31,81,31,147,31,84,31,84,30,116,31,198,31,125,31,125,30,110,31,154,31,42,31,104,31,200,31,181,31,18,31,18,30,218,31,218,30,29,31,29,30,162,31,220,31,224,31,214,31,225,31,46,31,39,31,64,31,231,31,231,30,137,31,11,31,195,31,195,30,110,31,246,31,95,31,77,31,62,31,220,31,79,31,30,31,79,31,166,31,166,30,166,29,201,31,194,31,180,31,248,31,144,31,168,31,93,31,221,31,221,30,221,29,221,28,23,31,178,31,178,30,178,29,87,31,218,31,207,31,142,31,41,31,104,31,104,30,19,31,188,31,118,31,211,31,183,31,183,30,249,31,249,30,189,31,179,31,128,31,106,31,203,31,228,31,45,31,146,31,168,31,189,31,196,31,186,31,209,31,222,31,41,31,150,31,124,31,179,31,179,30,169,31,212,31,137,31,251,31,110,31,71,31,71,30,216,31,57,31,40,31,40,30,34,31,34,30,64,31,154,31,154,30,57,31,129,31,129,30,128,31,56,31,39,31,186,31,71,31,139,31,82,31,1,31,67,31,198,31,147,31,234,31,227,31,227,30,227,29,129,31,197,31,52,31,67,31,67,30,25,31,171,31,27,31,164,31,152,31,236,31,133,31,92,31,170,31,217,31,45,31,45,30,45,29,3,31,29,31,135,31,138,31,138,30,246,31,204,31,207,31,170,31,170,30,170,29,190,31,217,31,217,30,78,31,78,30,89,31,89,30,89,29,113,31,248,31,149,31,254,31,17,31,251,31,175,31,4,31,60,31,91,31,63,31,83,31,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
