-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 304;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,221,0,81,0,8,0,113,0,107,0,225,0,154,0,191,0,29,0,22,0,207,0,118,0,0,0,155,0,0,0,0,0,179,0,78,0,254,0,214,0,10,0,100,0,106,0,97,0,249,0,106,0,147,0,125,0,148,0,207,0,200,0,120,0,0,0,134,0,215,0,219,0,0,0,0,0,255,0,159,0,0,0,76,0,8,0,34,0,0,0,10,0,217,0,0,0,130,0,237,0,159,0,66,0,119,0,195,0,160,0,77,0,104,0,151,0,229,0,228,0,58,0,149,0,29,0,161,0,0,0,0,0,187,0,97,0,35,0,0,0,89,0,0,0,0,0,25,0,0,0,184,0,182,0,88,0,84,0,225,0,0,0,111,0,145,0,240,0,97,0,163,0,68,0,63,0,173,0,0,0,0,0,49,0,43,0,62,0,96,0,207,0,72,0,0,0,115,0,0,0,151,0,190,0,85,0,166,0,212,0,161,0,16,0,246,0,120,0,209,0,0,0,101,0,131,0,219,0,191,0,134,0,246,0,116,0,8,0,112,0,193,0,9,0,0,0,3,0,165,0,161,0,142,0,62,0,222,0,20,0,11,0,42,0,209,0,242,0,54,0,238,0,219,0,178,0,241,0,0,0,7,0,165,0,218,0,220,0,129,0,0,0,105,0,138,0,0,0,51,0,198,0,214,0,76,0,170,0,168,0,0,0,132,0,150,0,111,0,167,0,0,0,50,0,161,0,82,0,137,0,98,0,229,0,223,0,151,0,10,0,168,0,204,0,64,0,195,0,170,0,0,0,29,0,56,0,5,0,125,0,144,0,180,0,0,0,243,0,225,0,0,0,145,0,112,0,0,0,216,0,16,0,222,0,125,0,0,0,0,0,0,0,0,0,219,0,172,0,0,0,0,0,141,0,106,0,46,0,199,0,201,0,26,0,165,0,247,0,54,0,76,0,181,0,216,0,0,0,166,0,0,0,74,0,0,0,22,0,144,0,32,0,175,0,20,0,252,0,215,0,63,0,243,0,0,0,0,0,141,0,87,0,215,0,230,0,10,0,220,0,197,0,0,0,0,0,154,0,255,0,86,0,37,0,0,0,246,0,63,0,192,0,173,0,234,0,180,0,0,0,0,0,44,0,3,0,245,0,206,0,171,0,0,0,0,0,69,0,7,0,189,0,134,0,47,0,240,0,41,0,47,0,110,0,133,0,117,0,0,0,0,0,0,0,223,0,154,0,146,0,250,0,39,0,118,0,0,0,55,0,247,0,150,0,110,0,225,0,0,0,3,0,92,0,129,0,83,0,227,0,0,0,31,0,0,0,240,0,203,0,0,0,207,0,59,0,7,0,167,0,176,0,64,0,184,0);
signal scenario_full  : scenario_type := (0,0,221,31,81,31,8,31,113,31,107,31,225,31,154,31,191,31,29,31,22,31,207,31,118,31,118,30,155,31,155,30,155,29,179,31,78,31,254,31,214,31,10,31,100,31,106,31,97,31,249,31,106,31,147,31,125,31,148,31,207,31,200,31,120,31,120,30,134,31,215,31,219,31,219,30,219,29,255,31,159,31,159,30,76,31,8,31,34,31,34,30,10,31,217,31,217,30,130,31,237,31,159,31,66,31,119,31,195,31,160,31,77,31,104,31,151,31,229,31,228,31,58,31,149,31,29,31,161,31,161,30,161,29,187,31,97,31,35,31,35,30,89,31,89,30,89,29,25,31,25,30,184,31,182,31,88,31,84,31,225,31,225,30,111,31,145,31,240,31,97,31,163,31,68,31,63,31,173,31,173,30,173,29,49,31,43,31,62,31,96,31,207,31,72,31,72,30,115,31,115,30,151,31,190,31,85,31,166,31,212,31,161,31,16,31,246,31,120,31,209,31,209,30,101,31,131,31,219,31,191,31,134,31,246,31,116,31,8,31,112,31,193,31,9,31,9,30,3,31,165,31,161,31,142,31,62,31,222,31,20,31,11,31,42,31,209,31,242,31,54,31,238,31,219,31,178,31,241,31,241,30,7,31,165,31,218,31,220,31,129,31,129,30,105,31,138,31,138,30,51,31,198,31,214,31,76,31,170,31,168,31,168,30,132,31,150,31,111,31,167,31,167,30,50,31,161,31,82,31,137,31,98,31,229,31,223,31,151,31,10,31,168,31,204,31,64,31,195,31,170,31,170,30,29,31,56,31,5,31,125,31,144,31,180,31,180,30,243,31,225,31,225,30,145,31,112,31,112,30,216,31,16,31,222,31,125,31,125,30,125,29,125,28,125,27,219,31,172,31,172,30,172,29,141,31,106,31,46,31,199,31,201,31,26,31,165,31,247,31,54,31,76,31,181,31,216,31,216,30,166,31,166,30,74,31,74,30,22,31,144,31,32,31,175,31,20,31,252,31,215,31,63,31,243,31,243,30,243,29,141,31,87,31,215,31,230,31,10,31,220,31,197,31,197,30,197,29,154,31,255,31,86,31,37,31,37,30,246,31,63,31,192,31,173,31,234,31,180,31,180,30,180,29,44,31,3,31,245,31,206,31,171,31,171,30,171,29,69,31,7,31,189,31,134,31,47,31,240,31,41,31,47,31,110,31,133,31,117,31,117,30,117,29,117,28,223,31,154,31,146,31,250,31,39,31,118,31,118,30,55,31,247,31,150,31,110,31,225,31,225,30,3,31,92,31,129,31,83,31,227,31,227,30,31,31,31,30,240,31,203,31,203,30,207,31,59,31,7,31,167,31,176,31,64,31,184,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
