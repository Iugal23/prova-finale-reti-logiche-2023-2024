-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_443 is
end project_tb_443;

architecture project_tb_arch_443 of project_tb_443 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 680;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,56,0,0,0,229,0,208,0,0,0,0,0,227,0,38,0,2,0,170,0,107,0,178,0,0,0,0,0,0,0,63,0,36,0,195,0,249,0,97,0,131,0,191,0,214,0,157,0,241,0,114,0,130,0,145,0,204,0,0,0,149,0,50,0,222,0,2,0,255,0,236,0,156,0,83,0,68,0,2,0,0,0,222,0,0,0,178,0,111,0,200,0,231,0,0,0,193,0,194,0,150,0,91,0,93,0,214,0,31,0,109,0,250,0,0,0,47,0,62,0,251,0,0,0,165,0,4,0,0,0,248,0,104,0,150,0,225,0,24,0,91,0,153,0,0,0,141,0,134,0,83,0,0,0,204,0,0,0,48,0,0,0,83,0,179,0,99,0,173,0,48,0,0,0,145,0,156,0,131,0,0,0,22,0,78,0,70,0,45,0,209,0,25,0,68,0,43,0,167,0,70,0,0,0,78,0,0,0,141,0,16,0,0,0,133,0,181,0,0,0,161,0,127,0,217,0,50,0,0,0,123,0,87,0,0,0,224,0,159,0,222,0,0,0,0,0,238,0,219,0,63,0,133,0,226,0,0,0,68,0,147,0,117,0,190,0,102,0,33,0,237,0,236,0,134,0,224,0,68,0,0,0,115,0,216,0,218,0,148,0,165,0,27,0,137,0,38,0,112,0,207,0,186,0,149,0,198,0,13,0,235,0,31,0,152,0,0,0,42,0,112,0,27,0,37,0,196,0,246,0,0,0,108,0,180,0,189,0,0,0,0,0,104,0,196,0,152,0,25,0,98,0,0,0,95,0,0,0,248,0,150,0,96,0,1,0,34,0,124,0,116,0,0,0,6,0,0,0,0,0,79,0,120,0,35,0,41,0,117,0,40,0,3,0,21,0,117,0,171,0,0,0,212,0,0,0,33,0,142,0,93,0,187,0,171,0,147,0,217,0,211,0,28,0,54,0,234,0,206,0,0,0,57,0,0,0,44,0,237,0,175,0,147,0,157,0,226,0,0,0,0,0,235,0,0,0,217,0,219,0,41,0,220,0,163,0,54,0,125,0,214,0,178,0,0,0,73,0,137,0,52,0,122,0,219,0,123,0,224,0,0,0,31,0,187,0,63,0,0,0,239,0,251,0,24,0,154,0,0,0,142,0,162,0,185,0,142,0,203,0,212,0,42,0,189,0,242,0,191,0,167,0,75,0,232,0,1,0,0,0,0,0,177,0,105,0,239,0,80,0,56,0,39,0,217,0,76,0,74,0,107,0,198,0,95,0,62,0,0,0,125,0,148,0,247,0,155,0,130,0,0,0,233,0,228,0,0,0,12,0,152,0,127,0,165,0,0,0,126,0,0,0,221,0,197,0,194,0,46,0,163,0,51,0,80,0,15,0,201,0,185,0,212,0,51,0,134,0,52,0,65,0,44,0,155,0,134,0,0,0,18,0,214,0,3,0,0,0,213,0,100,0,0,0,154,0,52,0,0,0,200,0,195,0,189,0,0,0,0,0,0,0,82,0,113,0,255,0,155,0,130,0,150,0,0,0,89,0,247,0,232,0,37,0,42,0,153,0,213,0,151,0,0,0,199,0,0,0,72,0,30,0,61,0,69,0,199,0,160,0,154,0,21,0,71,0,132,0,90,0,0,0,0,0,158,0,0,0,76,0,0,0,6,0,39,0,245,0,0,0,113,0,0,0,129,0,183,0,228,0,153,0,144,0,148,0,0,0,0,0,0,0,0,0,142,0,181,0,102,0,155,0,0,0,27,0,240,0,0,0,0,0,166,0,107,0,66,0,219,0,188,0,0,0,173,0,0,0,255,0,109,0,179,0,16,0,0,0,156,0,50,0,231,0,63,0,0,0,32,0,0,0,215,0,156,0,0,0,190,0,241,0,186,0,200,0,13,0,238,0,128,0,132,0,230,0,0,0,191,0,215,0,0,0,5,0,0,0,18,0,132,0,12,0,157,0,0,0,233,0,217,0,166,0,181,0,0,0,30,0,182,0,209,0,17,0,220,0,79,0,161,0,167,0,0,0,90,0,7,0,138,0,245,0,62,0,170,0,249,0,120,0,0,0,0,0,46,0,221,0,97,0,121,0,96,0,197,0,126,0,185,0,76,0,138,0,91,0,67,0,192,0,0,0,51,0,0,0,218,0,241,0,250,0,151,0,249,0,0,0,193,0,0,0,166,0,0,0,0,0,0,0,16,0,0,0,48,0,0,0,196,0,71,0,43,0,34,0,248,0,0,0,205,0,186,0,147,0,14,0,74,0,0,0,120,0,0,0,146,0,114,0,2,0,110,0,74,0,0,0,50,0,0,0,162,0,0,0,0,0,215,0,236,0,34,0,242,0,40,0,208,0,22,0,194,0,0,0,172,0,230,0,92,0,41,0,123,0,19,0,193,0,168,0,0,0,178,0,74,0,114,0,0,0,87,0,0,0,136,0,0,0,240,0,16,0,0,0,0,0,161,0,241,0,34,0,35,0,34,0,89,0,35,0,0,0,36,0,81,0,121,0,0,0,0,0,137,0,141,0,114,0,104,0,53,0,0,0,153,0,196,0,73,0,127,0,154,0,40,0,112,0,144,0,34,0,160,0,0,0,0,0,110,0,181,0,140,0,34,0,54,0,88,0,169,0,160,0,204,0,7,0,73,0,191,0,224,0,107,0,0,0,63,0,233,0,8,0,185,0,90,0,177,0,129,0,117,0,154,0,0,0,158,0,57,0,102,0,0,0,18,0,132,0,28,0,225,0,19,0,0,0,137,0,0,0,154,0,193,0,115,0,144,0,0,0,196,0,0,0,182,0,0,0,207,0,39,0,0,0,1,0,189,0,150,0,192,0,188,0,0,0,93,0,63,0,15,0,64,0,8,0,0,0,81,0,9,0,196,0,194,0,198,0,165,0,0,0,73,0,255,0,145,0,96,0,106,0,0,0,81,0,231,0,132,0,132,0,0,0,63,0,0,0,0,0,213,0,163,0,93,0,18,0,68,0,229,0,156,0,0,0,0,0,38,0,0,0,73,0,132,0,104,0,55,0,85,0);
signal scenario_full  : scenario_type := (0,0,56,31,56,30,229,31,208,31,208,30,208,29,227,31,38,31,2,31,170,31,107,31,178,31,178,30,178,29,178,28,63,31,36,31,195,31,249,31,97,31,131,31,191,31,214,31,157,31,241,31,114,31,130,31,145,31,204,31,204,30,149,31,50,31,222,31,2,31,255,31,236,31,156,31,83,31,68,31,2,31,2,30,222,31,222,30,178,31,111,31,200,31,231,31,231,30,193,31,194,31,150,31,91,31,93,31,214,31,31,31,109,31,250,31,250,30,47,31,62,31,251,31,251,30,165,31,4,31,4,30,248,31,104,31,150,31,225,31,24,31,91,31,153,31,153,30,141,31,134,31,83,31,83,30,204,31,204,30,48,31,48,30,83,31,179,31,99,31,173,31,48,31,48,30,145,31,156,31,131,31,131,30,22,31,78,31,70,31,45,31,209,31,25,31,68,31,43,31,167,31,70,31,70,30,78,31,78,30,141,31,16,31,16,30,133,31,181,31,181,30,161,31,127,31,217,31,50,31,50,30,123,31,87,31,87,30,224,31,159,31,222,31,222,30,222,29,238,31,219,31,63,31,133,31,226,31,226,30,68,31,147,31,117,31,190,31,102,31,33,31,237,31,236,31,134,31,224,31,68,31,68,30,115,31,216,31,218,31,148,31,165,31,27,31,137,31,38,31,112,31,207,31,186,31,149,31,198,31,13,31,235,31,31,31,152,31,152,30,42,31,112,31,27,31,37,31,196,31,246,31,246,30,108,31,180,31,189,31,189,30,189,29,104,31,196,31,152,31,25,31,98,31,98,30,95,31,95,30,248,31,150,31,96,31,1,31,34,31,124,31,116,31,116,30,6,31,6,30,6,29,79,31,120,31,35,31,41,31,117,31,40,31,3,31,21,31,117,31,171,31,171,30,212,31,212,30,33,31,142,31,93,31,187,31,171,31,147,31,217,31,211,31,28,31,54,31,234,31,206,31,206,30,57,31,57,30,44,31,237,31,175,31,147,31,157,31,226,31,226,30,226,29,235,31,235,30,217,31,219,31,41,31,220,31,163,31,54,31,125,31,214,31,178,31,178,30,73,31,137,31,52,31,122,31,219,31,123,31,224,31,224,30,31,31,187,31,63,31,63,30,239,31,251,31,24,31,154,31,154,30,142,31,162,31,185,31,142,31,203,31,212,31,42,31,189,31,242,31,191,31,167,31,75,31,232,31,1,31,1,30,1,29,177,31,105,31,239,31,80,31,56,31,39,31,217,31,76,31,74,31,107,31,198,31,95,31,62,31,62,30,125,31,148,31,247,31,155,31,130,31,130,30,233,31,228,31,228,30,12,31,152,31,127,31,165,31,165,30,126,31,126,30,221,31,197,31,194,31,46,31,163,31,51,31,80,31,15,31,201,31,185,31,212,31,51,31,134,31,52,31,65,31,44,31,155,31,134,31,134,30,18,31,214,31,3,31,3,30,213,31,100,31,100,30,154,31,52,31,52,30,200,31,195,31,189,31,189,30,189,29,189,28,82,31,113,31,255,31,155,31,130,31,150,31,150,30,89,31,247,31,232,31,37,31,42,31,153,31,213,31,151,31,151,30,199,31,199,30,72,31,30,31,61,31,69,31,199,31,160,31,154,31,21,31,71,31,132,31,90,31,90,30,90,29,158,31,158,30,76,31,76,30,6,31,39,31,245,31,245,30,113,31,113,30,129,31,183,31,228,31,153,31,144,31,148,31,148,30,148,29,148,28,148,27,142,31,181,31,102,31,155,31,155,30,27,31,240,31,240,30,240,29,166,31,107,31,66,31,219,31,188,31,188,30,173,31,173,30,255,31,109,31,179,31,16,31,16,30,156,31,50,31,231,31,63,31,63,30,32,31,32,30,215,31,156,31,156,30,190,31,241,31,186,31,200,31,13,31,238,31,128,31,132,31,230,31,230,30,191,31,215,31,215,30,5,31,5,30,18,31,132,31,12,31,157,31,157,30,233,31,217,31,166,31,181,31,181,30,30,31,182,31,209,31,17,31,220,31,79,31,161,31,167,31,167,30,90,31,7,31,138,31,245,31,62,31,170,31,249,31,120,31,120,30,120,29,46,31,221,31,97,31,121,31,96,31,197,31,126,31,185,31,76,31,138,31,91,31,67,31,192,31,192,30,51,31,51,30,218,31,241,31,250,31,151,31,249,31,249,30,193,31,193,30,166,31,166,30,166,29,166,28,16,31,16,30,48,31,48,30,196,31,71,31,43,31,34,31,248,31,248,30,205,31,186,31,147,31,14,31,74,31,74,30,120,31,120,30,146,31,114,31,2,31,110,31,74,31,74,30,50,31,50,30,162,31,162,30,162,29,215,31,236,31,34,31,242,31,40,31,208,31,22,31,194,31,194,30,172,31,230,31,92,31,41,31,123,31,19,31,193,31,168,31,168,30,178,31,74,31,114,31,114,30,87,31,87,30,136,31,136,30,240,31,16,31,16,30,16,29,161,31,241,31,34,31,35,31,34,31,89,31,35,31,35,30,36,31,81,31,121,31,121,30,121,29,137,31,141,31,114,31,104,31,53,31,53,30,153,31,196,31,73,31,127,31,154,31,40,31,112,31,144,31,34,31,160,31,160,30,160,29,110,31,181,31,140,31,34,31,54,31,88,31,169,31,160,31,204,31,7,31,73,31,191,31,224,31,107,31,107,30,63,31,233,31,8,31,185,31,90,31,177,31,129,31,117,31,154,31,154,30,158,31,57,31,102,31,102,30,18,31,132,31,28,31,225,31,19,31,19,30,137,31,137,30,154,31,193,31,115,31,144,31,144,30,196,31,196,30,182,31,182,30,207,31,39,31,39,30,1,31,189,31,150,31,192,31,188,31,188,30,93,31,63,31,15,31,64,31,8,31,8,30,81,31,9,31,196,31,194,31,198,31,165,31,165,30,73,31,255,31,145,31,96,31,106,31,106,30,81,31,231,31,132,31,132,31,132,30,63,31,63,30,63,29,213,31,163,31,93,31,18,31,68,31,229,31,156,31,156,30,156,29,38,31,38,30,73,31,132,31,104,31,55,31,85,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
