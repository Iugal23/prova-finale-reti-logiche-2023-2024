-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_765 is
end project_tb_765;

architecture project_tb_arch_765 of project_tb_765 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 324;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (144,0,230,0,0,0,0,0,153,0,193,0,55,0,0,0,108,0,62,0,205,0,76,0,147,0,89,0,72,0,88,0,104,0,51,0,105,0,0,0,0,0,0,0,102,0,179,0,169,0,17,0,21,0,140,0,0,0,47,0,0,0,174,0,97,0,102,0,193,0,0,0,0,0,197,0,0,0,169,0,0,0,93,0,253,0,145,0,221,0,71,0,0,0,253,0,149,0,72,0,0,0,59,0,46,0,152,0,146,0,59,0,34,0,0,0,0,0,203,0,149,0,165,0,135,0,99,0,106,0,0,0,25,0,213,0,143,0,141,0,232,0,0,0,209,0,236,0,0,0,0,0,41,0,0,0,109,0,26,0,0,0,106,0,162,0,155,0,195,0,28,0,57,0,200,0,121,0,233,0,46,0,176,0,125,0,81,0,33,0,143,0,46,0,116,0,192,0,118,0,170,0,184,0,174,0,0,0,10,0,68,0,148,0,93,0,159,0,193,0,164,0,136,0,0,0,136,0,0,0,46,0,83,0,174,0,0,0,127,0,0,0,55,0,236,0,155,0,33,0,106,0,94,0,202,0,0,0,0,0,93,0,0,0,0,0,125,0,60,0,0,0,161,0,203,0,16,0,63,0,186,0,233,0,58,0,161,0,104,0,0,0,250,0,143,0,24,0,151,0,103,0,47,0,0,0,119,0,143,0,211,0,240,0,0,0,250,0,0,0,225,0,53,0,236,0,35,0,208,0,192,0,106,0,126,0,0,0,0,0,248,0,59,0,239,0,188,0,56,0,174,0,97,0,237,0,137,0,253,0,138,0,0,0,75,0,0,0,36,0,33,0,65,0,0,0,0,0,183,0,108,0,248,0,0,0,159,0,0,0,63,0,246,0,212,0,151,0,0,0,0,0,221,0,0,0,75,0,243,0,144,0,156,0,120,0,252,0,167,0,72,0,104,0,158,0,0,0,112,0,37,0,154,0,130,0,254,0,169,0,10,0,201,0,204,0,160,0,168,0,76,0,123,0,155,0,18,0,232,0,228,0,217,0,0,0,0,0,247,0,125,0,35,0,0,0,237,0,242,0,217,0,0,0,12,0,8,0,204,0,0,0,72,0,198,0,217,0,187,0,230,0,17,0,196,0,102,0,84,0,147,0,114,0,165,0,99,0,46,0,79,0,117,0,165,0,77,0,195,0,4,0,223,0,86,0,39,0,35,0,44,0,243,0,0,0,130,0,0,0,134,0,203,0,61,0,52,0,31,0,122,0,102,0,151,0,130,0,13,0,145,0,68,0,224,0,0,0,0,0,0,0,124,0,0,0,118,0,4,0,135,0,251,0,92,0,59,0,139,0,99,0,234,0,133,0,118,0,1,0,89,0,230,0,0,0,181,0,143,0,3,0,37,0,248,0,181,0,109,0,161,0,170,0,170,0,156,0,129,0,91,0,142,0,97,0,222,0);
signal scenario_full  : scenario_type := (144,31,230,31,230,30,230,29,153,31,193,31,55,31,55,30,108,31,62,31,205,31,76,31,147,31,89,31,72,31,88,31,104,31,51,31,105,31,105,30,105,29,105,28,102,31,179,31,169,31,17,31,21,31,140,31,140,30,47,31,47,30,174,31,97,31,102,31,193,31,193,30,193,29,197,31,197,30,169,31,169,30,93,31,253,31,145,31,221,31,71,31,71,30,253,31,149,31,72,31,72,30,59,31,46,31,152,31,146,31,59,31,34,31,34,30,34,29,203,31,149,31,165,31,135,31,99,31,106,31,106,30,25,31,213,31,143,31,141,31,232,31,232,30,209,31,236,31,236,30,236,29,41,31,41,30,109,31,26,31,26,30,106,31,162,31,155,31,195,31,28,31,57,31,200,31,121,31,233,31,46,31,176,31,125,31,81,31,33,31,143,31,46,31,116,31,192,31,118,31,170,31,184,31,174,31,174,30,10,31,68,31,148,31,93,31,159,31,193,31,164,31,136,31,136,30,136,31,136,30,46,31,83,31,174,31,174,30,127,31,127,30,55,31,236,31,155,31,33,31,106,31,94,31,202,31,202,30,202,29,93,31,93,30,93,29,125,31,60,31,60,30,161,31,203,31,16,31,63,31,186,31,233,31,58,31,161,31,104,31,104,30,250,31,143,31,24,31,151,31,103,31,47,31,47,30,119,31,143,31,211,31,240,31,240,30,250,31,250,30,225,31,53,31,236,31,35,31,208,31,192,31,106,31,126,31,126,30,126,29,248,31,59,31,239,31,188,31,56,31,174,31,97,31,237,31,137,31,253,31,138,31,138,30,75,31,75,30,36,31,33,31,65,31,65,30,65,29,183,31,108,31,248,31,248,30,159,31,159,30,63,31,246,31,212,31,151,31,151,30,151,29,221,31,221,30,75,31,243,31,144,31,156,31,120,31,252,31,167,31,72,31,104,31,158,31,158,30,112,31,37,31,154,31,130,31,254,31,169,31,10,31,201,31,204,31,160,31,168,31,76,31,123,31,155,31,18,31,232,31,228,31,217,31,217,30,217,29,247,31,125,31,35,31,35,30,237,31,242,31,217,31,217,30,12,31,8,31,204,31,204,30,72,31,198,31,217,31,187,31,230,31,17,31,196,31,102,31,84,31,147,31,114,31,165,31,99,31,46,31,79,31,117,31,165,31,77,31,195,31,4,31,223,31,86,31,39,31,35,31,44,31,243,31,243,30,130,31,130,30,134,31,203,31,61,31,52,31,31,31,122,31,102,31,151,31,130,31,13,31,145,31,68,31,224,31,224,30,224,29,224,28,124,31,124,30,118,31,4,31,135,31,251,31,92,31,59,31,139,31,99,31,234,31,133,31,118,31,1,31,89,31,230,31,230,30,181,31,143,31,3,31,37,31,248,31,181,31,109,31,161,31,170,31,170,31,156,31,129,31,91,31,142,31,97,31,222,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
