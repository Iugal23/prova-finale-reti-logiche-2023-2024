-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1014;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (200,0,0,0,0,0,145,0,195,0,0,0,200,0,0,0,21,0,178,0,116,0,118,0,0,0,0,0,42,0,0,0,215,0,245,0,206,0,42,0,128,0,105,0,0,0,0,0,69,0,166,0,221,0,52,0,214,0,0,0,55,0,0,0,204,0,97,0,154,0,41,0,122,0,85,0,0,0,183,0,161,0,156,0,0,0,0,0,227,0,94,0,88,0,0,0,237,0,179,0,85,0,39,0,29,0,86,0,0,0,110,0,149,0,41,0,181,0,0,0,39,0,100,0,131,0,0,0,14,0,212,0,0,0,90,0,42,0,0,0,0,0,158,0,159,0,130,0,56,0,87,0,169,0,137,0,149,0,21,0,124,0,50,0,0,0,154,0,234,0,54,0,205,0,125,0,159,0,0,0,50,0,219,0,255,0,232,0,232,0,51,0,210,0,184,0,0,0,0,0,103,0,159,0,63,0,0,0,170,0,218,0,155,0,189,0,0,0,168,0,215,0,0,0,0,0,187,0,76,0,19,0,223,0,173,0,222,0,38,0,0,0,149,0,179,0,110,0,117,0,233,0,0,0,0,0,242,0,73,0,120,0,147,0,146,0,188,0,145,0,146,0,7,0,77,0,214,0,0,0,0,0,232,0,45,0,175,0,25,0,117,0,45,0,150,0,218,0,7,0,58,0,2,0,7,0,91,0,143,0,28,0,0,0,218,0,73,0,195,0,217,0,0,0,96,0,244,0,222,0,53,0,177,0,44,0,0,0,140,0,0,0,219,0,52,0,165,0,221,0,0,0,0,0,68,0,0,0,129,0,58,0,0,0,21,0,0,0,66,0,133,0,20,0,124,0,20,0,0,0,0,0,207,0,0,0,172,0,250,0,172,0,117,0,14,0,81,0,35,0,82,0,13,0,199,0,133,0,209,0,0,0,224,0,90,0,42,0,98,0,69,0,151,0,236,0,215,0,15,0,237,0,229,0,150,0,88,0,148,0,49,0,0,0,0,0,192,0,0,0,237,0,3,0,0,0,161,0,0,0,0,0,183,0,151,0,174,0,135,0,49,0,0,0,15,0,0,0,251,0,0,0,104,0,181,0,244,0,0,0,0,0,245,0,0,0,0,0,195,0,158,0,220,0,0,0,95,0,0,0,205,0,0,0,212,0,228,0,218,0,48,0,0,0,199,0,0,0,201,0,46,0,0,0,143,0,198,0,211,0,244,0,117,0,234,0,199,0,155,0,77,0,106,0,114,0,128,0,0,0,35,0,0,0,52,0,184,0,247,0,0,0,0,0,0,0,126,0,0,0,176,0,0,0,226,0,8,0,92,0,161,0,255,0,33,0,0,0,95,0,57,0,44,0,233,0,186,0,191,0,199,0,222,0,110,0,0,0,141,0,16,0,11,0,95,0,84,0,222,0,23,0,46,0,232,0,0,0,91,0,0,0,168,0,0,0,0,0,202,0,0,0,249,0,47,0,105,0,209,0,53,0,68,0,209,0,40,0,0,0,42,0,48,0,82,0,95,0,188,0,228,0,45,0,190,0,142,0,0,0,19,0,170,0,159,0,128,0,151,0,0,0,21,0,56,0,224,0,176,0,54,0,0,0,35,0,0,0,0,0,206,0,220,0,68,0,9,0,0,0,215,0,196,0,90,0,216,0,167,0,0,0,58,0,160,0,24,0,27,0,54,0,0,0,231,0,114,0,57,0,152,0,180,0,117,0,180,0,0,0,202,0,21,0,130,0,0,0,0,0,0,0,150,0,1,0,103,0,158,0,48,0,19,0,0,0,210,0,17,0,63,0,44,0,106,0,0,0,221,0,9,0,242,0,10,0,0,0,0,0,31,0,0,0,0,0,215,0,0,0,86,0,254,0,164,0,1,0,155,0,166,0,133,0,187,0,40,0,224,0,78,0,233,0,113,0,77,0,80,0,0,0,180,0,252,0,238,0,60,0,41,0,57,0,0,0,0,0,225,0,49,0,226,0,150,0,53,0,133,0,16,0,165,0,205,0,200,0,134,0,136,0,74,0,230,0,218,0,227,0,175,0,0,0,27,0,239,0,168,0,193,0,108,0,240,0,208,0,248,0,220,0,169,0,110,0,110,0,49,0,0,0,0,0,82,0,67,0,179,0,104,0,63,0,172,0,157,0,138,0,0,0,0,0,231,0,79,0,105,0,43,0,81,0,0,0,50,0,0,0,0,0,68,0,128,0,218,0,156,0,201,0,22,0,103,0,173,0,45,0,6,0,116,0,22,0,203,0,0,0,96,0,195,0,111,0,60,0,234,0,101,0,0,0,19,0,15,0,219,0,76,0,216,0,58,0,54,0,146,0,157,0,132,0,227,0,0,0,73,0,0,0,189,0,110,0,30,0,0,0,254,0,69,0,224,0,214,0,37,0,151,0,143,0,138,0,46,0,240,0,132,0,46,0,65,0,23,0,0,0,0,0,81,0,0,0,29,0,0,0,0,0,156,0,0,0,156,0,16,0,53,0,0,0,113,0,0,0,92,0,49,0,215,0,0,0,59,0,141,0,0,0,143,0,219,0,140,0,0,0,185,0,215,0,143,0,65,0,0,0,250,0,0,0,148,0,211,0,0,0,117,0,0,0,117,0,29,0,255,0,60,0,0,0,148,0,79,0,13,0,0,0,253,0,41,0,167,0,10,0,0,0,60,0,23,0,0,0,77,0,247,0,11,0,0,0,3,0,0,0,0,0,251,0,86,0,0,0,0,0,214,0,76,0,0,0,133,0,0,0,184,0,124,0,238,0,0,0,136,0,139,0,201,0,14,0,0,0,212,0,0,0,0,0,40,0,191,0,18,0,184,0,204,0,212,0,249,0,160,0,180,0,136,0,138,0,138,0,93,0,80,0,0,0,0,0,31,0,101,0,173,0,25,0,121,0,20,0,115,0,44,0,31,0,105,0,0,0,183,0,120,0,104,0,238,0,16,0,34,0,38,0,112,0,92,0,116,0,240,0,176,0,0,0,137,0,208,0,159,0,29,0,0,0,247,0,45,0,153,0,242,0,129,0,164,0,205,0,187,0,145,0,0,0,162,0,136,0,68,0,231,0,10,0,2,0,147,0,63,0,176,0,78,0,186,0,9,0,117,0,55,0,70,0,129,0,13,0,210,0,246,0,5,0,6,0,250,0,0,0,127,0,178,0,40,0,33,0,194,0,172,0,0,0,0,0,114,0,0,0,108,0,138,0,138,0,0,0,26,0,37,0,219,0,0,0,25,0,252,0,0,0,252,0,185,0,0,0,130,0,4,0,0,0,73,0,0,0,21,0,50,0,167,0,18,0,158,0,0,0,160,0,116,0,108,0,0,0,23,0,154,0,238,0,0,0,94,0,0,0,231,0,0,0,156,0,137,0,230,0,186,0,0,0,113,0,59,0,0,0,221,0,85,0,118,0,221,0,124,0,64,0,45,0,215,0,0,0,0,0,48,0,57,0,5,0,0,0,203,0,176,0,160,0,160,0,0,0,0,0,230,0,168,0,254,0,107,0,80,0,179,0,132,0,115,0,0,0,36,0,117,0,183,0,190,0,16,0,16,0,18,0,98,0,23,0,209,0,209,0,123,0,0,0,72,0,143,0,69,0,0,0,118,0,173,0,180,0,20,0,27,0,0,0,231,0,134,0,249,0,0,0,158,0,62,0,66,0,117,0,122,0,247,0,81,0,191,0,0,0,76,0,157,0,253,0,122,0,182,0,53,0,0,0,131,0,137,0,164,0,95,0,114,0,4,0,111,0,0,0,156,0,134,0,0,0,0,0,245,0,0,0,39,0,124,0,252,0,114,0,61,0,210,0,225,0,0,0,0,0,0,0,0,0,109,0,0,0,0,0,69,0,227,0,0,0,124,0,26,0,201,0,184,0,50,0,159,0,142,0,119,0,39,0,0,0,0,0,32,0,0,0,104,0,237,0,178,0,196,0,111,0,153,0,114,0,82,0,0,0,119,0,0,0,0,0,109,0,94,0,0,0,38,0,0,0,0,0,249,0,0,0,19,0,0,0,0,0,142,0,0,0,236,0,89,0,0,0,13,0,57,0,137,0,35,0,0,0,247,0,0,0,105,0,225,0,232,0,186,0,112,0,15,0,209,0,161,0,0,0,169,0,29,0,0,0,231,0,119,0,0,0,45,0,0,0,0,0,157,0,0,0,229,0,0,0,245,0,212,0,80,0,46,0,178,0,24,0,0,0,78,0,125,0,26,0,0,0,134,0,153,0,163,0,233,0,101,0,242,0,96,0,71,0,119,0,11,0,81,0,93,0,28,0,214,0,62,0,112,0,10,0,0,0,48,0,254,0,37,0,51,0,0,0,195,0,171,0,0,0,95,0,0,0,207,0,220,0,0,0,0,0,102,0,0,0,0,0,142,0,243,0,230,0,0,0,0,0,101,0,32,0,0,0,0,0,39,0,67,0,141,0,128,0,25,0,7,0,88,0,35,0,190,0,73,0,13,0,85,0,8,0,68,0,216,0,141,0,0,0,0,0,207,0,108,0,0,0,33,0,0,0,141,0,189,0,24,0);
signal scenario_full  : scenario_type := (200,31,200,30,200,29,145,31,195,31,195,30,200,31,200,30,21,31,178,31,116,31,118,31,118,30,118,29,42,31,42,30,215,31,245,31,206,31,42,31,128,31,105,31,105,30,105,29,69,31,166,31,221,31,52,31,214,31,214,30,55,31,55,30,204,31,97,31,154,31,41,31,122,31,85,31,85,30,183,31,161,31,156,31,156,30,156,29,227,31,94,31,88,31,88,30,237,31,179,31,85,31,39,31,29,31,86,31,86,30,110,31,149,31,41,31,181,31,181,30,39,31,100,31,131,31,131,30,14,31,212,31,212,30,90,31,42,31,42,30,42,29,158,31,159,31,130,31,56,31,87,31,169,31,137,31,149,31,21,31,124,31,50,31,50,30,154,31,234,31,54,31,205,31,125,31,159,31,159,30,50,31,219,31,255,31,232,31,232,31,51,31,210,31,184,31,184,30,184,29,103,31,159,31,63,31,63,30,170,31,218,31,155,31,189,31,189,30,168,31,215,31,215,30,215,29,187,31,76,31,19,31,223,31,173,31,222,31,38,31,38,30,149,31,179,31,110,31,117,31,233,31,233,30,233,29,242,31,73,31,120,31,147,31,146,31,188,31,145,31,146,31,7,31,77,31,214,31,214,30,214,29,232,31,45,31,175,31,25,31,117,31,45,31,150,31,218,31,7,31,58,31,2,31,7,31,91,31,143,31,28,31,28,30,218,31,73,31,195,31,217,31,217,30,96,31,244,31,222,31,53,31,177,31,44,31,44,30,140,31,140,30,219,31,52,31,165,31,221,31,221,30,221,29,68,31,68,30,129,31,58,31,58,30,21,31,21,30,66,31,133,31,20,31,124,31,20,31,20,30,20,29,207,31,207,30,172,31,250,31,172,31,117,31,14,31,81,31,35,31,82,31,13,31,199,31,133,31,209,31,209,30,224,31,90,31,42,31,98,31,69,31,151,31,236,31,215,31,15,31,237,31,229,31,150,31,88,31,148,31,49,31,49,30,49,29,192,31,192,30,237,31,3,31,3,30,161,31,161,30,161,29,183,31,151,31,174,31,135,31,49,31,49,30,15,31,15,30,251,31,251,30,104,31,181,31,244,31,244,30,244,29,245,31,245,30,245,29,195,31,158,31,220,31,220,30,95,31,95,30,205,31,205,30,212,31,228,31,218,31,48,31,48,30,199,31,199,30,201,31,46,31,46,30,143,31,198,31,211,31,244,31,117,31,234,31,199,31,155,31,77,31,106,31,114,31,128,31,128,30,35,31,35,30,52,31,184,31,247,31,247,30,247,29,247,28,126,31,126,30,176,31,176,30,226,31,8,31,92,31,161,31,255,31,33,31,33,30,95,31,57,31,44,31,233,31,186,31,191,31,199,31,222,31,110,31,110,30,141,31,16,31,11,31,95,31,84,31,222,31,23,31,46,31,232,31,232,30,91,31,91,30,168,31,168,30,168,29,202,31,202,30,249,31,47,31,105,31,209,31,53,31,68,31,209,31,40,31,40,30,42,31,48,31,82,31,95,31,188,31,228,31,45,31,190,31,142,31,142,30,19,31,170,31,159,31,128,31,151,31,151,30,21,31,56,31,224,31,176,31,54,31,54,30,35,31,35,30,35,29,206,31,220,31,68,31,9,31,9,30,215,31,196,31,90,31,216,31,167,31,167,30,58,31,160,31,24,31,27,31,54,31,54,30,231,31,114,31,57,31,152,31,180,31,117,31,180,31,180,30,202,31,21,31,130,31,130,30,130,29,130,28,150,31,1,31,103,31,158,31,48,31,19,31,19,30,210,31,17,31,63,31,44,31,106,31,106,30,221,31,9,31,242,31,10,31,10,30,10,29,31,31,31,30,31,29,215,31,215,30,86,31,254,31,164,31,1,31,155,31,166,31,133,31,187,31,40,31,224,31,78,31,233,31,113,31,77,31,80,31,80,30,180,31,252,31,238,31,60,31,41,31,57,31,57,30,57,29,225,31,49,31,226,31,150,31,53,31,133,31,16,31,165,31,205,31,200,31,134,31,136,31,74,31,230,31,218,31,227,31,175,31,175,30,27,31,239,31,168,31,193,31,108,31,240,31,208,31,248,31,220,31,169,31,110,31,110,31,49,31,49,30,49,29,82,31,67,31,179,31,104,31,63,31,172,31,157,31,138,31,138,30,138,29,231,31,79,31,105,31,43,31,81,31,81,30,50,31,50,30,50,29,68,31,128,31,218,31,156,31,201,31,22,31,103,31,173,31,45,31,6,31,116,31,22,31,203,31,203,30,96,31,195,31,111,31,60,31,234,31,101,31,101,30,19,31,15,31,219,31,76,31,216,31,58,31,54,31,146,31,157,31,132,31,227,31,227,30,73,31,73,30,189,31,110,31,30,31,30,30,254,31,69,31,224,31,214,31,37,31,151,31,143,31,138,31,46,31,240,31,132,31,46,31,65,31,23,31,23,30,23,29,81,31,81,30,29,31,29,30,29,29,156,31,156,30,156,31,16,31,53,31,53,30,113,31,113,30,92,31,49,31,215,31,215,30,59,31,141,31,141,30,143,31,219,31,140,31,140,30,185,31,215,31,143,31,65,31,65,30,250,31,250,30,148,31,211,31,211,30,117,31,117,30,117,31,29,31,255,31,60,31,60,30,148,31,79,31,13,31,13,30,253,31,41,31,167,31,10,31,10,30,60,31,23,31,23,30,77,31,247,31,11,31,11,30,3,31,3,30,3,29,251,31,86,31,86,30,86,29,214,31,76,31,76,30,133,31,133,30,184,31,124,31,238,31,238,30,136,31,139,31,201,31,14,31,14,30,212,31,212,30,212,29,40,31,191,31,18,31,184,31,204,31,212,31,249,31,160,31,180,31,136,31,138,31,138,31,93,31,80,31,80,30,80,29,31,31,101,31,173,31,25,31,121,31,20,31,115,31,44,31,31,31,105,31,105,30,183,31,120,31,104,31,238,31,16,31,34,31,38,31,112,31,92,31,116,31,240,31,176,31,176,30,137,31,208,31,159,31,29,31,29,30,247,31,45,31,153,31,242,31,129,31,164,31,205,31,187,31,145,31,145,30,162,31,136,31,68,31,231,31,10,31,2,31,147,31,63,31,176,31,78,31,186,31,9,31,117,31,55,31,70,31,129,31,13,31,210,31,246,31,5,31,6,31,250,31,250,30,127,31,178,31,40,31,33,31,194,31,172,31,172,30,172,29,114,31,114,30,108,31,138,31,138,31,138,30,26,31,37,31,219,31,219,30,25,31,252,31,252,30,252,31,185,31,185,30,130,31,4,31,4,30,73,31,73,30,21,31,50,31,167,31,18,31,158,31,158,30,160,31,116,31,108,31,108,30,23,31,154,31,238,31,238,30,94,31,94,30,231,31,231,30,156,31,137,31,230,31,186,31,186,30,113,31,59,31,59,30,221,31,85,31,118,31,221,31,124,31,64,31,45,31,215,31,215,30,215,29,48,31,57,31,5,31,5,30,203,31,176,31,160,31,160,31,160,30,160,29,230,31,168,31,254,31,107,31,80,31,179,31,132,31,115,31,115,30,36,31,117,31,183,31,190,31,16,31,16,31,18,31,98,31,23,31,209,31,209,31,123,31,123,30,72,31,143,31,69,31,69,30,118,31,173,31,180,31,20,31,27,31,27,30,231,31,134,31,249,31,249,30,158,31,62,31,66,31,117,31,122,31,247,31,81,31,191,31,191,30,76,31,157,31,253,31,122,31,182,31,53,31,53,30,131,31,137,31,164,31,95,31,114,31,4,31,111,31,111,30,156,31,134,31,134,30,134,29,245,31,245,30,39,31,124,31,252,31,114,31,61,31,210,31,225,31,225,30,225,29,225,28,225,27,109,31,109,30,109,29,69,31,227,31,227,30,124,31,26,31,201,31,184,31,50,31,159,31,142,31,119,31,39,31,39,30,39,29,32,31,32,30,104,31,237,31,178,31,196,31,111,31,153,31,114,31,82,31,82,30,119,31,119,30,119,29,109,31,94,31,94,30,38,31,38,30,38,29,249,31,249,30,19,31,19,30,19,29,142,31,142,30,236,31,89,31,89,30,13,31,57,31,137,31,35,31,35,30,247,31,247,30,105,31,225,31,232,31,186,31,112,31,15,31,209,31,161,31,161,30,169,31,29,31,29,30,231,31,119,31,119,30,45,31,45,30,45,29,157,31,157,30,229,31,229,30,245,31,212,31,80,31,46,31,178,31,24,31,24,30,78,31,125,31,26,31,26,30,134,31,153,31,163,31,233,31,101,31,242,31,96,31,71,31,119,31,11,31,81,31,93,31,28,31,214,31,62,31,112,31,10,31,10,30,48,31,254,31,37,31,51,31,51,30,195,31,171,31,171,30,95,31,95,30,207,31,220,31,220,30,220,29,102,31,102,30,102,29,142,31,243,31,230,31,230,30,230,29,101,31,32,31,32,30,32,29,39,31,67,31,141,31,128,31,25,31,7,31,88,31,35,31,190,31,73,31,13,31,85,31,8,31,68,31,216,31,141,31,141,30,141,29,207,31,108,31,108,30,33,31,33,30,141,31,189,31,24,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
