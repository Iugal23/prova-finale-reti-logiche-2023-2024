-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_439 is
end project_tb_439;

architecture project_tb_arch_439 of project_tb_439 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 522;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,144,0,70,0,254,0,82,0,243,0,99,0,237,0,84,0,232,0,179,0,102,0,32,0,248,0,150,0,137,0,203,0,0,0,0,0,109,0,0,0,152,0,0,0,78,0,46,0,212,0,219,0,73,0,167,0,11,0,27,0,225,0,0,0,16,0,59,0,228,0,242,0,247,0,0,0,227,0,0,0,167,0,0,0,174,0,124,0,7,0,91,0,78,0,82,0,54,0,0,0,224,0,106,0,75,0,0,0,0,0,151,0,223,0,104,0,0,0,79,0,0,0,141,0,17,0,236,0,8,0,113,0,217,0,117,0,41,0,94,0,221,0,43,0,119,0,52,0,53,0,178,0,112,0,154,0,0,0,239,0,192,0,204,0,237,0,239,0,98,0,65,0,0,0,0,0,18,0,0,0,65,0,192,0,243,0,215,0,0,0,0,0,128,0,84,0,0,0,125,0,89,0,188,0,235,0,55,0,220,0,40,0,95,0,19,0,244,0,212,0,97,0,77,0,0,0,0,0,181,0,58,0,0,0,119,0,0,0,131,0,14,0,163,0,243,0,255,0,25,0,170,0,76,0,139,0,0,0,103,0,0,0,232,0,165,0,37,0,106,0,186,0,0,0,175,0,0,0,0,0,65,0,155,0,18,0,161,0,216,0,0,0,47,0,36,0,0,0,212,0,0,0,198,0,192,0,107,0,226,0,0,0,126,0,79,0,0,0,136,0,79,0,81,0,103,0,99,0,131,0,138,0,84,0,43,0,154,0,136,0,120,0,14,0,0,0,0,0,96,0,24,0,135,0,158,0,53,0,140,0,242,0,15,0,56,0,185,0,245,0,14,0,226,0,233,0,44,0,86,0,0,0,140,0,74,0,0,0,169,0,108,0,160,0,129,0,0,0,108,0,27,0,0,0,180,0,30,0,0,0,0,0,141,0,0,0,0,0,57,0,106,0,160,0,218,0,171,0,0,0,0,0,117,0,74,0,229,0,205,0,205,0,2,0,246,0,165,0,120,0,244,0,84,0,179,0,247,0,37,0,51,0,0,0,0,0,224,0,182,0,66,0,67,0,0,0,247,0,162,0,42,0,152,0,166,0,42,0,191,0,33,0,147,0,59,0,164,0,0,0,90,0,27,0,208,0,159,0,205,0,180,0,231,0,172,0,212,0,245,0,0,0,191,0,140,0,26,0,60,0,138,0,21,0,87,0,0,0,187,0,0,0,254,0,44,0,70,0,225,0,0,0,105,0,212,0,56,0,70,0,138,0,247,0,0,0,0,0,0,0,255,0,105,0,90,0,60,0,180,0,162,0,0,0,0,0,201,0,0,0,0,0,208,0,74,0,4,0,193,0,116,0,30,0,142,0,88,0,202,0,121,0,69,0,0,0,0,0,253,0,10,0,155,0,168,0,12,0,84,0,175,0,36,0,35,0,243,0,127,0,252,0,117,0,99,0,0,0,10,0,0,0,0,0,0,0,237,0,215,0,132,0,152,0,0,0,51,0,27,0,2,0,0,0,105,0,0,0,74,0,229,0,97,0,136,0,78,0,189,0,20,0,73,0,255,0,55,0,177,0,41,0,238,0,72,0,156,0,32,0,0,0,31,0,178,0,215,0,176,0,143,0,207,0,70,0,0,0,216,0,47,0,201,0,79,0,105,0,159,0,0,0,0,0,152,0,236,0,12,0,228,0,108,0,56,0,0,0,105,0,60,0,0,0,0,0,57,0,163,0,153,0,245,0,150,0,0,0,0,0,188,0,28,0,24,0,0,0,114,0,123,0,0,0,191,0,117,0,228,0,202,0,53,0,182,0,0,0,49,0,104,0,54,0,70,0,78,0,0,0,188,0,179,0,130,0,7,0,0,0,0,0,0,0,42,0,104,0,133,0,2,0,132,0,210,0,0,0,247,0,28,0,197,0,0,0,0,0,81,0,207,0,95,0,154,0,139,0,0,0,89,0,158,0,251,0,0,0,244,0,113,0,0,0,69,0,186,0,0,0,43,0,18,0,181,0,47,0,131,0,69,0,238,0,9,0,11,0,117,0,169,0,178,0,63,0,154,0,26,0,55,0,145,0,173,0,92,0,139,0,0,0,89,0,227,0,0,0,84,0,170,0,243,0,77,0,233,0,0,0,0,0,198,0,123,0,0,0,214,0,32,0,36,0,59,0,67,0,0,0,108,0,216,0,85,0,0,0,85,0,169,0,65,0,46,0,184,0,162,0,0,0,0,0,67,0,0,0,163,0,0,0,0,0,180,0,123,0,242,0,0,0,0,0,4,0,207,0,248,0,100,0,64,0,126,0,16,0,153,0,117,0,216,0,105,0,24,0,156,0,237,0);
signal scenario_full  : scenario_type := (0,0,144,31,70,31,254,31,82,31,243,31,99,31,237,31,84,31,232,31,179,31,102,31,32,31,248,31,150,31,137,31,203,31,203,30,203,29,109,31,109,30,152,31,152,30,78,31,46,31,212,31,219,31,73,31,167,31,11,31,27,31,225,31,225,30,16,31,59,31,228,31,242,31,247,31,247,30,227,31,227,30,167,31,167,30,174,31,124,31,7,31,91,31,78,31,82,31,54,31,54,30,224,31,106,31,75,31,75,30,75,29,151,31,223,31,104,31,104,30,79,31,79,30,141,31,17,31,236,31,8,31,113,31,217,31,117,31,41,31,94,31,221,31,43,31,119,31,52,31,53,31,178,31,112,31,154,31,154,30,239,31,192,31,204,31,237,31,239,31,98,31,65,31,65,30,65,29,18,31,18,30,65,31,192,31,243,31,215,31,215,30,215,29,128,31,84,31,84,30,125,31,89,31,188,31,235,31,55,31,220,31,40,31,95,31,19,31,244,31,212,31,97,31,77,31,77,30,77,29,181,31,58,31,58,30,119,31,119,30,131,31,14,31,163,31,243,31,255,31,25,31,170,31,76,31,139,31,139,30,103,31,103,30,232,31,165,31,37,31,106,31,186,31,186,30,175,31,175,30,175,29,65,31,155,31,18,31,161,31,216,31,216,30,47,31,36,31,36,30,212,31,212,30,198,31,192,31,107,31,226,31,226,30,126,31,79,31,79,30,136,31,79,31,81,31,103,31,99,31,131,31,138,31,84,31,43,31,154,31,136,31,120,31,14,31,14,30,14,29,96,31,24,31,135,31,158,31,53,31,140,31,242,31,15,31,56,31,185,31,245,31,14,31,226,31,233,31,44,31,86,31,86,30,140,31,74,31,74,30,169,31,108,31,160,31,129,31,129,30,108,31,27,31,27,30,180,31,30,31,30,30,30,29,141,31,141,30,141,29,57,31,106,31,160,31,218,31,171,31,171,30,171,29,117,31,74,31,229,31,205,31,205,31,2,31,246,31,165,31,120,31,244,31,84,31,179,31,247,31,37,31,51,31,51,30,51,29,224,31,182,31,66,31,67,31,67,30,247,31,162,31,42,31,152,31,166,31,42,31,191,31,33,31,147,31,59,31,164,31,164,30,90,31,27,31,208,31,159,31,205,31,180,31,231,31,172,31,212,31,245,31,245,30,191,31,140,31,26,31,60,31,138,31,21,31,87,31,87,30,187,31,187,30,254,31,44,31,70,31,225,31,225,30,105,31,212,31,56,31,70,31,138,31,247,31,247,30,247,29,247,28,255,31,105,31,90,31,60,31,180,31,162,31,162,30,162,29,201,31,201,30,201,29,208,31,74,31,4,31,193,31,116,31,30,31,142,31,88,31,202,31,121,31,69,31,69,30,69,29,253,31,10,31,155,31,168,31,12,31,84,31,175,31,36,31,35,31,243,31,127,31,252,31,117,31,99,31,99,30,10,31,10,30,10,29,10,28,237,31,215,31,132,31,152,31,152,30,51,31,27,31,2,31,2,30,105,31,105,30,74,31,229,31,97,31,136,31,78,31,189,31,20,31,73,31,255,31,55,31,177,31,41,31,238,31,72,31,156,31,32,31,32,30,31,31,178,31,215,31,176,31,143,31,207,31,70,31,70,30,216,31,47,31,201,31,79,31,105,31,159,31,159,30,159,29,152,31,236,31,12,31,228,31,108,31,56,31,56,30,105,31,60,31,60,30,60,29,57,31,163,31,153,31,245,31,150,31,150,30,150,29,188,31,28,31,24,31,24,30,114,31,123,31,123,30,191,31,117,31,228,31,202,31,53,31,182,31,182,30,49,31,104,31,54,31,70,31,78,31,78,30,188,31,179,31,130,31,7,31,7,30,7,29,7,28,42,31,104,31,133,31,2,31,132,31,210,31,210,30,247,31,28,31,197,31,197,30,197,29,81,31,207,31,95,31,154,31,139,31,139,30,89,31,158,31,251,31,251,30,244,31,113,31,113,30,69,31,186,31,186,30,43,31,18,31,181,31,47,31,131,31,69,31,238,31,9,31,11,31,117,31,169,31,178,31,63,31,154,31,26,31,55,31,145,31,173,31,92,31,139,31,139,30,89,31,227,31,227,30,84,31,170,31,243,31,77,31,233,31,233,30,233,29,198,31,123,31,123,30,214,31,32,31,36,31,59,31,67,31,67,30,108,31,216,31,85,31,85,30,85,31,169,31,65,31,46,31,184,31,162,31,162,30,162,29,67,31,67,30,163,31,163,30,163,29,180,31,123,31,242,31,242,30,242,29,4,31,207,31,248,31,100,31,64,31,126,31,16,31,153,31,117,31,216,31,105,31,24,31,156,31,237,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
