-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_701 is
end project_tb_701;

architecture project_tb_arch_701 of project_tb_701 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 767;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (116,0,221,0,34,0,0,0,0,0,48,0,200,0,202,0,121,0,248,0,55,0,244,0,77,0,138,0,188,0,18,0,0,0,139,0,17,0,29,0,5,0,0,0,216,0,151,0,0,0,84,0,237,0,23,0,0,0,0,0,44,0,0,0,165,0,104,0,162,0,103,0,174,0,0,0,81,0,131,0,138,0,152,0,200,0,166,0,39,0,88,0,0,0,137,0,0,0,190,0,39,0,46,0,42,0,123,0,43,0,100,0,37,0,0,0,109,0,114,0,159,0,78,0,163,0,220,0,129,0,230,0,124,0,0,0,19,0,122,0,200,0,85,0,84,0,25,0,167,0,247,0,42,0,148,0,246,0,0,0,44,0,0,0,3,0,41,0,68,0,45,0,105,0,0,0,32,0,221,0,117,0,191,0,220,0,144,0,97,0,217,0,90,0,107,0,202,0,0,0,0,0,108,0,6,0,22,0,107,0,145,0,180,0,197,0,189,0,54,0,216,0,176,0,100,0,89,0,136,0,158,0,239,0,253,0,195,0,202,0,15,0,0,0,0,0,53,0,145,0,219,0,0,0,172,0,153,0,90,0,0,0,67,0,203,0,19,0,0,0,113,0,101,0,59,0,32,0,0,0,102,0,188,0,0,0,90,0,201,0,176,0,214,0,220,0,221,0,96,0,159,0,103,0,79,0,153,0,0,0,0,0,147,0,16,0,133,0,29,0,156,0,103,0,211,0,0,0,243,0,0,0,56,0,93,0,61,0,34,0,182,0,0,0,151,0,117,0,55,0,0,0,74,0,23,0,0,0,170,0,0,0,129,0,80,0,64,0,99,0,115,0,119,0,83,0,230,0,231,0,186,0,224,0,108,0,130,0,231,0,142,0,189,0,235,0,187,0,220,0,251,0,160,0,0,0,0,0,19,0,209,0,254,0,173,0,0,0,187,0,0,0,251,0,228,0,223,0,196,0,181,0,74,0,0,0,108,0,24,0,145,0,0,0,180,0,212,0,22,0,0,0,45,0,5,0,200,0,103,0,47,0,196,0,207,0,0,0,198,0,233,0,81,0,181,0,0,0,0,0,20,0,22,0,244,0,99,0,54,0,24,0,121,0,8,0,146,0,172,0,181,0,233,0,0,0,78,0,173,0,214,0,165,0,126,0,173,0,197,0,140,0,0,0,0,0,9,0,64,0,0,0,14,0,0,0,242,0,96,0,169,0,12,0,215,0,35,0,196,0,0,0,200,0,88,0,222,0,134,0,88,0,56,0,0,0,0,0,124,0,209,0,0,0,104,0,162,0,217,0,6,0,36,0,0,0,142,0,0,0,78,0,0,0,155,0,154,0,20,0,125,0,122,0,63,0,166,0,201,0,178,0,0,0,0,0,59,0,115,0,0,0,20,0,146,0,0,0,218,0,91,0,209,0,115,0,123,0,29,0,72,0,167,0,124,0,248,0,0,0,243,0,248,0,22,0,239,0,0,0,188,0,199,0,70,0,33,0,252,0,74,0,34,0,34,0,89,0,0,0,74,0,0,0,86,0,0,0,147,0,156,0,251,0,99,0,80,0,0,0,5,0,175,0,118,0,234,0,9,0,237,0,0,0,180,0,134,0,0,0,172,0,0,0,0,0,0,0,115,0,181,0,224,0,37,0,151,0,22,0,29,0,239,0,202,0,52,0,83,0,0,0,38,0,0,0,65,0,0,0,14,0,12,0,190,0,206,0,85,0,230,0,208,0,142,0,145,0,235,0,0,0,250,0,47,0,0,0,69,0,232,0,214,0,101,0,97,0,67,0,91,0,225,0,201,0,51,0,66,0,0,0,98,0,215,0,0,0,147,0,251,0,0,0,0,0,6,0,24,0,12,0,214,0,206,0,246,0,36,0,222,0,4,0,16,0,0,0,253,0,185,0,59,0,246,0,136,0,119,0,84,0,146,0,238,0,209,0,243,0,34,0,247,0,139,0,105,0,242,0,41,0,186,0,65,0,56,0,218,0,25,0,105,0,7,0,0,0,63,0,80,0,73,0,50,0,217,0,0,0,0,0,53,0,101,0,90,0,0,0,252,0,15,0,0,0,136,0,0,0,40,0,151,0,207,0,99,0,185,0,0,0,97,0,0,0,98,0,0,0,0,0,0,0,158,0,207,0,236,0,146,0,187,0,26,0,120,0,2,0,136,0,254,0,112,0,53,0,174,0,101,0,0,0,233,0,0,0,219,0,252,0,250,0,248,0,145,0,43,0,183,0,47,0,0,0,27,0,99,0,64,0,144,0,223,0,59,0,0,0,81,0,221,0,88,0,240,0,33,0,0,0,236,0,24,0,90,0,0,0,230,0,0,0,240,0,240,0,50,0,124,0,155,0,29,0,0,0,217,0,90,0,107,0,35,0,241,0,228,0,200,0,14,0,0,0,233,0,80,0,96,0,6,0,121,0,184,0,0,0,82,0,89,0,176,0,0,0,173,0,169,0,0,0,18,0,149,0,243,0,0,0,0,0,52,0,14,0,1,0,38,0,60,0,161,0,83,0,86,0,0,0,0,0,141,0,176,0,0,0,0,0,231,0,114,0,0,0,193,0,9,0,117,0,203,0,71,0,46,0,243,0,16,0,0,0,231,0,24,0,0,0,161,0,223,0,52,0,190,0,130,0,0,0,0,0,113,0,80,0,6,0,101,0,55,0,0,0,121,0,236,0,123,0,64,0,106,0,49,0,137,0,93,0,140,0,199,0,24,0,0,0,253,0,12,0,182,0,35,0,182,0,53,0,172,0,0,0,86,0,206,0,236,0,134,0,138,0,0,0,195,0,0,0,0,0,161,0,157,0,25,0,17,0,20,0,0,0,162,0,19,0,0,0,78,0,129,0,71,0,207,0,212,0,25,0,199,0,6,0,224,0,9,0,233,0,232,0,144,0,146,0,201,0,252,0,80,0,0,0,67,0,0,0,181,0,21,0,0,0,148,0,147,0,160,0,163,0,0,0,0,0,216,0,109,0,37,0,0,0,8,0,137,0,151,0,0,0,28,0,0,0,210,0,254,0,164,0,166,0,42,0,0,0,192,0,56,0,177,0,0,0,73,0,139,0,72,0,99,0,101,0,0,0,234,0,0,0,219,0,199,0,0,0,31,0,60,0,182,0,113,0,0,0,0,0,69,0,0,0,46,0,199,0,115,0,139,0,82,0,53,0,0,0,176,0,0,0,0,0,131,0,116,0,62,0,21,0,91,0,172,0,230,0,181,0,24,0,0,0,36,0,0,0,0,0,0,0,224,0,242,0,53,0,0,0,176,0,148,0,180,0,162,0,152,0,217,0,162,0,106,0,203,0,138,0,242,0,200,0,25,0,173,0,146,0,43,0,214,0,216,0,82,0,0,0,228,0,247,0,11,0,199,0,78,0,187,0,223,0,0,0,64,0,87,0,241,0,118,0,11,0,84,0);
signal scenario_full  : scenario_type := (116,31,221,31,34,31,34,30,34,29,48,31,200,31,202,31,121,31,248,31,55,31,244,31,77,31,138,31,188,31,18,31,18,30,139,31,17,31,29,31,5,31,5,30,216,31,151,31,151,30,84,31,237,31,23,31,23,30,23,29,44,31,44,30,165,31,104,31,162,31,103,31,174,31,174,30,81,31,131,31,138,31,152,31,200,31,166,31,39,31,88,31,88,30,137,31,137,30,190,31,39,31,46,31,42,31,123,31,43,31,100,31,37,31,37,30,109,31,114,31,159,31,78,31,163,31,220,31,129,31,230,31,124,31,124,30,19,31,122,31,200,31,85,31,84,31,25,31,167,31,247,31,42,31,148,31,246,31,246,30,44,31,44,30,3,31,41,31,68,31,45,31,105,31,105,30,32,31,221,31,117,31,191,31,220,31,144,31,97,31,217,31,90,31,107,31,202,31,202,30,202,29,108,31,6,31,22,31,107,31,145,31,180,31,197,31,189,31,54,31,216,31,176,31,100,31,89,31,136,31,158,31,239,31,253,31,195,31,202,31,15,31,15,30,15,29,53,31,145,31,219,31,219,30,172,31,153,31,90,31,90,30,67,31,203,31,19,31,19,30,113,31,101,31,59,31,32,31,32,30,102,31,188,31,188,30,90,31,201,31,176,31,214,31,220,31,221,31,96,31,159,31,103,31,79,31,153,31,153,30,153,29,147,31,16,31,133,31,29,31,156,31,103,31,211,31,211,30,243,31,243,30,56,31,93,31,61,31,34,31,182,31,182,30,151,31,117,31,55,31,55,30,74,31,23,31,23,30,170,31,170,30,129,31,80,31,64,31,99,31,115,31,119,31,83,31,230,31,231,31,186,31,224,31,108,31,130,31,231,31,142,31,189,31,235,31,187,31,220,31,251,31,160,31,160,30,160,29,19,31,209,31,254,31,173,31,173,30,187,31,187,30,251,31,228,31,223,31,196,31,181,31,74,31,74,30,108,31,24,31,145,31,145,30,180,31,212,31,22,31,22,30,45,31,5,31,200,31,103,31,47,31,196,31,207,31,207,30,198,31,233,31,81,31,181,31,181,30,181,29,20,31,22,31,244,31,99,31,54,31,24,31,121,31,8,31,146,31,172,31,181,31,233,31,233,30,78,31,173,31,214,31,165,31,126,31,173,31,197,31,140,31,140,30,140,29,9,31,64,31,64,30,14,31,14,30,242,31,96,31,169,31,12,31,215,31,35,31,196,31,196,30,200,31,88,31,222,31,134,31,88,31,56,31,56,30,56,29,124,31,209,31,209,30,104,31,162,31,217,31,6,31,36,31,36,30,142,31,142,30,78,31,78,30,155,31,154,31,20,31,125,31,122,31,63,31,166,31,201,31,178,31,178,30,178,29,59,31,115,31,115,30,20,31,146,31,146,30,218,31,91,31,209,31,115,31,123,31,29,31,72,31,167,31,124,31,248,31,248,30,243,31,248,31,22,31,239,31,239,30,188,31,199,31,70,31,33,31,252,31,74,31,34,31,34,31,89,31,89,30,74,31,74,30,86,31,86,30,147,31,156,31,251,31,99,31,80,31,80,30,5,31,175,31,118,31,234,31,9,31,237,31,237,30,180,31,134,31,134,30,172,31,172,30,172,29,172,28,115,31,181,31,224,31,37,31,151,31,22,31,29,31,239,31,202,31,52,31,83,31,83,30,38,31,38,30,65,31,65,30,14,31,12,31,190,31,206,31,85,31,230,31,208,31,142,31,145,31,235,31,235,30,250,31,47,31,47,30,69,31,232,31,214,31,101,31,97,31,67,31,91,31,225,31,201,31,51,31,66,31,66,30,98,31,215,31,215,30,147,31,251,31,251,30,251,29,6,31,24,31,12,31,214,31,206,31,246,31,36,31,222,31,4,31,16,31,16,30,253,31,185,31,59,31,246,31,136,31,119,31,84,31,146,31,238,31,209,31,243,31,34,31,247,31,139,31,105,31,242,31,41,31,186,31,65,31,56,31,218,31,25,31,105,31,7,31,7,30,63,31,80,31,73,31,50,31,217,31,217,30,217,29,53,31,101,31,90,31,90,30,252,31,15,31,15,30,136,31,136,30,40,31,151,31,207,31,99,31,185,31,185,30,97,31,97,30,98,31,98,30,98,29,98,28,158,31,207,31,236,31,146,31,187,31,26,31,120,31,2,31,136,31,254,31,112,31,53,31,174,31,101,31,101,30,233,31,233,30,219,31,252,31,250,31,248,31,145,31,43,31,183,31,47,31,47,30,27,31,99,31,64,31,144,31,223,31,59,31,59,30,81,31,221,31,88,31,240,31,33,31,33,30,236,31,24,31,90,31,90,30,230,31,230,30,240,31,240,31,50,31,124,31,155,31,29,31,29,30,217,31,90,31,107,31,35,31,241,31,228,31,200,31,14,31,14,30,233,31,80,31,96,31,6,31,121,31,184,31,184,30,82,31,89,31,176,31,176,30,173,31,169,31,169,30,18,31,149,31,243,31,243,30,243,29,52,31,14,31,1,31,38,31,60,31,161,31,83,31,86,31,86,30,86,29,141,31,176,31,176,30,176,29,231,31,114,31,114,30,193,31,9,31,117,31,203,31,71,31,46,31,243,31,16,31,16,30,231,31,24,31,24,30,161,31,223,31,52,31,190,31,130,31,130,30,130,29,113,31,80,31,6,31,101,31,55,31,55,30,121,31,236,31,123,31,64,31,106,31,49,31,137,31,93,31,140,31,199,31,24,31,24,30,253,31,12,31,182,31,35,31,182,31,53,31,172,31,172,30,86,31,206,31,236,31,134,31,138,31,138,30,195,31,195,30,195,29,161,31,157,31,25,31,17,31,20,31,20,30,162,31,19,31,19,30,78,31,129,31,71,31,207,31,212,31,25,31,199,31,6,31,224,31,9,31,233,31,232,31,144,31,146,31,201,31,252,31,80,31,80,30,67,31,67,30,181,31,21,31,21,30,148,31,147,31,160,31,163,31,163,30,163,29,216,31,109,31,37,31,37,30,8,31,137,31,151,31,151,30,28,31,28,30,210,31,254,31,164,31,166,31,42,31,42,30,192,31,56,31,177,31,177,30,73,31,139,31,72,31,99,31,101,31,101,30,234,31,234,30,219,31,199,31,199,30,31,31,60,31,182,31,113,31,113,30,113,29,69,31,69,30,46,31,199,31,115,31,139,31,82,31,53,31,53,30,176,31,176,30,176,29,131,31,116,31,62,31,21,31,91,31,172,31,230,31,181,31,24,31,24,30,36,31,36,30,36,29,36,28,224,31,242,31,53,31,53,30,176,31,148,31,180,31,162,31,152,31,217,31,162,31,106,31,203,31,138,31,242,31,200,31,25,31,173,31,146,31,43,31,214,31,216,31,82,31,82,30,228,31,247,31,11,31,199,31,78,31,187,31,223,31,223,30,64,31,87,31,241,31,118,31,11,31,84,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
