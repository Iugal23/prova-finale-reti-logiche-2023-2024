-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 333;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (224,0,0,0,176,0,0,0,127,0,183,0,85,0,3,0,47,0,209,0,195,0,247,0,0,0,199,0,12,0,25,0,133,0,146,0,24,0,173,0,66,0,198,0,108,0,128,0,0,0,114,0,38,0,0,0,223,0,131,0,7,0,254,0,210,0,0,0,77,0,243,0,9,0,98,0,40,0,101,0,143,0,108,0,210,0,217,0,0,0,220,0,12,0,29,0,142,0,176,0,180,0,0,0,117,0,87,0,141,0,177,0,0,0,0,0,3,0,0,0,203,0,0,0,183,0,187,0,228,0,19,0,97,0,23,0,0,0,147,0,178,0,173,0,228,0,115,0,21,0,90,0,57,0,132,0,180,0,163,0,165,0,141,0,112,0,140,0,236,0,118,0,79,0,24,0,93,0,251,0,158,0,200,0,85,0,0,0,0,0,243,0,141,0,175,0,207,0,0,0,202,0,119,0,103,0,15,0,64,0,19,0,160,0,174,0,3,0,154,0,0,0,0,0,0,0,0,0,47,0,173,0,24,0,68,0,0,0,137,0,155,0,84,0,138,0,222,0,195,0,136,0,169,0,30,0,223,0,110,0,126,0,97,0,0,0,192,0,162,0,226,0,181,0,0,0,0,0,165,0,243,0,132,0,0,0,155,0,4,0,89,0,193,0,226,0,172,0,146,0,121,0,132,0,61,0,77,0,88,0,114,0,0,0,116,0,96,0,225,0,0,0,217,0,70,0,111,0,0,0,103,0,255,0,123,0,217,0,106,0,94,0,0,0,204,0,0,0,100,0,57,0,202,0,61,0,70,0,149,0,107,0,0,0,0,0,176,0,0,0,0,0,168,0,242,0,33,0,253,0,0,0,1,0,0,0,0,0,174,0,85,0,119,0,160,0,0,0,51,0,0,0,106,0,0,0,25,0,98,0,247,0,8,0,0,0,73,0,174,0,0,0,113,0,57,0,155,0,116,0,0,0,10,0,181,0,179,0,218,0,122,0,191,0,40,0,0,0,216,0,121,0,100,0,0,0,242,0,0,0,0,0,88,0,163,0,151,0,248,0,130,0,62,0,239,0,70,0,63,0,156,0,189,0,60,0,0,0,204,0,183,0,196,0,0,0,249,0,168,0,0,0,213,0,0,0,139,0,192,0,74,0,154,0,0,0,199,0,65,0,250,0,234,0,146,0,97,0,84,0,74,0,114,0,188,0,81,0,183,0,133,0,96,0,210,0,100,0,1,0,51,0,136,0,103,0,123,0,105,0,78,0,134,0,207,0,53,0,98,0,0,0,45,0,52,0,52,0,36,0,21,0,136,0,169,0,87,0,91,0,172,0,0,0,156,0,76,0,106,0,251,0,40,0,88,0,211,0,206,0,73,0,78,0,156,0,0,0,87,0,0,0,0,0,43,0,35,0,0,0,180,0,117,0,115,0,49,0,110,0,200,0,88,0,0,0,221,0,0,0,0,0,248,0,0,0,66,0,105,0,145,0,0,0,202,0);
signal scenario_full  : scenario_type := (224,31,224,30,176,31,176,30,127,31,183,31,85,31,3,31,47,31,209,31,195,31,247,31,247,30,199,31,12,31,25,31,133,31,146,31,24,31,173,31,66,31,198,31,108,31,128,31,128,30,114,31,38,31,38,30,223,31,131,31,7,31,254,31,210,31,210,30,77,31,243,31,9,31,98,31,40,31,101,31,143,31,108,31,210,31,217,31,217,30,220,31,12,31,29,31,142,31,176,31,180,31,180,30,117,31,87,31,141,31,177,31,177,30,177,29,3,31,3,30,203,31,203,30,183,31,187,31,228,31,19,31,97,31,23,31,23,30,147,31,178,31,173,31,228,31,115,31,21,31,90,31,57,31,132,31,180,31,163,31,165,31,141,31,112,31,140,31,236,31,118,31,79,31,24,31,93,31,251,31,158,31,200,31,85,31,85,30,85,29,243,31,141,31,175,31,207,31,207,30,202,31,119,31,103,31,15,31,64,31,19,31,160,31,174,31,3,31,154,31,154,30,154,29,154,28,154,27,47,31,173,31,24,31,68,31,68,30,137,31,155,31,84,31,138,31,222,31,195,31,136,31,169,31,30,31,223,31,110,31,126,31,97,31,97,30,192,31,162,31,226,31,181,31,181,30,181,29,165,31,243,31,132,31,132,30,155,31,4,31,89,31,193,31,226,31,172,31,146,31,121,31,132,31,61,31,77,31,88,31,114,31,114,30,116,31,96,31,225,31,225,30,217,31,70,31,111,31,111,30,103,31,255,31,123,31,217,31,106,31,94,31,94,30,204,31,204,30,100,31,57,31,202,31,61,31,70,31,149,31,107,31,107,30,107,29,176,31,176,30,176,29,168,31,242,31,33,31,253,31,253,30,1,31,1,30,1,29,174,31,85,31,119,31,160,31,160,30,51,31,51,30,106,31,106,30,25,31,98,31,247,31,8,31,8,30,73,31,174,31,174,30,113,31,57,31,155,31,116,31,116,30,10,31,181,31,179,31,218,31,122,31,191,31,40,31,40,30,216,31,121,31,100,31,100,30,242,31,242,30,242,29,88,31,163,31,151,31,248,31,130,31,62,31,239,31,70,31,63,31,156,31,189,31,60,31,60,30,204,31,183,31,196,31,196,30,249,31,168,31,168,30,213,31,213,30,139,31,192,31,74,31,154,31,154,30,199,31,65,31,250,31,234,31,146,31,97,31,84,31,74,31,114,31,188,31,81,31,183,31,133,31,96,31,210,31,100,31,1,31,51,31,136,31,103,31,123,31,105,31,78,31,134,31,207,31,53,31,98,31,98,30,45,31,52,31,52,31,36,31,21,31,136,31,169,31,87,31,91,31,172,31,172,30,156,31,76,31,106,31,251,31,40,31,88,31,211,31,206,31,73,31,78,31,156,31,156,30,87,31,87,30,87,29,43,31,35,31,35,30,180,31,117,31,115,31,49,31,110,31,200,31,88,31,88,30,221,31,221,30,221,29,248,31,248,30,66,31,105,31,145,31,145,30,202,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
