-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_554 is
end project_tb_554;

architecture project_tb_arch_554 of project_tb_554 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 896;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (182,0,0,0,78,0,36,0,60,0,32,0,51,0,27,0,63,0,0,0,0,0,166,0,246,0,38,0,0,0,91,0,54,0,0,0,16,0,244,0,101,0,21,0,250,0,0,0,11,0,153,0,218,0,232,0,154,0,198,0,194,0,39,0,194,0,93,0,130,0,0,0,0,0,81,0,170,0,39,0,0,0,214,0,217,0,52,0,59,0,0,0,146,0,206,0,23,0,0,0,93,0,58,0,0,0,113,0,253,0,105,0,190,0,0,0,194,0,135,0,152,0,169,0,210,0,0,0,0,0,239,0,246,0,84,0,52,0,68,0,50,0,72,0,223,0,152,0,169,0,72,0,185,0,0,0,122,0,211,0,230,0,3,0,22,0,159,0,177,0,34,0,91,0,107,0,40,0,138,0,0,0,79,0,237,0,51,0,186,0,64,0,90,0,0,0,11,0,232,0,0,0,58,0,42,0,232,0,0,0,255,0,156,0,170,0,175,0,145,0,0,0,0,0,127,0,200,0,0,0,248,0,166,0,0,0,0,0,246,0,118,0,0,0,230,0,25,0,0,0,42,0,217,0,0,0,15,0,0,0,47,0,205,0,0,0,2,0,98,0,117,0,4,0,234,0,0,0,194,0,140,0,0,0,192,0,18,0,0,0,158,0,0,0,0,0,46,0,144,0,123,0,180,0,0,0,131,0,61,0,138,0,190,0,21,0,59,0,0,0,0,0,69,0,20,0,182,0,53,0,0,0,160,0,149,0,201,0,0,0,196,0,181,0,229,0,0,0,95,0,12,0,81,0,237,0,154,0,9,0,0,0,0,0,62,0,155,0,0,0,191,0,164,0,47,0,0,0,174,0,0,0,139,0,0,0,116,0,196,0,239,0,0,0,150,0,188,0,0,0,0,0,205,0,173,0,140,0,0,0,151,0,200,0,0,0,199,0,87,0,75,0,164,0,3,0,0,0,38,0,0,0,0,0,0,0,188,0,0,0,23,0,75,0,0,0,101,0,171,0,156,0,22,0,224,0,3,0,198,0,201,0,59,0,168,0,0,0,26,0,152,0,32,0,134,0,52,0,119,0,92,0,124,0,71,0,3,0,125,0,140,0,121,0,81,0,51,0,0,0,238,0,0,0,0,0,157,0,51,0,30,0,161,0,95,0,230,0,189,0,119,0,242,0,179,0,23,0,3,0,98,0,184,0,102,0,143,0,0,0,107,0,219,0,0,0,67,0,176,0,252,0,49,0,159,0,198,0,6,0,168,0,171,0,168,0,104,0,100,0,170,0,221,0,95,0,231,0,152,0,187,0,106,0,155,0,56,0,248,0,130,0,63,0,0,0,150,0,0,0,0,0,139,0,193,0,230,0,170,0,172,0,203,0,153,0,29,0,107,0,153,0,86,0,238,0,141,0,63,0,70,0,61,0,27,0,249,0,124,0,20,0,45,0,237,0,9,0,46,0,29,0,6,0,198,0,76,0,215,0,100,0,88,0,7,0,90,0,0,0,0,0,8,0,128,0,140,0,116,0,187,0,133,0,147,0,3,0,86,0,155,0,134,0,156,0,63,0,0,0,146,0,229,0,0,0,0,0,184,0,194,0,101,0,144,0,30,0,159,0,106,0,31,0,215,0,133,0,0,0,249,0,191,0,211,0,0,0,0,0,223,0,82,0,0,0,0,0,178,0,0,0,33,0,121,0,121,0,43,0,152,0,0,0,0,0,90,0,0,0,23,0,204,0,23,0,0,0,21,0,63,0,59,0,219,0,0,0,0,0,243,0,0,0,160,0,0,0,48,0,27,0,0,0,223,0,91,0,220,0,124,0,230,0,0,0,13,0,131,0,0,0,34,0,171,0,27,0,151,0,58,0,12,0,30,0,17,0,174,0,0,0,34,0,0,0,0,0,50,0,0,0,100,0,89,0,0,0,218,0,30,0,137,0,35,0,0,0,115,0,227,0,24,0,211,0,0,0,84,0,72,0,193,0,0,0,176,0,0,0,202,0,0,0,238,0,186,0,155,0,12,0,209,0,85,0,0,0,0,0,206,0,88,0,20,0,0,0,0,0,75,0,0,0,46,0,0,0,9,0,18,0,68,0,0,0,243,0,218,0,190,0,29,0,244,0,126,0,60,0,0,0,142,0,57,0,220,0,131,0,235,0,0,0,81,0,159,0,195,0,152,0,0,0,218,0,155,0,183,0,0,0,25,0,225,0,17,0,200,0,0,0,94,0,254,0,224,0,76,0,79,0,233,0,164,0,109,0,230,0,0,0,130,0,10,0,0,0,0,0,0,0,186,0,154,0,166,0,103,0,0,0,191,0,143,0,51,0,0,0,0,0,39,0,53,0,95,0,163,0,0,0,236,0,47,0,22,0,40,0,40,0,220,0,20,0,8,0,116,0,220,0,108,0,0,0,0,0,138,0,0,0,69,0,0,0,204,0,112,0,41,0,44,0,0,0,223,0,164,0,14,0,0,0,145,0,0,0,36,0,0,0,82,0,134,0,166,0,135,0,79,0,0,0,129,0,104,0,214,0,134,0,125,0,209,0,182,0,37,0,16,0,161,0,109,0,0,0,0,0,88,0,1,0,93,0,135,0,4,0,152,0,150,0,161,0,239,0,41,0,122,0,226,0,229,0,0,0,81,0,61,0,131,0,190,0,0,0,84,0,0,0,191,0,125,0,220,0,87,0,128,0,151,0,192,0,210,0,199,0,53,0,232,0,96,0,112,0,229,0,0,0,105,0,75,0,194,0,0,0,0,0,82,0,218,0,129,0,0,0,65,0,245,0,102,0,220,0,208,0,255,0,186,0,119,0,86,0,0,0,185,0,111,0,0,0,250,0,181,0,45,0,0,0,95,0,37,0,124,0,122,0,13,0,0,0,149,0,14,0,184,0,222,0,35,0,35,0,14,0,158,0,173,0,43,0,212,0,79,0,96,0,18,0,0,0,201,0,56,0,213,0,226,0,167,0,220,0,255,0,30,0,17,0,114,0,147,0,214,0,213,0,12,0,55,0,85,0,116,0,0,0,101,0,0,0,0,0,93,0,243,0,141,0,179,0,199,0,109,0,45,0,211,0,135,0,178,0,164,0,212,0,34,0,0,0,0,0,77,0,124,0,0,0,66,0,77,0,60,0,4,0,0,0,157,0,201,0,71,0,22,0,187,0,4,0,182,0,113,0,0,0,235,0,251,0,0,0,0,0,0,0,0,0,23,0,154,0,215,0,0,0,28,0,0,0,62,0,57,0,0,0,0,0,245,0,69,0,116,0,223,0,59,0,0,0,60,0,0,0,221,0,23,0,55,0,192,0,156,0,181,0,180,0,167,0,51,0,60,0,22,0,79,0,0,0,219,0,113,0,0,0,94,0,255,0,180,0,208,0,159,0,251,0,0,0,170,0,170,0,131,0,37,0,217,0,223,0,43,0,0,0,24,0,42,0,207,0,53,0,165,0,104,0,247,0,0,0,72,0,134,0,204,0,235,0,212,0,125,0,0,0,123,0,136,0,120,0,8,0,0,0,99,0,70,0,133,0,182,0,141,0,206,0,10,0,4,0,0,0,9,0,129,0,0,0,0,0,228,0,86,0,139,0,172,0,196,0,229,0,77,0,233,0,139,0,20,0,151,0,17,0,235,0,4,0,83,0,202,0,27,0,77,0,185,0,232,0,158,0,162,0,143,0,216,0,116,0,117,0,253,0,225,0,24,0,175,0,177,0,0,0,131,0,148,0,96,0,106,0,0,0,220,0,18,0,152,0,0,0,73,0,45,0,97,0,189,0,75,0,17,0,189,0,217,0,0,0,58,0,80,0,191,0,249,0,156,0,31,0,107,0,0,0,110,0,250,0,0,0,255,0,214,0,181,0,65,0,75,0,69,0,210,0,0,0,127,0,191,0,19,0,10,0,216,0,243,0,123,0,180,0,45,0,41,0,137,0,247,0,254,0,0,0,2,0,189,0,3,0,86,0,0,0,0,0,194,0,13,0,123,0,115,0,98,0,51,0,25,0,110,0);
signal scenario_full  : scenario_type := (182,31,182,30,78,31,36,31,60,31,32,31,51,31,27,31,63,31,63,30,63,29,166,31,246,31,38,31,38,30,91,31,54,31,54,30,16,31,244,31,101,31,21,31,250,31,250,30,11,31,153,31,218,31,232,31,154,31,198,31,194,31,39,31,194,31,93,31,130,31,130,30,130,29,81,31,170,31,39,31,39,30,214,31,217,31,52,31,59,31,59,30,146,31,206,31,23,31,23,30,93,31,58,31,58,30,113,31,253,31,105,31,190,31,190,30,194,31,135,31,152,31,169,31,210,31,210,30,210,29,239,31,246,31,84,31,52,31,68,31,50,31,72,31,223,31,152,31,169,31,72,31,185,31,185,30,122,31,211,31,230,31,3,31,22,31,159,31,177,31,34,31,91,31,107,31,40,31,138,31,138,30,79,31,237,31,51,31,186,31,64,31,90,31,90,30,11,31,232,31,232,30,58,31,42,31,232,31,232,30,255,31,156,31,170,31,175,31,145,31,145,30,145,29,127,31,200,31,200,30,248,31,166,31,166,30,166,29,246,31,118,31,118,30,230,31,25,31,25,30,42,31,217,31,217,30,15,31,15,30,47,31,205,31,205,30,2,31,98,31,117,31,4,31,234,31,234,30,194,31,140,31,140,30,192,31,18,31,18,30,158,31,158,30,158,29,46,31,144,31,123,31,180,31,180,30,131,31,61,31,138,31,190,31,21,31,59,31,59,30,59,29,69,31,20,31,182,31,53,31,53,30,160,31,149,31,201,31,201,30,196,31,181,31,229,31,229,30,95,31,12,31,81,31,237,31,154,31,9,31,9,30,9,29,62,31,155,31,155,30,191,31,164,31,47,31,47,30,174,31,174,30,139,31,139,30,116,31,196,31,239,31,239,30,150,31,188,31,188,30,188,29,205,31,173,31,140,31,140,30,151,31,200,31,200,30,199,31,87,31,75,31,164,31,3,31,3,30,38,31,38,30,38,29,38,28,188,31,188,30,23,31,75,31,75,30,101,31,171,31,156,31,22,31,224,31,3,31,198,31,201,31,59,31,168,31,168,30,26,31,152,31,32,31,134,31,52,31,119,31,92,31,124,31,71,31,3,31,125,31,140,31,121,31,81,31,51,31,51,30,238,31,238,30,238,29,157,31,51,31,30,31,161,31,95,31,230,31,189,31,119,31,242,31,179,31,23,31,3,31,98,31,184,31,102,31,143,31,143,30,107,31,219,31,219,30,67,31,176,31,252,31,49,31,159,31,198,31,6,31,168,31,171,31,168,31,104,31,100,31,170,31,221,31,95,31,231,31,152,31,187,31,106,31,155,31,56,31,248,31,130,31,63,31,63,30,150,31,150,30,150,29,139,31,193,31,230,31,170,31,172,31,203,31,153,31,29,31,107,31,153,31,86,31,238,31,141,31,63,31,70,31,61,31,27,31,249,31,124,31,20,31,45,31,237,31,9,31,46,31,29,31,6,31,198,31,76,31,215,31,100,31,88,31,7,31,90,31,90,30,90,29,8,31,128,31,140,31,116,31,187,31,133,31,147,31,3,31,86,31,155,31,134,31,156,31,63,31,63,30,146,31,229,31,229,30,229,29,184,31,194,31,101,31,144,31,30,31,159,31,106,31,31,31,215,31,133,31,133,30,249,31,191,31,211,31,211,30,211,29,223,31,82,31,82,30,82,29,178,31,178,30,33,31,121,31,121,31,43,31,152,31,152,30,152,29,90,31,90,30,23,31,204,31,23,31,23,30,21,31,63,31,59,31,219,31,219,30,219,29,243,31,243,30,160,31,160,30,48,31,27,31,27,30,223,31,91,31,220,31,124,31,230,31,230,30,13,31,131,31,131,30,34,31,171,31,27,31,151,31,58,31,12,31,30,31,17,31,174,31,174,30,34,31,34,30,34,29,50,31,50,30,100,31,89,31,89,30,218,31,30,31,137,31,35,31,35,30,115,31,227,31,24,31,211,31,211,30,84,31,72,31,193,31,193,30,176,31,176,30,202,31,202,30,238,31,186,31,155,31,12,31,209,31,85,31,85,30,85,29,206,31,88,31,20,31,20,30,20,29,75,31,75,30,46,31,46,30,9,31,18,31,68,31,68,30,243,31,218,31,190,31,29,31,244,31,126,31,60,31,60,30,142,31,57,31,220,31,131,31,235,31,235,30,81,31,159,31,195,31,152,31,152,30,218,31,155,31,183,31,183,30,25,31,225,31,17,31,200,31,200,30,94,31,254,31,224,31,76,31,79,31,233,31,164,31,109,31,230,31,230,30,130,31,10,31,10,30,10,29,10,28,186,31,154,31,166,31,103,31,103,30,191,31,143,31,51,31,51,30,51,29,39,31,53,31,95,31,163,31,163,30,236,31,47,31,22,31,40,31,40,31,220,31,20,31,8,31,116,31,220,31,108,31,108,30,108,29,138,31,138,30,69,31,69,30,204,31,112,31,41,31,44,31,44,30,223,31,164,31,14,31,14,30,145,31,145,30,36,31,36,30,82,31,134,31,166,31,135,31,79,31,79,30,129,31,104,31,214,31,134,31,125,31,209,31,182,31,37,31,16,31,161,31,109,31,109,30,109,29,88,31,1,31,93,31,135,31,4,31,152,31,150,31,161,31,239,31,41,31,122,31,226,31,229,31,229,30,81,31,61,31,131,31,190,31,190,30,84,31,84,30,191,31,125,31,220,31,87,31,128,31,151,31,192,31,210,31,199,31,53,31,232,31,96,31,112,31,229,31,229,30,105,31,75,31,194,31,194,30,194,29,82,31,218,31,129,31,129,30,65,31,245,31,102,31,220,31,208,31,255,31,186,31,119,31,86,31,86,30,185,31,111,31,111,30,250,31,181,31,45,31,45,30,95,31,37,31,124,31,122,31,13,31,13,30,149,31,14,31,184,31,222,31,35,31,35,31,14,31,158,31,173,31,43,31,212,31,79,31,96,31,18,31,18,30,201,31,56,31,213,31,226,31,167,31,220,31,255,31,30,31,17,31,114,31,147,31,214,31,213,31,12,31,55,31,85,31,116,31,116,30,101,31,101,30,101,29,93,31,243,31,141,31,179,31,199,31,109,31,45,31,211,31,135,31,178,31,164,31,212,31,34,31,34,30,34,29,77,31,124,31,124,30,66,31,77,31,60,31,4,31,4,30,157,31,201,31,71,31,22,31,187,31,4,31,182,31,113,31,113,30,235,31,251,31,251,30,251,29,251,28,251,27,23,31,154,31,215,31,215,30,28,31,28,30,62,31,57,31,57,30,57,29,245,31,69,31,116,31,223,31,59,31,59,30,60,31,60,30,221,31,23,31,55,31,192,31,156,31,181,31,180,31,167,31,51,31,60,31,22,31,79,31,79,30,219,31,113,31,113,30,94,31,255,31,180,31,208,31,159,31,251,31,251,30,170,31,170,31,131,31,37,31,217,31,223,31,43,31,43,30,24,31,42,31,207,31,53,31,165,31,104,31,247,31,247,30,72,31,134,31,204,31,235,31,212,31,125,31,125,30,123,31,136,31,120,31,8,31,8,30,99,31,70,31,133,31,182,31,141,31,206,31,10,31,4,31,4,30,9,31,129,31,129,30,129,29,228,31,86,31,139,31,172,31,196,31,229,31,77,31,233,31,139,31,20,31,151,31,17,31,235,31,4,31,83,31,202,31,27,31,77,31,185,31,232,31,158,31,162,31,143,31,216,31,116,31,117,31,253,31,225,31,24,31,175,31,177,31,177,30,131,31,148,31,96,31,106,31,106,30,220,31,18,31,152,31,152,30,73,31,45,31,97,31,189,31,75,31,17,31,189,31,217,31,217,30,58,31,80,31,191,31,249,31,156,31,31,31,107,31,107,30,110,31,250,31,250,30,255,31,214,31,181,31,65,31,75,31,69,31,210,31,210,30,127,31,191,31,19,31,10,31,216,31,243,31,123,31,180,31,45,31,41,31,137,31,247,31,254,31,254,30,2,31,189,31,3,31,86,31,86,30,86,29,194,31,13,31,123,31,115,31,98,31,51,31,25,31,110,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
