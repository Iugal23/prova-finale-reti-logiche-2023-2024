-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 859;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,117,0,175,0,110,0,241,0,111,0,0,0,226,0,49,0,110,0,80,0,182,0,0,0,149,0,0,0,65,0,143,0,48,0,0,0,0,0,14,0,137,0,199,0,140,0,0,0,102,0,228,0,16,0,158,0,111,0,105,0,194,0,127,0,142,0,0,0,48,0,0,0,177,0,0,0,225,0,0,0,120,0,32,0,160,0,216,0,0,0,102,0,165,0,184,0,222,0,50,0,114,0,88,0,0,0,95,0,118,0,24,0,168,0,208,0,224,0,213,0,108,0,161,0,115,0,184,0,135,0,0,0,95,0,246,0,88,0,91,0,131,0,231,0,41,0,34,0,56,0,194,0,141,0,11,0,177,0,0,0,202,0,93,0,89,0,159,0,189,0,0,0,98,0,71,0,222,0,91,0,56,0,39,0,127,0,86,0,0,0,152,0,50,0,57,0,194,0,0,0,0,0,90,0,59,0,233,0,179,0,115,0,104,0,0,0,173,0,202,0,3,0,199,0,46,0,0,0,79,0,107,0,32,0,0,0,5,0,0,0,239,0,93,0,62,0,251,0,83,0,129,0,15,0,85,0,197,0,156,0,215,0,121,0,75,0,137,0,199,0,215,0,62,0,0,0,0,0,65,0,0,0,0,0,77,0,14,0,39,0,154,0,131,0,48,0,0,0,119,0,36,0,0,0,0,0,42,0,0,0,0,0,0,0,51,0,0,0,0,0,67,0,42,0,63,0,0,0,120,0,0,0,172,0,158,0,72,0,210,0,170,0,251,0,45,0,35,0,0,0,163,0,194,0,0,0,63,0,215,0,24,0,0,0,137,0,140,0,64,0,115,0,0,0,226,0,161,0,61,0,210,0,152,0,191,0,136,0,52,0,199,0,91,0,0,0,0,0,0,0,216,0,19,0,0,0,89,0,36,0,144,0,249,0,0,0,62,0,28,0,88,0,244,0,225,0,131,0,65,0,213,0,252,0,0,0,53,0,176,0,0,0,45,0,189,0,36,0,0,0,137,0,84,0,254,0,43,0,238,0,0,0,205,0,47,0,100,0,145,0,0,0,7,0,17,0,0,0,67,0,119,0,0,0,115,0,0,0,102,0,171,0,10,0,234,0,168,0,123,0,18,0,117,0,27,0,0,0,0,0,0,0,0,0,0,0,0,0,194,0,149,0,0,0,90,0,108,0,240,0,0,0,0,0,114,0,33,0,146,0,73,0,0,0,58,0,171,0,218,0,0,0,160,0,0,0,27,0,12,0,200,0,208,0,0,0,9,0,61,0,23,0,21,0,78,0,0,0,0,0,136,0,10,0,95,0,0,0,18,0,216,0,152,0,127,0,234,0,219,0,148,0,172,0,150,0,84,0,71,0,0,0,148,0,144,0,0,0,58,0,165,0,114,0,0,0,246,0,145,0,130,0,0,0,64,0,101,0,65,0,50,0,228,0,215,0,238,0,146,0,0,0,0,0,83,0,246,0,0,0,0,0,240,0,232,0,55,0,131,0,221,0,159,0,39,0,20,0,186,0,53,0,220,0,243,0,226,0,0,0,22,0,178,0,0,0,104,0,154,0,11,0,244,0,0,0,187,0,126,0,0,0,186,0,57,0,139,0,0,0,0,0,0,0,32,0,0,0,163,0,152,0,86,0,124,0,51,0,128,0,54,0,150,0,177,0,187,0,253,0,154,0,38,0,167,0,183,0,185,0,124,0,87,0,124,0,165,0,100,0,0,0,199,0,240,0,59,0,92,0,191,0,140,0,138,0,68,0,129,0,0,0,250,0,0,0,226,0,12,0,119,0,4,0,0,0,173,0,163,0,16,0,66,0,121,0,0,0,97,0,211,0,57,0,207,0,248,0,120,0,111,0,0,0,96,0,171,0,141,0,103,0,148,0,0,0,0,0,175,0,83,0,60,0,136,0,34,0,0,0,119,0,97,0,0,0,31,0,0,0,0,0,58,0,226,0,121,0,111,0,223,0,104,0,218,0,117,0,249,0,243,0,0,0,78,0,125,0,16,0,0,0,198,0,0,0,134,0,249,0,233,0,0,0,0,0,39,0,202,0,81,0,175,0,0,0,54,0,41,0,0,0,157,0,43,0,249,0,47,0,0,0,44,0,245,0,157,0,91,0,0,0,14,0,74,0,58,0,93,0,0,0,5,0,222,0,121,0,0,0,0,0,94,0,0,0,48,0,248,0,113,0,113,0,100,0,0,0,255,0,57,0,191,0,92,0,0,0,157,0,217,0,0,0,138,0,0,0,238,0,57,0,133,0,0,0,244,0,197,0,145,0,6,0,141,0,186,0,235,0,113,0,42,0,0,0,217,0,7,0,210,0,133,0,200,0,29,0,202,0,0,0,241,0,253,0,0,0,107,0,16,0,138,0,0,0,10,0,237,0,208,0,64,0,213,0,103,0,199,0,89,0,70,0,214,0,223,0,133,0,33,0,0,0,210,0,0,0,63,0,201,0,132,0,237,0,0,0,0,0,31,0,58,0,0,0,119,0,69,0,207,0,0,0,0,0,0,0,0,0,64,0,206,0,14,0,32,0,109,0,88,0,215,0,20,0,63,0,96,0,0,0,80,0,222,0,67,0,108,0,120,0,0,0,32,0,175,0,249,0,0,0,119,0,25,0,0,0,100,0,243,0,157,0,107,0,0,0,49,0,10,0,0,0,80,0,0,0,128,0,10,0,167,0,52,0,78,0,188,0,81,0,89,0,51,0,153,0,240,0,0,0,139,0,58,0,51,0,170,0,104,0,91,0,164,0,0,0,106,0,49,0,198,0,136,0,252,0,161,0,70,0,188,0,194,0,0,0,138,0,200,0,68,0,64,0,0,0,187,0,211,0,132,0,0,0,0,0,195,0,43,0,0,0,58,0,35,0,0,0,235,0,0,0,67,0,82,0,22,0,81,0,0,0,47,0,180,0,7,0,50,0,102,0,205,0,0,0,22,0,244,0,0,0,164,0,222,0,0,0,74,0,0,0,152,0,0,0,231,0,118,0,62,0,157,0,0,0,193,0,168,0,97,0,234,0,109,0,104,0,147,0,82,0,240,0,145,0,204,0,231,0,83,0,0,0,0,0,0,0,149,0,140,0,237,0,168,0,229,0,127,0,213,0,0,0,0,0,38,0,102,0,112,0,81,0,157,0,0,0,77,0,165,0,149,0,18,0,207,0,5,0,248,0,240,0,54,0,61,0,17,0,203,0,0,0,0,0,0,0,220,0,64,0,0,0,175,0,0,0,251,0,169,0,19,0,0,0,213,0,159,0,6,0,7,0,0,0,117,0,130,0,156,0,30,0,62,0,194,0,156,0,0,0,135,0,143,0,12,0,234,0,195,0,208,0,71,0,88,0,212,0,185,0,42,0,122,0,198,0,7,0,0,0,115,0,90,0,177,0,25,0,25,0,29,0,198,0,0,0,0,0,70,0,242,0,48,0,0,0,48,0,250,0,118,0,57,0,111,0,149,0,109,0,141,0,0,0,41,0,180,0,0,0,122,0,90,0,87,0,153,0,208,0,9,0,0,0,172,0,103,0,128,0,107,0,246,0,9,0,191,0,12,0,0,0,179,0,147,0,207,0,20,0,138,0,0,0,217,0,0,0,247,0,0,0,0,0,160,0,0,0,230,0,38,0,133,0,222,0,201,0,242,0,0,0,13,0,208,0,200,0,74,0,85,0,235,0,92,0,232,0,159,0,0,0,0,0,0,0,170,0,175,0,0,0,126,0,128,0,175,0,248,0,0,0,191,0,0,0,252,0,178,0,0,0,232,0,143,0,109,0,38,0,189,0,170,0,142,0,82,0,0,0,70,0,77,0,0,0,28,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,117,31,175,31,110,31,241,31,111,31,111,30,226,31,49,31,110,31,80,31,182,31,182,30,149,31,149,30,65,31,143,31,48,31,48,30,48,29,14,31,137,31,199,31,140,31,140,30,102,31,228,31,16,31,158,31,111,31,105,31,194,31,127,31,142,31,142,30,48,31,48,30,177,31,177,30,225,31,225,30,120,31,32,31,160,31,216,31,216,30,102,31,165,31,184,31,222,31,50,31,114,31,88,31,88,30,95,31,118,31,24,31,168,31,208,31,224,31,213,31,108,31,161,31,115,31,184,31,135,31,135,30,95,31,246,31,88,31,91,31,131,31,231,31,41,31,34,31,56,31,194,31,141,31,11,31,177,31,177,30,202,31,93,31,89,31,159,31,189,31,189,30,98,31,71,31,222,31,91,31,56,31,39,31,127,31,86,31,86,30,152,31,50,31,57,31,194,31,194,30,194,29,90,31,59,31,233,31,179,31,115,31,104,31,104,30,173,31,202,31,3,31,199,31,46,31,46,30,79,31,107,31,32,31,32,30,5,31,5,30,239,31,93,31,62,31,251,31,83,31,129,31,15,31,85,31,197,31,156,31,215,31,121,31,75,31,137,31,199,31,215,31,62,31,62,30,62,29,65,31,65,30,65,29,77,31,14,31,39,31,154,31,131,31,48,31,48,30,119,31,36,31,36,30,36,29,42,31,42,30,42,29,42,28,51,31,51,30,51,29,67,31,42,31,63,31,63,30,120,31,120,30,172,31,158,31,72,31,210,31,170,31,251,31,45,31,35,31,35,30,163,31,194,31,194,30,63,31,215,31,24,31,24,30,137,31,140,31,64,31,115,31,115,30,226,31,161,31,61,31,210,31,152,31,191,31,136,31,52,31,199,31,91,31,91,30,91,29,91,28,216,31,19,31,19,30,89,31,36,31,144,31,249,31,249,30,62,31,28,31,88,31,244,31,225,31,131,31,65,31,213,31,252,31,252,30,53,31,176,31,176,30,45,31,189,31,36,31,36,30,137,31,84,31,254,31,43,31,238,31,238,30,205,31,47,31,100,31,145,31,145,30,7,31,17,31,17,30,67,31,119,31,119,30,115,31,115,30,102,31,171,31,10,31,234,31,168,31,123,31,18,31,117,31,27,31,27,30,27,29,27,28,27,27,27,26,27,25,194,31,149,31,149,30,90,31,108,31,240,31,240,30,240,29,114,31,33,31,146,31,73,31,73,30,58,31,171,31,218,31,218,30,160,31,160,30,27,31,12,31,200,31,208,31,208,30,9,31,61,31,23,31,21,31,78,31,78,30,78,29,136,31,10,31,95,31,95,30,18,31,216,31,152,31,127,31,234,31,219,31,148,31,172,31,150,31,84,31,71,31,71,30,148,31,144,31,144,30,58,31,165,31,114,31,114,30,246,31,145,31,130,31,130,30,64,31,101,31,65,31,50,31,228,31,215,31,238,31,146,31,146,30,146,29,83,31,246,31,246,30,246,29,240,31,232,31,55,31,131,31,221,31,159,31,39,31,20,31,186,31,53,31,220,31,243,31,226,31,226,30,22,31,178,31,178,30,104,31,154,31,11,31,244,31,244,30,187,31,126,31,126,30,186,31,57,31,139,31,139,30,139,29,139,28,32,31,32,30,163,31,152,31,86,31,124,31,51,31,128,31,54,31,150,31,177,31,187,31,253,31,154,31,38,31,167,31,183,31,185,31,124,31,87,31,124,31,165,31,100,31,100,30,199,31,240,31,59,31,92,31,191,31,140,31,138,31,68,31,129,31,129,30,250,31,250,30,226,31,12,31,119,31,4,31,4,30,173,31,163,31,16,31,66,31,121,31,121,30,97,31,211,31,57,31,207,31,248,31,120,31,111,31,111,30,96,31,171,31,141,31,103,31,148,31,148,30,148,29,175,31,83,31,60,31,136,31,34,31,34,30,119,31,97,31,97,30,31,31,31,30,31,29,58,31,226,31,121,31,111,31,223,31,104,31,218,31,117,31,249,31,243,31,243,30,78,31,125,31,16,31,16,30,198,31,198,30,134,31,249,31,233,31,233,30,233,29,39,31,202,31,81,31,175,31,175,30,54,31,41,31,41,30,157,31,43,31,249,31,47,31,47,30,44,31,245,31,157,31,91,31,91,30,14,31,74,31,58,31,93,31,93,30,5,31,222,31,121,31,121,30,121,29,94,31,94,30,48,31,248,31,113,31,113,31,100,31,100,30,255,31,57,31,191,31,92,31,92,30,157,31,217,31,217,30,138,31,138,30,238,31,57,31,133,31,133,30,244,31,197,31,145,31,6,31,141,31,186,31,235,31,113,31,42,31,42,30,217,31,7,31,210,31,133,31,200,31,29,31,202,31,202,30,241,31,253,31,253,30,107,31,16,31,138,31,138,30,10,31,237,31,208,31,64,31,213,31,103,31,199,31,89,31,70,31,214,31,223,31,133,31,33,31,33,30,210,31,210,30,63,31,201,31,132,31,237,31,237,30,237,29,31,31,58,31,58,30,119,31,69,31,207,31,207,30,207,29,207,28,207,27,64,31,206,31,14,31,32,31,109,31,88,31,215,31,20,31,63,31,96,31,96,30,80,31,222,31,67,31,108,31,120,31,120,30,32,31,175,31,249,31,249,30,119,31,25,31,25,30,100,31,243,31,157,31,107,31,107,30,49,31,10,31,10,30,80,31,80,30,128,31,10,31,167,31,52,31,78,31,188,31,81,31,89,31,51,31,153,31,240,31,240,30,139,31,58,31,51,31,170,31,104,31,91,31,164,31,164,30,106,31,49,31,198,31,136,31,252,31,161,31,70,31,188,31,194,31,194,30,138,31,200,31,68,31,64,31,64,30,187,31,211,31,132,31,132,30,132,29,195,31,43,31,43,30,58,31,35,31,35,30,235,31,235,30,67,31,82,31,22,31,81,31,81,30,47,31,180,31,7,31,50,31,102,31,205,31,205,30,22,31,244,31,244,30,164,31,222,31,222,30,74,31,74,30,152,31,152,30,231,31,118,31,62,31,157,31,157,30,193,31,168,31,97,31,234,31,109,31,104,31,147,31,82,31,240,31,145,31,204,31,231,31,83,31,83,30,83,29,83,28,149,31,140,31,237,31,168,31,229,31,127,31,213,31,213,30,213,29,38,31,102,31,112,31,81,31,157,31,157,30,77,31,165,31,149,31,18,31,207,31,5,31,248,31,240,31,54,31,61,31,17,31,203,31,203,30,203,29,203,28,220,31,64,31,64,30,175,31,175,30,251,31,169,31,19,31,19,30,213,31,159,31,6,31,7,31,7,30,117,31,130,31,156,31,30,31,62,31,194,31,156,31,156,30,135,31,143,31,12,31,234,31,195,31,208,31,71,31,88,31,212,31,185,31,42,31,122,31,198,31,7,31,7,30,115,31,90,31,177,31,25,31,25,31,29,31,198,31,198,30,198,29,70,31,242,31,48,31,48,30,48,31,250,31,118,31,57,31,111,31,149,31,109,31,141,31,141,30,41,31,180,31,180,30,122,31,90,31,87,31,153,31,208,31,9,31,9,30,172,31,103,31,128,31,107,31,246,31,9,31,191,31,12,31,12,30,179,31,147,31,207,31,20,31,138,31,138,30,217,31,217,30,247,31,247,30,247,29,160,31,160,30,230,31,38,31,133,31,222,31,201,31,242,31,242,30,13,31,208,31,200,31,74,31,85,31,235,31,92,31,232,31,159,31,159,30,159,29,159,28,170,31,175,31,175,30,126,31,128,31,175,31,248,31,248,30,191,31,191,30,252,31,178,31,178,30,232,31,143,31,109,31,38,31,189,31,170,31,142,31,82,31,82,30,70,31,77,31,77,30,28,31,28,30,28,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
