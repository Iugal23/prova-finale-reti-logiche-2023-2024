-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 651;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (91,0,39,0,149,0,51,0,245,0,178,0,110,0,164,0,217,0,0,0,165,0,124,0,251,0,194,0,1,0,182,0,176,0,96,0,0,0,94,0,86,0,0,0,0,0,105,0,16,0,72,0,175,0,30,0,39,0,0,0,141,0,167,0,0,0,32,0,160,0,154,0,0,0,0,0,238,0,0,0,200,0,176,0,215,0,255,0,59,0,233,0,199,0,0,0,240,0,59,0,150,0,71,0,178,0,11,0,203,0,32,0,0,0,157,0,0,0,140,0,91,0,206,0,249,0,149,0,0,0,183,0,0,0,44,0,18,0,0,0,255,0,0,0,170,0,8,0,205,0,221,0,54,0,15,0,181,0,59,0,148,0,42,0,0,0,246,0,134,0,49,0,56,0,57,0,24,0,0,0,0,0,144,0,158,0,173,0,215,0,110,0,250,0,132,0,148,0,133,0,228,0,245,0,0,0,0,0,216,0,0,0,209,0,127,0,159,0,218,0,0,0,234,0,253,0,192,0,52,0,238,0,222,0,10,0,167,0,241,0,219,0,56,0,210,0,226,0,155,0,249,0,250,0,233,0,19,0,52,0,251,0,0,0,126,0,0,0,0,0,38,0,173,0,23,0,239,0,61,0,68,0,0,0,0,0,216,0,0,0,0,0,212,0,241,0,41,0,76,0,222,0,114,0,4,0,0,0,235,0,60,0,213,0,56,0,183,0,200,0,37,0,84,0,175,0,202,0,49,0,72,0,123,0,0,0,184,0,117,0,199,0,207,0,0,0,143,0,35,0,0,0,12,0,60,0,244,0,76,0,25,0,201,0,176,0,127,0,0,0,174,0,214,0,217,0,72,0,87,0,1,0,149,0,78,0,109,0,0,0,111,0,170,0,0,0,160,0,81,0,203,0,52,0,151,0,129,0,253,0,78,0,0,0,169,0,102,0,0,0,188,0,23,0,158,0,21,0,98,0,40,0,131,0,0,0,246,0,109,0,120,0,249,0,8,0,22,0,245,0,76,0,0,0,0,0,22,0,176,0,196,0,220,0,74,0,8,0,156,0,177,0,61,0,28,0,188,0,190,0,135,0,0,0,0,0,145,0,131,0,111,0,96,0,69,0,0,0,0,0,136,0,124,0,119,0,177,0,0,0,157,0,192,0,177,0,61,0,243,0,0,0,0,0,213,0,209,0,11,0,0,0,242,0,242,0,29,0,60,0,120,0,94,0,60,0,87,0,170,0,92,0,109,0,10,0,219,0,72,0,144,0,33,0,13,0,165,0,8,0,147,0,35,0,44,0,0,0,26,0,0,0,23,0,228,0,175,0,189,0,184,0,191,0,90,0,0,0,0,0,64,0,28,0,72,0,94,0,0,0,183,0,38,0,65,0,0,0,0,0,17,0,47,0,171,0,148,0,67,0,0,0,184,0,0,0,0,0,154,0,146,0,206,0,0,0,91,0,0,0,0,0,85,0,203,0,41,0,233,0,35,0,249,0,202,0,216,0,196,0,185,0,199,0,105,0,183,0,103,0,139,0,90,0,6,0,228,0,26,0,111,0,93,0,174,0,105,0,36,0,193,0,248,0,0,0,0,0,109,0,8,0,192,0,0,0,74,0,0,0,0,0,4,0,58,0,0,0,203,0,0,0,145,0,0,0,47,0,184,0,47,0,0,0,28,0,0,0,221,0,13,0,232,0,158,0,192,0,193,0,214,0,0,0,190,0,139,0,116,0,125,0,62,0,146,0,217,0,77,0,132,0,212,0,61,0,122,0,176,0,247,0,76,0,23,0,0,0,0,0,170,0,243,0,0,0,0,0,127,0,0,0,0,0,0,0,80,0,0,0,69,0,90,0,0,0,23,0,232,0,109,0,0,0,94,0,0,0,126,0,0,0,248,0,178,0,100,0,172,0,176,0,0,0,43,0,200,0,116,0,243,0,100,0,139,0,16,0,137,0,35,0,28,0,180,0,90,0,0,0,203,0,43,0,218,0,0,0,214,0,165,0,60,0,82,0,77,0,226,0,126,0,0,0,0,0,179,0,222,0,122,0,160,0,0,0,187,0,0,0,151,0,0,0,214,0,0,0,82,0,190,0,0,0,91,0,57,0,126,0,75,0,60,0,189,0,132,0,62,0,15,0,0,0,116,0,21,0,111,0,234,0,0,0,0,0,201,0,200,0,216,0,9,0,24,0,29,0,201,0,152,0,39,0,139,0,15,0,64,0,170,0,0,0,125,0,0,0,0,0,163,0,0,0,146,0,56,0,114,0,47,0,173,0,190,0,40,0,131,0,0,0,0,0,249,0,198,0,139,0,30,0,139,0,34,0,41,0,92,0,0,0,110,0,136,0,0,0,77,0,197,0,192,0,236,0,0,0,0,0,0,0,0,0,56,0,82,0,188,0,0,0,141,0,44,0,82,0,212,0,97,0,45,0,0,0,174,0,160,0,98,0,46,0,20,0,196,0,254,0,247,0,59,0,55,0,134,0,70,0,0,0,0,0,154,0,65,0,192,0,0,0,225,0,246,0,231,0,225,0,195,0,103,0,221,0,54,0,187,0,4,0,130,0,232,0,0,0,161,0,222,0,98,0,0,0,145,0,76,0,20,0,108,0,21,0,0,0,133,0,0,0,0,0,143,0,145,0,173,0,22,0,0,0,24,0,231,0,216,0,0,0,0,0,254,0,106,0,88,0,89,0,211,0,11,0,232,0,73,0,0,0,2,0,0,0,0,0,111,0,0,0,138,0,0,0,0,0,133,0,59,0,156,0,69,0,164,0,29,0,57,0,66,0,161,0,59,0,200,0,39,0,158,0,69,0,0,0,63,0,0,0,5,0,15,0,167,0,0,0,17,0,134,0,220,0,152,0,172,0,10,0,76,0,236,0,235,0,97,0,251,0,187,0,92,0,107,0,102,0,86,0);
signal scenario_full  : scenario_type := (91,31,39,31,149,31,51,31,245,31,178,31,110,31,164,31,217,31,217,30,165,31,124,31,251,31,194,31,1,31,182,31,176,31,96,31,96,30,94,31,86,31,86,30,86,29,105,31,16,31,72,31,175,31,30,31,39,31,39,30,141,31,167,31,167,30,32,31,160,31,154,31,154,30,154,29,238,31,238,30,200,31,176,31,215,31,255,31,59,31,233,31,199,31,199,30,240,31,59,31,150,31,71,31,178,31,11,31,203,31,32,31,32,30,157,31,157,30,140,31,91,31,206,31,249,31,149,31,149,30,183,31,183,30,44,31,18,31,18,30,255,31,255,30,170,31,8,31,205,31,221,31,54,31,15,31,181,31,59,31,148,31,42,31,42,30,246,31,134,31,49,31,56,31,57,31,24,31,24,30,24,29,144,31,158,31,173,31,215,31,110,31,250,31,132,31,148,31,133,31,228,31,245,31,245,30,245,29,216,31,216,30,209,31,127,31,159,31,218,31,218,30,234,31,253,31,192,31,52,31,238,31,222,31,10,31,167,31,241,31,219,31,56,31,210,31,226,31,155,31,249,31,250,31,233,31,19,31,52,31,251,31,251,30,126,31,126,30,126,29,38,31,173,31,23,31,239,31,61,31,68,31,68,30,68,29,216,31,216,30,216,29,212,31,241,31,41,31,76,31,222,31,114,31,4,31,4,30,235,31,60,31,213,31,56,31,183,31,200,31,37,31,84,31,175,31,202,31,49,31,72,31,123,31,123,30,184,31,117,31,199,31,207,31,207,30,143,31,35,31,35,30,12,31,60,31,244,31,76,31,25,31,201,31,176,31,127,31,127,30,174,31,214,31,217,31,72,31,87,31,1,31,149,31,78,31,109,31,109,30,111,31,170,31,170,30,160,31,81,31,203,31,52,31,151,31,129,31,253,31,78,31,78,30,169,31,102,31,102,30,188,31,23,31,158,31,21,31,98,31,40,31,131,31,131,30,246,31,109,31,120,31,249,31,8,31,22,31,245,31,76,31,76,30,76,29,22,31,176,31,196,31,220,31,74,31,8,31,156,31,177,31,61,31,28,31,188,31,190,31,135,31,135,30,135,29,145,31,131,31,111,31,96,31,69,31,69,30,69,29,136,31,124,31,119,31,177,31,177,30,157,31,192,31,177,31,61,31,243,31,243,30,243,29,213,31,209,31,11,31,11,30,242,31,242,31,29,31,60,31,120,31,94,31,60,31,87,31,170,31,92,31,109,31,10,31,219,31,72,31,144,31,33,31,13,31,165,31,8,31,147,31,35,31,44,31,44,30,26,31,26,30,23,31,228,31,175,31,189,31,184,31,191,31,90,31,90,30,90,29,64,31,28,31,72,31,94,31,94,30,183,31,38,31,65,31,65,30,65,29,17,31,47,31,171,31,148,31,67,31,67,30,184,31,184,30,184,29,154,31,146,31,206,31,206,30,91,31,91,30,91,29,85,31,203,31,41,31,233,31,35,31,249,31,202,31,216,31,196,31,185,31,199,31,105,31,183,31,103,31,139,31,90,31,6,31,228,31,26,31,111,31,93,31,174,31,105,31,36,31,193,31,248,31,248,30,248,29,109,31,8,31,192,31,192,30,74,31,74,30,74,29,4,31,58,31,58,30,203,31,203,30,145,31,145,30,47,31,184,31,47,31,47,30,28,31,28,30,221,31,13,31,232,31,158,31,192,31,193,31,214,31,214,30,190,31,139,31,116,31,125,31,62,31,146,31,217,31,77,31,132,31,212,31,61,31,122,31,176,31,247,31,76,31,23,31,23,30,23,29,170,31,243,31,243,30,243,29,127,31,127,30,127,29,127,28,80,31,80,30,69,31,90,31,90,30,23,31,232,31,109,31,109,30,94,31,94,30,126,31,126,30,248,31,178,31,100,31,172,31,176,31,176,30,43,31,200,31,116,31,243,31,100,31,139,31,16,31,137,31,35,31,28,31,180,31,90,31,90,30,203,31,43,31,218,31,218,30,214,31,165,31,60,31,82,31,77,31,226,31,126,31,126,30,126,29,179,31,222,31,122,31,160,31,160,30,187,31,187,30,151,31,151,30,214,31,214,30,82,31,190,31,190,30,91,31,57,31,126,31,75,31,60,31,189,31,132,31,62,31,15,31,15,30,116,31,21,31,111,31,234,31,234,30,234,29,201,31,200,31,216,31,9,31,24,31,29,31,201,31,152,31,39,31,139,31,15,31,64,31,170,31,170,30,125,31,125,30,125,29,163,31,163,30,146,31,56,31,114,31,47,31,173,31,190,31,40,31,131,31,131,30,131,29,249,31,198,31,139,31,30,31,139,31,34,31,41,31,92,31,92,30,110,31,136,31,136,30,77,31,197,31,192,31,236,31,236,30,236,29,236,28,236,27,56,31,82,31,188,31,188,30,141,31,44,31,82,31,212,31,97,31,45,31,45,30,174,31,160,31,98,31,46,31,20,31,196,31,254,31,247,31,59,31,55,31,134,31,70,31,70,30,70,29,154,31,65,31,192,31,192,30,225,31,246,31,231,31,225,31,195,31,103,31,221,31,54,31,187,31,4,31,130,31,232,31,232,30,161,31,222,31,98,31,98,30,145,31,76,31,20,31,108,31,21,31,21,30,133,31,133,30,133,29,143,31,145,31,173,31,22,31,22,30,24,31,231,31,216,31,216,30,216,29,254,31,106,31,88,31,89,31,211,31,11,31,232,31,73,31,73,30,2,31,2,30,2,29,111,31,111,30,138,31,138,30,138,29,133,31,59,31,156,31,69,31,164,31,29,31,57,31,66,31,161,31,59,31,200,31,39,31,158,31,69,31,69,30,63,31,63,30,5,31,15,31,167,31,167,30,17,31,134,31,220,31,152,31,172,31,10,31,76,31,236,31,235,31,97,31,251,31,187,31,92,31,107,31,102,31,86,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
