-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_170 is
end project_tb_170;

architecture project_tb_arch_170 of project_tb_170 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 861;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,131,0,133,0,238,0,105,0,201,0,0,0,144,0,42,0,36,0,101,0,0,0,212,0,50,0,31,0,25,0,0,0,57,0,0,0,171,0,0,0,13,0,79,0,87,0,3,0,145,0,61,0,152,0,46,0,75,0,2,0,143,0,63,0,229,0,57,0,9,0,0,0,11,0,60,0,46,0,116,0,50,0,151,0,81,0,56,0,161,0,219,0,0,0,200,0,110,0,0,0,141,0,0,0,46,0,211,0,0,0,118,0,248,0,43,0,234,0,0,0,41,0,104,0,58,0,69,0,32,0,182,0,0,0,42,0,133,0,200,0,0,0,0,0,51,0,29,0,202,0,0,0,40,0,0,0,0,0,201,0,0,0,154,0,0,0,51,0,74,0,58,0,0,0,112,0,215,0,79,0,0,0,41,0,75,0,148,0,96,0,43,0,118,0,48,0,247,0,85,0,0,0,0,0,136,0,199,0,0,0,204,0,19,0,193,0,0,0,41,0,5,0,144,0,251,0,246,0,120,0,204,0,172,0,217,0,251,0,167,0,0,0,98,0,153,0,117,0,0,0,218,0,106,0,0,0,196,0,127,0,0,0,128,0,58,0,38,0,226,0,245,0,38,0,169,0,104,0,19,0,122,0,0,0,239,0,0,0,0,0,177,0,0,0,240,0,49,0,18,0,249,0,0,0,108,0,253,0,114,0,68,0,246,0,56,0,220,0,61,0,101,0,153,0,116,0,167,0,0,0,124,0,240,0,214,0,187,0,198,0,201,0,216,0,16,0,0,0,4,0,0,0,228,0,0,0,28,0,218,0,7,0,0,0,208,0,198,0,190,0,6,0,28,0,196,0,14,0,177,0,125,0,194,0,26,0,0,0,235,0,9,0,234,0,89,0,0,0,55,0,207,0,0,0,209,0,192,0,213,0,0,0,153,0,238,0,0,0,255,0,0,0,22,0,114,0,38,0,131,0,0,0,118,0,0,0,36,0,253,0,35,0,0,0,113,0,0,0,133,0,175,0,195,0,162,0,0,0,42,0,214,0,18,0,234,0,0,0,31,0,184,0,128,0,0,0,111,0,0,0,0,0,0,0,71,0,0,0,81,0,46,0,240,0,206,0,116,0,86,0,223,0,78,0,0,0,200,0,0,0,157,0,90,0,0,0,21,0,250,0,29,0,238,0,56,0,50,0,0,0,132,0,0,0,25,0,179,0,50,0,4,0,56,0,97,0,192,0,34,0,0,0,60,0,230,0,230,0,8,0,7,0,79,0,115,0,164,0,180,0,63,0,246,0,189,0,86,0,0,0,0,0,52,0,145,0,150,0,58,0,0,0,191,0,0,0,0,0,13,0,175,0,168,0,0,0,5,0,112,0,176,0,88,0,0,0,215,0,0,0,201,0,234,0,0,0,13,0,102,0,0,0,60,0,235,0,200,0,0,0,54,0,179,0,59,0,121,0,54,0,26,0,69,0,134,0,126,0,173,0,242,0,4,0,83,0,228,0,50,0,0,0,192,0,192,0,13,0,213,0,0,0,0,0,0,0,148,0,0,0,0,0,192,0,112,0,150,0,126,0,105,0,251,0,110,0,194,0,1,0,18,0,177,0,112,0,184,0,145,0,0,0,122,0,235,0,147,0,0,0,0,0,27,0,64,0,0,0,239,0,219,0,26,0,132,0,0,0,0,0,117,0,130,0,0,0,0,0,0,0,17,0,113,0,218,0,172,0,6,0,3,0,0,0,185,0,0,0,184,0,57,0,116,0,227,0,0,0,123,0,91,0,98,0,25,0,0,0,0,0,130,0,45,0,56,0,196,0,29,0,57,0,67,0,141,0,177,0,131,0,39,0,145,0,0,0,179,0,0,0,197,0,254,0,80,0,4,0,211,0,0,0,0,0,0,0,174,0,156,0,193,0,89,0,79,0,177,0,0,0,152,0,0,0,0,0,86,0,177,0,13,0,0,0,3,0,132,0,153,0,28,0,80,0,0,0,200,0,0,0,124,0,62,0,232,0,3,0,131,0,194,0,27,0,27,0,44,0,0,0,105,0,20,0,95,0,87,0,0,0,171,0,127,0,54,0,0,0,166,0,123,0,31,0,0,0,178,0,210,0,77,0,153,0,59,0,32,0,172,0,243,0,42,0,34,0,136,0,108,0,105,0,87,0,220,0,191,0,227,0,0,0,235,0,61,0,113,0,36,0,159,0,197,0,184,0,212,0,123,0,154,0,44,0,181,0,197,0,39,0,0,0,177,0,0,0,0,0,89,0,248,0,120,0,6,0,0,0,0,0,0,0,112,0,195,0,142,0,36,0,225,0,81,0,71,0,152,0,111,0,0,0,227,0,172,0,0,0,193,0,255,0,202,0,55,0,0,0,0,0,116,0,0,0,100,0,70,0,0,0,0,0,0,0,244,0,33,0,219,0,103,0,6,0,89,0,0,0,69,0,0,0,151,0,218,0,0,0,200,0,22,0,232,0,228,0,209,0,166,0,144,0,6,0,0,0,16,0,0,0,0,0,188,0,221,0,0,0,132,0,142,0,0,0,93,0,76,0,100,0,230,0,137,0,29,0,93,0,42,0,178,0,170,0,8,0,182,0,32,0,0,0,54,0,151,0,0,0,100,0,72,0,137,0,0,0,252,0,151,0,50,0,1,0,22,0,236,0,69,0,33,0,171,0,252,0,15,0,93,0,14,0,153,0,242,0,234,0,176,0,0,0,97,0,172,0,194,0,85,0,83,0,0,0,0,0,6,0,108,0,32,0,23,0,164,0,0,0,232,0,244,0,96,0,144,0,19,0,40,0,103,0,231,0,117,0,0,0,221,0,204,0,232,0,0,0,0,0,137,0,206,0,159,0,101,0,0,0,6,0,0,0,68,0,227,0,0,0,0,0,85,0,0,0,0,0,0,0,0,0,56,0,0,0,79,0,0,0,163,0,51,0,199,0,99,0,0,0,18,0,0,0,230,0,42,0,125,0,0,0,39,0,90,0,164,0,23,0,3,0,7,0,105,0,121,0,38,0,172,0,77,0,68,0,27,0,148,0,243,0,212,0,239,0,228,0,225,0,0,0,0,0,0,0,32,0,98,0,126,0,58,0,70,0,122,0,171,0,195,0,224,0,91,0,0,0,66,0,176,0,234,0,251,0,90,0,254,0,0,0,0,0,245,0,31,0,236,0,103,0,0,0,0,0,155,0,0,0,198,0,207,0,216,0,94,0,224,0,150,0,0,0,163,0,223,0,240,0,0,0,198,0,10,0,161,0,31,0,66,0,56,0,32,0,0,0,81,0,8,0,16,0,197,0,113,0,224,0,0,0,186,0,0,0,27,0,3,0,250,0,5,0,62,0,13,0,0,0,186,0,88,0,195,0,27,0,211,0,0,0,156,0,0,0,58,0,100,0,71,0,166,0,0,0,0,0,38,0,17,0,160,0,132,0,115,0,26,0,207,0,0,0,3,0,0,0,28,0,143,0,60,0,32,0,0,0,253,0,249,0,181,0,229,0,228,0,0,0,69,0,11,0,239,0,202,0,228,0,158,0,227,0,227,0,0,0,251,0,4,0,180,0,91,0,41,0,253,0,129,0,0,0,121,0,0,0,118,0,0,0,59,0,54,0,0,0,47,0,135,0,27,0,123,0,51,0,163,0,217,0,0,0,20,0,250,0,0,0,0,0,152,0,245,0,36,0,246,0,0,0,168,0,9,0,151,0,103,0,28,0,77,0,41,0,126,0,152,0,171,0,27,0,18,0,208,0,96,0,182,0,103,0,243,0,222,0,51,0,37,0,0,0,130,0,220,0,8,0,147,0,167,0,210,0,159,0,42,0,138,0,0,0,57,0,153,0,228,0,145,0);
signal scenario_full  : scenario_type := (189,31,131,31,133,31,238,31,105,31,201,31,201,30,144,31,42,31,36,31,101,31,101,30,212,31,50,31,31,31,25,31,25,30,57,31,57,30,171,31,171,30,13,31,79,31,87,31,3,31,145,31,61,31,152,31,46,31,75,31,2,31,143,31,63,31,229,31,57,31,9,31,9,30,11,31,60,31,46,31,116,31,50,31,151,31,81,31,56,31,161,31,219,31,219,30,200,31,110,31,110,30,141,31,141,30,46,31,211,31,211,30,118,31,248,31,43,31,234,31,234,30,41,31,104,31,58,31,69,31,32,31,182,31,182,30,42,31,133,31,200,31,200,30,200,29,51,31,29,31,202,31,202,30,40,31,40,30,40,29,201,31,201,30,154,31,154,30,51,31,74,31,58,31,58,30,112,31,215,31,79,31,79,30,41,31,75,31,148,31,96,31,43,31,118,31,48,31,247,31,85,31,85,30,85,29,136,31,199,31,199,30,204,31,19,31,193,31,193,30,41,31,5,31,144,31,251,31,246,31,120,31,204,31,172,31,217,31,251,31,167,31,167,30,98,31,153,31,117,31,117,30,218,31,106,31,106,30,196,31,127,31,127,30,128,31,58,31,38,31,226,31,245,31,38,31,169,31,104,31,19,31,122,31,122,30,239,31,239,30,239,29,177,31,177,30,240,31,49,31,18,31,249,31,249,30,108,31,253,31,114,31,68,31,246,31,56,31,220,31,61,31,101,31,153,31,116,31,167,31,167,30,124,31,240,31,214,31,187,31,198,31,201,31,216,31,16,31,16,30,4,31,4,30,228,31,228,30,28,31,218,31,7,31,7,30,208,31,198,31,190,31,6,31,28,31,196,31,14,31,177,31,125,31,194,31,26,31,26,30,235,31,9,31,234,31,89,31,89,30,55,31,207,31,207,30,209,31,192,31,213,31,213,30,153,31,238,31,238,30,255,31,255,30,22,31,114,31,38,31,131,31,131,30,118,31,118,30,36,31,253,31,35,31,35,30,113,31,113,30,133,31,175,31,195,31,162,31,162,30,42,31,214,31,18,31,234,31,234,30,31,31,184,31,128,31,128,30,111,31,111,30,111,29,111,28,71,31,71,30,81,31,46,31,240,31,206,31,116,31,86,31,223,31,78,31,78,30,200,31,200,30,157,31,90,31,90,30,21,31,250,31,29,31,238,31,56,31,50,31,50,30,132,31,132,30,25,31,179,31,50,31,4,31,56,31,97,31,192,31,34,31,34,30,60,31,230,31,230,31,8,31,7,31,79,31,115,31,164,31,180,31,63,31,246,31,189,31,86,31,86,30,86,29,52,31,145,31,150,31,58,31,58,30,191,31,191,30,191,29,13,31,175,31,168,31,168,30,5,31,112,31,176,31,88,31,88,30,215,31,215,30,201,31,234,31,234,30,13,31,102,31,102,30,60,31,235,31,200,31,200,30,54,31,179,31,59,31,121,31,54,31,26,31,69,31,134,31,126,31,173,31,242,31,4,31,83,31,228,31,50,31,50,30,192,31,192,31,13,31,213,31,213,30,213,29,213,28,148,31,148,30,148,29,192,31,112,31,150,31,126,31,105,31,251,31,110,31,194,31,1,31,18,31,177,31,112,31,184,31,145,31,145,30,122,31,235,31,147,31,147,30,147,29,27,31,64,31,64,30,239,31,219,31,26,31,132,31,132,30,132,29,117,31,130,31,130,30,130,29,130,28,17,31,113,31,218,31,172,31,6,31,3,31,3,30,185,31,185,30,184,31,57,31,116,31,227,31,227,30,123,31,91,31,98,31,25,31,25,30,25,29,130,31,45,31,56,31,196,31,29,31,57,31,67,31,141,31,177,31,131,31,39,31,145,31,145,30,179,31,179,30,197,31,254,31,80,31,4,31,211,31,211,30,211,29,211,28,174,31,156,31,193,31,89,31,79,31,177,31,177,30,152,31,152,30,152,29,86,31,177,31,13,31,13,30,3,31,132,31,153,31,28,31,80,31,80,30,200,31,200,30,124,31,62,31,232,31,3,31,131,31,194,31,27,31,27,31,44,31,44,30,105,31,20,31,95,31,87,31,87,30,171,31,127,31,54,31,54,30,166,31,123,31,31,31,31,30,178,31,210,31,77,31,153,31,59,31,32,31,172,31,243,31,42,31,34,31,136,31,108,31,105,31,87,31,220,31,191,31,227,31,227,30,235,31,61,31,113,31,36,31,159,31,197,31,184,31,212,31,123,31,154,31,44,31,181,31,197,31,39,31,39,30,177,31,177,30,177,29,89,31,248,31,120,31,6,31,6,30,6,29,6,28,112,31,195,31,142,31,36,31,225,31,81,31,71,31,152,31,111,31,111,30,227,31,172,31,172,30,193,31,255,31,202,31,55,31,55,30,55,29,116,31,116,30,100,31,70,31,70,30,70,29,70,28,244,31,33,31,219,31,103,31,6,31,89,31,89,30,69,31,69,30,151,31,218,31,218,30,200,31,22,31,232,31,228,31,209,31,166,31,144,31,6,31,6,30,16,31,16,30,16,29,188,31,221,31,221,30,132,31,142,31,142,30,93,31,76,31,100,31,230,31,137,31,29,31,93,31,42,31,178,31,170,31,8,31,182,31,32,31,32,30,54,31,151,31,151,30,100,31,72,31,137,31,137,30,252,31,151,31,50,31,1,31,22,31,236,31,69,31,33,31,171,31,252,31,15,31,93,31,14,31,153,31,242,31,234,31,176,31,176,30,97,31,172,31,194,31,85,31,83,31,83,30,83,29,6,31,108,31,32,31,23,31,164,31,164,30,232,31,244,31,96,31,144,31,19,31,40,31,103,31,231,31,117,31,117,30,221,31,204,31,232,31,232,30,232,29,137,31,206,31,159,31,101,31,101,30,6,31,6,30,68,31,227,31,227,30,227,29,85,31,85,30,85,29,85,28,85,27,56,31,56,30,79,31,79,30,163,31,51,31,199,31,99,31,99,30,18,31,18,30,230,31,42,31,125,31,125,30,39,31,90,31,164,31,23,31,3,31,7,31,105,31,121,31,38,31,172,31,77,31,68,31,27,31,148,31,243,31,212,31,239,31,228,31,225,31,225,30,225,29,225,28,32,31,98,31,126,31,58,31,70,31,122,31,171,31,195,31,224,31,91,31,91,30,66,31,176,31,234,31,251,31,90,31,254,31,254,30,254,29,245,31,31,31,236,31,103,31,103,30,103,29,155,31,155,30,198,31,207,31,216,31,94,31,224,31,150,31,150,30,163,31,223,31,240,31,240,30,198,31,10,31,161,31,31,31,66,31,56,31,32,31,32,30,81,31,8,31,16,31,197,31,113,31,224,31,224,30,186,31,186,30,27,31,3,31,250,31,5,31,62,31,13,31,13,30,186,31,88,31,195,31,27,31,211,31,211,30,156,31,156,30,58,31,100,31,71,31,166,31,166,30,166,29,38,31,17,31,160,31,132,31,115,31,26,31,207,31,207,30,3,31,3,30,28,31,143,31,60,31,32,31,32,30,253,31,249,31,181,31,229,31,228,31,228,30,69,31,11,31,239,31,202,31,228,31,158,31,227,31,227,31,227,30,251,31,4,31,180,31,91,31,41,31,253,31,129,31,129,30,121,31,121,30,118,31,118,30,59,31,54,31,54,30,47,31,135,31,27,31,123,31,51,31,163,31,217,31,217,30,20,31,250,31,250,30,250,29,152,31,245,31,36,31,246,31,246,30,168,31,9,31,151,31,103,31,28,31,77,31,41,31,126,31,152,31,171,31,27,31,18,31,208,31,96,31,182,31,103,31,243,31,222,31,51,31,37,31,37,30,130,31,220,31,8,31,147,31,167,31,210,31,159,31,42,31,138,31,138,30,57,31,153,31,228,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
