-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 821;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,8,0,228,0,194,0,71,0,250,0,0,0,109,0,0,0,189,0,0,0,17,0,158,0,19,0,206,0,28,0,227,0,20,0,248,0,217,0,8,0,240,0,252,0,89,0,0,0,0,0,0,0,0,0,33,0,0,0,244,0,99,0,10,0,72,0,0,0,0,0,230,0,93,0,0,0,51,0,0,0,105,0,98,0,197,0,105,0,0,0,189,0,59,0,169,0,245,0,173,0,137,0,24,0,144,0,247,0,219,0,185,0,153,0,175,0,64,0,138,0,141,0,212,0,0,0,244,0,75,0,0,0,230,0,195,0,144,0,21,0,179,0,0,0,0,0,135,0,239,0,44,0,60,0,14,0,46,0,57,0,140,0,112,0,0,0,130,0,11,0,193,0,206,0,0,0,93,0,39,0,233,0,127,0,0,0,203,0,164,0,68,0,0,0,8,0,189,0,0,0,57,0,69,0,69,0,46,0,162,0,0,0,133,0,146,0,153,0,133,0,0,0,78,0,66,0,113,0,254,0,52,0,200,0,13,0,217,0,35,0,91,0,156,0,67,0,151,0,127,0,94,0,208,0,0,0,167,0,60,0,83,0,76,0,3,0,0,0,0,0,211,0,0,0,17,0,0,0,47,0,69,0,0,0,178,0,174,0,242,0,201,0,0,0,0,0,212,0,104,0,168,0,35,0,162,0,2,0,153,0,93,0,230,0,58,0,159,0,236,0,181,0,210,0,158,0,0,0,0,0,0,0,255,0,188,0,182,0,138,0,76,0,246,0,235,0,143,0,135,0,29,0,228,0,0,0,78,0,105,0,221,0,122,0,0,0,103,0,0,0,17,0,195,0,229,0,0,0,156,0,0,0,176,0,0,0,133,0,37,0,136,0,240,0,156,0,0,0,0,0,150,0,27,0,53,0,0,0,179,0,138,0,88,0,243,0,51,0,27,0,133,0,4,0,244,0,5,0,0,0,186,0,67,0,25,0,63,0,214,0,0,0,107,0,166,0,0,0,127,0,110,0,254,0,4,0,176,0,141,0,61,0,202,0,0,0,0,0,236,0,142,0,245,0,127,0,69,0,0,0,222,0,0,0,128,0,0,0,0,0,75,0,65,0,50,0,162,0,183,0,37,0,0,0,0,0,99,0,0,0,202,0,152,0,26,0,0,0,28,0,101,0,0,0,44,0,0,0,0,0,26,0,0,0,202,0,94,0,191,0,0,0,253,0,0,0,48,0,239,0,0,0,169,0,0,0,56,0,46,0,134,0,107,0,0,0,80,0,150,0,4,0,88,0,161,0,57,0,0,0,86,0,0,0,122,0,0,0,3,0,90,0,75,0,156,0,0,0,0,0,133,0,253,0,0,0,0,0,0,0,74,0,23,0,246,0,115,0,41,0,0,0,96,0,156,0,44,0,102,0,0,0,119,0,149,0,114,0,0,0,0,0,53,0,36,0,2,0,133,0,62,0,132,0,219,0,0,0,0,0,0,0,105,0,0,0,95,0,157,0,0,0,149,0,252,0,39,0,0,0,2,0,88,0,129,0,0,0,28,0,114,0,219,0,221,0,0,0,103,0,7,0,211,0,197,0,179,0,119,0,0,0,6,0,124,0,32,0,14,0,0,0,92,0,1,0,183,0,37,0,14,0,23,0,0,0,177,0,22,0,216,0,217,0,0,0,137,0,95,0,0,0,64,0,135,0,70,0,188,0,106,0,0,0,0,0,198,0,73,0,61,0,149,0,0,0,0,0,36,0,0,0,77,0,174,0,163,0,0,0,0,0,16,0,48,0,210,0,242,0,21,0,18,0,147,0,57,0,0,0,186,0,171,0,9,0,232,0,15,0,239,0,0,0,94,0,93,0,57,0,149,0,17,0,28,0,209,0,209,0,37,0,62,0,25,0,143,0,0,0,33,0,192,0,110,0,215,0,170,0,201,0,0,0,253,0,0,0,81,0,246,0,56,0,158,0,132,0,136,0,43,0,116,0,177,0,0,0,235,0,0,0,74,0,200,0,185,0,169,0,68,0,252,0,196,0,0,0,0,0,114,0,0,0,193,0,249,0,143,0,139,0,63,0,236,0,232,0,54,0,247,0,0,0,140,0,69,0,50,0,0,0,0,0,0,0,253,0,0,0,151,0,7,0,164,0,180,0,15,0,26,0,237,0,130,0,131,0,22,0,101,0,38,0,176,0,131,0,0,0,95,0,163,0,115,0,133,0,90,0,0,0,232,0,4,0,101,0,99,0,37,0,213,0,124,0,0,0,0,0,80,0,50,0,215,0,175,0,38,0,51,0,220,0,231,0,177,0,156,0,91,0,8,0,0,0,167,0,232,0,123,0,18,0,217,0,7,0,106,0,32,0,247,0,107,0,26,0,147,0,9,0,111,0,57,0,235,0,0,0,190,0,30,0,129,0,10,0,254,0,100,0,2,0,226,0,0,0,39,0,50,0,250,0,216,0,74,0,1,0,118,0,64,0,142,0,194,0,176,0,11,0,60,0,67,0,25,0,190,0,25,0,51,0,237,0,29,0,48,0,179,0,39,0,28,0,233,0,21,0,45,0,0,0,73,0,0,0,0,0,191,0,0,0,149,0,229,0,184,0,160,0,179,0,7,0,201,0,114,0,203,0,204,0,156,0,199,0,182,0,0,0,140,0,151,0,11,0,41,0,220,0,0,0,103,0,142,0,0,0,218,0,7,0,89,0,0,0,83,0,0,0,80,0,58,0,191,0,0,0,55,0,0,0,205,0,186,0,60,0,255,0,0,0,87,0,0,0,169,0,251,0,90,0,86,0,171,0,0,0,40,0,175,0,20,0,0,0,151,0,114,0,0,0,6,0,246,0,174,0,0,0,213,0,214,0,216,0,164,0,207,0,26,0,61,0,41,0,0,0,0,0,0,0,115,0,0,0,183,0,8,0,0,0,40,0,0,0,0,0,239,0,41,0,45,0,0,0,197,0,148,0,163,0,112,0,14,0,252,0,241,0,86,0,63,0,25,0,141,0,171,0,143,0,94,0,90,0,178,0,225,0,14,0,141,0,160,0,202,0,255,0,82,0,201,0,128,0,143,0,31,0,124,0,193,0,0,0,0,0,29,0,20,0,200,0,0,0,64,0,95,0,99,0,58,0,232,0,0,0,0,0,0,0,158,0,0,0,92,0,88,0,2,0,155,0,23,0,28,0,80,0,57,0,136,0,115,0,0,0,236,0,0,0,195,0,0,0,157,0,8,0,60,0,0,0,229,0,95,0,0,0,178,0,247,0,162,0,142,0,43,0,243,0,175,0,139,0,44,0,101,0,245,0,73,0,153,0,156,0,0,0,0,0,182,0,162,0,219,0,222,0,222,0,217,0,34,0,207,0,0,0,236,0,0,0,0,0,8,0,137,0,134,0,15,0,0,0,47,0,249,0,58,0,250,0,14,0,20,0,0,0,249,0,0,0,247,0,252,0,65,0,65,0,78,0,0,0,98,0,128,0,223,0,117,0,215,0,84,0,110,0,84,0,116,0,174,0,62,0,159,0,0,0,1,0,164,0,0,0,147,0,101,0,195,0,149,0,0,0,0,0,56,0,5,0,39,0,98,0,0,0,0,0,53,0,68,0,133,0,0,0,224,0,127,0,215,0,181,0,33,0,0,0,119,0,96,0,139,0,0,0,182,0,0,0,28,0,118,0);
signal scenario_full  : scenario_type := (24,31,8,31,228,31,194,31,71,31,250,31,250,30,109,31,109,30,189,31,189,30,17,31,158,31,19,31,206,31,28,31,227,31,20,31,248,31,217,31,8,31,240,31,252,31,89,31,89,30,89,29,89,28,89,27,33,31,33,30,244,31,99,31,10,31,72,31,72,30,72,29,230,31,93,31,93,30,51,31,51,30,105,31,98,31,197,31,105,31,105,30,189,31,59,31,169,31,245,31,173,31,137,31,24,31,144,31,247,31,219,31,185,31,153,31,175,31,64,31,138,31,141,31,212,31,212,30,244,31,75,31,75,30,230,31,195,31,144,31,21,31,179,31,179,30,179,29,135,31,239,31,44,31,60,31,14,31,46,31,57,31,140,31,112,31,112,30,130,31,11,31,193,31,206,31,206,30,93,31,39,31,233,31,127,31,127,30,203,31,164,31,68,31,68,30,8,31,189,31,189,30,57,31,69,31,69,31,46,31,162,31,162,30,133,31,146,31,153,31,133,31,133,30,78,31,66,31,113,31,254,31,52,31,200,31,13,31,217,31,35,31,91,31,156,31,67,31,151,31,127,31,94,31,208,31,208,30,167,31,60,31,83,31,76,31,3,31,3,30,3,29,211,31,211,30,17,31,17,30,47,31,69,31,69,30,178,31,174,31,242,31,201,31,201,30,201,29,212,31,104,31,168,31,35,31,162,31,2,31,153,31,93,31,230,31,58,31,159,31,236,31,181,31,210,31,158,31,158,30,158,29,158,28,255,31,188,31,182,31,138,31,76,31,246,31,235,31,143,31,135,31,29,31,228,31,228,30,78,31,105,31,221,31,122,31,122,30,103,31,103,30,17,31,195,31,229,31,229,30,156,31,156,30,176,31,176,30,133,31,37,31,136,31,240,31,156,31,156,30,156,29,150,31,27,31,53,31,53,30,179,31,138,31,88,31,243,31,51,31,27,31,133,31,4,31,244,31,5,31,5,30,186,31,67,31,25,31,63,31,214,31,214,30,107,31,166,31,166,30,127,31,110,31,254,31,4,31,176,31,141,31,61,31,202,31,202,30,202,29,236,31,142,31,245,31,127,31,69,31,69,30,222,31,222,30,128,31,128,30,128,29,75,31,65,31,50,31,162,31,183,31,37,31,37,30,37,29,99,31,99,30,202,31,152,31,26,31,26,30,28,31,101,31,101,30,44,31,44,30,44,29,26,31,26,30,202,31,94,31,191,31,191,30,253,31,253,30,48,31,239,31,239,30,169,31,169,30,56,31,46,31,134,31,107,31,107,30,80,31,150,31,4,31,88,31,161,31,57,31,57,30,86,31,86,30,122,31,122,30,3,31,90,31,75,31,156,31,156,30,156,29,133,31,253,31,253,30,253,29,253,28,74,31,23,31,246,31,115,31,41,31,41,30,96,31,156,31,44,31,102,31,102,30,119,31,149,31,114,31,114,30,114,29,53,31,36,31,2,31,133,31,62,31,132,31,219,31,219,30,219,29,219,28,105,31,105,30,95,31,157,31,157,30,149,31,252,31,39,31,39,30,2,31,88,31,129,31,129,30,28,31,114,31,219,31,221,31,221,30,103,31,7,31,211,31,197,31,179,31,119,31,119,30,6,31,124,31,32,31,14,31,14,30,92,31,1,31,183,31,37,31,14,31,23,31,23,30,177,31,22,31,216,31,217,31,217,30,137,31,95,31,95,30,64,31,135,31,70,31,188,31,106,31,106,30,106,29,198,31,73,31,61,31,149,31,149,30,149,29,36,31,36,30,77,31,174,31,163,31,163,30,163,29,16,31,48,31,210,31,242,31,21,31,18,31,147,31,57,31,57,30,186,31,171,31,9,31,232,31,15,31,239,31,239,30,94,31,93,31,57,31,149,31,17,31,28,31,209,31,209,31,37,31,62,31,25,31,143,31,143,30,33,31,192,31,110,31,215,31,170,31,201,31,201,30,253,31,253,30,81,31,246,31,56,31,158,31,132,31,136,31,43,31,116,31,177,31,177,30,235,31,235,30,74,31,200,31,185,31,169,31,68,31,252,31,196,31,196,30,196,29,114,31,114,30,193,31,249,31,143,31,139,31,63,31,236,31,232,31,54,31,247,31,247,30,140,31,69,31,50,31,50,30,50,29,50,28,253,31,253,30,151,31,7,31,164,31,180,31,15,31,26,31,237,31,130,31,131,31,22,31,101,31,38,31,176,31,131,31,131,30,95,31,163,31,115,31,133,31,90,31,90,30,232,31,4,31,101,31,99,31,37,31,213,31,124,31,124,30,124,29,80,31,50,31,215,31,175,31,38,31,51,31,220,31,231,31,177,31,156,31,91,31,8,31,8,30,167,31,232,31,123,31,18,31,217,31,7,31,106,31,32,31,247,31,107,31,26,31,147,31,9,31,111,31,57,31,235,31,235,30,190,31,30,31,129,31,10,31,254,31,100,31,2,31,226,31,226,30,39,31,50,31,250,31,216,31,74,31,1,31,118,31,64,31,142,31,194,31,176,31,11,31,60,31,67,31,25,31,190,31,25,31,51,31,237,31,29,31,48,31,179,31,39,31,28,31,233,31,21,31,45,31,45,30,73,31,73,30,73,29,191,31,191,30,149,31,229,31,184,31,160,31,179,31,7,31,201,31,114,31,203,31,204,31,156,31,199,31,182,31,182,30,140,31,151,31,11,31,41,31,220,31,220,30,103,31,142,31,142,30,218,31,7,31,89,31,89,30,83,31,83,30,80,31,58,31,191,31,191,30,55,31,55,30,205,31,186,31,60,31,255,31,255,30,87,31,87,30,169,31,251,31,90,31,86,31,171,31,171,30,40,31,175,31,20,31,20,30,151,31,114,31,114,30,6,31,246,31,174,31,174,30,213,31,214,31,216,31,164,31,207,31,26,31,61,31,41,31,41,30,41,29,41,28,115,31,115,30,183,31,8,31,8,30,40,31,40,30,40,29,239,31,41,31,45,31,45,30,197,31,148,31,163,31,112,31,14,31,252,31,241,31,86,31,63,31,25,31,141,31,171,31,143,31,94,31,90,31,178,31,225,31,14,31,141,31,160,31,202,31,255,31,82,31,201,31,128,31,143,31,31,31,124,31,193,31,193,30,193,29,29,31,20,31,200,31,200,30,64,31,95,31,99,31,58,31,232,31,232,30,232,29,232,28,158,31,158,30,92,31,88,31,2,31,155,31,23,31,28,31,80,31,57,31,136,31,115,31,115,30,236,31,236,30,195,31,195,30,157,31,8,31,60,31,60,30,229,31,95,31,95,30,178,31,247,31,162,31,142,31,43,31,243,31,175,31,139,31,44,31,101,31,245,31,73,31,153,31,156,31,156,30,156,29,182,31,162,31,219,31,222,31,222,31,217,31,34,31,207,31,207,30,236,31,236,30,236,29,8,31,137,31,134,31,15,31,15,30,47,31,249,31,58,31,250,31,14,31,20,31,20,30,249,31,249,30,247,31,252,31,65,31,65,31,78,31,78,30,98,31,128,31,223,31,117,31,215,31,84,31,110,31,84,31,116,31,174,31,62,31,159,31,159,30,1,31,164,31,164,30,147,31,101,31,195,31,149,31,149,30,149,29,56,31,5,31,39,31,98,31,98,30,98,29,53,31,68,31,133,31,133,30,224,31,127,31,215,31,181,31,33,31,33,30,119,31,96,31,139,31,139,30,182,31,182,30,28,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
