-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 425;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,0,0,200,0,166,0,97,0,250,0,95,0,82,0,0,0,234,0,0,0,165,0,0,0,44,0,83,0,69,0,209,0,154,0,244,0,86,0,0,0,0,0,10,0,138,0,49,0,224,0,0,0,0,0,23,0,0,0,0,0,31,0,64,0,25,0,34,0,18,0,46,0,111,0,201,0,235,0,213,0,72,0,16,0,113,0,0,0,0,0,18,0,14,0,138,0,252,0,34,0,116,0,174,0,254,0,140,0,94,0,0,0,36,0,121,0,142,0,98,0,200,0,0,0,222,0,22,0,79,0,156,0,0,0,167,0,196,0,191,0,166,0,232,0,124,0,87,0,129,0,58,0,117,0,212,0,245,0,60,0,18,0,0,0,178,0,54,0,160,0,0,0,49,0,45,0,0,0,237,0,144,0,136,0,125,0,186,0,199,0,30,0,134,0,118,0,157,0,133,0,122,0,95,0,254,0,46,0,180,0,1,0,244,0,28,0,124,0,196,0,207,0,0,0,127,0,250,0,94,0,201,0,175,0,36,0,150,0,235,0,118,0,47,0,147,0,54,0,0,0,116,0,6,0,14,0,187,0,242,0,63,0,13,0,181,0,192,0,126,0,0,0,100,0,142,0,0,0,88,0,208,0,200,0,187,0,0,0,173,0,65,0,95,0,249,0,241,0,191,0,216,0,192,0,66,0,237,0,250,0,255,0,188,0,233,0,88,0,205,0,0,0,160,0,15,0,81,0,157,0,139,0,248,0,17,0,0,0,0,0,91,0,8,0,90,0,13,0,210,0,34,0,251,0,86,0,0,0,216,0,95,0,202,0,0,0,213,0,0,0,75,0,219,0,0,0,200,0,247,0,94,0,0,0,158,0,39,0,219,0,0,0,225,0,101,0,19,0,193,0,255,0,217,0,140,0,199,0,187,0,237,0,123,0,52,0,149,0,86,0,0,0,135,0,0,0,229,0,0,0,30,0,12,0,154,0,231,0,0,0,133,0,215,0,67,0,33,0,36,0,118,0,211,0,4,0,0,0,0,0,104,0,251,0,51,0,243,0,102,0,160,0,0,0,167,0,190,0,225,0,215,0,118,0,11,0,0,0,166,0,90,0,254,0,163,0,127,0,158,0,173,0,0,0,4,0,213,0,0,0,150,0,65,0,0,0,159,0,186,0,184,0,68,0,92,0,252,0,129,0,184,0,0,0,96,0,0,0,209,0,0,0,144,0,129,0,114,0,10,0,252,0,33,0,0,0,188,0,129,0,159,0,158,0,201,0,229,0,84,0,0,0,28,0,3,0,225,0,122,0,116,0,86,0,105,0,140,0,15,0,169,0,0,0,252,0,123,0,95,0,46,0,7,0,125,0,202,0,122,0,0,0,219,0,27,0,0,0,188,0,110,0,0,0,18,0,0,0,43,0,109,0,63,0,173,0,176,0,183,0,34,0,169,0,29,0,41,0,28,0,0,0,19,0,212,0,51,0,248,0,210,0,215,0,244,0,110,0,0,0,176,0,44,0,0,0,174,0,0,0,19,0,84,0,254,0,0,0,78,0,33,0,0,0,0,0,0,0,104,0,154,0,0,0,0,0,0,0,0,0,228,0,0,0,248,0,210,0,71,0,153,0,112,0,0,0,0,0,22,0,244,0,233,0,45,0,0,0,242,0,132,0,195,0,204,0,16,0,160,0,145,0,115,0,0,0,0,0,89,0,90,0,51,0,0,0,9,0,212,0,151,0,0,0,0,0,19,0,61,0,0,0,251,0,110,0,13,0,169,0,0,0,0,0,0,0,56,0,50,0,0,0,186,0,155,0,0,0,32,0,23,0,157,0,197,0,193,0,0,0,155,0,247,0,147,0,181,0,91,0,17,0,109,0,0,0,237,0,242,0,119,0,0,0,65,0,116,0);
signal scenario_full  : scenario_type := (36,31,36,30,200,31,166,31,97,31,250,31,95,31,82,31,82,30,234,31,234,30,165,31,165,30,44,31,83,31,69,31,209,31,154,31,244,31,86,31,86,30,86,29,10,31,138,31,49,31,224,31,224,30,224,29,23,31,23,30,23,29,31,31,64,31,25,31,34,31,18,31,46,31,111,31,201,31,235,31,213,31,72,31,16,31,113,31,113,30,113,29,18,31,14,31,138,31,252,31,34,31,116,31,174,31,254,31,140,31,94,31,94,30,36,31,121,31,142,31,98,31,200,31,200,30,222,31,22,31,79,31,156,31,156,30,167,31,196,31,191,31,166,31,232,31,124,31,87,31,129,31,58,31,117,31,212,31,245,31,60,31,18,31,18,30,178,31,54,31,160,31,160,30,49,31,45,31,45,30,237,31,144,31,136,31,125,31,186,31,199,31,30,31,134,31,118,31,157,31,133,31,122,31,95,31,254,31,46,31,180,31,1,31,244,31,28,31,124,31,196,31,207,31,207,30,127,31,250,31,94,31,201,31,175,31,36,31,150,31,235,31,118,31,47,31,147,31,54,31,54,30,116,31,6,31,14,31,187,31,242,31,63,31,13,31,181,31,192,31,126,31,126,30,100,31,142,31,142,30,88,31,208,31,200,31,187,31,187,30,173,31,65,31,95,31,249,31,241,31,191,31,216,31,192,31,66,31,237,31,250,31,255,31,188,31,233,31,88,31,205,31,205,30,160,31,15,31,81,31,157,31,139,31,248,31,17,31,17,30,17,29,91,31,8,31,90,31,13,31,210,31,34,31,251,31,86,31,86,30,216,31,95,31,202,31,202,30,213,31,213,30,75,31,219,31,219,30,200,31,247,31,94,31,94,30,158,31,39,31,219,31,219,30,225,31,101,31,19,31,193,31,255,31,217,31,140,31,199,31,187,31,237,31,123,31,52,31,149,31,86,31,86,30,135,31,135,30,229,31,229,30,30,31,12,31,154,31,231,31,231,30,133,31,215,31,67,31,33,31,36,31,118,31,211,31,4,31,4,30,4,29,104,31,251,31,51,31,243,31,102,31,160,31,160,30,167,31,190,31,225,31,215,31,118,31,11,31,11,30,166,31,90,31,254,31,163,31,127,31,158,31,173,31,173,30,4,31,213,31,213,30,150,31,65,31,65,30,159,31,186,31,184,31,68,31,92,31,252,31,129,31,184,31,184,30,96,31,96,30,209,31,209,30,144,31,129,31,114,31,10,31,252,31,33,31,33,30,188,31,129,31,159,31,158,31,201,31,229,31,84,31,84,30,28,31,3,31,225,31,122,31,116,31,86,31,105,31,140,31,15,31,169,31,169,30,252,31,123,31,95,31,46,31,7,31,125,31,202,31,122,31,122,30,219,31,27,31,27,30,188,31,110,31,110,30,18,31,18,30,43,31,109,31,63,31,173,31,176,31,183,31,34,31,169,31,29,31,41,31,28,31,28,30,19,31,212,31,51,31,248,31,210,31,215,31,244,31,110,31,110,30,176,31,44,31,44,30,174,31,174,30,19,31,84,31,254,31,254,30,78,31,33,31,33,30,33,29,33,28,104,31,154,31,154,30,154,29,154,28,154,27,228,31,228,30,248,31,210,31,71,31,153,31,112,31,112,30,112,29,22,31,244,31,233,31,45,31,45,30,242,31,132,31,195,31,204,31,16,31,160,31,145,31,115,31,115,30,115,29,89,31,90,31,51,31,51,30,9,31,212,31,151,31,151,30,151,29,19,31,61,31,61,30,251,31,110,31,13,31,169,31,169,30,169,29,169,28,56,31,50,31,50,30,186,31,155,31,155,30,32,31,23,31,157,31,197,31,193,31,193,30,155,31,247,31,147,31,181,31,91,31,17,31,109,31,109,30,237,31,242,31,119,31,119,30,65,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
