-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_267 is
end project_tb_267;

architecture project_tb_arch_267 of project_tb_267 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 752;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (161,0,229,0,0,0,0,0,110,0,0,0,25,0,0,0,151,0,210,0,0,0,90,0,90,0,64,0,215,0,154,0,0,0,236,0,0,0,42,0,46,0,235,0,4,0,150,0,0,0,0,0,0,0,98,0,88,0,191,0,0,0,237,0,0,0,0,0,190,0,83,0,210,0,150,0,206,0,80,0,212,0,204,0,0,0,0,0,134,0,231,0,0,0,79,0,170,0,59,0,2,0,91,0,36,0,44,0,219,0,233,0,249,0,126,0,180,0,0,0,29,0,1,0,187,0,0,0,228,0,0,0,73,0,204,0,0,0,128,0,130,0,194,0,0,0,2,0,218,0,59,0,178,0,240,0,0,0,205,0,249,0,111,0,145,0,209,0,159,0,60,0,0,0,82,0,186,0,161,0,62,0,42,0,224,0,81,0,117,0,0,0,64,0,251,0,0,0,69,0,0,0,177,0,109,0,81,0,132,0,69,0,171,0,57,0,137,0,0,0,0,0,0,0,0,0,76,0,0,0,230,0,65,0,33,0,0,0,48,0,162,0,129,0,52,0,226,0,0,0,106,0,0,0,224,0,150,0,2,0,48,0,189,0,0,0,58,0,141,0,106,0,23,0,113,0,0,0,165,0,197,0,218,0,0,0,116,0,0,0,66,0,0,0,0,0,205,0,52,0,0,0,177,0,75,0,39,0,0,0,158,0,38,0,0,0,230,0,2,0,173,0,29,0,0,0,74,0,128,0,143,0,0,0,58,0,73,0,0,0,67,0,0,0,53,0,50,0,42,0,20,0,148,0,39,0,6,0,0,0,108,0,153,0,19,0,0,0,92,0,217,0,0,0,164,0,86,0,0,0,33,0,62,0,201,0,143,0,0,0,108,0,78,0,0,0,186,0,57,0,0,0,0,0,210,0,205,0,0,0,28,0,232,0,190,0,0,0,149,0,115,0,35,0,249,0,226,0,171,0,206,0,246,0,90,0,131,0,246,0,184,0,203,0,0,0,0,0,170,0,41,0,183,0,0,0,0,0,0,0,213,0,108,0,193,0,14,0,189,0,191,0,0,0,0,0,0,0,78,0,86,0,134,0,72,0,0,0,166,0,117,0,196,0,99,0,214,0,0,0,81,0,164,0,242,0,146,0,111,0,15,0,224,0,198,0,163,0,0,0,169,0,169,0,218,0,21,0,0,0,155,0,0,0,0,0,227,0,122,0,80,0,95,0,10,0,137,0,0,0,76,0,232,0,0,0,4,0,153,0,107,0,0,0,0,0,185,0,121,0,247,0,141,0,15,0,219,0,0,0,0,0,30,0,102,0,68,0,29,0,109,0,252,0,179,0,240,0,224,0,224,0,1,0,80,0,234,0,80,0,191,0,23,0,165,0,146,0,94,0,207,0,51,0,0,0,27,0,5,0,237,0,168,0,0,0,71,0,200,0,214,0,84,0,33,0,254,0,46,0,0,0,33,0,222,0,233,0,0,0,247,0,227,0,254,0,0,0,143,0,238,0,127,0,37,0,0,0,227,0,147,0,32,0,61,0,132,0,53,0,114,0,54,0,0,0,189,0,240,0,109,0,221,0,141,0,0,0,186,0,0,0,0,0,74,0,1,0,0,0,57,0,152,0,0,0,224,0,144,0,65,0,118,0,0,0,177,0,0,0,0,0,195,0,174,0,186,0,82,0,62,0,62,0,0,0,67,0,0,0,167,0,0,0,130,0,119,0,88,0,125,0,58,0,203,0,169,0,105,0,237,0,5,0,51,0,192,0,218,0,147,0,233,0,0,0,155,0,238,0,133,0,73,0,111,0,0,0,6,0,203,0,76,0,119,0,0,0,0,0,26,0,59,0,0,0,212,0,188,0,59,0,234,0,151,0,70,0,123,0,0,0,45,0,0,0,8,0,0,0,121,0,208,0,37,0,212,0,0,0,0,0,0,0,44,0,186,0,64,0,0,0,146,0,158,0,0,0,0,0,72,0,220,0,19,0,53,0,236,0,0,0,27,0,211,0,134,0,0,0,240,0,168,0,34,0,100,0,20,0,51,0,73,0,0,0,122,0,150,0,103,0,4,0,38,0,113,0,187,0,136,0,187,0,107,0,0,0,12,0,45,0,0,0,108,0,106,0,0,0,135,0,166,0,161,0,162,0,0,0,0,0,203,0,45,0,0,0,122,0,140,0,122,0,218,0,128,0,110,0,69,0,238,0,195,0,244,0,185,0,22,0,31,0,0,0,190,0,0,0,179,0,61,0,112,0,178,0,80,0,130,0,108,0,109,0,0,0,70,0,116,0,172,0,0,0,0,0,174,0,118,0,110,0,0,0,147,0,0,0,98,0,70,0,105,0,241,0,206,0,141,0,198,0,3,0,39,0,215,0,126,0,26,0,139,0,228,0,74,0,125,0,131,0,67,0,183,0,32,0,208,0,128,0,242,0,0,0,77,0,239,0,87,0,58,0,154,0,134,0,0,0,65,0,243,0,0,0,0,0,255,0,0,0,27,0,19,0,214,0,191,0,119,0,170,0,71,0,0,0,47,0,187,0,0,0,232,0,97,0,81,0,211,0,4,0,85,0,0,0,37,0,0,0,77,0,53,0,105,0,36,0,120,0,80,0,94,0,150,0,0,0,83,0,0,0,191,0,0,0,247,0,189,0,113,0,239,0,0,0,246,0,28,0,0,0,191,0,205,0,178,0,0,0,44,0,36,0,63,0,0,0,228,0,0,0,206,0,163,0,83,0,0,0,151,0,247,0,75,0,137,0,0,0,0,0,196,0,194,0,0,0,113,0,0,0,0,0,79,0,78,0,0,0,56,0,204,0,41,0,0,0,153,0,159,0,92,0,32,0,149,0,0,0,86,0,12,0,23,0,59,0,92,0,134,0,59,0,233,0,197,0,35,0,61,0,142,0,119,0,163,0,236,0,16,0,74,0,201,0,184,0,221,0,105,0,45,0,116,0,80,0,25,0,171,0,123,0,0,0,12,0,172,0,139,0,0,0,140,0,0,0,117,0,128,0,0,0,0,0,176,0,127,0,66,0,175,0,37,0,24,0,247,0,0,0,131,0,0,0,234,0,49,0,162,0,234,0,0,0,222,0,212,0,131,0,235,0,1,0,5,0,163,0,0,0,78,0,0,0,21,0,34,0,69,0,23,0,200,0,0,0,0,0,147,0,154,0,93,0,124,0,64,0,224,0,147,0,0,0,227,0,137,0,250,0,58,0,130,0,245,0,55,0,77,0,224,0,69,0,48,0,9,0,218,0,40,0,110,0,20,0,74,0,78,0,44,0,156,0,207,0,210,0,235,0,91,0,191,0,222,0,84,0,40,0,125,0,213,0,20,0,0,0,0,0,105,0,0,0,0,0,202,0);
signal scenario_full  : scenario_type := (161,31,229,31,229,30,229,29,110,31,110,30,25,31,25,30,151,31,210,31,210,30,90,31,90,31,64,31,215,31,154,31,154,30,236,31,236,30,42,31,46,31,235,31,4,31,150,31,150,30,150,29,150,28,98,31,88,31,191,31,191,30,237,31,237,30,237,29,190,31,83,31,210,31,150,31,206,31,80,31,212,31,204,31,204,30,204,29,134,31,231,31,231,30,79,31,170,31,59,31,2,31,91,31,36,31,44,31,219,31,233,31,249,31,126,31,180,31,180,30,29,31,1,31,187,31,187,30,228,31,228,30,73,31,204,31,204,30,128,31,130,31,194,31,194,30,2,31,218,31,59,31,178,31,240,31,240,30,205,31,249,31,111,31,145,31,209,31,159,31,60,31,60,30,82,31,186,31,161,31,62,31,42,31,224,31,81,31,117,31,117,30,64,31,251,31,251,30,69,31,69,30,177,31,109,31,81,31,132,31,69,31,171,31,57,31,137,31,137,30,137,29,137,28,137,27,76,31,76,30,230,31,65,31,33,31,33,30,48,31,162,31,129,31,52,31,226,31,226,30,106,31,106,30,224,31,150,31,2,31,48,31,189,31,189,30,58,31,141,31,106,31,23,31,113,31,113,30,165,31,197,31,218,31,218,30,116,31,116,30,66,31,66,30,66,29,205,31,52,31,52,30,177,31,75,31,39,31,39,30,158,31,38,31,38,30,230,31,2,31,173,31,29,31,29,30,74,31,128,31,143,31,143,30,58,31,73,31,73,30,67,31,67,30,53,31,50,31,42,31,20,31,148,31,39,31,6,31,6,30,108,31,153,31,19,31,19,30,92,31,217,31,217,30,164,31,86,31,86,30,33,31,62,31,201,31,143,31,143,30,108,31,78,31,78,30,186,31,57,31,57,30,57,29,210,31,205,31,205,30,28,31,232,31,190,31,190,30,149,31,115,31,35,31,249,31,226,31,171,31,206,31,246,31,90,31,131,31,246,31,184,31,203,31,203,30,203,29,170,31,41,31,183,31,183,30,183,29,183,28,213,31,108,31,193,31,14,31,189,31,191,31,191,30,191,29,191,28,78,31,86,31,134,31,72,31,72,30,166,31,117,31,196,31,99,31,214,31,214,30,81,31,164,31,242,31,146,31,111,31,15,31,224,31,198,31,163,31,163,30,169,31,169,31,218,31,21,31,21,30,155,31,155,30,155,29,227,31,122,31,80,31,95,31,10,31,137,31,137,30,76,31,232,31,232,30,4,31,153,31,107,31,107,30,107,29,185,31,121,31,247,31,141,31,15,31,219,31,219,30,219,29,30,31,102,31,68,31,29,31,109,31,252,31,179,31,240,31,224,31,224,31,1,31,80,31,234,31,80,31,191,31,23,31,165,31,146,31,94,31,207,31,51,31,51,30,27,31,5,31,237,31,168,31,168,30,71,31,200,31,214,31,84,31,33,31,254,31,46,31,46,30,33,31,222,31,233,31,233,30,247,31,227,31,254,31,254,30,143,31,238,31,127,31,37,31,37,30,227,31,147,31,32,31,61,31,132,31,53,31,114,31,54,31,54,30,189,31,240,31,109,31,221,31,141,31,141,30,186,31,186,30,186,29,74,31,1,31,1,30,57,31,152,31,152,30,224,31,144,31,65,31,118,31,118,30,177,31,177,30,177,29,195,31,174,31,186,31,82,31,62,31,62,31,62,30,67,31,67,30,167,31,167,30,130,31,119,31,88,31,125,31,58,31,203,31,169,31,105,31,237,31,5,31,51,31,192,31,218,31,147,31,233,31,233,30,155,31,238,31,133,31,73,31,111,31,111,30,6,31,203,31,76,31,119,31,119,30,119,29,26,31,59,31,59,30,212,31,188,31,59,31,234,31,151,31,70,31,123,31,123,30,45,31,45,30,8,31,8,30,121,31,208,31,37,31,212,31,212,30,212,29,212,28,44,31,186,31,64,31,64,30,146,31,158,31,158,30,158,29,72,31,220,31,19,31,53,31,236,31,236,30,27,31,211,31,134,31,134,30,240,31,168,31,34,31,100,31,20,31,51,31,73,31,73,30,122,31,150,31,103,31,4,31,38,31,113,31,187,31,136,31,187,31,107,31,107,30,12,31,45,31,45,30,108,31,106,31,106,30,135,31,166,31,161,31,162,31,162,30,162,29,203,31,45,31,45,30,122,31,140,31,122,31,218,31,128,31,110,31,69,31,238,31,195,31,244,31,185,31,22,31,31,31,31,30,190,31,190,30,179,31,61,31,112,31,178,31,80,31,130,31,108,31,109,31,109,30,70,31,116,31,172,31,172,30,172,29,174,31,118,31,110,31,110,30,147,31,147,30,98,31,70,31,105,31,241,31,206,31,141,31,198,31,3,31,39,31,215,31,126,31,26,31,139,31,228,31,74,31,125,31,131,31,67,31,183,31,32,31,208,31,128,31,242,31,242,30,77,31,239,31,87,31,58,31,154,31,134,31,134,30,65,31,243,31,243,30,243,29,255,31,255,30,27,31,19,31,214,31,191,31,119,31,170,31,71,31,71,30,47,31,187,31,187,30,232,31,97,31,81,31,211,31,4,31,85,31,85,30,37,31,37,30,77,31,53,31,105,31,36,31,120,31,80,31,94,31,150,31,150,30,83,31,83,30,191,31,191,30,247,31,189,31,113,31,239,31,239,30,246,31,28,31,28,30,191,31,205,31,178,31,178,30,44,31,36,31,63,31,63,30,228,31,228,30,206,31,163,31,83,31,83,30,151,31,247,31,75,31,137,31,137,30,137,29,196,31,194,31,194,30,113,31,113,30,113,29,79,31,78,31,78,30,56,31,204,31,41,31,41,30,153,31,159,31,92,31,32,31,149,31,149,30,86,31,12,31,23,31,59,31,92,31,134,31,59,31,233,31,197,31,35,31,61,31,142,31,119,31,163,31,236,31,16,31,74,31,201,31,184,31,221,31,105,31,45,31,116,31,80,31,25,31,171,31,123,31,123,30,12,31,172,31,139,31,139,30,140,31,140,30,117,31,128,31,128,30,128,29,176,31,127,31,66,31,175,31,37,31,24,31,247,31,247,30,131,31,131,30,234,31,49,31,162,31,234,31,234,30,222,31,212,31,131,31,235,31,1,31,5,31,163,31,163,30,78,31,78,30,21,31,34,31,69,31,23,31,200,31,200,30,200,29,147,31,154,31,93,31,124,31,64,31,224,31,147,31,147,30,227,31,137,31,250,31,58,31,130,31,245,31,55,31,77,31,224,31,69,31,48,31,9,31,218,31,40,31,110,31,20,31,74,31,78,31,44,31,156,31,207,31,210,31,235,31,91,31,191,31,222,31,84,31,40,31,125,31,213,31,20,31,20,30,20,29,105,31,105,30,105,29,202,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
