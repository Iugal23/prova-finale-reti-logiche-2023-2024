-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_777 is
end project_tb_777;

architecture project_tb_arch_777 of project_tb_777 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 636;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (193,0,74,0,0,0,227,0,254,0,0,0,31,0,0,0,112,0,32,0,18,0,137,0,0,0,45,0,107,0,245,0,41,0,103,0,40,0,74,0,5,0,0,0,0,0,100,0,87,0,102,0,0,0,255,0,0,0,63,0,121,0,211,0,165,0,227,0,0,0,48,0,0,0,3,0,102,0,15,0,243,0,0,0,234,0,139,0,102,0,0,0,136,0,0,0,0,0,0,0,135,0,120,0,28,0,4,0,100,0,0,0,0,0,165,0,11,0,140,0,221,0,188,0,7,0,7,0,141,0,75,0,174,0,0,0,182,0,111,0,42,0,0,0,72,0,166,0,114,0,5,0,242,0,174,0,139,0,92,0,38,0,0,0,141,0,112,0,120,0,0,0,0,0,0,0,0,0,1,0,126,0,120,0,76,0,14,0,0,0,63,0,152,0,0,0,82,0,1,0,82,0,177,0,244,0,162,0,156,0,242,0,0,0,129,0,98,0,4,0,100,0,9,0,90,0,10,0,18,0,199,0,160,0,142,0,0,0,51,0,227,0,54,0,47,0,123,0,0,0,203,0,120,0,48,0,113,0,204,0,170,0,114,0,152,0,0,0,0,0,45,0,80,0,154,0,214,0,0,0,178,0,163,0,20,0,189,0,52,0,155,0,153,0,129,0,0,0,41,0,233,0,151,0,151,0,202,0,169,0,118,0,232,0,0,0,0,0,212,0,0,0,133,0,249,0,152,0,112,0,134,0,120,0,0,0,236,0,223,0,0,0,141,0,0,0,229,0,119,0,0,0,244,0,0,0,0,0,133,0,255,0,165,0,0,0,56,0,250,0,223,0,37,0,190,0,11,0,0,0,39,0,0,0,49,0,191,0,104,0,36,0,151,0,0,0,0,0,233,0,0,0,250,0,29,0,160,0,190,0,92,0,9,0,160,0,14,0,0,0,171,0,137,0,38,0,82,0,76,0,198,0,76,0,201,0,225,0,39,0,206,0,104,0,22,0,9,0,239,0,193,0,168,0,221,0,0,0,154,0,0,0,0,0,189,0,0,0,0,0,0,0,172,0,183,0,0,0,105,0,141,0,126,0,53,0,139,0,31,0,47,0,111,0,0,0,36,0,0,0,28,0,251,0,191,0,113,0,0,0,0,0,129,0,0,0,52,0,39,0,1,0,0,0,119,0,0,0,153,0,167,0,69,0,40,0,76,0,151,0,220,0,0,0,245,0,4,0,231,0,0,0,170,0,62,0,205,0,46,0,0,0,37,0,0,0,28,0,0,0,50,0,0,0,178,0,181,0,62,0,119,0,65,0,155,0,247,0,0,0,236,0,0,0,83,0,130,0,243,0,176,0,165,0,208,0,235,0,139,0,11,0,125,0,69,0,0,0,206,0,0,0,0,0,142,0,110,0,36,0,141,0,151,0,239,0,228,0,0,0,234,0,142,0,90,0,0,0,98,0,117,0,168,0,171,0,11,0,236,0,129,0,0,0,0,0,127,0,0,0,38,0,33,0,92,0,0,0,194,0,220,0,248,0,108,0,32,0,231,0,81,0,137,0,82,0,0,0,0,0,0,0,67,0,217,0,0,0,117,0,107,0,61,0,151,0,116,0,254,0,118,0,179,0,104,0,16,0,52,0,209,0,238,0,51,0,208,0,185,0,230,0,159,0,149,0,40,0,133,0,83,0,0,0,118,0,78,0,59,0,28,0,91,0,133,0,143,0,135,0,158,0,212,0,144,0,14,0,91,0,121,0,75,0,0,0,181,0,143,0,145,0,147,0,224,0,215,0,68,0,29,0,19,0,0,0,160,0,107,0,66,0,0,0,0,0,164,0,236,0,64,0,156,0,159,0,176,0,197,0,199,0,123,0,58,0,240,0,18,0,0,0,138,0,115,0,146,0,76,0,0,0,94,0,223,0,0,0,208,0,135,0,169,0,0,0,90,0,68,0,104,0,117,0,136,0,21,0,76,0,50,0,210,0,200,0,189,0,148,0,89,0,196,0,129,0,205,0,146,0,77,0,0,0,154,0,17,0,230,0,213,0,114,0,0,0,0,0,134,0,17,0,0,0,191,0,0,0,77,0,172,0,101,0,254,0,182,0,178,0,217,0,0,0,16,0,48,0,253,0,0,0,255,0,0,0,0,0,147,0,0,0,4,0,169,0,126,0,0,0,23,0,14,0,0,0,46,0,149,0,231,0,34,0,153,0,26,0,209,0,220,0,191,0,238,0,253,0,0,0,129,0,163,0,172,0,126,0,59,0,0,0,159,0,73,0,146,0,20,0,27,0,0,0,180,0,202,0,0,0,192,0,0,0,0,0,197,0,70,0,221,0,241,0,156,0,0,0,33,0,81,0,236,0,48,0,0,0,198,0,43,0,0,0,31,0,224,0,101,0,142,0,239,0,216,0,217,0,74,0,0,0,0,0,0,0,232,0,211,0,110,0,129,0,185,0,198,0,89,0,145,0,103,0,35,0,149,0,0,0,90,0,230,0,0,0,80,0,248,0,101,0,116,0,0,0,236,0,232,0,110,0,76,0,0,0,0,0,121,0,239,0,135,0,5,0,124,0,215,0,31,0,203,0,189,0,9,0,24,0,179,0,142,0,212,0,30,0,203,0,126,0,116,0,221,0,0,0,82,0,57,0,50,0,76,0,36,0,237,0,0,0,215,0,130,0,191,0,137,0,0,0,218,0,166,0,23,0,180,0,174,0,56,0,240,0,0,0,48,0,128,0,79,0,16,0,154,0,102,0,106,0,0,0,64,0,181,0,191,0,54,0,11,0,199,0,108,0,54,0,126,0,74,0,0,0,200,0,21,0,125,0,226,0,181,0,89,0,194,0,179,0);
signal scenario_full  : scenario_type := (193,31,74,31,74,30,227,31,254,31,254,30,31,31,31,30,112,31,32,31,18,31,137,31,137,30,45,31,107,31,245,31,41,31,103,31,40,31,74,31,5,31,5,30,5,29,100,31,87,31,102,31,102,30,255,31,255,30,63,31,121,31,211,31,165,31,227,31,227,30,48,31,48,30,3,31,102,31,15,31,243,31,243,30,234,31,139,31,102,31,102,30,136,31,136,30,136,29,136,28,135,31,120,31,28,31,4,31,100,31,100,30,100,29,165,31,11,31,140,31,221,31,188,31,7,31,7,31,141,31,75,31,174,31,174,30,182,31,111,31,42,31,42,30,72,31,166,31,114,31,5,31,242,31,174,31,139,31,92,31,38,31,38,30,141,31,112,31,120,31,120,30,120,29,120,28,120,27,1,31,126,31,120,31,76,31,14,31,14,30,63,31,152,31,152,30,82,31,1,31,82,31,177,31,244,31,162,31,156,31,242,31,242,30,129,31,98,31,4,31,100,31,9,31,90,31,10,31,18,31,199,31,160,31,142,31,142,30,51,31,227,31,54,31,47,31,123,31,123,30,203,31,120,31,48,31,113,31,204,31,170,31,114,31,152,31,152,30,152,29,45,31,80,31,154,31,214,31,214,30,178,31,163,31,20,31,189,31,52,31,155,31,153,31,129,31,129,30,41,31,233,31,151,31,151,31,202,31,169,31,118,31,232,31,232,30,232,29,212,31,212,30,133,31,249,31,152,31,112,31,134,31,120,31,120,30,236,31,223,31,223,30,141,31,141,30,229,31,119,31,119,30,244,31,244,30,244,29,133,31,255,31,165,31,165,30,56,31,250,31,223,31,37,31,190,31,11,31,11,30,39,31,39,30,49,31,191,31,104,31,36,31,151,31,151,30,151,29,233,31,233,30,250,31,29,31,160,31,190,31,92,31,9,31,160,31,14,31,14,30,171,31,137,31,38,31,82,31,76,31,198,31,76,31,201,31,225,31,39,31,206,31,104,31,22,31,9,31,239,31,193,31,168,31,221,31,221,30,154,31,154,30,154,29,189,31,189,30,189,29,189,28,172,31,183,31,183,30,105,31,141,31,126,31,53,31,139,31,31,31,47,31,111,31,111,30,36,31,36,30,28,31,251,31,191,31,113,31,113,30,113,29,129,31,129,30,52,31,39,31,1,31,1,30,119,31,119,30,153,31,167,31,69,31,40,31,76,31,151,31,220,31,220,30,245,31,4,31,231,31,231,30,170,31,62,31,205,31,46,31,46,30,37,31,37,30,28,31,28,30,50,31,50,30,178,31,181,31,62,31,119,31,65,31,155,31,247,31,247,30,236,31,236,30,83,31,130,31,243,31,176,31,165,31,208,31,235,31,139,31,11,31,125,31,69,31,69,30,206,31,206,30,206,29,142,31,110,31,36,31,141,31,151,31,239,31,228,31,228,30,234,31,142,31,90,31,90,30,98,31,117,31,168,31,171,31,11,31,236,31,129,31,129,30,129,29,127,31,127,30,38,31,33,31,92,31,92,30,194,31,220,31,248,31,108,31,32,31,231,31,81,31,137,31,82,31,82,30,82,29,82,28,67,31,217,31,217,30,117,31,107,31,61,31,151,31,116,31,254,31,118,31,179,31,104,31,16,31,52,31,209,31,238,31,51,31,208,31,185,31,230,31,159,31,149,31,40,31,133,31,83,31,83,30,118,31,78,31,59,31,28,31,91,31,133,31,143,31,135,31,158,31,212,31,144,31,14,31,91,31,121,31,75,31,75,30,181,31,143,31,145,31,147,31,224,31,215,31,68,31,29,31,19,31,19,30,160,31,107,31,66,31,66,30,66,29,164,31,236,31,64,31,156,31,159,31,176,31,197,31,199,31,123,31,58,31,240,31,18,31,18,30,138,31,115,31,146,31,76,31,76,30,94,31,223,31,223,30,208,31,135,31,169,31,169,30,90,31,68,31,104,31,117,31,136,31,21,31,76,31,50,31,210,31,200,31,189,31,148,31,89,31,196,31,129,31,205,31,146,31,77,31,77,30,154,31,17,31,230,31,213,31,114,31,114,30,114,29,134,31,17,31,17,30,191,31,191,30,77,31,172,31,101,31,254,31,182,31,178,31,217,31,217,30,16,31,48,31,253,31,253,30,255,31,255,30,255,29,147,31,147,30,4,31,169,31,126,31,126,30,23,31,14,31,14,30,46,31,149,31,231,31,34,31,153,31,26,31,209,31,220,31,191,31,238,31,253,31,253,30,129,31,163,31,172,31,126,31,59,31,59,30,159,31,73,31,146,31,20,31,27,31,27,30,180,31,202,31,202,30,192,31,192,30,192,29,197,31,70,31,221,31,241,31,156,31,156,30,33,31,81,31,236,31,48,31,48,30,198,31,43,31,43,30,31,31,224,31,101,31,142,31,239,31,216,31,217,31,74,31,74,30,74,29,74,28,232,31,211,31,110,31,129,31,185,31,198,31,89,31,145,31,103,31,35,31,149,31,149,30,90,31,230,31,230,30,80,31,248,31,101,31,116,31,116,30,236,31,232,31,110,31,76,31,76,30,76,29,121,31,239,31,135,31,5,31,124,31,215,31,31,31,203,31,189,31,9,31,24,31,179,31,142,31,212,31,30,31,203,31,126,31,116,31,221,31,221,30,82,31,57,31,50,31,76,31,36,31,237,31,237,30,215,31,130,31,191,31,137,31,137,30,218,31,166,31,23,31,180,31,174,31,56,31,240,31,240,30,48,31,128,31,79,31,16,31,154,31,102,31,106,31,106,30,64,31,181,31,191,31,54,31,11,31,199,31,108,31,54,31,126,31,74,31,74,30,200,31,21,31,125,31,226,31,181,31,89,31,194,31,179,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
