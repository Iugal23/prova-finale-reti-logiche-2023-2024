-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_42 is
end project_tb_42;

architecture project_tb_arch_42 of project_tb_42 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 380;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,189,0,110,0,245,0,66,0,217,0,107,0,163,0,42,0,38,0,0,0,101,0,0,0,0,0,255,0,0,0,28,0,141,0,131,0,139,0,104,0,0,0,110,0,36,0,103,0,0,0,0,0,0,0,204,0,0,0,75,0,0,0,0,0,0,0,237,0,57,0,244,0,155,0,0,0,0,0,103,0,107,0,176,0,39,0,166,0,34,0,215,0,115,0,103,0,18,0,193,0,193,0,39,0,133,0,17,0,182,0,0,0,0,0,147,0,203,0,54,0,85,0,203,0,1,0,187,0,241,0,24,0,32,0,10,0,208,0,0,0,0,0,222,0,46,0,109,0,238,0,7,0,244,0,166,0,0,0,197,0,218,0,13,0,251,0,92,0,29,0,0,0,82,0,128,0,102,0,0,0,94,0,202,0,0,0,73,0,185,0,84,0,0,0,156,0,164,0,1,0,46,0,122,0,0,0,50,0,224,0,19,0,0,0,0,0,28,0,194,0,0,0,0,0,233,0,166,0,240,0,0,0,178,0,0,0,0,0,0,0,183,0,91,0,233,0,0,0,0,0,249,0,208,0,162,0,0,0,208,0,0,0,127,0,0,0,108,0,4,0,216,0,232,0,0,0,114,0,68,0,0,0,148,0,55,0,0,0,97,0,37,0,2,0,157,0,159,0,0,0,203,0,99,0,61,0,0,0,145,0,252,0,0,0,245,0,187,0,241,0,231,0,0,0,132,0,60,0,0,0,140,0,171,0,165,0,1,0,94,0,90,0,41,0,19,0,39,0,0,0,252,0,170,0,149,0,58,0,202,0,161,0,158,0,160,0,253,0,113,0,189,0,169,0,242,0,131,0,195,0,0,0,156,0,188,0,239,0,174,0,0,0,59,0,246,0,115,0,160,0,243,0,223,0,148,0,21,0,237,0,191,0,0,0,60,0,22,0,80,0,170,0,0,0,138,0,220,0,159,0,225,0,180,0,225,0,88,0,253,0,45,0,46,0,111,0,90,0,21,0,0,0,13,0,215,0,179,0,18,0,76,0,32,0,66,0,66,0,0,0,208,0,130,0,0,0,0,0,0,0,65,0,18,0,170,0,102,0,249,0,0,0,82,0,117,0,0,0,54,0,112,0,30,0,198,0,57,0,181,0,55,0,225,0,73,0,204,0,0,0,218,0,104,0,0,0,108,0,31,0,128,0,0,0,242,0,151,0,196,0,0,0,56,0,106,0,148,0,0,0,104,0,242,0,205,0,238,0,116,0,70,0,161,0,123,0,18,0,19,0,202,0,251,0,0,0,0,0,91,0,218,0,116,0,91,0,112,0,246,0,199,0,5,0,0,0,58,0,175,0,98,0,245,0,0,0,117,0,192,0,170,0,0,0,13,0,158,0,57,0,208,0,66,0,32,0,53,0,0,0,240,0,99,0,0,0,0,0,0,0,206,0,178,0,0,0,170,0,115,0,20,0,168,0,186,0,109,0,214,0,118,0,132,0,208,0,154,0,41,0,57,0,58,0,15,0,237,0,125,0,118,0,71,0,0,0,138,0,165,0,29,0,64,0,28,0,148,0,23,0,150,0,101,0,129,0,61,0,44,0,51,0,255,0,2,0,132,0,0,0,33,0,33,0,109,0,96,0,99,0,175,0,49,0,0,0,30,0,84,0,109,0,153,0,0,0,126,0,86,0,84,0,2,0,141,0,250,0);
signal scenario_full  : scenario_type := (1,31,189,31,110,31,245,31,66,31,217,31,107,31,163,31,42,31,38,31,38,30,101,31,101,30,101,29,255,31,255,30,28,31,141,31,131,31,139,31,104,31,104,30,110,31,36,31,103,31,103,30,103,29,103,28,204,31,204,30,75,31,75,30,75,29,75,28,237,31,57,31,244,31,155,31,155,30,155,29,103,31,107,31,176,31,39,31,166,31,34,31,215,31,115,31,103,31,18,31,193,31,193,31,39,31,133,31,17,31,182,31,182,30,182,29,147,31,203,31,54,31,85,31,203,31,1,31,187,31,241,31,24,31,32,31,10,31,208,31,208,30,208,29,222,31,46,31,109,31,238,31,7,31,244,31,166,31,166,30,197,31,218,31,13,31,251,31,92,31,29,31,29,30,82,31,128,31,102,31,102,30,94,31,202,31,202,30,73,31,185,31,84,31,84,30,156,31,164,31,1,31,46,31,122,31,122,30,50,31,224,31,19,31,19,30,19,29,28,31,194,31,194,30,194,29,233,31,166,31,240,31,240,30,178,31,178,30,178,29,178,28,183,31,91,31,233,31,233,30,233,29,249,31,208,31,162,31,162,30,208,31,208,30,127,31,127,30,108,31,4,31,216,31,232,31,232,30,114,31,68,31,68,30,148,31,55,31,55,30,97,31,37,31,2,31,157,31,159,31,159,30,203,31,99,31,61,31,61,30,145,31,252,31,252,30,245,31,187,31,241,31,231,31,231,30,132,31,60,31,60,30,140,31,171,31,165,31,1,31,94,31,90,31,41,31,19,31,39,31,39,30,252,31,170,31,149,31,58,31,202,31,161,31,158,31,160,31,253,31,113,31,189,31,169,31,242,31,131,31,195,31,195,30,156,31,188,31,239,31,174,31,174,30,59,31,246,31,115,31,160,31,243,31,223,31,148,31,21,31,237,31,191,31,191,30,60,31,22,31,80,31,170,31,170,30,138,31,220,31,159,31,225,31,180,31,225,31,88,31,253,31,45,31,46,31,111,31,90,31,21,31,21,30,13,31,215,31,179,31,18,31,76,31,32,31,66,31,66,31,66,30,208,31,130,31,130,30,130,29,130,28,65,31,18,31,170,31,102,31,249,31,249,30,82,31,117,31,117,30,54,31,112,31,30,31,198,31,57,31,181,31,55,31,225,31,73,31,204,31,204,30,218,31,104,31,104,30,108,31,31,31,128,31,128,30,242,31,151,31,196,31,196,30,56,31,106,31,148,31,148,30,104,31,242,31,205,31,238,31,116,31,70,31,161,31,123,31,18,31,19,31,202,31,251,31,251,30,251,29,91,31,218,31,116,31,91,31,112,31,246,31,199,31,5,31,5,30,58,31,175,31,98,31,245,31,245,30,117,31,192,31,170,31,170,30,13,31,158,31,57,31,208,31,66,31,32,31,53,31,53,30,240,31,99,31,99,30,99,29,99,28,206,31,178,31,178,30,170,31,115,31,20,31,168,31,186,31,109,31,214,31,118,31,132,31,208,31,154,31,41,31,57,31,58,31,15,31,237,31,125,31,118,31,71,31,71,30,138,31,165,31,29,31,64,31,28,31,148,31,23,31,150,31,101,31,129,31,61,31,44,31,51,31,255,31,2,31,132,31,132,30,33,31,33,31,109,31,96,31,99,31,175,31,49,31,49,30,30,31,84,31,109,31,153,31,153,30,126,31,86,31,84,31,2,31,141,31,250,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
