-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_178 is
end project_tb_178;

architecture project_tb_arch_178 of project_tb_178 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 203;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,55,0,0,0,72,0,222,0,0,0,19,0,206,0,228,0,245,0,119,0,123,0,90,0,72,0,220,0,199,0,0,0,152,0,79,0,137,0,75,0,0,0,20,0,100,0,0,0,63,0,237,0,16,0,31,0,0,0,112,0,23,0,157,0,41,0,197,0,152,0,0,0,107,0,173,0,19,0,91,0,41,0,239,0,252,0,0,0,239,0,53,0,57,0,78,0,196,0,0,0,160,0,2,0,65,0,1,0,31,0,0,0,31,0,74,0,191,0,0,0,227,0,126,0,51,0,89,0,192,0,85,0,19,0,7,0,0,0,61,0,0,0,64,0,79,0,0,0,87,0,132,0,121,0,0,0,145,0,119,0,124,0,62,0,109,0,135,0,128,0,135,0,248,0,15,0,15,0,3,0,0,0,79,0,0,0,129,0,27,0,227,0,23,0,26,0,0,0,1,0,0,0,84,0,219,0,0,0,167,0,0,0,0,0,0,0,117,0,136,0,0,0,232,0,0,0,0,0,0,0,94,0,84,0,38,0,98,0,224,0,101,0,122,0,231,0,8,0,0,0,229,0,0,0,62,0,99,0,58,0,22,0,183,0,227,0,250,0,217,0,200,0,155,0,109,0,48,0,0,0,100,0,102,0,206,0,111,0,35,0,108,0,247,0,204,0,214,0,198,0,63,0,232,0,173,0,79,0,170,0,158,0,48,0,0,0,0,0,112,0,0,0,18,0,0,0,23,0,253,0,114,0,121,0,19,0,213,0,0,0,229,0,46,0,154,0,217,0,207,0,204,0,161,0,157,0,134,0,0,0,0,0,0,0,216,0,93,0,234,0,21,0,99,0,46,0,0,0,27,0,203,0,167,0,65,0,55,0,204,0,240,0,203,0,83,0,226,0,160,0,233,0,215,0);
signal scenario_full  : scenario_type := (0,0,55,31,55,30,72,31,222,31,222,30,19,31,206,31,228,31,245,31,119,31,123,31,90,31,72,31,220,31,199,31,199,30,152,31,79,31,137,31,75,31,75,30,20,31,100,31,100,30,63,31,237,31,16,31,31,31,31,30,112,31,23,31,157,31,41,31,197,31,152,31,152,30,107,31,173,31,19,31,91,31,41,31,239,31,252,31,252,30,239,31,53,31,57,31,78,31,196,31,196,30,160,31,2,31,65,31,1,31,31,31,31,30,31,31,74,31,191,31,191,30,227,31,126,31,51,31,89,31,192,31,85,31,19,31,7,31,7,30,61,31,61,30,64,31,79,31,79,30,87,31,132,31,121,31,121,30,145,31,119,31,124,31,62,31,109,31,135,31,128,31,135,31,248,31,15,31,15,31,3,31,3,30,79,31,79,30,129,31,27,31,227,31,23,31,26,31,26,30,1,31,1,30,84,31,219,31,219,30,167,31,167,30,167,29,167,28,117,31,136,31,136,30,232,31,232,30,232,29,232,28,94,31,84,31,38,31,98,31,224,31,101,31,122,31,231,31,8,31,8,30,229,31,229,30,62,31,99,31,58,31,22,31,183,31,227,31,250,31,217,31,200,31,155,31,109,31,48,31,48,30,100,31,102,31,206,31,111,31,35,31,108,31,247,31,204,31,214,31,198,31,63,31,232,31,173,31,79,31,170,31,158,31,48,31,48,30,48,29,112,31,112,30,18,31,18,30,23,31,253,31,114,31,121,31,19,31,213,31,213,30,229,31,46,31,154,31,217,31,207,31,204,31,161,31,157,31,134,31,134,30,134,29,134,28,216,31,93,31,234,31,21,31,99,31,46,31,46,30,27,31,203,31,167,31,65,31,55,31,204,31,240,31,203,31,83,31,226,31,160,31,233,31,215,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
