-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_116 is
end project_tb_116;

architecture project_tb_arch_116 of project_tb_116 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 341;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (81,0,0,0,209,0,208,0,255,0,157,0,141,0,0,0,206,0,0,0,141,0,172,0,188,0,238,0,37,0,222,0,212,0,11,0,123,0,207,0,67,0,72,0,187,0,0,0,140,0,239,0,113,0,217,0,0,0,77,0,53,0,37,0,229,0,142,0,0,0,69,0,31,0,77,0,0,0,18,0,48,0,56,0,33,0,231,0,192,0,181,0,0,0,125,0,48,0,162,0,237,0,77,0,134,0,100,0,137,0,223,0,174,0,148,0,60,0,158,0,98,0,152,0,175,0,184,0,194,0,239,0,202,0,0,0,214,0,0,0,237,0,220,0,0,0,253,0,43,0,111,0,101,0,0,0,45,0,0,0,22,0,122,0,211,0,1,0,0,0,44,0,15,0,221,0,179,0,202,0,83,0,218,0,0,0,157,0,189,0,88,0,245,0,107,0,60,0,52,0,4,0,111,0,193,0,169,0,51,0,134,0,49,0,10,0,150,0,226,0,94,0,70,0,147,0,60,0,29,0,196,0,8,0,63,0,0,0,149,0,129,0,71,0,128,0,0,0,69,0,163,0,181,0,0,0,120,0,203,0,0,0,0,0,159,0,121,0,216,0,35,0,0,0,0,0,75,0,126,0,0,0,166,0,0,0,219,0,240,0,0,0,0,0,42,0,211,0,183,0,210,0,183,0,114,0,244,0,35,0,33,0,14,0,0,0,0,0,183,0,0,0,254,0,78,0,163,0,244,0,17,0,237,0,21,0,183,0,0,0,23,0,0,0,227,0,0,0,152,0,0,0,0,0,95,0,180,0,115,0,0,0,220,0,0,0,213,0,0,0,0,0,92,0,58,0,227,0,0,0,49,0,0,0,52,0,204,0,74,0,230,0,52,0,0,0,30,0,0,0,220,0,11,0,16,0,0,0,22,0,48,0,230,0,142,0,0,0,207,0,0,0,187,0,149,0,152,0,213,0,77,0,28,0,0,0,0,0,189,0,0,0,10,0,89,0,214,0,111,0,13,0,0,0,176,0,172,0,206,0,125,0,35,0,0,0,56,0,120,0,168,0,239,0,207,0,0,0,65,0,38,0,216,0,114,0,199,0,0,0,0,0,0,0,187,0,214,0,35,0,0,0,77,0,118,0,126,0,134,0,11,0,74,0,127,0,40,0,200,0,26,0,0,0,136,0,215,0,0,0,223,0,51,0,241,0,44,0,151,0,172,0,70,0,193,0,102,0,235,0,238,0,21,0,0,0,245,0,165,0,38,0,155,0,214,0,215,0,6,0,211,0,15,0,185,0,154,0,242,0,198,0,0,0,192,0,206,0,47,0,79,0,144,0,69,0,49,0,0,0,132,0,103,0,58,0,166,0,31,0,217,0,152,0,184,0,223,0,211,0,99,0,17,0,210,0,119,0,225,0,148,0,29,0,230,0,182,0,70,0,70,0,193,0,245,0,0,0,200,0,109,0,78,0,4,0,98,0,5,0,0,0,50,0,86,0,120,0,24,0,52,0,6,0,125,0,227,0,86,0,0,0);
signal scenario_full  : scenario_type := (81,31,81,30,209,31,208,31,255,31,157,31,141,31,141,30,206,31,206,30,141,31,172,31,188,31,238,31,37,31,222,31,212,31,11,31,123,31,207,31,67,31,72,31,187,31,187,30,140,31,239,31,113,31,217,31,217,30,77,31,53,31,37,31,229,31,142,31,142,30,69,31,31,31,77,31,77,30,18,31,48,31,56,31,33,31,231,31,192,31,181,31,181,30,125,31,48,31,162,31,237,31,77,31,134,31,100,31,137,31,223,31,174,31,148,31,60,31,158,31,98,31,152,31,175,31,184,31,194,31,239,31,202,31,202,30,214,31,214,30,237,31,220,31,220,30,253,31,43,31,111,31,101,31,101,30,45,31,45,30,22,31,122,31,211,31,1,31,1,30,44,31,15,31,221,31,179,31,202,31,83,31,218,31,218,30,157,31,189,31,88,31,245,31,107,31,60,31,52,31,4,31,111,31,193,31,169,31,51,31,134,31,49,31,10,31,150,31,226,31,94,31,70,31,147,31,60,31,29,31,196,31,8,31,63,31,63,30,149,31,129,31,71,31,128,31,128,30,69,31,163,31,181,31,181,30,120,31,203,31,203,30,203,29,159,31,121,31,216,31,35,31,35,30,35,29,75,31,126,31,126,30,166,31,166,30,219,31,240,31,240,30,240,29,42,31,211,31,183,31,210,31,183,31,114,31,244,31,35,31,33,31,14,31,14,30,14,29,183,31,183,30,254,31,78,31,163,31,244,31,17,31,237,31,21,31,183,31,183,30,23,31,23,30,227,31,227,30,152,31,152,30,152,29,95,31,180,31,115,31,115,30,220,31,220,30,213,31,213,30,213,29,92,31,58,31,227,31,227,30,49,31,49,30,52,31,204,31,74,31,230,31,52,31,52,30,30,31,30,30,220,31,11,31,16,31,16,30,22,31,48,31,230,31,142,31,142,30,207,31,207,30,187,31,149,31,152,31,213,31,77,31,28,31,28,30,28,29,189,31,189,30,10,31,89,31,214,31,111,31,13,31,13,30,176,31,172,31,206,31,125,31,35,31,35,30,56,31,120,31,168,31,239,31,207,31,207,30,65,31,38,31,216,31,114,31,199,31,199,30,199,29,199,28,187,31,214,31,35,31,35,30,77,31,118,31,126,31,134,31,11,31,74,31,127,31,40,31,200,31,26,31,26,30,136,31,215,31,215,30,223,31,51,31,241,31,44,31,151,31,172,31,70,31,193,31,102,31,235,31,238,31,21,31,21,30,245,31,165,31,38,31,155,31,214,31,215,31,6,31,211,31,15,31,185,31,154,31,242,31,198,31,198,30,192,31,206,31,47,31,79,31,144,31,69,31,49,31,49,30,132,31,103,31,58,31,166,31,31,31,217,31,152,31,184,31,223,31,211,31,99,31,17,31,210,31,119,31,225,31,148,31,29,31,230,31,182,31,70,31,70,31,193,31,245,31,245,30,200,31,109,31,78,31,4,31,98,31,5,31,5,30,50,31,86,31,120,31,24,31,52,31,6,31,125,31,227,31,86,31,86,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
