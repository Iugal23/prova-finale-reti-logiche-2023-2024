-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 758;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (234,0,179,0,31,0,188,0,146,0,2,0,108,0,0,0,64,0,201,0,96,0,0,0,112,0,48,0,218,0,54,0,77,0,99,0,35,0,0,0,66,0,0,0,19,0,63,0,0,0,44,0,218,0,191,0,103,0,39,0,128,0,0,0,141,0,136,0,135,0,0,0,80,0,40,0,218,0,85,0,126,0,0,0,84,0,131,0,0,0,0,0,215,0,231,0,16,0,226,0,0,0,73,0,0,0,176,0,232,0,173,0,0,0,186,0,125,0,147,0,80,0,255,0,33,0,197,0,33,0,0,0,0,0,0,0,200,0,0,0,0,0,151,0,21,0,190,0,0,0,68,0,171,0,177,0,6,0,250,0,72,0,224,0,210,0,43,0,157,0,153,0,56,0,51,0,240,0,59,0,220,0,13,0,162,0,230,0,41,0,82,0,112,0,1,0,41,0,251,0,64,0,0,0,18,0,23,0,22,0,137,0,123,0,118,0,206,0,42,0,132,0,146,0,53,0,0,0,184,0,0,0,109,0,184,0,6,0,0,0,51,0,10,0,168,0,245,0,202,0,254,0,45,0,133,0,76,0,233,0,174,0,0,0,0,0,195,0,0,0,188,0,39,0,215,0,109,0,130,0,0,0,0,0,36,0,204,0,51,0,22,0,134,0,0,0,123,0,0,0,118,0,134,0,203,0,12,0,217,0,138,0,232,0,91,0,235,0,203,0,210,0,124,0,167,0,166,0,53,0,222,0,13,0,0,0,255,0,182,0,42,0,0,0,0,0,207,0,0,0,101,0,145,0,0,0,170,0,48,0,76,0,119,0,0,0,177,0,62,0,0,0,227,0,42,0,43,0,123,0,0,0,91,0,0,0,170,0,243,0,114,0,0,0,77,0,0,0,0,0,215,0,93,0,133,0,0,0,156,0,190,0,0,0,193,0,107,0,114,0,161,0,234,0,48,0,0,0,7,0,236,0,20,0,255,0,0,0,54,0,157,0,0,0,175,0,41,0,112,0,186,0,152,0,120,0,202,0,150,0,21,0,203,0,175,0,254,0,0,0,243,0,238,0,63,0,0,0,0,0,3,0,11,0,190,0,0,0,161,0,150,0,235,0,0,0,0,0,239,0,215,0,0,0,84,0,217,0,167,0,187,0,237,0,19,0,146,0,0,0,167,0,99,0,0,0,50,0,42,0,65,0,6,0,37,0,143,0,93,0,30,0,5,0,204,0,223,0,131,0,83,0,51,0,0,0,223,0,0,0,0,0,155,0,222,0,58,0,0,0,174,0,61,0,57,0,186,0,125,0,1,0,173,0,19,0,60,0,163,0,0,0,112,0,188,0,240,0,235,0,0,0,221,0,0,0,0,0,0,0,227,0,0,0,150,0,40,0,221,0,144,0,2,0,76,0,245,0,0,0,0,0,170,0,138,0,184,0,78,0,4,0,135,0,239,0,100,0,253,0,167,0,139,0,1,0,118,0,104,0,216,0,248,0,87,0,102,0,191,0,0,0,181,0,235,0,173,0,207,0,170,0,248,0,183,0,0,0,140,0,116,0,204,0,71,0,45,0,13,0,112,0,66,0,61,0,180,0,135,0,182,0,106,0,121,0,208,0,124,0,0,0,0,0,137,0,127,0,179,0,115,0,122,0,0,0,249,0,0,0,40,0,138,0,118,0,235,0,65,0,196,0,80,0,75,0,142,0,136,0,0,0,88,0,181,0,174,0,48,0,105,0,195,0,0,0,0,0,68,0,133,0,189,0,0,0,154,0,244,0,0,0,189,0,95,0,52,0,0,0,158,0,117,0,144,0,242,0,57,0,0,0,51,0,145,0,157,0,56,0,253,0,198,0,197,0,99,0,86,0,191,0,46,0,249,0,81,0,113,0,28,0,0,0,232,0,0,0,54,0,91,0,0,0,186,0,74,0,0,0,242,0,0,0,124,0,30,0,157,0,0,0,168,0,214,0,193,0,0,0,218,0,33,0,203,0,0,0,235,0,132,0,181,0,163,0,211,0,16,0,162,0,0,0,52,0,234,0,80,0,0,0,0,0,102,0,0,0,127,0,0,0,0,0,225,0,24,0,213,0,106,0,0,0,247,0,113,0,204,0,253,0,184,0,238,0,25,0,42,0,0,0,0,0,154,0,172,0,215,0,24,0,221,0,0,0,233,0,218,0,168,0,229,0,188,0,0,0,51,0,152,0,141,0,89,0,232,0,86,0,124,0,103,0,72,0,244,0,226,0,0,0,137,0,0,0,194,0,123,0,110,0,86,0,139,0,12,0,80,0,131,0,84,0,175,0,133,0,0,0,0,0,175,0,37,0,19,0,108,0,64,0,117,0,204,0,46,0,12,0,114,0,0,0,237,0,179,0,0,0,123,0,74,0,221,0,0,0,0,0,179,0,212,0,120,0,0,0,153,0,73,0,162,0,2,0,44,0,143,0,254,0,212,0,229,0,254,0,145,0,224,0,212,0,60,0,0,0,52,0,93,0,102,0,241,0,168,0,89,0,118,0,11,0,3,0,0,0,150,0,150,0,71,0,179,0,0,0,62,0,0,0,201,0,245,0,228,0,55,0,237,0,66,0,162,0,251,0,12,0,58,0,100,0,100,0,56,0,0,0,89,0,0,0,172,0,70,0,177,0,66,0,0,0,188,0,0,0,221,0,87,0,167,0,132,0,135,0,71,0,250,0,205,0,239,0,2,0,0,0,19,0,73,0,99,0,31,0,103,0,188,0,145,0,183,0,0,0,154,0,193,0,144,0,0,0,6,0,167,0,0,0,182,0,230,0,0,0,213,0,241,0,173,0,160,0,177,0,110,0,0,0,139,0,82,0,194,0,23,0,151,0,0,0,81,0,138,0,76,0,206,0,167,0,152,0,0,0,53,0,251,0,193,0,246,0,82,0,50,0,14,0,0,0,0,0,190,0,76,0,237,0,250,0,0,0,218,0,235,0,140,0,102,0,179,0,232,0,0,0,215,0,0,0,12,0,112,0,0,0,0,0,131,0,57,0,87,0,0,0,57,0,220,0,0,0,0,0,52,0,10,0,31,0,159,0,171,0,237,0,19,0,2,0,85,0,180,0,235,0,103,0,122,0,102,0,48,0,17,0,175,0,141,0,84,0,0,0,110,0,195,0,38,0,210,0,141,0,97,0,0,0,88,0,113,0,121,0,0,0,201,0,8,0,0,0,0,0,213,0,0,0,65,0,56,0,241,0,0,0,0,0,177,0,169,0,2,0,232,0,247,0,14,0,148,0,103,0,0,0,192,0,88,0,14,0,237,0,237,0,0,0,180,0,102,0,236,0,0,0,46,0,188,0,47,0,154,0,211,0,220,0,173,0,114,0,169,0,85,0,176,0,90,0,25,0,135,0,145,0,78,0,7,0,244,0);
signal scenario_full  : scenario_type := (234,31,179,31,31,31,188,31,146,31,2,31,108,31,108,30,64,31,201,31,96,31,96,30,112,31,48,31,218,31,54,31,77,31,99,31,35,31,35,30,66,31,66,30,19,31,63,31,63,30,44,31,218,31,191,31,103,31,39,31,128,31,128,30,141,31,136,31,135,31,135,30,80,31,40,31,218,31,85,31,126,31,126,30,84,31,131,31,131,30,131,29,215,31,231,31,16,31,226,31,226,30,73,31,73,30,176,31,232,31,173,31,173,30,186,31,125,31,147,31,80,31,255,31,33,31,197,31,33,31,33,30,33,29,33,28,200,31,200,30,200,29,151,31,21,31,190,31,190,30,68,31,171,31,177,31,6,31,250,31,72,31,224,31,210,31,43,31,157,31,153,31,56,31,51,31,240,31,59,31,220,31,13,31,162,31,230,31,41,31,82,31,112,31,1,31,41,31,251,31,64,31,64,30,18,31,23,31,22,31,137,31,123,31,118,31,206,31,42,31,132,31,146,31,53,31,53,30,184,31,184,30,109,31,184,31,6,31,6,30,51,31,10,31,168,31,245,31,202,31,254,31,45,31,133,31,76,31,233,31,174,31,174,30,174,29,195,31,195,30,188,31,39,31,215,31,109,31,130,31,130,30,130,29,36,31,204,31,51,31,22,31,134,31,134,30,123,31,123,30,118,31,134,31,203,31,12,31,217,31,138,31,232,31,91,31,235,31,203,31,210,31,124,31,167,31,166,31,53,31,222,31,13,31,13,30,255,31,182,31,42,31,42,30,42,29,207,31,207,30,101,31,145,31,145,30,170,31,48,31,76,31,119,31,119,30,177,31,62,31,62,30,227,31,42,31,43,31,123,31,123,30,91,31,91,30,170,31,243,31,114,31,114,30,77,31,77,30,77,29,215,31,93,31,133,31,133,30,156,31,190,31,190,30,193,31,107,31,114,31,161,31,234,31,48,31,48,30,7,31,236,31,20,31,255,31,255,30,54,31,157,31,157,30,175,31,41,31,112,31,186,31,152,31,120,31,202,31,150,31,21,31,203,31,175,31,254,31,254,30,243,31,238,31,63,31,63,30,63,29,3,31,11,31,190,31,190,30,161,31,150,31,235,31,235,30,235,29,239,31,215,31,215,30,84,31,217,31,167,31,187,31,237,31,19,31,146,31,146,30,167,31,99,31,99,30,50,31,42,31,65,31,6,31,37,31,143,31,93,31,30,31,5,31,204,31,223,31,131,31,83,31,51,31,51,30,223,31,223,30,223,29,155,31,222,31,58,31,58,30,174,31,61,31,57,31,186,31,125,31,1,31,173,31,19,31,60,31,163,31,163,30,112,31,188,31,240,31,235,31,235,30,221,31,221,30,221,29,221,28,227,31,227,30,150,31,40,31,221,31,144,31,2,31,76,31,245,31,245,30,245,29,170,31,138,31,184,31,78,31,4,31,135,31,239,31,100,31,253,31,167,31,139,31,1,31,118,31,104,31,216,31,248,31,87,31,102,31,191,31,191,30,181,31,235,31,173,31,207,31,170,31,248,31,183,31,183,30,140,31,116,31,204,31,71,31,45,31,13,31,112,31,66,31,61,31,180,31,135,31,182,31,106,31,121,31,208,31,124,31,124,30,124,29,137,31,127,31,179,31,115,31,122,31,122,30,249,31,249,30,40,31,138,31,118,31,235,31,65,31,196,31,80,31,75,31,142,31,136,31,136,30,88,31,181,31,174,31,48,31,105,31,195,31,195,30,195,29,68,31,133,31,189,31,189,30,154,31,244,31,244,30,189,31,95,31,52,31,52,30,158,31,117,31,144,31,242,31,57,31,57,30,51,31,145,31,157,31,56,31,253,31,198,31,197,31,99,31,86,31,191,31,46,31,249,31,81,31,113,31,28,31,28,30,232,31,232,30,54,31,91,31,91,30,186,31,74,31,74,30,242,31,242,30,124,31,30,31,157,31,157,30,168,31,214,31,193,31,193,30,218,31,33,31,203,31,203,30,235,31,132,31,181,31,163,31,211,31,16,31,162,31,162,30,52,31,234,31,80,31,80,30,80,29,102,31,102,30,127,31,127,30,127,29,225,31,24,31,213,31,106,31,106,30,247,31,113,31,204,31,253,31,184,31,238,31,25,31,42,31,42,30,42,29,154,31,172,31,215,31,24,31,221,31,221,30,233,31,218,31,168,31,229,31,188,31,188,30,51,31,152,31,141,31,89,31,232,31,86,31,124,31,103,31,72,31,244,31,226,31,226,30,137,31,137,30,194,31,123,31,110,31,86,31,139,31,12,31,80,31,131,31,84,31,175,31,133,31,133,30,133,29,175,31,37,31,19,31,108,31,64,31,117,31,204,31,46,31,12,31,114,31,114,30,237,31,179,31,179,30,123,31,74,31,221,31,221,30,221,29,179,31,212,31,120,31,120,30,153,31,73,31,162,31,2,31,44,31,143,31,254,31,212,31,229,31,254,31,145,31,224,31,212,31,60,31,60,30,52,31,93,31,102,31,241,31,168,31,89,31,118,31,11,31,3,31,3,30,150,31,150,31,71,31,179,31,179,30,62,31,62,30,201,31,245,31,228,31,55,31,237,31,66,31,162,31,251,31,12,31,58,31,100,31,100,31,56,31,56,30,89,31,89,30,172,31,70,31,177,31,66,31,66,30,188,31,188,30,221,31,87,31,167,31,132,31,135,31,71,31,250,31,205,31,239,31,2,31,2,30,19,31,73,31,99,31,31,31,103,31,188,31,145,31,183,31,183,30,154,31,193,31,144,31,144,30,6,31,167,31,167,30,182,31,230,31,230,30,213,31,241,31,173,31,160,31,177,31,110,31,110,30,139,31,82,31,194,31,23,31,151,31,151,30,81,31,138,31,76,31,206,31,167,31,152,31,152,30,53,31,251,31,193,31,246,31,82,31,50,31,14,31,14,30,14,29,190,31,76,31,237,31,250,31,250,30,218,31,235,31,140,31,102,31,179,31,232,31,232,30,215,31,215,30,12,31,112,31,112,30,112,29,131,31,57,31,87,31,87,30,57,31,220,31,220,30,220,29,52,31,10,31,31,31,159,31,171,31,237,31,19,31,2,31,85,31,180,31,235,31,103,31,122,31,102,31,48,31,17,31,175,31,141,31,84,31,84,30,110,31,195,31,38,31,210,31,141,31,97,31,97,30,88,31,113,31,121,31,121,30,201,31,8,31,8,30,8,29,213,31,213,30,65,31,56,31,241,31,241,30,241,29,177,31,169,31,2,31,232,31,247,31,14,31,148,31,103,31,103,30,192,31,88,31,14,31,237,31,237,31,237,30,180,31,102,31,236,31,236,30,46,31,188,31,47,31,154,31,211,31,220,31,173,31,114,31,169,31,85,31,176,31,90,31,25,31,135,31,145,31,78,31,7,31,244,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
