-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 674;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,0,0,0,0,0,0,101,0,202,0,89,0,0,0,0,0,0,0,154,0,231,0,211,0,223,0,58,0,132,0,107,0,87,0,42,0,81,0,0,0,118,0,135,0,193,0,222,0,226,0,249,0,20,0,132,0,84,0,0,0,180,0,84,0,158,0,114,0,35,0,0,0,42,0,181,0,119,0,0,0,35,0,158,0,0,0,0,0,0,0,145,0,13,0,251,0,98,0,250,0,225,0,0,0,26,0,0,0,75,0,29,0,65,0,110,0,236,0,103,0,197,0,49,0,79,0,22,0,0,0,0,0,139,0,159,0,219,0,176,0,0,0,13,0,77,0,0,0,216,0,62,0,2,0,0,0,97,0,163,0,0,0,5,0,54,0,41,0,0,0,9,0,96,0,200,0,215,0,227,0,86,0,225,0,241,0,208,0,37,0,49,0,228,0,156,0,11,0,222,0,64,0,197,0,0,0,36,0,171,0,86,0,59,0,200,0,229,0,112,0,79,0,101,0,229,0,25,0,184,0,0,0,200,0,42,0,161,0,22,0,115,0,0,0,180,0,16,0,72,0,113,0,74,0,171,0,5,0,66,0,0,0,60,0,159,0,248,0,212,0,69,0,119,0,50,0,239,0,128,0,190,0,94,0,118,0,206,0,119,0,22,0,0,0,12,0,4,0,236,0,221,0,75,0,69,0,0,0,0,0,244,0,156,0,0,0,128,0,74,0,0,0,138,0,134,0,72,0,0,0,82,0,90,0,113,0,231,0,0,0,49,0,177,0,55,0,14,0,150,0,70,0,111,0,158,0,37,0,215,0,9,0,43,0,154,0,229,0,43,0,162,0,218,0,72,0,160,0,0,0,186,0,126,0,59,0,145,0,137,0,71,0,232,0,226,0,174,0,35,0,192,0,0,0,155,0,38,0,247,0,160,0,1,0,0,0,76,0,33,0,247,0,148,0,113,0,31,0,140,0,21,0,82,0,0,0,14,0,230,0,7,0,28,0,99,0,54,0,1,0,146,0,160,0,120,0,0,0,0,0,0,0,9,0,32,0,176,0,0,0,79,0,139,0,32,0,4,0,0,0,184,0,53,0,190,0,150,0,213,0,26,0,76,0,108,0,85,0,254,0,0,0,64,0,201,0,132,0,73,0,153,0,109,0,200,0,168,0,0,0,20,0,0,0,113,0,212,0,145,0,241,0,72,0,170,0,150,0,144,0,130,0,10,0,25,0,0,0,167,0,156,0,225,0,0,0,208,0,38,0,0,0,0,0,140,0,145,0,238,0,74,0,126,0,246,0,18,0,109,0,0,0,7,0,98,0,43,0,7,0,172,0,45,0,28,0,102,0,74,0,14,0,133,0,13,0,139,0,0,0,138,0,0,0,202,0,150,0,177,0,193,0,229,0,87,0,18,0,49,0,215,0,50,0,241,0,183,0,0,0,167,0,22,0,227,0,97,0,0,0,189,0,130,0,0,0,133,0,196,0,0,0,174,0,231,0,166,0,226,0,30,0,245,0,184,0,0,0,102,0,0,0,65,0,234,0,241,0,0,0,154,0,0,0,241,0,216,0,219,0,46,0,125,0,133,0,173,0,180,0,0,0,103,0,94,0,235,0,47,0,62,0,163,0,132,0,243,0,0,0,239,0,204,0,243,0,116,0,0,0,0,0,42,0,192,0,7,0,202,0,50,0,0,0,235,0,66,0,194,0,0,0,245,0,90,0,100,0,0,0,0,0,105,0,79,0,217,0,153,0,151,0,177,0,231,0,25,0,59,0,166,0,129,0,134,0,10,0,65,0,0,0,186,0,199,0,100,0,0,0,69,0,135,0,157,0,49,0,181,0,48,0,0,0,38,0,253,0,107,0,56,0,97,0,120,0,13,0,74,0,154,0,119,0,211,0,45,0,56,0,0,0,43,0,9,0,188,0,0,0,2,0,0,0,128,0,28,0,0,0,83,0,131,0,211,0,140,0,103,0,216,0,24,0,0,0,183,0,173,0,108,0,0,0,204,0,87,0,167,0,0,0,0,0,63,0,246,0,7,0,195,0,200,0,156,0,0,0,204,0,230,0,53,0,127,0,148,0,227,0,251,0,253,0,31,0,22,0,114,0,0,0,98,0,85,0,187,0,105,0,0,0,28,0,103,0,204,0,0,0,101,0,0,0,53,0,221,0,145,0,0,0,231,0,247,0,53,0,69,0,171,0,0,0,0,0,91,0,8,0,0,0,225,0,130,0,104,0,253,0,206,0,0,0,245,0,113,0,83,0,173,0,0,0,29,0,84,0,222,0,172,0,121,0,216,0,64,0,223,0,0,0,245,0,161,0,0,0,241,0,29,0,0,0,111,0,56,0,0,0,104,0,2,0,60,0,88,0,250,0,177,0,101,0,187,0,0,0,59,0,161,0,64,0,0,0,255,0,105,0,76,0,0,0,40,0,94,0,138,0,116,0,81,0,0,0,95,0,0,0,0,0,24,0,28,0,105,0,182,0,0,0,180,0,55,0,233,0,0,0,0,0,108,0,108,0,215,0,67,0,193,0,122,0,0,0,179,0,0,0,230,0,235,0,159,0,34,0,117,0,157,0,0,0,14,0,0,0,0,0,220,0,56,0,111,0,207,0,123,0,51,0,0,0,9,0,0,0,125,0,65,0,51,0,151,0,193,0,17,0,89,0,171,0,11,0,39,0,234,0,0,0,31,0,49,0,0,0,83,0,20,0,97,0,0,0,190,0,160,0,123,0,229,0,163,0,241,0,191,0,175,0,2,0,26,0,0,0,198,0,22,0,210,0,65,0,198,0,0,0,92,0,94,0,203,0,229,0,0,0,0,0,191,0,161,0,2,0,0,0,70,0,26,0,0,0,0,0,158,0,161,0,158,0,190,0,114,0,0,0,0,0,158,0,0,0,10,0,0,0,89,0,222,0,0,0,217,0,61,0,100,0,181,0,32,0,8,0,185,0,24,0,41,0,193,0,7,0,81,0,0,0,150,0,122,0,25,0,170,0,229,0,142,0,188,0);
signal scenario_full  : scenario_type := (83,31,83,30,83,29,83,28,101,31,202,31,89,31,89,30,89,29,89,28,154,31,231,31,211,31,223,31,58,31,132,31,107,31,87,31,42,31,81,31,81,30,118,31,135,31,193,31,222,31,226,31,249,31,20,31,132,31,84,31,84,30,180,31,84,31,158,31,114,31,35,31,35,30,42,31,181,31,119,31,119,30,35,31,158,31,158,30,158,29,158,28,145,31,13,31,251,31,98,31,250,31,225,31,225,30,26,31,26,30,75,31,29,31,65,31,110,31,236,31,103,31,197,31,49,31,79,31,22,31,22,30,22,29,139,31,159,31,219,31,176,31,176,30,13,31,77,31,77,30,216,31,62,31,2,31,2,30,97,31,163,31,163,30,5,31,54,31,41,31,41,30,9,31,96,31,200,31,215,31,227,31,86,31,225,31,241,31,208,31,37,31,49,31,228,31,156,31,11,31,222,31,64,31,197,31,197,30,36,31,171,31,86,31,59,31,200,31,229,31,112,31,79,31,101,31,229,31,25,31,184,31,184,30,200,31,42,31,161,31,22,31,115,31,115,30,180,31,16,31,72,31,113,31,74,31,171,31,5,31,66,31,66,30,60,31,159,31,248,31,212,31,69,31,119,31,50,31,239,31,128,31,190,31,94,31,118,31,206,31,119,31,22,31,22,30,12,31,4,31,236,31,221,31,75,31,69,31,69,30,69,29,244,31,156,31,156,30,128,31,74,31,74,30,138,31,134,31,72,31,72,30,82,31,90,31,113,31,231,31,231,30,49,31,177,31,55,31,14,31,150,31,70,31,111,31,158,31,37,31,215,31,9,31,43,31,154,31,229,31,43,31,162,31,218,31,72,31,160,31,160,30,186,31,126,31,59,31,145,31,137,31,71,31,232,31,226,31,174,31,35,31,192,31,192,30,155,31,38,31,247,31,160,31,1,31,1,30,76,31,33,31,247,31,148,31,113,31,31,31,140,31,21,31,82,31,82,30,14,31,230,31,7,31,28,31,99,31,54,31,1,31,146,31,160,31,120,31,120,30,120,29,120,28,9,31,32,31,176,31,176,30,79,31,139,31,32,31,4,31,4,30,184,31,53,31,190,31,150,31,213,31,26,31,76,31,108,31,85,31,254,31,254,30,64,31,201,31,132,31,73,31,153,31,109,31,200,31,168,31,168,30,20,31,20,30,113,31,212,31,145,31,241,31,72,31,170,31,150,31,144,31,130,31,10,31,25,31,25,30,167,31,156,31,225,31,225,30,208,31,38,31,38,30,38,29,140,31,145,31,238,31,74,31,126,31,246,31,18,31,109,31,109,30,7,31,98,31,43,31,7,31,172,31,45,31,28,31,102,31,74,31,14,31,133,31,13,31,139,31,139,30,138,31,138,30,202,31,150,31,177,31,193,31,229,31,87,31,18,31,49,31,215,31,50,31,241,31,183,31,183,30,167,31,22,31,227,31,97,31,97,30,189,31,130,31,130,30,133,31,196,31,196,30,174,31,231,31,166,31,226,31,30,31,245,31,184,31,184,30,102,31,102,30,65,31,234,31,241,31,241,30,154,31,154,30,241,31,216,31,219,31,46,31,125,31,133,31,173,31,180,31,180,30,103,31,94,31,235,31,47,31,62,31,163,31,132,31,243,31,243,30,239,31,204,31,243,31,116,31,116,30,116,29,42,31,192,31,7,31,202,31,50,31,50,30,235,31,66,31,194,31,194,30,245,31,90,31,100,31,100,30,100,29,105,31,79,31,217,31,153,31,151,31,177,31,231,31,25,31,59,31,166,31,129,31,134,31,10,31,65,31,65,30,186,31,199,31,100,31,100,30,69,31,135,31,157,31,49,31,181,31,48,31,48,30,38,31,253,31,107,31,56,31,97,31,120,31,13,31,74,31,154,31,119,31,211,31,45,31,56,31,56,30,43,31,9,31,188,31,188,30,2,31,2,30,128,31,28,31,28,30,83,31,131,31,211,31,140,31,103,31,216,31,24,31,24,30,183,31,173,31,108,31,108,30,204,31,87,31,167,31,167,30,167,29,63,31,246,31,7,31,195,31,200,31,156,31,156,30,204,31,230,31,53,31,127,31,148,31,227,31,251,31,253,31,31,31,22,31,114,31,114,30,98,31,85,31,187,31,105,31,105,30,28,31,103,31,204,31,204,30,101,31,101,30,53,31,221,31,145,31,145,30,231,31,247,31,53,31,69,31,171,31,171,30,171,29,91,31,8,31,8,30,225,31,130,31,104,31,253,31,206,31,206,30,245,31,113,31,83,31,173,31,173,30,29,31,84,31,222,31,172,31,121,31,216,31,64,31,223,31,223,30,245,31,161,31,161,30,241,31,29,31,29,30,111,31,56,31,56,30,104,31,2,31,60,31,88,31,250,31,177,31,101,31,187,31,187,30,59,31,161,31,64,31,64,30,255,31,105,31,76,31,76,30,40,31,94,31,138,31,116,31,81,31,81,30,95,31,95,30,95,29,24,31,28,31,105,31,182,31,182,30,180,31,55,31,233,31,233,30,233,29,108,31,108,31,215,31,67,31,193,31,122,31,122,30,179,31,179,30,230,31,235,31,159,31,34,31,117,31,157,31,157,30,14,31,14,30,14,29,220,31,56,31,111,31,207,31,123,31,51,31,51,30,9,31,9,30,125,31,65,31,51,31,151,31,193,31,17,31,89,31,171,31,11,31,39,31,234,31,234,30,31,31,49,31,49,30,83,31,20,31,97,31,97,30,190,31,160,31,123,31,229,31,163,31,241,31,191,31,175,31,2,31,26,31,26,30,198,31,22,31,210,31,65,31,198,31,198,30,92,31,94,31,203,31,229,31,229,30,229,29,191,31,161,31,2,31,2,30,70,31,26,31,26,30,26,29,158,31,161,31,158,31,190,31,114,31,114,30,114,29,158,31,158,30,10,31,10,30,89,31,222,31,222,30,217,31,61,31,100,31,181,31,32,31,8,31,185,31,24,31,41,31,193,31,7,31,81,31,81,30,150,31,122,31,25,31,170,31,229,31,142,31,188,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
