-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 412;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,176,0,144,0,160,0,171,0,170,0,222,0,166,0,78,0,0,0,6,0,0,0,185,0,88,0,217,0,77,0,87,0,149,0,0,0,149,0,0,0,96,0,0,0,137,0,0,0,213,0,0,0,5,0,61,0,142,0,64,0,218,0,159,0,182,0,229,0,120,0,0,0,116,0,247,0,152,0,0,0,81,0,135,0,143,0,154,0,0,0,252,0,191,0,26,0,42,0,0,0,0,0,0,0,13,0,86,0,141,0,191,0,23,0,160,0,0,0,95,0,78,0,147,0,231,0,0,0,78,0,98,0,31,0,176,0,121,0,31,0,0,0,80,0,146,0,69,0,125,0,206,0,205,0,76,0,111,0,16,0,217,0,82,0,168,0,145,0,0,0,0,0,74,0,30,0,202,0,187,0,16,0,0,0,250,0,112,0,203,0,240,0,235,0,106,0,70,0,205,0,64,0,70,0,216,0,6,0,175,0,157,0,0,0,224,0,71,0,248,0,254,0,0,0,52,0,168,0,0,0,21,0,139,0,162,0,43,0,203,0,0,0,181,0,147,0,124,0,0,0,8,0,108,0,71,0,135,0,6,0,204,0,221,0,0,0,107,0,34,0,69,0,118,0,110,0,173,0,0,0,58,0,221,0,0,0,242,0,0,0,185,0,174,0,130,0,0,0,31,0,211,0,68,0,0,0,0,0,176,0,55,0,187,0,28,0,107,0,251,0,78,0,54,0,3,0,0,0,236,0,240,0,47,0,0,0,0,0,34,0,0,0,116,0,0,0,210,0,46,0,206,0,234,0,251,0,176,0,124,0,231,0,0,0,162,0,247,0,211,0,158,0,224,0,90,0,85,0,32,0,176,0,168,0,79,0,181,0,147,0,244,0,154,0,37,0,15,0,57,0,174,0,84,0,38,0,163,0,195,0,0,0,0,0,0,0,0,0,79,0,186,0,233,0,251,0,122,0,0,0,0,0,5,0,78,0,239,0,171,0,41,0,166,0,240,0,247,0,0,0,0,0,218,0,223,0,217,0,183,0,182,0,187,0,155,0,0,0,169,0,0,0,202,0,118,0,31,0,222,0,85,0,0,0,89,0,31,0,217,0,49,0,126,0,207,0,93,0,186,0,41,0,0,0,138,0,143,0,0,0,27,0,0,0,69,0,165,0,0,0,133,0,0,0,140,0,233,0,80,0,31,0,188,0,20,0,212,0,0,0,0,0,145,0,173,0,94,0,0,0,0,0,199,0,0,0,0,0,0,0,0,0,82,0,216,0,0,0,0,0,0,0,35,0,103,0,243,0,0,0,0,0,38,0,192,0,0,0,0,0,0,0,138,0,230,0,0,0,249,0,0,0,33,0,0,0,63,0,222,0,105,0,5,0,249,0,237,0,27,0,0,0,172,0,225,0,123,0,168,0,204,0,110,0,29,0,88,0,153,0,0,0,108,0,0,0,0,0,6,0,250,0,138,0,93,0,31,0,234,0,88,0,209,0,87,0,107,0,0,0,18,0,0,0,85,0,74,0,46,0,163,0,0,0,60,0,96,0,235,0,86,0,0,0,58,0,206,0,179,0,206,0,252,0,236,0,231,0,0,0,197,0,181,0,178,0,181,0,81,0,253,0,51,0,33,0,39,0,253,0,0,0,161,0,161,0,132,0,0,0,49,0,166,0,131,0,0,0,98,0,105,0,249,0,6,0,190,0,33,0,32,0,0,0,107,0,22,0,148,0,1,0,177,0,155,0,116,0,0,0,0,0,189,0,0,0,114,0,36,0,26,0,199,0,0,0,102,0,84,0,128,0,91,0,79,0,200,0,210,0,77,0,43,0,10,0,70,0,249,0,135,0);
signal scenario_full  : scenario_type := (0,0,176,31,144,31,160,31,171,31,170,31,222,31,166,31,78,31,78,30,6,31,6,30,185,31,88,31,217,31,77,31,87,31,149,31,149,30,149,31,149,30,96,31,96,30,137,31,137,30,213,31,213,30,5,31,61,31,142,31,64,31,218,31,159,31,182,31,229,31,120,31,120,30,116,31,247,31,152,31,152,30,81,31,135,31,143,31,154,31,154,30,252,31,191,31,26,31,42,31,42,30,42,29,42,28,13,31,86,31,141,31,191,31,23,31,160,31,160,30,95,31,78,31,147,31,231,31,231,30,78,31,98,31,31,31,176,31,121,31,31,31,31,30,80,31,146,31,69,31,125,31,206,31,205,31,76,31,111,31,16,31,217,31,82,31,168,31,145,31,145,30,145,29,74,31,30,31,202,31,187,31,16,31,16,30,250,31,112,31,203,31,240,31,235,31,106,31,70,31,205,31,64,31,70,31,216,31,6,31,175,31,157,31,157,30,224,31,71,31,248,31,254,31,254,30,52,31,168,31,168,30,21,31,139,31,162,31,43,31,203,31,203,30,181,31,147,31,124,31,124,30,8,31,108,31,71,31,135,31,6,31,204,31,221,31,221,30,107,31,34,31,69,31,118,31,110,31,173,31,173,30,58,31,221,31,221,30,242,31,242,30,185,31,174,31,130,31,130,30,31,31,211,31,68,31,68,30,68,29,176,31,55,31,187,31,28,31,107,31,251,31,78,31,54,31,3,31,3,30,236,31,240,31,47,31,47,30,47,29,34,31,34,30,116,31,116,30,210,31,46,31,206,31,234,31,251,31,176,31,124,31,231,31,231,30,162,31,247,31,211,31,158,31,224,31,90,31,85,31,32,31,176,31,168,31,79,31,181,31,147,31,244,31,154,31,37,31,15,31,57,31,174,31,84,31,38,31,163,31,195,31,195,30,195,29,195,28,195,27,79,31,186,31,233,31,251,31,122,31,122,30,122,29,5,31,78,31,239,31,171,31,41,31,166,31,240,31,247,31,247,30,247,29,218,31,223,31,217,31,183,31,182,31,187,31,155,31,155,30,169,31,169,30,202,31,118,31,31,31,222,31,85,31,85,30,89,31,31,31,217,31,49,31,126,31,207,31,93,31,186,31,41,31,41,30,138,31,143,31,143,30,27,31,27,30,69,31,165,31,165,30,133,31,133,30,140,31,233,31,80,31,31,31,188,31,20,31,212,31,212,30,212,29,145,31,173,31,94,31,94,30,94,29,199,31,199,30,199,29,199,28,199,27,82,31,216,31,216,30,216,29,216,28,35,31,103,31,243,31,243,30,243,29,38,31,192,31,192,30,192,29,192,28,138,31,230,31,230,30,249,31,249,30,33,31,33,30,63,31,222,31,105,31,5,31,249,31,237,31,27,31,27,30,172,31,225,31,123,31,168,31,204,31,110,31,29,31,88,31,153,31,153,30,108,31,108,30,108,29,6,31,250,31,138,31,93,31,31,31,234,31,88,31,209,31,87,31,107,31,107,30,18,31,18,30,85,31,74,31,46,31,163,31,163,30,60,31,96,31,235,31,86,31,86,30,58,31,206,31,179,31,206,31,252,31,236,31,231,31,231,30,197,31,181,31,178,31,181,31,81,31,253,31,51,31,33,31,39,31,253,31,253,30,161,31,161,31,132,31,132,30,49,31,166,31,131,31,131,30,98,31,105,31,249,31,6,31,190,31,33,31,32,31,32,30,107,31,22,31,148,31,1,31,177,31,155,31,116,31,116,30,116,29,189,31,189,30,114,31,36,31,26,31,199,31,199,30,102,31,84,31,128,31,91,31,79,31,200,31,210,31,77,31,43,31,10,31,70,31,249,31,135,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
