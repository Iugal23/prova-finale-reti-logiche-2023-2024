-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 705;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (63,0,0,0,50,0,128,0,82,0,32,0,0,0,0,0,112,0,87,0,182,0,106,0,0,0,10,0,78,0,164,0,197,0,24,0,190,0,43,0,26,0,195,0,154,0,0,0,0,0,216,0,121,0,0,0,71,0,80,0,147,0,232,0,126,0,58,0,6,0,170,0,238,0,0,0,232,0,0,0,167,0,231,0,27,0,248,0,109,0,0,0,109,0,59,0,254,0,160,0,48,0,63,0,90,0,93,0,113,0,118,0,39,0,155,0,246,0,121,0,0,0,108,0,5,0,84,0,126,0,190,0,124,0,28,0,149,0,74,0,149,0,188,0,37,0,0,0,236,0,103,0,139,0,36,0,181,0,233,0,138,0,0,0,22,0,254,0,182,0,244,0,149,0,64,0,239,0,146,0,189,0,152,0,197,0,91,0,0,0,238,0,60,0,54,0,223,0,64,0,0,0,233,0,6,0,223,0,0,0,254,0,197,0,228,0,116,0,177,0,107,0,28,0,58,0,40,0,156,0,220,0,51,0,242,0,100,0,0,0,132,0,0,0,143,0,239,0,106,0,223,0,52,0,66,0,224,0,0,0,72,0,82,0,0,0,219,0,166,0,209,0,0,0,3,0,184,0,164,0,65,0,166,0,87,0,173,0,237,0,219,0,0,0,169,0,0,0,214,0,0,0,165,0,122,0,172,0,24,0,235,0,51,0,79,0,26,0,161,0,192,0,154,0,78,0,195,0,112,0,30,0,209,0,0,0,136,0,0,0,0,0,52,0,33,0,87,0,229,0,104,0,155,0,0,0,46,0,103,0,80,0,123,0,12,0,106,0,35,0,44,0,107,0,76,0,115,0,241,0,163,0,231,0,213,0,6,0,61,0,110,0,110,0,135,0,228,0,0,0,33,0,233,0,122,0,94,0,0,0,122,0,187,0,20,0,0,0,125,0,240,0,215,0,248,0,18,0,201,0,40,0,230,0,0,0,196,0,0,0,163,0,84,0,245,0,140,0,147,0,150,0,0,0,0,0,0,0,112,0,93,0,255,0,170,0,18,0,143,0,112,0,61,0,156,0,203,0,195,0,191,0,20,0,210,0,189,0,81,0,203,0,81,0,4,0,238,0,0,0,0,0,198,0,20,0,0,0,31,0,235,0,224,0,237,0,162,0,60,0,138,0,127,0,0,0,0,0,179,0,72,0,73,0,150,0,241,0,164,0,0,0,242,0,61,0,244,0,0,0,0,0,0,0,102,0,14,0,166,0,52,0,108,0,61,0,118,0,168,0,215,0,0,0,79,0,0,0,131,0,7,0,0,0,15,0,198,0,0,0,30,0,0,0,168,0,217,0,142,0,149,0,0,0,220,0,151,0,55,0,0,0,231,0,21,0,0,0,0,0,165,0,0,0,10,0,153,0,4,0,241,0,93,0,0,0,0,0,198,0,206,0,38,0,151,0,40,0,147,0,76,0,43,0,0,0,200,0,0,0,0,0,0,0,242,0,28,0,5,0,128,0,182,0,205,0,162,0,191,0,196,0,199,0,253,0,0,0,0,0,120,0,220,0,0,0,15,0,21,0,118,0,0,0,246,0,221,0,47,0,0,0,41,0,206,0,35,0,239,0,91,0,165,0,0,0,0,0,31,0,246,0,105,0,164,0,0,0,247,0,0,0,6,0,21,0,55,0,5,0,133,0,192,0,111,0,120,0,213,0,71,0,59,0,11,0,254,0,49,0,229,0,2,0,96,0,200,0,250,0,113,0,35,0,136,0,225,0,160,0,158,0,132,0,218,0,31,0,0,0,201,0,0,0,50,0,209,0,139,0,0,0,244,0,196,0,174,0,0,0,132,0,202,0,164,0,80,0,201,0,215,0,134,0,206,0,75,0,93,0,144,0,69,0,69,0,18,0,248,0,125,0,252,0,225,0,81,0,63,0,113,0,0,0,108,0,29,0,160,0,0,0,194,0,235,0,187,0,222,0,34,0,160,0,0,0,0,0,232,0,52,0,27,0,80,0,185,0,206,0,28,0,105,0,8,0,0,0,0,0,0,0,247,0,179,0,7,0,217,0,194,0,132,0,67,0,190,0,237,0,12,0,251,0,91,0,179,0,212,0,0,0,30,0,59,0,245,0,242,0,143,0,10,0,218,0,0,0,230,0,154,0,156,0,114,0,151,0,226,0,26,0,88,0,216,0,155,0,230,0,0,0,188,0,142,0,75,0,207,0,205,0,0,0,86,0,92,0,106,0,133,0,30,0,0,0,99,0,93,0,168,0,0,0,185,0,233,0,59,0,12,0,50,0,251,0,46,0,26,0,0,0,0,0,226,0,31,0,143,0,75,0,0,0,182,0,130,0,0,0,99,0,103,0,21,0,7,0,116,0,141,0,0,0,10,0,141,0,57,0,247,0,0,0,85,0,201,0,124,0,15,0,254,0,91,0,46,0,242,0,132,0,0,0,24,0,0,0,111,0,0,0,54,0,22,0,234,0,145,0,182,0,248,0,157,0,100,0,108,0,29,0,64,0,0,0,30,0,29,0,222,0,107,0,76,0,146,0,223,0,194,0,126,0,20,0,133,0,91,0,117,0,196,0,165,0,110,0,0,0,78,0,108,0,163,0,147,0,0,0,96,0,164,0,0,0,25,0,0,0,139,0,214,0,67,0,123,0,15,0,117,0,75,0,0,0,0,0,242,0,68,0,0,0,7,0,101,0,0,0,0,0,212,0,137,0,182,0,131,0,0,0,208,0,160,0,135,0,199,0,210,0,133,0,163,0,67,0,0,0,24,0,80,0,97,0,12,0,109,0,133,0,74,0,2,0,191,0,0,0,0,0,177,0,68,0,195,0,27,0,233,0,19,0,3,0,94,0,52,0,227,0,184,0,228,0,91,0,24,0,0,0,224,0,109,0,239,0,0,0,0,0,0,0,130,0,156,0,148,0,0,0,0,0,65,0,70,0,44,0,0,0,16,0,0,0,0,0,79,0,171,0,26,0,123,0,123,0,161,0,0,0,0,0,115,0,49,0,205,0,254,0,22,0,138,0,234,0,0,0,19,0,59,0,82,0,33,0,17,0,246,0,0,0,0,0,0,0,167,0,231,0,241,0,159,0,100,0,72,0,85,0,6,0,246,0,0,0,163,0,3,0,0,0,0,0,170,0,136,0);
signal scenario_full  : scenario_type := (63,31,63,30,50,31,128,31,82,31,32,31,32,30,32,29,112,31,87,31,182,31,106,31,106,30,10,31,78,31,164,31,197,31,24,31,190,31,43,31,26,31,195,31,154,31,154,30,154,29,216,31,121,31,121,30,71,31,80,31,147,31,232,31,126,31,58,31,6,31,170,31,238,31,238,30,232,31,232,30,167,31,231,31,27,31,248,31,109,31,109,30,109,31,59,31,254,31,160,31,48,31,63,31,90,31,93,31,113,31,118,31,39,31,155,31,246,31,121,31,121,30,108,31,5,31,84,31,126,31,190,31,124,31,28,31,149,31,74,31,149,31,188,31,37,31,37,30,236,31,103,31,139,31,36,31,181,31,233,31,138,31,138,30,22,31,254,31,182,31,244,31,149,31,64,31,239,31,146,31,189,31,152,31,197,31,91,31,91,30,238,31,60,31,54,31,223,31,64,31,64,30,233,31,6,31,223,31,223,30,254,31,197,31,228,31,116,31,177,31,107,31,28,31,58,31,40,31,156,31,220,31,51,31,242,31,100,31,100,30,132,31,132,30,143,31,239,31,106,31,223,31,52,31,66,31,224,31,224,30,72,31,82,31,82,30,219,31,166,31,209,31,209,30,3,31,184,31,164,31,65,31,166,31,87,31,173,31,237,31,219,31,219,30,169,31,169,30,214,31,214,30,165,31,122,31,172,31,24,31,235,31,51,31,79,31,26,31,161,31,192,31,154,31,78,31,195,31,112,31,30,31,209,31,209,30,136,31,136,30,136,29,52,31,33,31,87,31,229,31,104,31,155,31,155,30,46,31,103,31,80,31,123,31,12,31,106,31,35,31,44,31,107,31,76,31,115,31,241,31,163,31,231,31,213,31,6,31,61,31,110,31,110,31,135,31,228,31,228,30,33,31,233,31,122,31,94,31,94,30,122,31,187,31,20,31,20,30,125,31,240,31,215,31,248,31,18,31,201,31,40,31,230,31,230,30,196,31,196,30,163,31,84,31,245,31,140,31,147,31,150,31,150,30,150,29,150,28,112,31,93,31,255,31,170,31,18,31,143,31,112,31,61,31,156,31,203,31,195,31,191,31,20,31,210,31,189,31,81,31,203,31,81,31,4,31,238,31,238,30,238,29,198,31,20,31,20,30,31,31,235,31,224,31,237,31,162,31,60,31,138,31,127,31,127,30,127,29,179,31,72,31,73,31,150,31,241,31,164,31,164,30,242,31,61,31,244,31,244,30,244,29,244,28,102,31,14,31,166,31,52,31,108,31,61,31,118,31,168,31,215,31,215,30,79,31,79,30,131,31,7,31,7,30,15,31,198,31,198,30,30,31,30,30,168,31,217,31,142,31,149,31,149,30,220,31,151,31,55,31,55,30,231,31,21,31,21,30,21,29,165,31,165,30,10,31,153,31,4,31,241,31,93,31,93,30,93,29,198,31,206,31,38,31,151,31,40,31,147,31,76,31,43,31,43,30,200,31,200,30,200,29,200,28,242,31,28,31,5,31,128,31,182,31,205,31,162,31,191,31,196,31,199,31,253,31,253,30,253,29,120,31,220,31,220,30,15,31,21,31,118,31,118,30,246,31,221,31,47,31,47,30,41,31,206,31,35,31,239,31,91,31,165,31,165,30,165,29,31,31,246,31,105,31,164,31,164,30,247,31,247,30,6,31,21,31,55,31,5,31,133,31,192,31,111,31,120,31,213,31,71,31,59,31,11,31,254,31,49,31,229,31,2,31,96,31,200,31,250,31,113,31,35,31,136,31,225,31,160,31,158,31,132,31,218,31,31,31,31,30,201,31,201,30,50,31,209,31,139,31,139,30,244,31,196,31,174,31,174,30,132,31,202,31,164,31,80,31,201,31,215,31,134,31,206,31,75,31,93,31,144,31,69,31,69,31,18,31,248,31,125,31,252,31,225,31,81,31,63,31,113,31,113,30,108,31,29,31,160,31,160,30,194,31,235,31,187,31,222,31,34,31,160,31,160,30,160,29,232,31,52,31,27,31,80,31,185,31,206,31,28,31,105,31,8,31,8,30,8,29,8,28,247,31,179,31,7,31,217,31,194,31,132,31,67,31,190,31,237,31,12,31,251,31,91,31,179,31,212,31,212,30,30,31,59,31,245,31,242,31,143,31,10,31,218,31,218,30,230,31,154,31,156,31,114,31,151,31,226,31,26,31,88,31,216,31,155,31,230,31,230,30,188,31,142,31,75,31,207,31,205,31,205,30,86,31,92,31,106,31,133,31,30,31,30,30,99,31,93,31,168,31,168,30,185,31,233,31,59,31,12,31,50,31,251,31,46,31,26,31,26,30,26,29,226,31,31,31,143,31,75,31,75,30,182,31,130,31,130,30,99,31,103,31,21,31,7,31,116,31,141,31,141,30,10,31,141,31,57,31,247,31,247,30,85,31,201,31,124,31,15,31,254,31,91,31,46,31,242,31,132,31,132,30,24,31,24,30,111,31,111,30,54,31,22,31,234,31,145,31,182,31,248,31,157,31,100,31,108,31,29,31,64,31,64,30,30,31,29,31,222,31,107,31,76,31,146,31,223,31,194,31,126,31,20,31,133,31,91,31,117,31,196,31,165,31,110,31,110,30,78,31,108,31,163,31,147,31,147,30,96,31,164,31,164,30,25,31,25,30,139,31,214,31,67,31,123,31,15,31,117,31,75,31,75,30,75,29,242,31,68,31,68,30,7,31,101,31,101,30,101,29,212,31,137,31,182,31,131,31,131,30,208,31,160,31,135,31,199,31,210,31,133,31,163,31,67,31,67,30,24,31,80,31,97,31,12,31,109,31,133,31,74,31,2,31,191,31,191,30,191,29,177,31,68,31,195,31,27,31,233,31,19,31,3,31,94,31,52,31,227,31,184,31,228,31,91,31,24,31,24,30,224,31,109,31,239,31,239,30,239,29,239,28,130,31,156,31,148,31,148,30,148,29,65,31,70,31,44,31,44,30,16,31,16,30,16,29,79,31,171,31,26,31,123,31,123,31,161,31,161,30,161,29,115,31,49,31,205,31,254,31,22,31,138,31,234,31,234,30,19,31,59,31,82,31,33,31,17,31,246,31,246,30,246,29,246,28,167,31,231,31,241,31,159,31,100,31,72,31,85,31,6,31,246,31,246,30,163,31,3,31,3,30,3,29,170,31,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
