-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 937;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,131,0,50,0,191,0,196,0,41,0,188,0,81,0,100,0,244,0,137,0,56,0,236,0,159,0,46,0,76,0,88,0,190,0,82,0,104,0,36,0,133,0,161,0,0,0,158,0,89,0,203,0,112,0,119,0,173,0,31,0,0,0,109,0,0,0,247,0,0,0,67,0,164,0,0,0,0,0,0,0,219,0,89,0,50,0,218,0,105,0,231,0,186,0,53,0,0,0,140,0,210,0,198,0,152,0,78,0,100,0,27,0,0,0,93,0,156,0,60,0,118,0,0,0,219,0,0,0,133,0,105,0,0,0,0,0,35,0,0,0,255,0,227,0,0,0,79,0,31,0,182,0,0,0,53,0,1,0,45,0,239,0,113,0,59,0,87,0,0,0,201,0,0,0,58,0,0,0,218,0,246,0,161,0,106,0,199,0,179,0,246,0,63,0,22,0,98,0,182,0,226,0,222,0,158,0,17,0,99,0,0,0,0,0,0,0,0,0,251,0,219,0,35,0,24,0,72,0,185,0,54,0,197,0,240,0,34,0,97,0,0,0,63,0,195,0,0,0,184,0,80,0,65,0,83,0,251,0,39,0,0,0,207,0,225,0,128,0,101,0,35,0,215,0,111,0,64,0,82,0,18,0,158,0,41,0,25,0,237,0,99,0,59,0,57,0,0,0,0,0,104,0,213,0,241,0,117,0,235,0,0,0,81,0,152,0,26,0,253,0,119,0,18,0,2,0,52,0,63,0,0,0,0,0,180,0,216,0,241,0,166,0,120,0,0,0,196,0,91,0,227,0,183,0,34,0,47,0,154,0,34,0,218,0,93,0,6,0,233,0,211,0,178,0,177,0,141,0,33,0,143,0,135,0,235,0,101,0,211,0,13,0,0,0,243,0,67,0,0,0,0,0,95,0,0,0,22,0,0,0,166,0,188,0,22,0,0,0,164,0,49,0,215,0,118,0,152,0,107,0,0,0,0,0,0,0,235,0,117,0,234,0,217,0,196,0,12,0,125,0,148,0,172,0,199,0,220,0,217,0,179,0,0,0,129,0,0,0,149,0,39,0,51,0,230,0,243,0,205,0,55,0,53,0,170,0,254,0,85,0,44,0,120,0,192,0,252,0,228,0,117,0,197,0,157,0,213,0,244,0,0,0,0,0,1,0,0,0,42,0,219,0,243,0,0,0,51,0,25,0,87,0,76,0,55,0,167,0,238,0,222,0,0,0,212,0,165,0,72,0,148,0,227,0,77,0,0,0,145,0,79,0,131,0,0,0,234,0,69,0,45,0,55,0,68,0,90,0,142,0,223,0,113,0,174,0,65,0,128,0,37,0,145,0,151,0,36,0,189,0,241,0,0,0,0,0,0,0,0,0,246,0,0,0,0,0,229,0,106,0,148,0,93,0,151,0,144,0,0,0,27,0,184,0,88,0,44,0,251,0,70,0,172,0,19,0,197,0,68,0,213,0,57,0,173,0,123,0,34,0,70,0,198,0,0,0,73,0,0,0,134,0,6,0,110,0,154,0,193,0,25,0,173,0,39,0,236,0,3,0,4,0,197,0,209,0,27,0,101,0,9,0,193,0,1,0,195,0,0,0,211,0,252,0,0,0,251,0,196,0,133,0,236,0,0,0,181,0,63,0,167,0,67,0,0,0,35,0,59,0,201,0,229,0,166,0,38,0,92,0,154,0,156,0,140,0,25,0,31,0,145,0,237,0,0,0,172,0,204,0,78,0,0,0,0,0,80,0,115,0,112,0,113,0,157,0,252,0,21,0,236,0,0,0,144,0,0,0,0,0,18,0,153,0,138,0,0,0,0,0,78,0,0,0,241,0,160,0,206,0,33,0,239,0,144,0,214,0,74,0,0,0,65,0,213,0,229,0,186,0,0,0,83,0,0,0,228,0,217,0,63,0,25,0,44,0,106,0,0,0,194,0,46,0,0,0,0,0,40,0,0,0,0,0,89,0,167,0,0,0,0,0,25,0,162,0,0,0,19,0,226,0,0,0,0,0,136,0,174,0,127,0,73,0,24,0,227,0,125,0,178,0,211,0,0,0,0,0,0,0,12,0,0,0,148,0,55,0,100,0,84,0,71,0,58,0,0,0,0,0,0,0,64,0,164,0,188,0,167,0,228,0,25,0,71,0,37,0,220,0,51,0,46,0,140,0,0,0,203,0,22,0,13,0,180,0,0,0,247,0,93,0,201,0,0,0,30,0,62,0,126,0,0,0,163,0,149,0,0,0,173,0,100,0,55,0,200,0,43,0,112,0,29,0,98,0,254,0,0,0,212,0,244,0,185,0,56,0,82,0,180,0,0,0,71,0,226,0,0,0,218,0,117,0,31,0,1,0,183,0,231,0,239,0,62,0,101,0,33,0,0,0,0,0,120,0,89,0,54,0,200,0,82,0,0,0,0,0,87,0,40,0,0,0,0,0,225,0,0,0,0,0,66,0,134,0,124,0,0,0,0,0,10,0,41,0,0,0,186,0,175,0,0,0,212,0,165,0,71,0,38,0,0,0,252,0,75,0,235,0,25,0,171,0,141,0,240,0,189,0,18,0,214,0,167,0,210,0,33,0,115,0,0,0,0,0,191,0,245,0,101,0,188,0,72,0,238,0,185,0,15,0,124,0,53,0,122,0,205,0,187,0,0,0,254,0,0,0,0,0,152,0,0,0,161,0,118,0,67,0,159,0,163,0,0,0,0,0,0,0,22,0,117,0,182,0,92,0,233,0,5,0,20,0,76,0,212,0,75,0,99,0,0,0,177,0,254,0,247,0,127,0,0,0,0,0,186,0,190,0,45,0,126,0,30,0,0,0,163,0,110,0,0,0,190,0,104,0,113,0,62,0,211,0,26,0,218,0,53,0,229,0,0,0,203,0,187,0,42,0,63,0,133,0,103,0,108,0,120,0,98,0,119,0,216,0,238,0,95,0,190,0,46,0,56,0,145,0,113,0,16,0,0,0,190,0,103,0,0,0,143,0,196,0,160,0,16,0,102,0,150,0,96,0,0,0,24,0,138,0,35,0,31,0,12,0,0,0,0,0,199,0,141,0,145,0,0,0,254,0,0,0,0,0,183,0,95,0,116,0,226,0,0,0,39,0,0,0,62,0,205,0,0,0,78,0,241,0,0,0,37,0,28,0,15,0,4,0,0,0,69,0,244,0,5,0,223,0,25,0,249,0,2,0,200,0,140,0,229,0,92,0,234,0,248,0,149,0,234,0,123,0,18,0,24,0,5,0,109,0,140,0,108,0,0,0,79,0,13,0,0,0,191,0,18,0,30,0,100,0,169,0,80,0,229,0,164,0,0,0,10,0,220,0,218,0,63,0,106,0,0,0,253,0,44,0,0,0,0,0,25,0,12,0,199,0,40,0,199,0,10,0,0,0,54,0,189,0,185,0,0,0,109,0,112,0,0,0,0,0,135,0,135,0,242,0,152,0,0,0,107,0,65,0,136,0,107,0,0,0,0,0,199,0,0,0,112,0,134,0,0,0,52,0,232,0,8,0,181,0,0,0,0,0,0,0,151,0,215,0,156,0,61,0,12,0,0,0,32,0,229,0,190,0,71,0,28,0,245,0,94,0,3,0,0,0,133,0,0,0,166,0,185,0,178,0,108,0,0,0,93,0,142,0,0,0,129,0,127,0,0,0,182,0,0,0,0,0,87,0,133,0,146,0,110,0,68,0,1,0,102,0,95,0,176,0,5,0,246,0,145,0,0,0,233,0,99,0,0,0,22,0,3,0,45,0,197,0,122,0,206,0,37,0,86,0,18,0,213,0,22,0,18,0,0,0,0,0,0,0,0,0,159,0,88,0,235,0,162,0,97,0,21,0,48,0,23,0,30,0,182,0,0,0,0,0,85,0,16,0,234,0,65,0,222,0,192,0,198,0,214,0,94,0,0,0,0,0,19,0,0,0,190,0,196,0,184,0,0,0,221,0,39,0,252,0,99,0,178,0,140,0,113,0,166,0,252,0,66,0,0,0,185,0,0,0,6,0,98,0,239,0,206,0,58,0,220,0,13,0,192,0,35,0,60,0,0,0,30,0,128,0,133,0,0,0,148,0,55,0,178,0,184,0,90,0,254,0,0,0,29,0,0,0,58,0,0,0,181,0,0,0,247,0,0,0,21,0,185,0,70,0,37,0,28,0,1,0,239,0,228,0,19,0,0,0,0,0,0,0,105,0);
signal scenario_full  : scenario_type := (0,0,131,31,50,31,191,31,196,31,41,31,188,31,81,31,100,31,244,31,137,31,56,31,236,31,159,31,46,31,76,31,88,31,190,31,82,31,104,31,36,31,133,31,161,31,161,30,158,31,89,31,203,31,112,31,119,31,173,31,31,31,31,30,109,31,109,30,247,31,247,30,67,31,164,31,164,30,164,29,164,28,219,31,89,31,50,31,218,31,105,31,231,31,186,31,53,31,53,30,140,31,210,31,198,31,152,31,78,31,100,31,27,31,27,30,93,31,156,31,60,31,118,31,118,30,219,31,219,30,133,31,105,31,105,30,105,29,35,31,35,30,255,31,227,31,227,30,79,31,31,31,182,31,182,30,53,31,1,31,45,31,239,31,113,31,59,31,87,31,87,30,201,31,201,30,58,31,58,30,218,31,246,31,161,31,106,31,199,31,179,31,246,31,63,31,22,31,98,31,182,31,226,31,222,31,158,31,17,31,99,31,99,30,99,29,99,28,99,27,251,31,219,31,35,31,24,31,72,31,185,31,54,31,197,31,240,31,34,31,97,31,97,30,63,31,195,31,195,30,184,31,80,31,65,31,83,31,251,31,39,31,39,30,207,31,225,31,128,31,101,31,35,31,215,31,111,31,64,31,82,31,18,31,158,31,41,31,25,31,237,31,99,31,59,31,57,31,57,30,57,29,104,31,213,31,241,31,117,31,235,31,235,30,81,31,152,31,26,31,253,31,119,31,18,31,2,31,52,31,63,31,63,30,63,29,180,31,216,31,241,31,166,31,120,31,120,30,196,31,91,31,227,31,183,31,34,31,47,31,154,31,34,31,218,31,93,31,6,31,233,31,211,31,178,31,177,31,141,31,33,31,143,31,135,31,235,31,101,31,211,31,13,31,13,30,243,31,67,31,67,30,67,29,95,31,95,30,22,31,22,30,166,31,188,31,22,31,22,30,164,31,49,31,215,31,118,31,152,31,107,31,107,30,107,29,107,28,235,31,117,31,234,31,217,31,196,31,12,31,125,31,148,31,172,31,199,31,220,31,217,31,179,31,179,30,129,31,129,30,149,31,39,31,51,31,230,31,243,31,205,31,55,31,53,31,170,31,254,31,85,31,44,31,120,31,192,31,252,31,228,31,117,31,197,31,157,31,213,31,244,31,244,30,244,29,1,31,1,30,42,31,219,31,243,31,243,30,51,31,25,31,87,31,76,31,55,31,167,31,238,31,222,31,222,30,212,31,165,31,72,31,148,31,227,31,77,31,77,30,145,31,79,31,131,31,131,30,234,31,69,31,45,31,55,31,68,31,90,31,142,31,223,31,113,31,174,31,65,31,128,31,37,31,145,31,151,31,36,31,189,31,241,31,241,30,241,29,241,28,241,27,246,31,246,30,246,29,229,31,106,31,148,31,93,31,151,31,144,31,144,30,27,31,184,31,88,31,44,31,251,31,70,31,172,31,19,31,197,31,68,31,213,31,57,31,173,31,123,31,34,31,70,31,198,31,198,30,73,31,73,30,134,31,6,31,110,31,154,31,193,31,25,31,173,31,39,31,236,31,3,31,4,31,197,31,209,31,27,31,101,31,9,31,193,31,1,31,195,31,195,30,211,31,252,31,252,30,251,31,196,31,133,31,236,31,236,30,181,31,63,31,167,31,67,31,67,30,35,31,59,31,201,31,229,31,166,31,38,31,92,31,154,31,156,31,140,31,25,31,31,31,145,31,237,31,237,30,172,31,204,31,78,31,78,30,78,29,80,31,115,31,112,31,113,31,157,31,252,31,21,31,236,31,236,30,144,31,144,30,144,29,18,31,153,31,138,31,138,30,138,29,78,31,78,30,241,31,160,31,206,31,33,31,239,31,144,31,214,31,74,31,74,30,65,31,213,31,229,31,186,31,186,30,83,31,83,30,228,31,217,31,63,31,25,31,44,31,106,31,106,30,194,31,46,31,46,30,46,29,40,31,40,30,40,29,89,31,167,31,167,30,167,29,25,31,162,31,162,30,19,31,226,31,226,30,226,29,136,31,174,31,127,31,73,31,24,31,227,31,125,31,178,31,211,31,211,30,211,29,211,28,12,31,12,30,148,31,55,31,100,31,84,31,71,31,58,31,58,30,58,29,58,28,64,31,164,31,188,31,167,31,228,31,25,31,71,31,37,31,220,31,51,31,46,31,140,31,140,30,203,31,22,31,13,31,180,31,180,30,247,31,93,31,201,31,201,30,30,31,62,31,126,31,126,30,163,31,149,31,149,30,173,31,100,31,55,31,200,31,43,31,112,31,29,31,98,31,254,31,254,30,212,31,244,31,185,31,56,31,82,31,180,31,180,30,71,31,226,31,226,30,218,31,117,31,31,31,1,31,183,31,231,31,239,31,62,31,101,31,33,31,33,30,33,29,120,31,89,31,54,31,200,31,82,31,82,30,82,29,87,31,40,31,40,30,40,29,225,31,225,30,225,29,66,31,134,31,124,31,124,30,124,29,10,31,41,31,41,30,186,31,175,31,175,30,212,31,165,31,71,31,38,31,38,30,252,31,75,31,235,31,25,31,171,31,141,31,240,31,189,31,18,31,214,31,167,31,210,31,33,31,115,31,115,30,115,29,191,31,245,31,101,31,188,31,72,31,238,31,185,31,15,31,124,31,53,31,122,31,205,31,187,31,187,30,254,31,254,30,254,29,152,31,152,30,161,31,118,31,67,31,159,31,163,31,163,30,163,29,163,28,22,31,117,31,182,31,92,31,233,31,5,31,20,31,76,31,212,31,75,31,99,31,99,30,177,31,254,31,247,31,127,31,127,30,127,29,186,31,190,31,45,31,126,31,30,31,30,30,163,31,110,31,110,30,190,31,104,31,113,31,62,31,211,31,26,31,218,31,53,31,229,31,229,30,203,31,187,31,42,31,63,31,133,31,103,31,108,31,120,31,98,31,119,31,216,31,238,31,95,31,190,31,46,31,56,31,145,31,113,31,16,31,16,30,190,31,103,31,103,30,143,31,196,31,160,31,16,31,102,31,150,31,96,31,96,30,24,31,138,31,35,31,31,31,12,31,12,30,12,29,199,31,141,31,145,31,145,30,254,31,254,30,254,29,183,31,95,31,116,31,226,31,226,30,39,31,39,30,62,31,205,31,205,30,78,31,241,31,241,30,37,31,28,31,15,31,4,31,4,30,69,31,244,31,5,31,223,31,25,31,249,31,2,31,200,31,140,31,229,31,92,31,234,31,248,31,149,31,234,31,123,31,18,31,24,31,5,31,109,31,140,31,108,31,108,30,79,31,13,31,13,30,191,31,18,31,30,31,100,31,169,31,80,31,229,31,164,31,164,30,10,31,220,31,218,31,63,31,106,31,106,30,253,31,44,31,44,30,44,29,25,31,12,31,199,31,40,31,199,31,10,31,10,30,54,31,189,31,185,31,185,30,109,31,112,31,112,30,112,29,135,31,135,31,242,31,152,31,152,30,107,31,65,31,136,31,107,31,107,30,107,29,199,31,199,30,112,31,134,31,134,30,52,31,232,31,8,31,181,31,181,30,181,29,181,28,151,31,215,31,156,31,61,31,12,31,12,30,32,31,229,31,190,31,71,31,28,31,245,31,94,31,3,31,3,30,133,31,133,30,166,31,185,31,178,31,108,31,108,30,93,31,142,31,142,30,129,31,127,31,127,30,182,31,182,30,182,29,87,31,133,31,146,31,110,31,68,31,1,31,102,31,95,31,176,31,5,31,246,31,145,31,145,30,233,31,99,31,99,30,22,31,3,31,45,31,197,31,122,31,206,31,37,31,86,31,18,31,213,31,22,31,18,31,18,30,18,29,18,28,18,27,159,31,88,31,235,31,162,31,97,31,21,31,48,31,23,31,30,31,182,31,182,30,182,29,85,31,16,31,234,31,65,31,222,31,192,31,198,31,214,31,94,31,94,30,94,29,19,31,19,30,190,31,196,31,184,31,184,30,221,31,39,31,252,31,99,31,178,31,140,31,113,31,166,31,252,31,66,31,66,30,185,31,185,30,6,31,98,31,239,31,206,31,58,31,220,31,13,31,192,31,35,31,60,31,60,30,30,31,128,31,133,31,133,30,148,31,55,31,178,31,184,31,90,31,254,31,254,30,29,31,29,30,58,31,58,30,181,31,181,30,247,31,247,30,21,31,185,31,70,31,37,31,28,31,1,31,239,31,228,31,19,31,19,30,19,29,19,28,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
