-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_245 is
end project_tb_245;

architecture project_tb_arch_245 of project_tb_245 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (175,0,113,0,186,0,158,0,162,0,130,0,12,0,133,0,83,0,247,0,88,0,122,0,128,0,0,0,98,0,43,0,11,0,96,0,0,0,0,0,5,0,44,0,129,0,0,0,0,0,249,0,81,0,155,0,105,0,0,0,0,0,68,0,0,0,205,0,144,0,73,0,20,0,125,0,0,0,39,0,84,0,174,0,167,0,0,0,0,0,0,0,0,0,0,0,119,0,190,0,100,0,92,0,89,0,223,0,147,0,245,0,102,0,41,0,44,0,140,0,253,0,198,0,0,0,203,0,106,0,0,0,55,0,12,0,188,0,201,0,173,0,0,0,0,0,0,0,148,0,118,0,158,0,0,0,170,0,91,0,45,0,24,0,0,0,248,0,231,0,178,0,55,0,162,0,45,0,43,0,147,0,0,0,251,0,115,0,151,0,64,0,237,0,1,0,198,0,154,0,90,0,11,0,131,0,0,0,214,0,144,0,170,0,87,0,145,0,98,0,24,0,194,0,47,0,43,0,179,0,251,0,165,0,170,0,0,0,56,0,67,0,205,0,104,0,105,0,0,0,210,0,250,0,77,0,194,0,11,0,0,0,0,0,64,0,93,0,42,0,35,0,0,0,90,0,226,0,125,0,181,0,87,0,99,0,100,0,102,0,10,0,51,0,21,0,0,0,0,0,5,0,114,0,46,0,7,0,31,0,106,0,3,0,118,0,53,0,158,0,9,0,154,0,0,0,255,0,214,0,126,0,106,0,74,0,211,0,135,0,27,0,241,0,216,0,180,0,41,0,0,0,60,0,251,0,217,0,0,0,179,0,22,0,72,0,125,0,0,0,16,0,0,0,38,0,126,0,139,0,145,0,114,0,206,0,221,0,202,0,177,0,195,0,44,0,26,0,108,0,25,0,17,0,10,0,19,0,124,0,200,0,28,0,0,0,78,0,94,0,249,0,139,0,0,0,46,0,108,0,154,0,249,0,0,0,27,0,58,0,82,0,30,0,0,0,0,0,134,0,31,0,126,0,98,0,136,0,22,0,33,0,0,0,0,0,87,0,105,0,144,0,0,0,0,0,0,0,221,0,187,0,242,0,130,0,125,0,20,0,147,0,38,0,255,0,33,0,78,0,19,0,0,0,0,0,88,0,160,0,81,0,7,0,34,0,0,0,136,0,11,0,56,0,75,0,0,0,26,0,104,0,204,0,84,0,171,0,209,0,196,0,152,0,118,0,67,0,59,0,199,0,174,0,106,0,0,0,186,0,125,0,173,0,155,0,111,0,34,0,172,0,20,0,99,0,233,0,0,0,177,0,90,0,249,0,59,0,0,0,244,0,190,0,93,0,96,0,157,0,155,0,253,0,125,0,36,0,226,0,97,0,131,0,109,0,184,0,192,0,236,0,5,0,225,0,133,0,115,0,43,0,0,0,134,0,26,0,123,0,196,0,0,0,0,0,9,0,107,0,0,0,254,0,165,0,120,0,76,0,172,0,0,0,228,0,0,0,238,0,148,0,252,0,106,0,0,0,245,0,144,0,93,0,0,0,95,0,54,0,35,0,100,0,0,0,82,0,238,0,29,0,133,0,235,0,49,0,0,0,152,0,213,0,172,0,127,0,50,0,28,0,21,0,4,0,111,0,0,0,165,0,195,0,102,0,90,0,236,0,5,0,0,0,189,0,144,0,234,0,147,0,0,0,0,0,188,0,119,0,213,0,249,0,17,0,0,0,222,0,182,0,12,0,155,0,244,0,211,0,0,0,186,0,92,0,231,0,179,0,92,0,46,0,7,0,78,0,105,0,159,0,105,0,30,0,38,0,41,0,0,0,0,0,238,0,111,0,234,0,0,0,0,0,0,0,0,0,144,0,100,0,43,0,0,0,232,0,0,0,22,0,230,0,100,0,0,0,0,0,76,0,0,0,0,0,140,0,114,0,234,0,0,0,122,0,107,0,146,0,180,0,225,0,94,0,0,0,182,0,169,0,4,0,215,0,94,0,151,0,246,0,68,0,0,0,206,0,83,0,20,0,228,0,189,0,171,0,0,0,142,0,145,0,128,0,0,0,0,0,75,0,199,0,203,0,0,0,0,0,0,0,120,0,174,0,99,0,237,0,102,0,169,0,0,0,239,0,0,0,234,0,0,0,109,0,133,0,0,0,0,0,196,0,16,0,121,0,50,0,0,0,11,0,116,0,160,0,192,0,0,0,105,0,62,0,3,0,157,0,65,0,70,0,163,0,133,0,140,0,84,0,216,0,64,0,0,0,221,0,0,0,215,0,0,0,0,0,87,0,209,0,201,0,87,0,42,0,17,0,13,0,2,0,32,0,8,0,0,0,16,0,117,0,229,0,218,0,36,0,253,0,117,0,250,0,169,0,0,0,35,0,190,0,0,0,78,0,74,0,185,0,94,0,48,0,42,0,39,0,197,0,88,0,191,0,197,0,118,0,167,0,0,0,0,0,0,0,57,0,0,0,0,0,201,0,87,0,170,0,64,0,178,0,196,0,182,0,95,0,72,0,82,0,229,0,0,0,189,0,0,0,88,0,143,0,0,0,0,0,78,0,11,0,137,0,1,0,252,0,56,0,143,0,193,0,0,0,124,0,79,0,163,0,10,0,214,0,217,0,49,0,95,0,20,0,39,0,253,0,0,0,192,0,212,0,191,0,90,0,119,0,38,0,205,0,0,0,209,0,0,0,35,0,187,0,1,0,111,0,129,0,169,0,151,0,99,0,0,0,180,0,120,0,169,0,145,0,136,0,154,0,73,0,54,0,18,0,68,0,0,0,6,0,109,0,94,0,160,0,66,0,15,0,100,0,181,0,91,0,0,0,159,0,116,0,0,0,19,0,196,0,211,0,0,0,0,0,247,0,8,0,147,0,7,0,17,0,236,0,54,0,180,0,47,0,0,0,68,0,94,0,21,0,87,0,211,0,0,0,0,0,106,0,65,0,148,0,26,0,79,0,0,0,170,0,66,0,19,0,242,0,0,0,216,0,142,0,175,0,205,0,86,0,0,0,0,0,36,0,216,0,161,0,62,0,0,0,213,0,211,0,247,0,102,0,239,0,46,0,213,0,38,0,0,0,14,0,119,0,96,0,67,0,0,0,213,0,163,0,74,0,56,0,147,0,142,0,171,0,138,0,2,0,136,0,192,0,0,0,133,0,232,0,0,0,73,0,0,0,248,0,187,0,138,0,72,0,146,0,0,0,0,0,165,0,207,0,29,0,58,0,59,0,148,0,228,0,78,0,241,0,0,0,255,0,172,0,98,0,100,0,0,0,116,0,154,0,0,0,3,0,167,0,175,0,149,0,71,0,224,0,72,0,16,0,185,0,0,0,200,0,0,0,133,0,51,0,0,0,0,0,151,0,70,0,248,0,112,0,31,0,69,0,158,0,0,0,165,0,0,0,190,0,0,0,178,0,223,0,59,0,43,0,252,0,59,0,155,0,55,0,96,0,66,0,233,0,0,0,185,0,134,0,0,0,247,0,188,0,197,0,0,0,2,0,234,0,129,0,150,0,134,0,243,0,77,0,234,0,0,0,0,0,18,0,70,0,178,0,212,0,117,0,227,0,46,0,120,0,216,0,12,0,28,0,150,0,230,0,148,0,63,0,0,0,19,0,0,0,0,0,182,0,196,0,155,0,255,0,244,0,238,0,22,0,179,0,167,0,210,0,100,0,244,0,242,0,166,0,175,0,79,0,28,0,246,0,140,0,0,0,156,0,0,0,0,0,33,0,0,0,224,0,0,0,87,0,83,0,38,0,20,0,75,0,0,0,0,0,5,0,76,0,0,0,197,0,244,0,60,0,117,0,255,0,0,0,192,0,194,0,175,0,103,0,215,0,210,0,0,0,35,0,158,0,253,0,85,0,74,0,36,0,0,0,0,0,14,0,197,0,207,0,253,0,125,0,130,0,60,0,70,0,56,0,0,0,140,0,60,0,45,0,2,0,249,0,40,0,240,0,250,0,0,0,63,0,0,0,0,0,125,0,248,0,0,0,8,0,119,0,0,0,196,0,53,0,233,0,193,0,0,0,160,0,89,0,151,0,0,0,33,0,212,0,81,0,20,0,11,0,179,0,205,0,173,0,192,0,64,0,139,0,0,0,99,0,0,0,40,0,233,0,205,0,255,0,131,0,86,0,19,0,65,0,165,0,41,0,55,0,104,0,110,0,121,0,163,0,224,0,0,0,143,0,189,0,244,0,0,0,174,0,0,0,151,0,32,0,186,0,244,0,17,0,0,0,231,0,163,0,70,0,0,0,62,0,48,0,98,0,241,0,0,0,115,0,0,0,116,0,126,0,0,0,101,0,6,0,168,0,0,0,0,0,95,0,44,0,161,0,185,0,246,0,255,0,0,0);
signal scenario_full  : scenario_type := (175,31,113,31,186,31,158,31,162,31,130,31,12,31,133,31,83,31,247,31,88,31,122,31,128,31,128,30,98,31,43,31,11,31,96,31,96,30,96,29,5,31,44,31,129,31,129,30,129,29,249,31,81,31,155,31,105,31,105,30,105,29,68,31,68,30,205,31,144,31,73,31,20,31,125,31,125,30,39,31,84,31,174,31,167,31,167,30,167,29,167,28,167,27,167,26,119,31,190,31,100,31,92,31,89,31,223,31,147,31,245,31,102,31,41,31,44,31,140,31,253,31,198,31,198,30,203,31,106,31,106,30,55,31,12,31,188,31,201,31,173,31,173,30,173,29,173,28,148,31,118,31,158,31,158,30,170,31,91,31,45,31,24,31,24,30,248,31,231,31,178,31,55,31,162,31,45,31,43,31,147,31,147,30,251,31,115,31,151,31,64,31,237,31,1,31,198,31,154,31,90,31,11,31,131,31,131,30,214,31,144,31,170,31,87,31,145,31,98,31,24,31,194,31,47,31,43,31,179,31,251,31,165,31,170,31,170,30,56,31,67,31,205,31,104,31,105,31,105,30,210,31,250,31,77,31,194,31,11,31,11,30,11,29,64,31,93,31,42,31,35,31,35,30,90,31,226,31,125,31,181,31,87,31,99,31,100,31,102,31,10,31,51,31,21,31,21,30,21,29,5,31,114,31,46,31,7,31,31,31,106,31,3,31,118,31,53,31,158,31,9,31,154,31,154,30,255,31,214,31,126,31,106,31,74,31,211,31,135,31,27,31,241,31,216,31,180,31,41,31,41,30,60,31,251,31,217,31,217,30,179,31,22,31,72,31,125,31,125,30,16,31,16,30,38,31,126,31,139,31,145,31,114,31,206,31,221,31,202,31,177,31,195,31,44,31,26,31,108,31,25,31,17,31,10,31,19,31,124,31,200,31,28,31,28,30,78,31,94,31,249,31,139,31,139,30,46,31,108,31,154,31,249,31,249,30,27,31,58,31,82,31,30,31,30,30,30,29,134,31,31,31,126,31,98,31,136,31,22,31,33,31,33,30,33,29,87,31,105,31,144,31,144,30,144,29,144,28,221,31,187,31,242,31,130,31,125,31,20,31,147,31,38,31,255,31,33,31,78,31,19,31,19,30,19,29,88,31,160,31,81,31,7,31,34,31,34,30,136,31,11,31,56,31,75,31,75,30,26,31,104,31,204,31,84,31,171,31,209,31,196,31,152,31,118,31,67,31,59,31,199,31,174,31,106,31,106,30,186,31,125,31,173,31,155,31,111,31,34,31,172,31,20,31,99,31,233,31,233,30,177,31,90,31,249,31,59,31,59,30,244,31,190,31,93,31,96,31,157,31,155,31,253,31,125,31,36,31,226,31,97,31,131,31,109,31,184,31,192,31,236,31,5,31,225,31,133,31,115,31,43,31,43,30,134,31,26,31,123,31,196,31,196,30,196,29,9,31,107,31,107,30,254,31,165,31,120,31,76,31,172,31,172,30,228,31,228,30,238,31,148,31,252,31,106,31,106,30,245,31,144,31,93,31,93,30,95,31,54,31,35,31,100,31,100,30,82,31,238,31,29,31,133,31,235,31,49,31,49,30,152,31,213,31,172,31,127,31,50,31,28,31,21,31,4,31,111,31,111,30,165,31,195,31,102,31,90,31,236,31,5,31,5,30,189,31,144,31,234,31,147,31,147,30,147,29,188,31,119,31,213,31,249,31,17,31,17,30,222,31,182,31,12,31,155,31,244,31,211,31,211,30,186,31,92,31,231,31,179,31,92,31,46,31,7,31,78,31,105,31,159,31,105,31,30,31,38,31,41,31,41,30,41,29,238,31,111,31,234,31,234,30,234,29,234,28,234,27,144,31,100,31,43,31,43,30,232,31,232,30,22,31,230,31,100,31,100,30,100,29,76,31,76,30,76,29,140,31,114,31,234,31,234,30,122,31,107,31,146,31,180,31,225,31,94,31,94,30,182,31,169,31,4,31,215,31,94,31,151,31,246,31,68,31,68,30,206,31,83,31,20,31,228,31,189,31,171,31,171,30,142,31,145,31,128,31,128,30,128,29,75,31,199,31,203,31,203,30,203,29,203,28,120,31,174,31,99,31,237,31,102,31,169,31,169,30,239,31,239,30,234,31,234,30,109,31,133,31,133,30,133,29,196,31,16,31,121,31,50,31,50,30,11,31,116,31,160,31,192,31,192,30,105,31,62,31,3,31,157,31,65,31,70,31,163,31,133,31,140,31,84,31,216,31,64,31,64,30,221,31,221,30,215,31,215,30,215,29,87,31,209,31,201,31,87,31,42,31,17,31,13,31,2,31,32,31,8,31,8,30,16,31,117,31,229,31,218,31,36,31,253,31,117,31,250,31,169,31,169,30,35,31,190,31,190,30,78,31,74,31,185,31,94,31,48,31,42,31,39,31,197,31,88,31,191,31,197,31,118,31,167,31,167,30,167,29,167,28,57,31,57,30,57,29,201,31,87,31,170,31,64,31,178,31,196,31,182,31,95,31,72,31,82,31,229,31,229,30,189,31,189,30,88,31,143,31,143,30,143,29,78,31,11,31,137,31,1,31,252,31,56,31,143,31,193,31,193,30,124,31,79,31,163,31,10,31,214,31,217,31,49,31,95,31,20,31,39,31,253,31,253,30,192,31,212,31,191,31,90,31,119,31,38,31,205,31,205,30,209,31,209,30,35,31,187,31,1,31,111,31,129,31,169,31,151,31,99,31,99,30,180,31,120,31,169,31,145,31,136,31,154,31,73,31,54,31,18,31,68,31,68,30,6,31,109,31,94,31,160,31,66,31,15,31,100,31,181,31,91,31,91,30,159,31,116,31,116,30,19,31,196,31,211,31,211,30,211,29,247,31,8,31,147,31,7,31,17,31,236,31,54,31,180,31,47,31,47,30,68,31,94,31,21,31,87,31,211,31,211,30,211,29,106,31,65,31,148,31,26,31,79,31,79,30,170,31,66,31,19,31,242,31,242,30,216,31,142,31,175,31,205,31,86,31,86,30,86,29,36,31,216,31,161,31,62,31,62,30,213,31,211,31,247,31,102,31,239,31,46,31,213,31,38,31,38,30,14,31,119,31,96,31,67,31,67,30,213,31,163,31,74,31,56,31,147,31,142,31,171,31,138,31,2,31,136,31,192,31,192,30,133,31,232,31,232,30,73,31,73,30,248,31,187,31,138,31,72,31,146,31,146,30,146,29,165,31,207,31,29,31,58,31,59,31,148,31,228,31,78,31,241,31,241,30,255,31,172,31,98,31,100,31,100,30,116,31,154,31,154,30,3,31,167,31,175,31,149,31,71,31,224,31,72,31,16,31,185,31,185,30,200,31,200,30,133,31,51,31,51,30,51,29,151,31,70,31,248,31,112,31,31,31,69,31,158,31,158,30,165,31,165,30,190,31,190,30,178,31,223,31,59,31,43,31,252,31,59,31,155,31,55,31,96,31,66,31,233,31,233,30,185,31,134,31,134,30,247,31,188,31,197,31,197,30,2,31,234,31,129,31,150,31,134,31,243,31,77,31,234,31,234,30,234,29,18,31,70,31,178,31,212,31,117,31,227,31,46,31,120,31,216,31,12,31,28,31,150,31,230,31,148,31,63,31,63,30,19,31,19,30,19,29,182,31,196,31,155,31,255,31,244,31,238,31,22,31,179,31,167,31,210,31,100,31,244,31,242,31,166,31,175,31,79,31,28,31,246,31,140,31,140,30,156,31,156,30,156,29,33,31,33,30,224,31,224,30,87,31,83,31,38,31,20,31,75,31,75,30,75,29,5,31,76,31,76,30,197,31,244,31,60,31,117,31,255,31,255,30,192,31,194,31,175,31,103,31,215,31,210,31,210,30,35,31,158,31,253,31,85,31,74,31,36,31,36,30,36,29,14,31,197,31,207,31,253,31,125,31,130,31,60,31,70,31,56,31,56,30,140,31,60,31,45,31,2,31,249,31,40,31,240,31,250,31,250,30,63,31,63,30,63,29,125,31,248,31,248,30,8,31,119,31,119,30,196,31,53,31,233,31,193,31,193,30,160,31,89,31,151,31,151,30,33,31,212,31,81,31,20,31,11,31,179,31,205,31,173,31,192,31,64,31,139,31,139,30,99,31,99,30,40,31,233,31,205,31,255,31,131,31,86,31,19,31,65,31,165,31,41,31,55,31,104,31,110,31,121,31,163,31,224,31,224,30,143,31,189,31,244,31,244,30,174,31,174,30,151,31,32,31,186,31,244,31,17,31,17,30,231,31,163,31,70,31,70,30,62,31,48,31,98,31,241,31,241,30,115,31,115,30,116,31,126,31,126,30,101,31,6,31,168,31,168,30,168,29,95,31,44,31,161,31,185,31,246,31,255,31,255,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
