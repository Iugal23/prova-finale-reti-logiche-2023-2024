-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 373;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (210,0,171,0,228,0,0,0,0,0,214,0,0,0,93,0,0,0,0,0,124,0,91,0,138,0,28,0,197,0,147,0,88,0,218,0,0,0,128,0,170,0,113,0,45,0,0,0,151,0,123,0,102,0,52,0,50,0,165,0,0,0,2,0,0,0,113,0,63,0,69,0,0,0,4,0,224,0,210,0,132,0,196,0,34,0,252,0,196,0,137,0,192,0,85,0,243,0,236,0,237,0,0,0,76,0,0,0,0,0,81,0,85,0,142,0,0,0,143,0,36,0,38,0,143,0,113,0,0,0,219,0,17,0,67,0,255,0,0,0,0,0,18,0,227,0,97,0,253,0,0,0,0,0,183,0,86,0,220,0,0,0,0,0,146,0,48,0,128,0,0,0,7,0,47,0,170,0,38,0,202,0,0,0,0,0,110,0,207,0,162,0,90,0,239,0,36,0,88,0,215,0,111,0,1,0,0,0,241,0,227,0,21,0,0,0,211,0,19,0,166,0,23,0,199,0,243,0,116,0,7,0,167,0,105,0,88,0,100,0,0,0,0,0,92,0,163,0,9,0,0,0,0,0,0,0,123,0,0,0,191,0,89,0,82,0,251,0,202,0,193,0,0,0,25,0,110,0,0,0,0,0,146,0,30,0,156,0,7,0,200,0,166,0,152,0,56,0,197,0,133,0,176,0,123,0,135,0,202,0,171,0,0,0,97,0,143,0,151,0,198,0,74,0,122,0,167,0,24,0,182,0,18,0,54,0,40,0,170,0,228,0,8,0,217,0,52,0,0,0,140,0,231,0,0,0,63,0,145,0,136,0,202,0,129,0,169,0,147,0,189,0,175,0,100,0,3,0,157,0,139,0,1,0,139,0,0,0,166,0,239,0,0,0,183,0,66,0,241,0,159,0,115,0,0,0,31,0,0,0,0,0,0,0,208,0,130,0,85,0,255,0,236,0,9,0,0,0,83,0,56,0,10,0,158,0,114,0,0,0,0,0,73,0,113,0,138,0,0,0,129,0,99,0,142,0,65,0,0,0,88,0,0,0,102,0,206,0,0,0,110,0,113,0,163,0,181,0,97,0,88,0,0,0,8,0,214,0,0,0,142,0,225,0,98,0,179,0,0,0,3,0,176,0,118,0,0,0,142,0,32,0,0,0,62,0,0,0,212,0,6,0,209,0,0,0,140,0,108,0,237,0,76,0,0,0,89,0,84,0,5,0,0,0,65,0,61,0,17,0,122,0,73,0,45,0,0,0,167,0,3,0,0,0,57,0,240,0,244,0,92,0,116,0,0,0,251,0,107,0,0,0,116,0,135,0,0,0,0,0,47,0,200,0,222,0,226,0,179,0,127,0,255,0,201,0,152,0,111,0,0,0,0,0,107,0,113,0,242,0,0,0,54,0,15,0,17,0,56,0,49,0,152,0,233,0,10,0,246,0,254,0,0,0,144,0,222,0,68,0,33,0,72,0,230,0,0,0,0,0,50,0,184,0,176,0,0,0,78,0,71,0,170,0,147,0,223,0,61,0,26,0,49,0,12,0,108,0,114,0,16,0,1,0,133,0,207,0,32,0,239,0,211,0,79,0,103,0,21,0,0,0,177,0,0,0,132,0,0,0,151,0,115,0,55,0,158,0,14,0,8,0,0,0,13,0,144,0,226,0,16,0,107,0,219,0);
signal scenario_full  : scenario_type := (210,31,171,31,228,31,228,30,228,29,214,31,214,30,93,31,93,30,93,29,124,31,91,31,138,31,28,31,197,31,147,31,88,31,218,31,218,30,128,31,170,31,113,31,45,31,45,30,151,31,123,31,102,31,52,31,50,31,165,31,165,30,2,31,2,30,113,31,63,31,69,31,69,30,4,31,224,31,210,31,132,31,196,31,34,31,252,31,196,31,137,31,192,31,85,31,243,31,236,31,237,31,237,30,76,31,76,30,76,29,81,31,85,31,142,31,142,30,143,31,36,31,38,31,143,31,113,31,113,30,219,31,17,31,67,31,255,31,255,30,255,29,18,31,227,31,97,31,253,31,253,30,253,29,183,31,86,31,220,31,220,30,220,29,146,31,48,31,128,31,128,30,7,31,47,31,170,31,38,31,202,31,202,30,202,29,110,31,207,31,162,31,90,31,239,31,36,31,88,31,215,31,111,31,1,31,1,30,241,31,227,31,21,31,21,30,211,31,19,31,166,31,23,31,199,31,243,31,116,31,7,31,167,31,105,31,88,31,100,31,100,30,100,29,92,31,163,31,9,31,9,30,9,29,9,28,123,31,123,30,191,31,89,31,82,31,251,31,202,31,193,31,193,30,25,31,110,31,110,30,110,29,146,31,30,31,156,31,7,31,200,31,166,31,152,31,56,31,197,31,133,31,176,31,123,31,135,31,202,31,171,31,171,30,97,31,143,31,151,31,198,31,74,31,122,31,167,31,24,31,182,31,18,31,54,31,40,31,170,31,228,31,8,31,217,31,52,31,52,30,140,31,231,31,231,30,63,31,145,31,136,31,202,31,129,31,169,31,147,31,189,31,175,31,100,31,3,31,157,31,139,31,1,31,139,31,139,30,166,31,239,31,239,30,183,31,66,31,241,31,159,31,115,31,115,30,31,31,31,30,31,29,31,28,208,31,130,31,85,31,255,31,236,31,9,31,9,30,83,31,56,31,10,31,158,31,114,31,114,30,114,29,73,31,113,31,138,31,138,30,129,31,99,31,142,31,65,31,65,30,88,31,88,30,102,31,206,31,206,30,110,31,113,31,163,31,181,31,97,31,88,31,88,30,8,31,214,31,214,30,142,31,225,31,98,31,179,31,179,30,3,31,176,31,118,31,118,30,142,31,32,31,32,30,62,31,62,30,212,31,6,31,209,31,209,30,140,31,108,31,237,31,76,31,76,30,89,31,84,31,5,31,5,30,65,31,61,31,17,31,122,31,73,31,45,31,45,30,167,31,3,31,3,30,57,31,240,31,244,31,92,31,116,31,116,30,251,31,107,31,107,30,116,31,135,31,135,30,135,29,47,31,200,31,222,31,226,31,179,31,127,31,255,31,201,31,152,31,111,31,111,30,111,29,107,31,113,31,242,31,242,30,54,31,15,31,17,31,56,31,49,31,152,31,233,31,10,31,246,31,254,31,254,30,144,31,222,31,68,31,33,31,72,31,230,31,230,30,230,29,50,31,184,31,176,31,176,30,78,31,71,31,170,31,147,31,223,31,61,31,26,31,49,31,12,31,108,31,114,31,16,31,1,31,133,31,207,31,32,31,239,31,211,31,79,31,103,31,21,31,21,30,177,31,177,30,132,31,132,30,151,31,115,31,55,31,158,31,14,31,8,31,8,30,13,31,144,31,226,31,16,31,107,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
