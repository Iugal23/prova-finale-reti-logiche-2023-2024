-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 668;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (111,0,5,0,29,0,64,0,100,0,163,0,216,0,147,0,27,0,0,0,133,0,151,0,226,0,7,0,48,0,176,0,39,0,249,0,125,0,24,0,160,0,0,0,212,0,207,0,178,0,79,0,197,0,77,0,8,0,0,0,213,0,3,0,175,0,0,0,120,0,0,0,0,0,131,0,66,0,180,0,247,0,2,0,115,0,182,0,160,0,96,0,0,0,162,0,110,0,74,0,0,0,228,0,176,0,85,0,246,0,165,0,0,0,14,0,186,0,65,0,0,0,241,0,83,0,38,0,128,0,64,0,62,0,104,0,179,0,187,0,0,0,189,0,100,0,107,0,122,0,179,0,115,0,209,0,0,0,240,0,0,0,0,0,26,0,10,0,193,0,89,0,172,0,83,0,37,0,175,0,0,0,106,0,151,0,0,0,0,0,60,0,106,0,18,0,0,0,0,0,0,0,93,0,247,0,55,0,43,0,10,0,134,0,17,0,166,0,6,0,0,0,255,0,0,0,72,0,90,0,0,0,220,0,19,0,67,0,46,0,74,0,22,0,0,0,129,0,0,0,26,0,7,0,0,0,87,0,118,0,231,0,62,0,55,0,197,0,71,0,251,0,183,0,22,0,0,0,128,0,0,0,0,0,116,0,109,0,230,0,178,0,24,0,96,0,148,0,140,0,0,0,0,0,132,0,56,0,164,0,55,0,0,0,149,0,109,0,203,0,0,0,119,0,228,0,121,0,191,0,0,0,192,0,95,0,16,0,40,0,8,0,0,0,7,0,198,0,57,0,68,0,114,0,190,0,0,0,124,0,214,0,137,0,58,0,33,0,88,0,255,0,79,0,0,0,158,0,0,0,135,0,204,0,243,0,35,0,54,0,27,0,0,0,8,0,171,0,127,0,0,0,0,0,175,0,9,0,173,0,58,0,210,0,0,0,228,0,231,0,0,0,137,0,46,0,142,0,230,0,52,0,156,0,44,0,72,0,170,0,245,0,188,0,156,0,142,0,0,0,161,0,136,0,215,0,251,0,137,0,55,0,32,0,174,0,1,0,64,0,166,0,0,0,56,0,109,0,64,0,18,0,255,0,14,0,139,0,203,0,0,0,244,0,184,0,124,0,0,0,205,0,130,0,163,0,2,0,140,0,10,0,0,0,61,0,0,0,0,0,51,0,60,0,0,0,170,0,183,0,184,0,7,0,172,0,243,0,227,0,145,0,0,0,199,0,0,0,93,0,124,0,116,0,55,0,45,0,62,0,52,0,8,0,110,0,0,0,173,0,196,0,0,0,0,0,37,0,25,0,0,0,132,0,209,0,10,0,71,0,0,0,153,0,0,0,237,0,0,0,147,0,232,0,117,0,214,0,0,0,0,0,0,0,146,0,229,0,78,0,98,0,179,0,0,0,95,0,79,0,0,0,123,0,73,0,90,0,16,0,29,0,101,0,188,0,42,0,234,0,195,0,246,0,255,0,0,0,0,0,184,0,158,0,241,0,173,0,41,0,63,0,141,0,186,0,192,0,109,0,246,0,115,0,75,0,114,0,155,0,234,0,20,0,34,0,0,0,121,0,44,0,129,0,0,0,0,0,43,0,3,0,12,0,189,0,124,0,128,0,116,0,42,0,0,0,33,0,166,0,20,0,0,0,39,0,182,0,238,0,83,0,141,0,223,0,0,0,222,0,136,0,156,0,58,0,0,0,0,0,66,0,0,0,12,0,194,0,9,0,0,0,0,0,0,0,0,0,220,0,221,0,191,0,210,0,187,0,244,0,0,0,65,0,55,0,75,0,0,0,160,0,14,0,128,0,123,0,0,0,163,0,0,0,0,0,59,0,141,0,0,0,102,0,113,0,213,0,222,0,57,0,233,0,122,0,92,0,150,0,212,0,250,0,45,0,117,0,223,0,218,0,25,0,106,0,135,0,218,0,109,0,184,0,84,0,104,0,232,0,39,0,155,0,0,0,193,0,117,0,0,0,239,0,72,0,135,0,36,0,254,0,242,0,73,0,0,0,221,0,0,0,13,0,132,0,187,0,149,0,71,0,169,0,94,0,0,0,136,0,163,0,22,0,68,0,244,0,211,0,51,0,37,0,178,0,71,0,0,0,0,0,14,0,218,0,213,0,0,0,0,0,132,0,0,0,0,0,136,0,72,0,126,0,187,0,50,0,0,0,162,0,56,0,5,0,0,0,0,0,235,0,6,0,0,0,66,0,0,0,12,0,84,0,68,0,238,0,1,0,162,0,0,0,0,0,10,0,167,0,218,0,42,0,43,0,74,0,13,0,8,0,137,0,248,0,7,0,214,0,171,0,0,0,167,0,176,0,205,0,82,0,0,0,174,0,101,0,32,0,221,0,200,0,42,0,163,0,93,0,244,0,221,0,243,0,180,0,44,0,107,0,217,0,186,0,170,0,10,0,33,0,152,0,101,0,249,0,25,0,193,0,73,0,46,0,0,0,0,0,0,0,46,0,230,0,0,0,155,0,88,0,44,0,253,0,184,0,177,0,134,0,102,0,0,0,82,0,160,0,191,0,73,0,215,0,0,0,208,0,252,0,0,0,250,0,89,0,138,0,228,0,239,0,36,0,168,0,64,0,0,0,146,0,69,0,8,0,53,0,147,0,112,0,226,0,183,0,171,0,8,0,92,0,0,0,56,0,57,0,0,0,0,0,78,0,0,0,33,0,178,0,56,0,198,0,153,0,83,0,0,0,42,0,122,0,125,0,0,0,59,0,156,0,0,0,103,0,0,0,187,0,58,0,0,0,190,0,0,0,0,0,115,0,138,0,0,0,219,0,0,0,0,0,0,0,112,0,234,0,0,0,130,0,33,0,197,0,236,0,154,0,0,0,223,0,128,0,0,0,242,0,157,0,0,0,166,0,0,0,172,0,255,0,98,0,78,0,108,0,146,0,119,0,83,0,124,0,0,0,0,0,0,0,126,0,0,0,99,0,2,0,110,0,177,0,0,0,64,0,12,0,138,0,172,0);
signal scenario_full  : scenario_type := (111,31,5,31,29,31,64,31,100,31,163,31,216,31,147,31,27,31,27,30,133,31,151,31,226,31,7,31,48,31,176,31,39,31,249,31,125,31,24,31,160,31,160,30,212,31,207,31,178,31,79,31,197,31,77,31,8,31,8,30,213,31,3,31,175,31,175,30,120,31,120,30,120,29,131,31,66,31,180,31,247,31,2,31,115,31,182,31,160,31,96,31,96,30,162,31,110,31,74,31,74,30,228,31,176,31,85,31,246,31,165,31,165,30,14,31,186,31,65,31,65,30,241,31,83,31,38,31,128,31,64,31,62,31,104,31,179,31,187,31,187,30,189,31,100,31,107,31,122,31,179,31,115,31,209,31,209,30,240,31,240,30,240,29,26,31,10,31,193,31,89,31,172,31,83,31,37,31,175,31,175,30,106,31,151,31,151,30,151,29,60,31,106,31,18,31,18,30,18,29,18,28,93,31,247,31,55,31,43,31,10,31,134,31,17,31,166,31,6,31,6,30,255,31,255,30,72,31,90,31,90,30,220,31,19,31,67,31,46,31,74,31,22,31,22,30,129,31,129,30,26,31,7,31,7,30,87,31,118,31,231,31,62,31,55,31,197,31,71,31,251,31,183,31,22,31,22,30,128,31,128,30,128,29,116,31,109,31,230,31,178,31,24,31,96,31,148,31,140,31,140,30,140,29,132,31,56,31,164,31,55,31,55,30,149,31,109,31,203,31,203,30,119,31,228,31,121,31,191,31,191,30,192,31,95,31,16,31,40,31,8,31,8,30,7,31,198,31,57,31,68,31,114,31,190,31,190,30,124,31,214,31,137,31,58,31,33,31,88,31,255,31,79,31,79,30,158,31,158,30,135,31,204,31,243,31,35,31,54,31,27,31,27,30,8,31,171,31,127,31,127,30,127,29,175,31,9,31,173,31,58,31,210,31,210,30,228,31,231,31,231,30,137,31,46,31,142,31,230,31,52,31,156,31,44,31,72,31,170,31,245,31,188,31,156,31,142,31,142,30,161,31,136,31,215,31,251,31,137,31,55,31,32,31,174,31,1,31,64,31,166,31,166,30,56,31,109,31,64,31,18,31,255,31,14,31,139,31,203,31,203,30,244,31,184,31,124,31,124,30,205,31,130,31,163,31,2,31,140,31,10,31,10,30,61,31,61,30,61,29,51,31,60,31,60,30,170,31,183,31,184,31,7,31,172,31,243,31,227,31,145,31,145,30,199,31,199,30,93,31,124,31,116,31,55,31,45,31,62,31,52,31,8,31,110,31,110,30,173,31,196,31,196,30,196,29,37,31,25,31,25,30,132,31,209,31,10,31,71,31,71,30,153,31,153,30,237,31,237,30,147,31,232,31,117,31,214,31,214,30,214,29,214,28,146,31,229,31,78,31,98,31,179,31,179,30,95,31,79,31,79,30,123,31,73,31,90,31,16,31,29,31,101,31,188,31,42,31,234,31,195,31,246,31,255,31,255,30,255,29,184,31,158,31,241,31,173,31,41,31,63,31,141,31,186,31,192,31,109,31,246,31,115,31,75,31,114,31,155,31,234,31,20,31,34,31,34,30,121,31,44,31,129,31,129,30,129,29,43,31,3,31,12,31,189,31,124,31,128,31,116,31,42,31,42,30,33,31,166,31,20,31,20,30,39,31,182,31,238,31,83,31,141,31,223,31,223,30,222,31,136,31,156,31,58,31,58,30,58,29,66,31,66,30,12,31,194,31,9,31,9,30,9,29,9,28,9,27,220,31,221,31,191,31,210,31,187,31,244,31,244,30,65,31,55,31,75,31,75,30,160,31,14,31,128,31,123,31,123,30,163,31,163,30,163,29,59,31,141,31,141,30,102,31,113,31,213,31,222,31,57,31,233,31,122,31,92,31,150,31,212,31,250,31,45,31,117,31,223,31,218,31,25,31,106,31,135,31,218,31,109,31,184,31,84,31,104,31,232,31,39,31,155,31,155,30,193,31,117,31,117,30,239,31,72,31,135,31,36,31,254,31,242,31,73,31,73,30,221,31,221,30,13,31,132,31,187,31,149,31,71,31,169,31,94,31,94,30,136,31,163,31,22,31,68,31,244,31,211,31,51,31,37,31,178,31,71,31,71,30,71,29,14,31,218,31,213,31,213,30,213,29,132,31,132,30,132,29,136,31,72,31,126,31,187,31,50,31,50,30,162,31,56,31,5,31,5,30,5,29,235,31,6,31,6,30,66,31,66,30,12,31,84,31,68,31,238,31,1,31,162,31,162,30,162,29,10,31,167,31,218,31,42,31,43,31,74,31,13,31,8,31,137,31,248,31,7,31,214,31,171,31,171,30,167,31,176,31,205,31,82,31,82,30,174,31,101,31,32,31,221,31,200,31,42,31,163,31,93,31,244,31,221,31,243,31,180,31,44,31,107,31,217,31,186,31,170,31,10,31,33,31,152,31,101,31,249,31,25,31,193,31,73,31,46,31,46,30,46,29,46,28,46,31,230,31,230,30,155,31,88,31,44,31,253,31,184,31,177,31,134,31,102,31,102,30,82,31,160,31,191,31,73,31,215,31,215,30,208,31,252,31,252,30,250,31,89,31,138,31,228,31,239,31,36,31,168,31,64,31,64,30,146,31,69,31,8,31,53,31,147,31,112,31,226,31,183,31,171,31,8,31,92,31,92,30,56,31,57,31,57,30,57,29,78,31,78,30,33,31,178,31,56,31,198,31,153,31,83,31,83,30,42,31,122,31,125,31,125,30,59,31,156,31,156,30,103,31,103,30,187,31,58,31,58,30,190,31,190,30,190,29,115,31,138,31,138,30,219,31,219,30,219,29,219,28,112,31,234,31,234,30,130,31,33,31,197,31,236,31,154,31,154,30,223,31,128,31,128,30,242,31,157,31,157,30,166,31,166,30,172,31,255,31,98,31,78,31,108,31,146,31,119,31,83,31,124,31,124,30,124,29,124,28,126,31,126,30,99,31,2,31,110,31,177,31,177,30,64,31,12,31,138,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
