-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_819 is
end project_tb_819;

architecture project_tb_arch_819 of project_tb_819 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 830;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (208,0,194,0,0,0,0,0,175,0,25,0,41,0,0,0,118,0,134,0,77,0,240,0,0,0,6,0,0,0,219,0,133,0,20,0,0,0,144,0,0,0,25,0,147,0,47,0,179,0,0,0,62,0,151,0,205,0,0,0,174,0,49,0,12,0,0,0,112,0,203,0,20,0,0,0,0,0,169,0,0,0,0,0,231,0,27,0,164,0,152,0,194,0,50,0,96,0,233,0,224,0,180,0,0,0,240,0,252,0,229,0,53,0,224,0,0,0,6,0,35,0,159,0,48,0,18,0,67,0,91,0,128,0,0,0,150,0,238,0,241,0,0,0,107,0,62,0,223,0,84,0,93,0,108,0,31,0,146,0,217,0,83,0,73,0,60,0,37,0,218,0,183,0,211,0,99,0,0,0,204,0,95,0,0,0,0,0,107,0,25,0,233,0,119,0,54,0,215,0,22,0,0,0,57,0,0,0,189,0,185,0,181,0,219,0,156,0,70,0,0,0,111,0,187,0,250,0,153,0,57,0,206,0,213,0,0,0,101,0,0,0,63,0,78,0,180,0,65,0,27,0,0,0,254,0,21,0,178,0,237,0,84,0,28,0,90,0,6,0,45,0,250,0,79,0,141,0,198,0,127,0,8,0,0,0,0,0,213,0,138,0,0,0,50,0,220,0,0,0,49,0,40,0,82,0,138,0,7,0,35,0,69,0,0,0,90,0,186,0,61,0,18,0,231,0,0,0,143,0,239,0,1,0,221,0,105,0,24,0,86,0,0,0,254,0,249,0,156,0,34,0,19,0,134,0,133,0,101,0,222,0,0,0,35,0,226,0,28,0,164,0,49,0,157,0,0,0,149,0,76,0,0,0,0,0,0,0,24,0,132,0,100,0,210,0,176,0,239,0,66,0,242,0,200,0,131,0,53,0,49,0,26,0,105,0,140,0,87,0,133,0,29,0,105,0,191,0,212,0,25,0,0,0,185,0,0,0,53,0,3,0,7,0,14,0,0,0,219,0,221,0,19,0,158,0,175,0,28,0,95,0,85,0,0,0,142,0,198,0,0,0,0,0,220,0,23,0,77,0,81,0,216,0,167,0,55,0,240,0,124,0,122,0,42,0,229,0,98,0,65,0,194,0,0,0,142,0,92,0,0,0,0,0,96,0,11,0,149,0,35,0,115,0,0,0,117,0,0,0,0,0,175,0,81,0,61,0,207,0,58,0,0,0,29,0,110,0,190,0,155,0,0,0,0,0,0,0,141,0,0,0,101,0,250,0,25,0,84,0,230,0,233,0,0,0,106,0,0,0,36,0,32,0,113,0,251,0,136,0,0,0,155,0,201,0,156,0,15,0,67,0,116,0,56,0,0,0,0,0,206,0,69,0,111,0,87,0,252,0,246,0,200,0,194,0,0,0,105,0,194,0,38,0,1,0,117,0,0,0,225,0,243,0,227,0,39,0,0,0,178,0,124,0,25,0,160,0,0,0,213,0,95,0,72,0,68,0,148,0,116,0,0,0,104,0,253,0,170,0,0,0,97,0,63,0,0,0,42,0,83,0,80,0,190,0,30,0,72,0,115,0,89,0,89,0,114,0,0,0,231,0,130,0,197,0,0,0,30,0,145,0,14,0,155,0,172,0,0,0,211,0,191,0,96,0,26,0,72,0,0,0,84,0,13,0,0,0,174,0,0,0,5,0,142,0,163,0,0,0,160,0,30,0,61,0,0,0,120,0,94,0,63,0,0,0,72,0,109,0,131,0,116,0,105,0,156,0,7,0,55,0,19,0,95,0,216,0,0,0,245,0,82,0,7,0,174,0,197,0,179,0,136,0,128,0,170,0,89,0,178,0,80,0,241,0,32,0,165,0,18,0,0,0,0,0,24,0,200,0,0,0,0,0,22,0,90,0,169,0,69,0,205,0,30,0,7,0,76,0,129,0,87,0,41,0,170,0,150,0,208,0,233,0,57,0,171,0,229,0,0,0,28,0,117,0,0,0,101,0,143,0,137,0,222,0,220,0,164,0,56,0,0,0,74,0,0,0,254,0,140,0,241,0,86,0,193,0,98,0,0,0,0,0,82,0,171,0,205,0,216,0,77,0,0,0,165,0,74,0,42,0,0,0,127,0,181,0,178,0,48,0,195,0,87,0,0,0,0,0,170,0,99,0,95,0,164,0,123,0,61,0,85,0,111,0,178,0,126,0,192,0,58,0,36,0,160,0,0,0,32,0,180,0,0,0,95,0,221,0,219,0,115,0,0,0,190,0,0,0,0,0,72,0,0,0,0,0,223,0,254,0,175,0,139,0,180,0,0,0,57,0,196,0,0,0,0,0,97,0,193,0,193,0,0,0,161,0,204,0,150,0,253,0,171,0,50,0,103,0,123,0,10,0,210,0,201,0,0,0,28,0,187,0,155,0,105,0,122,0,160,0,240,0,63,0,232,0,35,0,210,0,46,0,39,0,7,0,179,0,176,0,97,0,87,0,23,0,0,0,20,0,146,0,0,0,6,0,67,0,242,0,12,0,2,0,90,0,150,0,0,0,0,0,148,0,79,0,40,0,44,0,254,0,0,0,100,0,205,0,68,0,0,0,76,0,62,0,190,0,12,0,24,0,0,0,231,0,186,0,33,0,117,0,197,0,193,0,0,0,7,0,190,0,40,0,238,0,131,0,57,0,55,0,226,0,96,0,194,0,117,0,239,0,0,0,58,0,145,0,162,0,99,0,118,0,161,0,209,0,36,0,54,0,0,0,0,0,69,0,216,0,240,0,166,0,53,0,0,0,0,0,73,0,162,0,130,0,132,0,50,0,0,0,0,0,246,0,115,0,16,0,55,0,189,0,0,0,0,0,85,0,0,0,182,0,129,0,127,0,202,0,135,0,144,0,85,0,59,0,246,0,212,0,0,0,46,0,37,0,156,0,250,0,0,0,177,0,0,0,121,0,14,0,0,0,201,0,0,0,85,0,236,0,35,0,69,0,29,0,28,0,200,0,0,0,49,0,255,0,90,0,233,0,84,0,173,0,147,0,152,0,0,0,144,0,199,0,73,0,184,0,190,0,221,0,162,0,25,0,132,0,246,0,103,0,93,0,160,0,0,0,211,0,0,0,93,0,116,0,87,0,0,0,95,0,122,0,111,0,200,0,137,0,214,0,100,0,249,0,169,0,0,0,47,0,110,0,210,0,143,0,156,0,0,0,0,0,0,0,218,0,233,0,37,0,0,0,150,0,45,0,91,0,246,0,187,0,35,0,171,0,0,0,222,0,158,0,94,0,132,0,100,0,0,0,77,0,0,0,239,0,0,0,38,0,126,0,0,0,164,0,130,0,0,0,0,0,22,0,93,0,100,0,188,0,55,0,0,0,120,0,2,0,14,0,66,0,3,0,229,0,93,0,162,0,0,0,44,0,0,0,192,0,40,0,0,0,92,0,125,0,151,0,144,0,0,0,245,0,79,0,135,0,221,0,0,0,38,0,155,0,56,0,140,0,0,0,163,0,0,0,101,0,245,0,238,0,161,0,19,0,132,0,77,0,192,0,187,0,252,0,221,0,68,0,212,0,163,0,48,0,0,0,132,0,19,0,0,0,234,0,0,0,185,0,195,0,97,0,169,0,98,0,224,0,12,0,0,0,214,0,133,0,0,0,130,0,205,0,50,0,89,0,242,0,0,0,0,0,177,0,3,0,106,0,106,0,48,0,241,0,131,0,239,0,117,0,168,0);
signal scenario_full  : scenario_type := (208,31,194,31,194,30,194,29,175,31,25,31,41,31,41,30,118,31,134,31,77,31,240,31,240,30,6,31,6,30,219,31,133,31,20,31,20,30,144,31,144,30,25,31,147,31,47,31,179,31,179,30,62,31,151,31,205,31,205,30,174,31,49,31,12,31,12,30,112,31,203,31,20,31,20,30,20,29,169,31,169,30,169,29,231,31,27,31,164,31,152,31,194,31,50,31,96,31,233,31,224,31,180,31,180,30,240,31,252,31,229,31,53,31,224,31,224,30,6,31,35,31,159,31,48,31,18,31,67,31,91,31,128,31,128,30,150,31,238,31,241,31,241,30,107,31,62,31,223,31,84,31,93,31,108,31,31,31,146,31,217,31,83,31,73,31,60,31,37,31,218,31,183,31,211,31,99,31,99,30,204,31,95,31,95,30,95,29,107,31,25,31,233,31,119,31,54,31,215,31,22,31,22,30,57,31,57,30,189,31,185,31,181,31,219,31,156,31,70,31,70,30,111,31,187,31,250,31,153,31,57,31,206,31,213,31,213,30,101,31,101,30,63,31,78,31,180,31,65,31,27,31,27,30,254,31,21,31,178,31,237,31,84,31,28,31,90,31,6,31,45,31,250,31,79,31,141,31,198,31,127,31,8,31,8,30,8,29,213,31,138,31,138,30,50,31,220,31,220,30,49,31,40,31,82,31,138,31,7,31,35,31,69,31,69,30,90,31,186,31,61,31,18,31,231,31,231,30,143,31,239,31,1,31,221,31,105,31,24,31,86,31,86,30,254,31,249,31,156,31,34,31,19,31,134,31,133,31,101,31,222,31,222,30,35,31,226,31,28,31,164,31,49,31,157,31,157,30,149,31,76,31,76,30,76,29,76,28,24,31,132,31,100,31,210,31,176,31,239,31,66,31,242,31,200,31,131,31,53,31,49,31,26,31,105,31,140,31,87,31,133,31,29,31,105,31,191,31,212,31,25,31,25,30,185,31,185,30,53,31,3,31,7,31,14,31,14,30,219,31,221,31,19,31,158,31,175,31,28,31,95,31,85,31,85,30,142,31,198,31,198,30,198,29,220,31,23,31,77,31,81,31,216,31,167,31,55,31,240,31,124,31,122,31,42,31,229,31,98,31,65,31,194,31,194,30,142,31,92,31,92,30,92,29,96,31,11,31,149,31,35,31,115,31,115,30,117,31,117,30,117,29,175,31,81,31,61,31,207,31,58,31,58,30,29,31,110,31,190,31,155,31,155,30,155,29,155,28,141,31,141,30,101,31,250,31,25,31,84,31,230,31,233,31,233,30,106,31,106,30,36,31,32,31,113,31,251,31,136,31,136,30,155,31,201,31,156,31,15,31,67,31,116,31,56,31,56,30,56,29,206,31,69,31,111,31,87,31,252,31,246,31,200,31,194,31,194,30,105,31,194,31,38,31,1,31,117,31,117,30,225,31,243,31,227,31,39,31,39,30,178,31,124,31,25,31,160,31,160,30,213,31,95,31,72,31,68,31,148,31,116,31,116,30,104,31,253,31,170,31,170,30,97,31,63,31,63,30,42,31,83,31,80,31,190,31,30,31,72,31,115,31,89,31,89,31,114,31,114,30,231,31,130,31,197,31,197,30,30,31,145,31,14,31,155,31,172,31,172,30,211,31,191,31,96,31,26,31,72,31,72,30,84,31,13,31,13,30,174,31,174,30,5,31,142,31,163,31,163,30,160,31,30,31,61,31,61,30,120,31,94,31,63,31,63,30,72,31,109,31,131,31,116,31,105,31,156,31,7,31,55,31,19,31,95,31,216,31,216,30,245,31,82,31,7,31,174,31,197,31,179,31,136,31,128,31,170,31,89,31,178,31,80,31,241,31,32,31,165,31,18,31,18,30,18,29,24,31,200,31,200,30,200,29,22,31,90,31,169,31,69,31,205,31,30,31,7,31,76,31,129,31,87,31,41,31,170,31,150,31,208,31,233,31,57,31,171,31,229,31,229,30,28,31,117,31,117,30,101,31,143,31,137,31,222,31,220,31,164,31,56,31,56,30,74,31,74,30,254,31,140,31,241,31,86,31,193,31,98,31,98,30,98,29,82,31,171,31,205,31,216,31,77,31,77,30,165,31,74,31,42,31,42,30,127,31,181,31,178,31,48,31,195,31,87,31,87,30,87,29,170,31,99,31,95,31,164,31,123,31,61,31,85,31,111,31,178,31,126,31,192,31,58,31,36,31,160,31,160,30,32,31,180,31,180,30,95,31,221,31,219,31,115,31,115,30,190,31,190,30,190,29,72,31,72,30,72,29,223,31,254,31,175,31,139,31,180,31,180,30,57,31,196,31,196,30,196,29,97,31,193,31,193,31,193,30,161,31,204,31,150,31,253,31,171,31,50,31,103,31,123,31,10,31,210,31,201,31,201,30,28,31,187,31,155,31,105,31,122,31,160,31,240,31,63,31,232,31,35,31,210,31,46,31,39,31,7,31,179,31,176,31,97,31,87,31,23,31,23,30,20,31,146,31,146,30,6,31,67,31,242,31,12,31,2,31,90,31,150,31,150,30,150,29,148,31,79,31,40,31,44,31,254,31,254,30,100,31,205,31,68,31,68,30,76,31,62,31,190,31,12,31,24,31,24,30,231,31,186,31,33,31,117,31,197,31,193,31,193,30,7,31,190,31,40,31,238,31,131,31,57,31,55,31,226,31,96,31,194,31,117,31,239,31,239,30,58,31,145,31,162,31,99,31,118,31,161,31,209,31,36,31,54,31,54,30,54,29,69,31,216,31,240,31,166,31,53,31,53,30,53,29,73,31,162,31,130,31,132,31,50,31,50,30,50,29,246,31,115,31,16,31,55,31,189,31,189,30,189,29,85,31,85,30,182,31,129,31,127,31,202,31,135,31,144,31,85,31,59,31,246,31,212,31,212,30,46,31,37,31,156,31,250,31,250,30,177,31,177,30,121,31,14,31,14,30,201,31,201,30,85,31,236,31,35,31,69,31,29,31,28,31,200,31,200,30,49,31,255,31,90,31,233,31,84,31,173,31,147,31,152,31,152,30,144,31,199,31,73,31,184,31,190,31,221,31,162,31,25,31,132,31,246,31,103,31,93,31,160,31,160,30,211,31,211,30,93,31,116,31,87,31,87,30,95,31,122,31,111,31,200,31,137,31,214,31,100,31,249,31,169,31,169,30,47,31,110,31,210,31,143,31,156,31,156,30,156,29,156,28,218,31,233,31,37,31,37,30,150,31,45,31,91,31,246,31,187,31,35,31,171,31,171,30,222,31,158,31,94,31,132,31,100,31,100,30,77,31,77,30,239,31,239,30,38,31,126,31,126,30,164,31,130,31,130,30,130,29,22,31,93,31,100,31,188,31,55,31,55,30,120,31,2,31,14,31,66,31,3,31,229,31,93,31,162,31,162,30,44,31,44,30,192,31,40,31,40,30,92,31,125,31,151,31,144,31,144,30,245,31,79,31,135,31,221,31,221,30,38,31,155,31,56,31,140,31,140,30,163,31,163,30,101,31,245,31,238,31,161,31,19,31,132,31,77,31,192,31,187,31,252,31,221,31,68,31,212,31,163,31,48,31,48,30,132,31,19,31,19,30,234,31,234,30,185,31,195,31,97,31,169,31,98,31,224,31,12,31,12,30,214,31,133,31,133,30,130,31,205,31,50,31,89,31,242,31,242,30,242,29,177,31,3,31,106,31,106,31,48,31,241,31,131,31,239,31,117,31,168,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
