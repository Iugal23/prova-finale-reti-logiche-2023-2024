-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_216 is
end project_tb_216;

architecture project_tb_arch_216 of project_tb_216 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (38,0,158,0,0,0,174,0,211,0,107,0,133,0,166,0,152,0,25,0,120,0,0,0,4,0,132,0,30,0,103,0,7,0,231,0,220,0,189,0,48,0,207,0,181,0,248,0,50,0,220,0,149,0,160,0,54,0,216,0,31,0,190,0,155,0,59,0,131,0,187,0,191,0,252,0,233,0,6,0,219,0,187,0,56,0,27,0,94,0,0,0,143,0,18,0,252,0,0,0,12,0,0,0,171,0,29,0,122,0,169,0,213,0,0,0,73,0,199,0,0,0,72,0,125,0,63,0,199,0,12,0,209,0,205,0,41,0,132,0,159,0,53,0,127,0,109,0,50,0,0,0,183,0,161,0,162,0,59,0,115,0,2,0,50,0,0,0,88,0,208,0,25,0,31,0,87,0,172,0,0,0,137,0,155,0,7,0,0,0,196,0,168,0,82,0,134,0,241,0,160,0,184,0,92,0,145,0,163,0,34,0,0,0,86,0,0,0,0,0,19,0,41,0,106,0,129,0,11,0,210,0,92,0,38,0,69,0,0,0,126,0,75,0,181,0,18,0,102,0,0,0,110,0,90,0,181,0,0,0,128,0,6,0,50,0,179,0,7,0,3,0,234,0,14,0,96,0,0,0,116,0,0,0,37,0,88,0,16,0,30,0,160,0,158,0,104,0,0,0,143,0,20,0,162,0,130,0,0,0,0,0,8,0,216,0,164,0,212,0,222,0,0,0,153,0,66,0,69,0,0,0,0,0,232,0,85,0,63,0,10,0,113,0,49,0,195,0,37,0,0,0,56,0,0,0,64,0,116,0,0,0,92,0,0,0,136,0,237,0,125,0,55,0,0,0,0,0,236,0,134,0,0,0,18,0,120,0,0,0,205,0,109,0,32,0,215,0,0,0,91,0,36,0,169,0,169,0,162,0,146,0,103,0,0,0,0,0,0,0,116,0,0,0,0,0,229,0,71,0,234,0,203,0,35,0,200,0,240,0,0,0,39,0,227,0,0,0,46,0,179,0,126,0,56,0,255,0,62,0,38,0,28,0,10,0,111,0,85,0,55,0,22,0,147,0,176,0,136,0,42,0,0,0,229,0,94,0,2,0,162,0,0,0,80,0,207,0,130,0,0,0,46,0,0,0,187,0,0,0,0,0,95,0,253,0,78,0,0,0,0,0,0,0,225,0,194,0,104,0,75,0,134,0,212,0,142,0,11,0,227,0,154,0,158,0,174,0,60,0,113,0,252,0,63,0,0,0,95,0,0,0,252,0,0,0,80,0,25,0,220,0,237,0,17,0,139,0,36,0,126,0,132,0,0,0,177,0,98,0,134,0,115,0,0,0,0,0,0,0,0,0,54,0,207,0,226,0,205,0,68,0,29,0,240,0,226,0,33,0,175,0,237,0,64,0,0,0,146,0,228,0,36,0,113,0,232,0,18,0,178,0,192,0,227,0,95,0,193,0,18,0,0,0,189,0,107,0,245,0,30,0,112,0,69,0,0,0,241,0,29,0,148,0,111,0,107,0,95,0,101,0,0,0,21,0,125,0,0,0,0,0,124,0,251,0,185,0,0,0,0,0,0,0,172,0,93,0,253,0,183,0,72,0,0,0,0,0,136,0,129,0,156,0,50,0,0,0,225,0,16,0,51,0,244,0,111,0,135,0,134,0,225,0,46,0,87,0,132,0,141,0,202,0,197,0,251,0,233,0,65,0,0,0,0,0,253,0,96,0,242,0,170,0,74,0,188,0,212,0,0,0,213,0,100,0,89,0,22,0,86,0,10,0,7,0,13,0,81,0,39,0,97,0,234,0,176,0,100,0,178,0,207,0,0,0,132,0,163,0,140,0,69,0,163,0,183,0,233,0,122,0,12,0,172,0,179,0,173,0,133,0,0,0,174,0,57,0,126,0,96,0,0,0,65,0,197,0,217,0,132,0,54,0,245,0,122,0,12,0,54,0,78,0,59,0,146,0,231,0,180,0,121,0,37,0,0,0,0,0,247,0,174,0,218,0,0,0,0,0,42,0,0,0,231,0,127,0,36,0,22,0,0,0,60,0,75,0,122,0,81,0,125,0,168,0,95,0,199,0,156,0,32,0,0,0,103,0,251,0,123,0,125,0,0,0,141,0,0,0,255,0,70,0,60,0,176,0,0,0,128,0,221,0,85,0,222,0,162,0,0,0,75,0,112,0,132,0,0,0,207,0,45,0,115,0,203,0,235,0,0,0,89,0,0,0,0,0,0,0,120,0,113,0,44,0,0,0,144,0,242,0,169,0,84,0,18,0,61,0,26,0,80,0,0,0,0,0,233,0,181,0,121,0,201,0,230,0,13,0,158,0,239,0,13,0,0,0,0,0,25,0,218,0,0,0,246,0,207,0,122,0,201,0,30,0,0,0,124,0,102,0,0,0,0,0,105,0,153,0,92,0,0,0,205,0,137,0,214,0,70,0,127,0,221,0,214,0,241,0,135,0,228,0,119,0,8,0,0,0,254,0,83,0,47,0,23,0,123,0,34,0,154,0,89,0,0,0,24,0,102,0,54,0,125,0,114,0,173,0,191,0,6,0,172,0,224,0,191,0,184,0,170,0,23,0,132,0,74,0,246,0,217,0,0,0,229,0,115,0,0,0,17,0,229,0,0,0,179,0,112,0,142,0,0,0,167,0,30,0,46,0,0,0,82,0,173,0,234,0,0,0,91,0,195,0,172,0,128,0,157,0,0,0,176,0,106,0,21,0,0,0,185,0,195,0,0,0,71,0,157,0,163,0,172,0,0,0,70,0,0,0,46,0,215,0,170,0,182,0,0,0,181,0,0,0,220,0,0,0,29,0,0,0,202,0,27,0,244,0,85,0,0,0,0,0,209,0,0,0,68,0,51,0,60,0,81,0,100,0,0,0);
signal scenario_full  : scenario_type := (38,31,158,31,158,30,174,31,211,31,107,31,133,31,166,31,152,31,25,31,120,31,120,30,4,31,132,31,30,31,103,31,7,31,231,31,220,31,189,31,48,31,207,31,181,31,248,31,50,31,220,31,149,31,160,31,54,31,216,31,31,31,190,31,155,31,59,31,131,31,187,31,191,31,252,31,233,31,6,31,219,31,187,31,56,31,27,31,94,31,94,30,143,31,18,31,252,31,252,30,12,31,12,30,171,31,29,31,122,31,169,31,213,31,213,30,73,31,199,31,199,30,72,31,125,31,63,31,199,31,12,31,209,31,205,31,41,31,132,31,159,31,53,31,127,31,109,31,50,31,50,30,183,31,161,31,162,31,59,31,115,31,2,31,50,31,50,30,88,31,208,31,25,31,31,31,87,31,172,31,172,30,137,31,155,31,7,31,7,30,196,31,168,31,82,31,134,31,241,31,160,31,184,31,92,31,145,31,163,31,34,31,34,30,86,31,86,30,86,29,19,31,41,31,106,31,129,31,11,31,210,31,92,31,38,31,69,31,69,30,126,31,75,31,181,31,18,31,102,31,102,30,110,31,90,31,181,31,181,30,128,31,6,31,50,31,179,31,7,31,3,31,234,31,14,31,96,31,96,30,116,31,116,30,37,31,88,31,16,31,30,31,160,31,158,31,104,31,104,30,143,31,20,31,162,31,130,31,130,30,130,29,8,31,216,31,164,31,212,31,222,31,222,30,153,31,66,31,69,31,69,30,69,29,232,31,85,31,63,31,10,31,113,31,49,31,195,31,37,31,37,30,56,31,56,30,64,31,116,31,116,30,92,31,92,30,136,31,237,31,125,31,55,31,55,30,55,29,236,31,134,31,134,30,18,31,120,31,120,30,205,31,109,31,32,31,215,31,215,30,91,31,36,31,169,31,169,31,162,31,146,31,103,31,103,30,103,29,103,28,116,31,116,30,116,29,229,31,71,31,234,31,203,31,35,31,200,31,240,31,240,30,39,31,227,31,227,30,46,31,179,31,126,31,56,31,255,31,62,31,38,31,28,31,10,31,111,31,85,31,55,31,22,31,147,31,176,31,136,31,42,31,42,30,229,31,94,31,2,31,162,31,162,30,80,31,207,31,130,31,130,30,46,31,46,30,187,31,187,30,187,29,95,31,253,31,78,31,78,30,78,29,78,28,225,31,194,31,104,31,75,31,134,31,212,31,142,31,11,31,227,31,154,31,158,31,174,31,60,31,113,31,252,31,63,31,63,30,95,31,95,30,252,31,252,30,80,31,25,31,220,31,237,31,17,31,139,31,36,31,126,31,132,31,132,30,177,31,98,31,134,31,115,31,115,30,115,29,115,28,115,27,54,31,207,31,226,31,205,31,68,31,29,31,240,31,226,31,33,31,175,31,237,31,64,31,64,30,146,31,228,31,36,31,113,31,232,31,18,31,178,31,192,31,227,31,95,31,193,31,18,31,18,30,189,31,107,31,245,31,30,31,112,31,69,31,69,30,241,31,29,31,148,31,111,31,107,31,95,31,101,31,101,30,21,31,125,31,125,30,125,29,124,31,251,31,185,31,185,30,185,29,185,28,172,31,93,31,253,31,183,31,72,31,72,30,72,29,136,31,129,31,156,31,50,31,50,30,225,31,16,31,51,31,244,31,111,31,135,31,134,31,225,31,46,31,87,31,132,31,141,31,202,31,197,31,251,31,233,31,65,31,65,30,65,29,253,31,96,31,242,31,170,31,74,31,188,31,212,31,212,30,213,31,100,31,89,31,22,31,86,31,10,31,7,31,13,31,81,31,39,31,97,31,234,31,176,31,100,31,178,31,207,31,207,30,132,31,163,31,140,31,69,31,163,31,183,31,233,31,122,31,12,31,172,31,179,31,173,31,133,31,133,30,174,31,57,31,126,31,96,31,96,30,65,31,197,31,217,31,132,31,54,31,245,31,122,31,12,31,54,31,78,31,59,31,146,31,231,31,180,31,121,31,37,31,37,30,37,29,247,31,174,31,218,31,218,30,218,29,42,31,42,30,231,31,127,31,36,31,22,31,22,30,60,31,75,31,122,31,81,31,125,31,168,31,95,31,199,31,156,31,32,31,32,30,103,31,251,31,123,31,125,31,125,30,141,31,141,30,255,31,70,31,60,31,176,31,176,30,128,31,221,31,85,31,222,31,162,31,162,30,75,31,112,31,132,31,132,30,207,31,45,31,115,31,203,31,235,31,235,30,89,31,89,30,89,29,89,28,120,31,113,31,44,31,44,30,144,31,242,31,169,31,84,31,18,31,61,31,26,31,80,31,80,30,80,29,233,31,181,31,121,31,201,31,230,31,13,31,158,31,239,31,13,31,13,30,13,29,25,31,218,31,218,30,246,31,207,31,122,31,201,31,30,31,30,30,124,31,102,31,102,30,102,29,105,31,153,31,92,31,92,30,205,31,137,31,214,31,70,31,127,31,221,31,214,31,241,31,135,31,228,31,119,31,8,31,8,30,254,31,83,31,47,31,23,31,123,31,34,31,154,31,89,31,89,30,24,31,102,31,54,31,125,31,114,31,173,31,191,31,6,31,172,31,224,31,191,31,184,31,170,31,23,31,132,31,74,31,246,31,217,31,217,30,229,31,115,31,115,30,17,31,229,31,229,30,179,31,112,31,142,31,142,30,167,31,30,31,46,31,46,30,82,31,173,31,234,31,234,30,91,31,195,31,172,31,128,31,157,31,157,30,176,31,106,31,21,31,21,30,185,31,195,31,195,30,71,31,157,31,163,31,172,31,172,30,70,31,70,30,46,31,215,31,170,31,182,31,182,30,181,31,181,30,220,31,220,30,29,31,29,30,202,31,27,31,244,31,85,31,85,30,85,29,209,31,209,30,68,31,51,31,60,31,81,31,100,31,100,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
