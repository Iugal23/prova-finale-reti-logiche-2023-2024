-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_751 is
end project_tb_751;

architecture project_tb_arch_751 of project_tb_751 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 932;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,0,0,249,0,201,0,68,0,160,0,55,0,89,0,119,0,45,0,32,0,161,0,254,0,0,0,194,0,174,0,202,0,173,0,51,0,175,0,66,0,74,0,43,0,83,0,92,0,0,0,86,0,0,0,42,0,130,0,179,0,0,0,6,0,0,0,154,0,228,0,0,0,48,0,224,0,0,0,162,0,100,0,4,0,79,0,76,0,202,0,144,0,209,0,146,0,0,0,157,0,47,0,25,0,191,0,91,0,65,0,251,0,0,0,152,0,222,0,0,0,90,0,187,0,215,0,166,0,122,0,211,0,215,0,251,0,187,0,67,0,80,0,140,0,34,0,159,0,254,0,191,0,143,0,39,0,231,0,25,0,161,0,92,0,0,0,145,0,0,0,36,0,0,0,58,0,67,0,166,0,222,0,86,0,45,0,192,0,0,0,243,0,0,0,189,0,139,0,0,0,0,0,150,0,201,0,106,0,140,0,0,0,189,0,48,0,108,0,210,0,20,0,236,0,250,0,21,0,117,0,243,0,68,0,53,0,0,0,228,0,0,0,122,0,33,0,170,0,0,0,60,0,217,0,0,0,213,0,207,0,134,0,104,0,0,0,135,0,48,0,0,0,52,0,35,0,0,0,0,0,187,0,220,0,0,0,134,0,37,0,150,0,73,0,222,0,242,0,25,0,21,0,0,0,0,0,139,0,192,0,217,0,0,0,67,0,96,0,251,0,0,0,30,0,34,0,0,0,0,0,0,0,0,0,94,0,213,0,38,0,144,0,245,0,0,0,0,0,97,0,230,0,37,0,31,0,0,0,229,0,37,0,108,0,0,0,141,0,239,0,202,0,85,0,46,0,84,0,178,0,221,0,0,0,37,0,162,0,179,0,149,0,205,0,0,0,0,0,0,0,163,0,157,0,93,0,0,0,0,0,0,0,210,0,0,0,0,0,245,0,111,0,193,0,125,0,0,0,117,0,71,0,203,0,209,0,135,0,169,0,0,0,45,0,167,0,0,0,94,0,5,0,227,0,249,0,161,0,0,0,0,0,223,0,220,0,28,0,217,0,232,0,0,0,230,0,178,0,189,0,234,0,0,0,183,0,145,0,21,0,231,0,123,0,80,0,209,0,227,0,47,0,2,0,220,0,226,0,49,0,213,0,45,0,78,0,0,0,169,0,200,0,157,0,193,0,111,0,157,0,0,0,173,0,231,0,119,0,110,0,102,0,181,0,162,0,61,0,2,0,0,0,4,0,76,0,116,0,165,0,0,0,0,0,3,0,111,0,49,0,141,0,79,0,49,0,228,0,74,0,201,0,190,0,34,0,249,0,0,0,0,0,126,0,39,0,104,0,39,0,246,0,0,0,37,0,98,0,59,0,142,0,73,0,59,0,37,0,217,0,72,0,0,0,227,0,9,0,0,0,0,0,0,0,0,0,35,0,152,0,78,0,223,0,131,0,41,0,132,0,6,0,152,0,103,0,0,0,20,0,0,0,0,0,214,0,81,0,142,0,253,0,68,0,62,0,100,0,21,0,191,0,222,0,149,0,28,0,162,0,209,0,49,0,69,0,247,0,0,0,182,0,2,0,0,0,0,0,197,0,102,0,0,0,42,0,128,0,131,0,63,0,61,0,84,0,0,0,0,0,172,0,86,0,0,0,83,0,242,0,246,0,51,0,120,0,156,0,0,0,243,0,151,0,183,0,91,0,244,0,5,0,220,0,194,0,69,0,84,0,125,0,215,0,231,0,245,0,120,0,73,0,188,0,124,0,25,0,92,0,117,0,49,0,146,0,211,0,0,0,18,0,5,0,0,0,136,0,171,0,0,0,195,0,109,0,187,0,202,0,112,0,212,0,221,0,15,0,56,0,161,0,202,0,0,0,27,0,236,0,0,0,221,0,172,0,214,0,120,0,37,0,206,0,0,0,182,0,251,0,92,0,204,0,44,0,135,0,95,0,0,0,0,0,0,0,0,0,17,0,100,0,160,0,29,0,224,0,34,0,87,0,173,0,87,0,4,0,15,0,114,0,0,0,193,0,246,0,0,0,0,0,109,0,132,0,0,0,14,0,31,0,17,0,0,0,197,0,0,0,111,0,134,0,254,0,0,0,57,0,127,0,166,0,134,0,201,0,30,0,69,0,157,0,55,0,169,0,66,0,16,0,189,0,0,0,0,0,22,0,243,0,82,0,184,0,0,0,238,0,221,0,0,0,231,0,230,0,4,0,49,0,83,0,0,0,0,0,184,0,203,0,166,0,160,0,181,0,68,0,0,0,0,0,236,0,0,0,152,0,0,0,254,0,104,0,8,0,234,0,189,0,18,0,68,0,192,0,55,0,134,0,0,0,19,0,93,0,35,0,240,0,139,0,163,0,123,0,9,0,7,0,0,0,82,0,0,0,184,0,202,0,150,0,195,0,147,0,81,0,140,0,54,0,0,0,9,0,0,0,141,0,129,0,250,0,11,0,247,0,0,0,66,0,0,0,188,0,207,0,42,0,194,0,0,0,105,0,213,0,0,0,107,0,198,0,0,0,220,0,249,0,135,0,164,0,14,0,120,0,211,0,207,0,220,0,45,0,129,0,38,0,102,0,155,0,0,0,192,0,197,0,45,0,0,0,196,0,100,0,125,0,237,0,214,0,181,0,51,0,132,0,3,0,179,0,137,0,0,0,166,0,247,0,116,0,235,0,96,0,107,0,42,0,0,0,13,0,0,0,0,0,6,0,164,0,208,0,140,0,231,0,44,0,80,0,178,0,0,0,229,0,171,0,3,0,197,0,13,0,55,0,0,0,0,0,175,0,161,0,235,0,0,0,175,0,72,0,154,0,219,0,183,0,171,0,141,0,207,0,115,0,20,0,229,0,181,0,158,0,30,0,0,0,254,0,0,0,38,0,163,0,95,0,131,0,123,0,25,0,0,0,203,0,118,0,105,0,208,0,12,0,0,0,40,0,36,0,214,0,0,0,239,0,69,0,0,0,0,0,77,0,68,0,0,0,87,0,0,0,42,0,67,0,75,0,0,0,134,0,0,0,113,0,118,0,0,0,151,0,59,0,157,0,0,0,0,0,0,0,192,0,71,0,62,0,242,0,20,0,0,0,197,0,81,0,218,0,141,0,170,0,223,0,131,0,177,0,241,0,84,0,243,0,200,0,108,0,119,0,134,0,255,0,163,0,235,0,17,0,139,0,115,0,0,0,94,0,150,0,138,0,0,0,0,0,230,0,191,0,0,0,212,0,143,0,0,0,33,0,146,0,0,0,233,0,0,0,253,0,90,0,101,0,142,0,86,0,154,0,209,0,212,0,24,0,247,0,230,0,0,0,231,0,110,0,0,0,200,0,0,0,173,0,0,0,64,0,20,0,0,0,168,0,0,0,221,0,132,0,75,0,28,0,161,0,0,0,116,0,0,0,193,0,209,0,99,0,181,0,0,0,151,0,104,0,166,0,185,0,0,0,246,0,193,0,0,0,239,0,231,0,85,0,252,0,50,0,192,0,68,0,248,0,176,0,0,0,157,0,41,0,95,0,79,0,0,0,11,0,112,0,244,0,0,0,78,0,168,0,184,0,229,0,66,0,200,0,209,0,235,0,223,0,180,0,0,0,0,0,0,0,0,0,129,0,34,0,244,0,31,0,51,0,22,0,0,0,53,0,0,0,191,0,112,0,213,0,0,0,0,0,0,0,0,0,84,0,225,0,27,0,0,0,115,0,186,0,192,0,0,0,0,0,91,0,103,0,218,0,229,0,247,0,31,0,0,0,110,0,78,0,0,0,252,0,177,0,63,0,5,0,216,0,13,0,243,0,123,0,229,0,0,0,142,0,0,0,232,0,225,0,14,0,0,0,115,0,31,0,224,0,101,0,66,0,68,0,17,0,0,0,89,0,177,0,45,0,144,0,42,0,56,0,97,0,139,0,23,0,143,0,0,0,0,0,150,0,224,0,143,0,193,0,73,0,22,0,171,0,143,0,0,0,223,0,147,0,64,0,0,0,51,0,14,0,227,0,0,0,32,0,39,0,158,0,65,0,224,0,165,0,64,0,221,0,160,0,49,0,0,0,109,0,25,0,232,0,143,0,79,0,173,0,21,0,172,0,97,0,61,0,247,0,0,0,201,0,223,0,140,0,59,0,23,0,81,0,162,0,57,0,118,0,0,0,25,0,247,0,181,0);
signal scenario_full  : scenario_type := (102,31,102,30,249,31,201,31,68,31,160,31,55,31,89,31,119,31,45,31,32,31,161,31,254,31,254,30,194,31,174,31,202,31,173,31,51,31,175,31,66,31,74,31,43,31,83,31,92,31,92,30,86,31,86,30,42,31,130,31,179,31,179,30,6,31,6,30,154,31,228,31,228,30,48,31,224,31,224,30,162,31,100,31,4,31,79,31,76,31,202,31,144,31,209,31,146,31,146,30,157,31,47,31,25,31,191,31,91,31,65,31,251,31,251,30,152,31,222,31,222,30,90,31,187,31,215,31,166,31,122,31,211,31,215,31,251,31,187,31,67,31,80,31,140,31,34,31,159,31,254,31,191,31,143,31,39,31,231,31,25,31,161,31,92,31,92,30,145,31,145,30,36,31,36,30,58,31,67,31,166,31,222,31,86,31,45,31,192,31,192,30,243,31,243,30,189,31,139,31,139,30,139,29,150,31,201,31,106,31,140,31,140,30,189,31,48,31,108,31,210,31,20,31,236,31,250,31,21,31,117,31,243,31,68,31,53,31,53,30,228,31,228,30,122,31,33,31,170,31,170,30,60,31,217,31,217,30,213,31,207,31,134,31,104,31,104,30,135,31,48,31,48,30,52,31,35,31,35,30,35,29,187,31,220,31,220,30,134,31,37,31,150,31,73,31,222,31,242,31,25,31,21,31,21,30,21,29,139,31,192,31,217,31,217,30,67,31,96,31,251,31,251,30,30,31,34,31,34,30,34,29,34,28,34,27,94,31,213,31,38,31,144,31,245,31,245,30,245,29,97,31,230,31,37,31,31,31,31,30,229,31,37,31,108,31,108,30,141,31,239,31,202,31,85,31,46,31,84,31,178,31,221,31,221,30,37,31,162,31,179,31,149,31,205,31,205,30,205,29,205,28,163,31,157,31,93,31,93,30,93,29,93,28,210,31,210,30,210,29,245,31,111,31,193,31,125,31,125,30,117,31,71,31,203,31,209,31,135,31,169,31,169,30,45,31,167,31,167,30,94,31,5,31,227,31,249,31,161,31,161,30,161,29,223,31,220,31,28,31,217,31,232,31,232,30,230,31,178,31,189,31,234,31,234,30,183,31,145,31,21,31,231,31,123,31,80,31,209,31,227,31,47,31,2,31,220,31,226,31,49,31,213,31,45,31,78,31,78,30,169,31,200,31,157,31,193,31,111,31,157,31,157,30,173,31,231,31,119,31,110,31,102,31,181,31,162,31,61,31,2,31,2,30,4,31,76,31,116,31,165,31,165,30,165,29,3,31,111,31,49,31,141,31,79,31,49,31,228,31,74,31,201,31,190,31,34,31,249,31,249,30,249,29,126,31,39,31,104,31,39,31,246,31,246,30,37,31,98,31,59,31,142,31,73,31,59,31,37,31,217,31,72,31,72,30,227,31,9,31,9,30,9,29,9,28,9,27,35,31,152,31,78,31,223,31,131,31,41,31,132,31,6,31,152,31,103,31,103,30,20,31,20,30,20,29,214,31,81,31,142,31,253,31,68,31,62,31,100,31,21,31,191,31,222,31,149,31,28,31,162,31,209,31,49,31,69,31,247,31,247,30,182,31,2,31,2,30,2,29,197,31,102,31,102,30,42,31,128,31,131,31,63,31,61,31,84,31,84,30,84,29,172,31,86,31,86,30,83,31,242,31,246,31,51,31,120,31,156,31,156,30,243,31,151,31,183,31,91,31,244,31,5,31,220,31,194,31,69,31,84,31,125,31,215,31,231,31,245,31,120,31,73,31,188,31,124,31,25,31,92,31,117,31,49,31,146,31,211,31,211,30,18,31,5,31,5,30,136,31,171,31,171,30,195,31,109,31,187,31,202,31,112,31,212,31,221,31,15,31,56,31,161,31,202,31,202,30,27,31,236,31,236,30,221,31,172,31,214,31,120,31,37,31,206,31,206,30,182,31,251,31,92,31,204,31,44,31,135,31,95,31,95,30,95,29,95,28,95,27,17,31,100,31,160,31,29,31,224,31,34,31,87,31,173,31,87,31,4,31,15,31,114,31,114,30,193,31,246,31,246,30,246,29,109,31,132,31,132,30,14,31,31,31,17,31,17,30,197,31,197,30,111,31,134,31,254,31,254,30,57,31,127,31,166,31,134,31,201,31,30,31,69,31,157,31,55,31,169,31,66,31,16,31,189,31,189,30,189,29,22,31,243,31,82,31,184,31,184,30,238,31,221,31,221,30,231,31,230,31,4,31,49,31,83,31,83,30,83,29,184,31,203,31,166,31,160,31,181,31,68,31,68,30,68,29,236,31,236,30,152,31,152,30,254,31,104,31,8,31,234,31,189,31,18,31,68,31,192,31,55,31,134,31,134,30,19,31,93,31,35,31,240,31,139,31,163,31,123,31,9,31,7,31,7,30,82,31,82,30,184,31,202,31,150,31,195,31,147,31,81,31,140,31,54,31,54,30,9,31,9,30,141,31,129,31,250,31,11,31,247,31,247,30,66,31,66,30,188,31,207,31,42,31,194,31,194,30,105,31,213,31,213,30,107,31,198,31,198,30,220,31,249,31,135,31,164,31,14,31,120,31,211,31,207,31,220,31,45,31,129,31,38,31,102,31,155,31,155,30,192,31,197,31,45,31,45,30,196,31,100,31,125,31,237,31,214,31,181,31,51,31,132,31,3,31,179,31,137,31,137,30,166,31,247,31,116,31,235,31,96,31,107,31,42,31,42,30,13,31,13,30,13,29,6,31,164,31,208,31,140,31,231,31,44,31,80,31,178,31,178,30,229,31,171,31,3,31,197,31,13,31,55,31,55,30,55,29,175,31,161,31,235,31,235,30,175,31,72,31,154,31,219,31,183,31,171,31,141,31,207,31,115,31,20,31,229,31,181,31,158,31,30,31,30,30,254,31,254,30,38,31,163,31,95,31,131,31,123,31,25,31,25,30,203,31,118,31,105,31,208,31,12,31,12,30,40,31,36,31,214,31,214,30,239,31,69,31,69,30,69,29,77,31,68,31,68,30,87,31,87,30,42,31,67,31,75,31,75,30,134,31,134,30,113,31,118,31,118,30,151,31,59,31,157,31,157,30,157,29,157,28,192,31,71,31,62,31,242,31,20,31,20,30,197,31,81,31,218,31,141,31,170,31,223,31,131,31,177,31,241,31,84,31,243,31,200,31,108,31,119,31,134,31,255,31,163,31,235,31,17,31,139,31,115,31,115,30,94,31,150,31,138,31,138,30,138,29,230,31,191,31,191,30,212,31,143,31,143,30,33,31,146,31,146,30,233,31,233,30,253,31,90,31,101,31,142,31,86,31,154,31,209,31,212,31,24,31,247,31,230,31,230,30,231,31,110,31,110,30,200,31,200,30,173,31,173,30,64,31,20,31,20,30,168,31,168,30,221,31,132,31,75,31,28,31,161,31,161,30,116,31,116,30,193,31,209,31,99,31,181,31,181,30,151,31,104,31,166,31,185,31,185,30,246,31,193,31,193,30,239,31,231,31,85,31,252,31,50,31,192,31,68,31,248,31,176,31,176,30,157,31,41,31,95,31,79,31,79,30,11,31,112,31,244,31,244,30,78,31,168,31,184,31,229,31,66,31,200,31,209,31,235,31,223,31,180,31,180,30,180,29,180,28,180,27,129,31,34,31,244,31,31,31,51,31,22,31,22,30,53,31,53,30,191,31,112,31,213,31,213,30,213,29,213,28,213,27,84,31,225,31,27,31,27,30,115,31,186,31,192,31,192,30,192,29,91,31,103,31,218,31,229,31,247,31,31,31,31,30,110,31,78,31,78,30,252,31,177,31,63,31,5,31,216,31,13,31,243,31,123,31,229,31,229,30,142,31,142,30,232,31,225,31,14,31,14,30,115,31,31,31,224,31,101,31,66,31,68,31,17,31,17,30,89,31,177,31,45,31,144,31,42,31,56,31,97,31,139,31,23,31,143,31,143,30,143,29,150,31,224,31,143,31,193,31,73,31,22,31,171,31,143,31,143,30,223,31,147,31,64,31,64,30,51,31,14,31,227,31,227,30,32,31,39,31,158,31,65,31,224,31,165,31,64,31,221,31,160,31,49,31,49,30,109,31,25,31,232,31,143,31,79,31,173,31,21,31,172,31,97,31,61,31,247,31,247,30,201,31,223,31,140,31,59,31,23,31,81,31,162,31,57,31,118,31,118,30,25,31,247,31,181,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
