-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_784 is
end project_tb_784;

architecture project_tb_arch_784 of project_tb_784 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 800;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (236,0,0,0,201,0,107,0,126,0,54,0,148,0,221,0,201,0,0,0,121,0,0,0,218,0,76,0,0,0,90,0,202,0,70,0,180,0,5,0,0,0,8,0,0,0,39,0,208,0,142,0,0,0,2,0,164,0,57,0,48,0,0,0,253,0,61,0,181,0,217,0,118,0,246,0,216,0,166,0,218,0,198,0,0,0,0,0,2,0,116,0,0,0,171,0,0,0,114,0,207,0,183,0,48,0,133,0,229,0,0,0,192,0,0,0,12,0,198,0,196,0,69,0,33,0,156,0,90,0,2,0,0,0,0,0,0,0,67,0,246,0,185,0,21,0,252,0,130,0,82,0,21,0,0,0,236,0,0,0,220,0,189,0,167,0,124,0,0,0,192,0,205,0,203,0,193,0,89,0,104,0,57,0,147,0,123,0,132,0,98,0,154,0,198,0,146,0,0,0,180,0,177,0,210,0,0,0,0,0,57,0,159,0,66,0,209,0,97,0,171,0,37,0,73,0,86,0,238,0,229,0,233,0,0,0,149,0,47,0,226,0,0,0,0,0,254,0,203,0,196,0,0,0,48,0,0,0,111,0,0,0,0,0,250,0,114,0,90,0,195,0,55,0,0,0,61,0,0,0,0,0,168,0,0,0,41,0,110,0,59,0,0,0,0,0,56,0,159,0,200,0,160,0,134,0,0,0,14,0,0,0,82,0,119,0,167,0,87,0,134,0,119,0,0,0,0,0,71,0,37,0,127,0,0,0,0,0,135,0,52,0,66,0,191,0,0,0,218,0,11,0,97,0,42,0,110,0,0,0,193,0,184,0,133,0,105,0,9,0,0,0,33,0,147,0,0,0,96,0,6,0,33,0,85,0,132,0,63,0,3,0,121,0,167,0,250,0,233,0,123,0,224,0,49,0,225,0,50,0,252,0,145,0,0,0,15,0,229,0,222,0,145,0,148,0,121,0,0,0,249,0,249,0,15,0,206,0,101,0,191,0,42,0,9,0,128,0,0,0,0,0,36,0,151,0,116,0,103,0,0,0,0,0,130,0,36,0,0,0,151,0,0,0,0,0,84,0,34,0,0,0,59,0,39,0,0,0,0,0,109,0,212,0,192,0,0,0,232,0,110,0,155,0,147,0,197,0,152,0,97,0,38,0,167,0,207,0,114,0,246,0,0,0,163,0,85,0,143,0,140,0,0,0,102,0,220,0,0,0,134,0,214,0,211,0,237,0,252,0,1,0,0,0,134,0,250,0,51,0,204,0,11,0,46,0,107,0,152,0,32,0,136,0,45,0,0,0,0,0,0,0,43,0,0,0,75,0,10,0,210,0,99,0,0,0,199,0,250,0,33,0,0,0,162,0,11,0,232,0,0,0,199,0,60,0,0,0,0,0,0,0,237,0,105,0,181,0,248,0,252,0,215,0,0,0,139,0,105,0,159,0,28,0,159,0,113,0,78,0,13,0,227,0,99,0,59,0,222,0,27,0,0,0,9,0,132,0,166,0,35,0,0,0,135,0,36,0,54,0,53,0,110,0,190,0,124,0,109,0,128,0,235,0,33,0,0,0,39,0,58,0,244,0,132,0,80,0,182,0,0,0,0,0,0,0,0,0,237,0,85,0,3,0,196,0,25,0,37,0,247,0,211,0,82,0,194,0,0,0,0,0,160,0,127,0,171,0,34,0,0,0,49,0,211,0,41,0,130,0,216,0,176,0,18,0,255,0,115,0,249,0,0,0,253,0,49,0,15,0,113,0,224,0,0,0,151,0,208,0,122,0,0,0,80,0,254,0,0,0,186,0,0,0,54,0,145,0,13,0,192,0,41,0,140,0,0,0,147,0,105,0,18,0,2,0,37,0,42,0,71,0,0,0,237,0,183,0,203,0,0,0,57,0,248,0,119,0,0,0,112,0,122,0,93,0,17,0,83,0,78,0,157,0,217,0,0,0,173,0,104,0,38,0,0,0,26,0,103,0,190,0,234,0,76,0,125,0,223,0,176,0,65,0,28,0,232,0,42,0,80,0,128,0,81,0,181,0,130,0,65,0,226,0,81,0,141,0,118,0,177,0,245,0,174,0,234,0,97,0,30,0,176,0,138,0,125,0,63,0,198,0,98,0,32,0,62,0,232,0,87,0,222,0,61,0,178,0,80,0,0,0,31,0,148,0,17,0,3,0,0,0,47,0,133,0,163,0,0,0,247,0,54,0,116,0,177,0,208,0,82,0,173,0,11,0,41,0,53,0,13,0,160,0,94,0,0,0,116,0,129,0,85,0,94,0,0,0,230,0,22,0,102,0,151,0,13,0,131,0,62,0,52,0,20,0,120,0,76,0,202,0,207,0,227,0,0,0,2,0,17,0,177,0,215,0,91,0,103,0,16,0,7,0,66,0,0,0,177,0,129,0,22,0,115,0,0,0,0,0,0,0,0,0,116,0,172,0,178,0,142,0,177,0,189,0,103,0,171,0,248,0,3,0,189,0,18,0,0,0,95,0,158,0,0,0,11,0,53,0,144,0,20,0,0,0,30,0,82,0,25,0,172,0,235,0,0,0,148,0,0,0,243,0,66,0,2,0,48,0,217,0,131,0,169,0,0,0,0,0,233,0,94,0,0,0,255,0,16,0,181,0,0,0,0,0,112,0,0,0,0,0,0,0,0,0,245,0,131,0,17,0,100,0,21,0,212,0,145,0,158,0,175,0,219,0,251,0,103,0,73,0,0,0,13,0,0,0,165,0,106,0,79,0,0,0,136,0,240,0,251,0,233,0,57,0,211,0,90,0,21,0,187,0,0,0,201,0,227,0,250,0,6,0,216,0,213,0,125,0,0,0,94,0,223,0,0,0,0,0,73,0,251,0,89,0,36,0,184,0,252,0,251,0,210,0,166,0,175,0,0,0,0,0,123,0,245,0,117,0,174,0,143,0,156,0,114,0,96,0,0,0,0,0,117,0,0,0,15,0,56,0,160,0,0,0,239,0,6,0,139,0,37,0,0,0,44,0,0,0,217,0,0,0,0,0,10,0,0,0,53,0,0,0,33,0,41,0,8,0,46,0,79,0,47,0,129,0,66,0,119,0,138,0,96,0,158,0,138,0,65,0,230,0,0,0,7,0,116,0,105,0,127,0,33,0,247,0,216,0,214,0,10,0,0,0,151,0,176,0,73,0,0,0,172,0,189,0,0,0,83,0,0,0,211,0,116,0,167,0,0,0,93,0,168,0,103,0,40,0,134,0,219,0,27,0,0,0,221,0,0,0,101,0,202,0,140,0,20,0,250,0,95,0,3,0,206,0,246,0,115,0,120,0,135,0,2,0,253,0,103,0,0,0,175,0,1,0,32,0,150,0,0,0,244,0,76,0,0,0,55,0,0,0,209,0,0,0,8,0,41,0,30,0,6,0,94,0,199,0,0,0,24,0,50,0,171,0,113,0,77,0,0,0,251,0,64,0,13,0,168,0,155,0,226,0,32,0,63,0,19,0,103,0,17,0,113,0,125,0,8,0,164,0,0,0,0,0,63,0,245,0,110,0,191,0,82,0,68,0,56,0,191,0,159,0,238,0,105,0,90,0,220,0,0,0,111,0,77,0);
signal scenario_full  : scenario_type := (236,31,236,30,201,31,107,31,126,31,54,31,148,31,221,31,201,31,201,30,121,31,121,30,218,31,76,31,76,30,90,31,202,31,70,31,180,31,5,31,5,30,8,31,8,30,39,31,208,31,142,31,142,30,2,31,164,31,57,31,48,31,48,30,253,31,61,31,181,31,217,31,118,31,246,31,216,31,166,31,218,31,198,31,198,30,198,29,2,31,116,31,116,30,171,31,171,30,114,31,207,31,183,31,48,31,133,31,229,31,229,30,192,31,192,30,12,31,198,31,196,31,69,31,33,31,156,31,90,31,2,31,2,30,2,29,2,28,67,31,246,31,185,31,21,31,252,31,130,31,82,31,21,31,21,30,236,31,236,30,220,31,189,31,167,31,124,31,124,30,192,31,205,31,203,31,193,31,89,31,104,31,57,31,147,31,123,31,132,31,98,31,154,31,198,31,146,31,146,30,180,31,177,31,210,31,210,30,210,29,57,31,159,31,66,31,209,31,97,31,171,31,37,31,73,31,86,31,238,31,229,31,233,31,233,30,149,31,47,31,226,31,226,30,226,29,254,31,203,31,196,31,196,30,48,31,48,30,111,31,111,30,111,29,250,31,114,31,90,31,195,31,55,31,55,30,61,31,61,30,61,29,168,31,168,30,41,31,110,31,59,31,59,30,59,29,56,31,159,31,200,31,160,31,134,31,134,30,14,31,14,30,82,31,119,31,167,31,87,31,134,31,119,31,119,30,119,29,71,31,37,31,127,31,127,30,127,29,135,31,52,31,66,31,191,31,191,30,218,31,11,31,97,31,42,31,110,31,110,30,193,31,184,31,133,31,105,31,9,31,9,30,33,31,147,31,147,30,96,31,6,31,33,31,85,31,132,31,63,31,3,31,121,31,167,31,250,31,233,31,123,31,224,31,49,31,225,31,50,31,252,31,145,31,145,30,15,31,229,31,222,31,145,31,148,31,121,31,121,30,249,31,249,31,15,31,206,31,101,31,191,31,42,31,9,31,128,31,128,30,128,29,36,31,151,31,116,31,103,31,103,30,103,29,130,31,36,31,36,30,151,31,151,30,151,29,84,31,34,31,34,30,59,31,39,31,39,30,39,29,109,31,212,31,192,31,192,30,232,31,110,31,155,31,147,31,197,31,152,31,97,31,38,31,167,31,207,31,114,31,246,31,246,30,163,31,85,31,143,31,140,31,140,30,102,31,220,31,220,30,134,31,214,31,211,31,237,31,252,31,1,31,1,30,134,31,250,31,51,31,204,31,11,31,46,31,107,31,152,31,32,31,136,31,45,31,45,30,45,29,45,28,43,31,43,30,75,31,10,31,210,31,99,31,99,30,199,31,250,31,33,31,33,30,162,31,11,31,232,31,232,30,199,31,60,31,60,30,60,29,60,28,237,31,105,31,181,31,248,31,252,31,215,31,215,30,139,31,105,31,159,31,28,31,159,31,113,31,78,31,13,31,227,31,99,31,59,31,222,31,27,31,27,30,9,31,132,31,166,31,35,31,35,30,135,31,36,31,54,31,53,31,110,31,190,31,124,31,109,31,128,31,235,31,33,31,33,30,39,31,58,31,244,31,132,31,80,31,182,31,182,30,182,29,182,28,182,27,237,31,85,31,3,31,196,31,25,31,37,31,247,31,211,31,82,31,194,31,194,30,194,29,160,31,127,31,171,31,34,31,34,30,49,31,211,31,41,31,130,31,216,31,176,31,18,31,255,31,115,31,249,31,249,30,253,31,49,31,15,31,113,31,224,31,224,30,151,31,208,31,122,31,122,30,80,31,254,31,254,30,186,31,186,30,54,31,145,31,13,31,192,31,41,31,140,31,140,30,147,31,105,31,18,31,2,31,37,31,42,31,71,31,71,30,237,31,183,31,203,31,203,30,57,31,248,31,119,31,119,30,112,31,122,31,93,31,17,31,83,31,78,31,157,31,217,31,217,30,173,31,104,31,38,31,38,30,26,31,103,31,190,31,234,31,76,31,125,31,223,31,176,31,65,31,28,31,232,31,42,31,80,31,128,31,81,31,181,31,130,31,65,31,226,31,81,31,141,31,118,31,177,31,245,31,174,31,234,31,97,31,30,31,176,31,138,31,125,31,63,31,198,31,98,31,32,31,62,31,232,31,87,31,222,31,61,31,178,31,80,31,80,30,31,31,148,31,17,31,3,31,3,30,47,31,133,31,163,31,163,30,247,31,54,31,116,31,177,31,208,31,82,31,173,31,11,31,41,31,53,31,13,31,160,31,94,31,94,30,116,31,129,31,85,31,94,31,94,30,230,31,22,31,102,31,151,31,13,31,131,31,62,31,52,31,20,31,120,31,76,31,202,31,207,31,227,31,227,30,2,31,17,31,177,31,215,31,91,31,103,31,16,31,7,31,66,31,66,30,177,31,129,31,22,31,115,31,115,30,115,29,115,28,115,27,116,31,172,31,178,31,142,31,177,31,189,31,103,31,171,31,248,31,3,31,189,31,18,31,18,30,95,31,158,31,158,30,11,31,53,31,144,31,20,31,20,30,30,31,82,31,25,31,172,31,235,31,235,30,148,31,148,30,243,31,66,31,2,31,48,31,217,31,131,31,169,31,169,30,169,29,233,31,94,31,94,30,255,31,16,31,181,31,181,30,181,29,112,31,112,30,112,29,112,28,112,27,245,31,131,31,17,31,100,31,21,31,212,31,145,31,158,31,175,31,219,31,251,31,103,31,73,31,73,30,13,31,13,30,165,31,106,31,79,31,79,30,136,31,240,31,251,31,233,31,57,31,211,31,90,31,21,31,187,31,187,30,201,31,227,31,250,31,6,31,216,31,213,31,125,31,125,30,94,31,223,31,223,30,223,29,73,31,251,31,89,31,36,31,184,31,252,31,251,31,210,31,166,31,175,31,175,30,175,29,123,31,245,31,117,31,174,31,143,31,156,31,114,31,96,31,96,30,96,29,117,31,117,30,15,31,56,31,160,31,160,30,239,31,6,31,139,31,37,31,37,30,44,31,44,30,217,31,217,30,217,29,10,31,10,30,53,31,53,30,33,31,41,31,8,31,46,31,79,31,47,31,129,31,66,31,119,31,138,31,96,31,158,31,138,31,65,31,230,31,230,30,7,31,116,31,105,31,127,31,33,31,247,31,216,31,214,31,10,31,10,30,151,31,176,31,73,31,73,30,172,31,189,31,189,30,83,31,83,30,211,31,116,31,167,31,167,30,93,31,168,31,103,31,40,31,134,31,219,31,27,31,27,30,221,31,221,30,101,31,202,31,140,31,20,31,250,31,95,31,3,31,206,31,246,31,115,31,120,31,135,31,2,31,253,31,103,31,103,30,175,31,1,31,32,31,150,31,150,30,244,31,76,31,76,30,55,31,55,30,209,31,209,30,8,31,41,31,30,31,6,31,94,31,199,31,199,30,24,31,50,31,171,31,113,31,77,31,77,30,251,31,64,31,13,31,168,31,155,31,226,31,32,31,63,31,19,31,103,31,17,31,113,31,125,31,8,31,164,31,164,30,164,29,63,31,245,31,110,31,191,31,82,31,68,31,56,31,191,31,159,31,238,31,105,31,90,31,220,31,220,30,111,31,77,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
