-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 847;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,139,0,77,0,2,0,86,0,11,0,201,0,92,0,164,0,0,0,0,0,118,0,0,0,16,0,8,0,10,0,191,0,36,0,42,0,32,0,0,0,25,0,238,0,202,0,8,0,0,0,208,0,72,0,33,0,85,0,34,0,0,0,131,0,0,0,12,0,155,0,5,0,41,0,108,0,104,0,4,0,114,0,205,0,248,0,0,0,0,0,249,0,87,0,0,0,131,0,0,0,129,0,34,0,0,0,25,0,0,0,94,0,194,0,99,0,186,0,160,0,145,0,219,0,226,0,33,0,0,0,0,0,227,0,63,0,0,0,221,0,0,0,32,0,46,0,215,0,181,0,0,0,0,0,96,0,170,0,203,0,246,0,138,0,34,0,123,0,44,0,0,0,0,0,0,0,0,0,28,0,40,0,199,0,47,0,91,0,0,0,8,0,228,0,0,0,135,0,203,0,55,0,197,0,81,0,0,0,175,0,59,0,232,0,96,0,135,0,0,0,241,0,49,0,0,0,64,0,197,0,210,0,63,0,146,0,0,0,250,0,254,0,149,0,92,0,111,0,61,0,148,0,68,0,10,0,79,0,147,0,120,0,158,0,219,0,208,0,10,0,44,0,0,0,184,0,0,0,173,0,228,0,9,0,158,0,252,0,164,0,44,0,55,0,238,0,33,0,107,0,199,0,0,0,134,0,117,0,15,0,246,0,2,0,0,0,57,0,233,0,0,0,80,0,18,0,34,0,83,0,0,0,105,0,0,0,101,0,229,0,0,0,122,0,32,0,0,0,58,0,36,0,0,0,224,0,0,0,93,0,0,0,0,0,95,0,210,0,250,0,133,0,174,0,0,0,0,0,210,0,118,0,167,0,0,0,65,0,173,0,140,0,62,0,94,0,17,0,148,0,0,0,0,0,214,0,189,0,209,0,0,0,18,0,55,0,229,0,142,0,9,0,216,0,228,0,46,0,93,0,171,0,124,0,65,0,164,0,0,0,199,0,238,0,0,0,63,0,179,0,0,0,25,0,60,0,0,0,185,0,18,0,57,0,52,0,237,0,49,0,102,0,0,0,116,0,28,0,0,0,0,0,252,0,139,0,68,0,194,0,173,0,88,0,0,0,61,0,68,0,204,0,23,0,0,0,21,0,228,0,231,0,119,0,121,0,38,0,78,0,101,0,188,0,67,0,74,0,131,0,243,0,231,0,106,0,0,0,0,0,238,0,122,0,2,0,198,0,234,0,86,0,254,0,122,0,229,0,0,0,52,0,36,0,0,0,0,0,0,0,73,0,109,0,43,0,218,0,249,0,197,0,132,0,74,0,32,0,163,0,202,0,40,0,189,0,66,0,145,0,198,0,244,0,0,0,247,0,68,0,0,0,0,0,0,0,250,0,0,0,0,0,99,0,98,0,81,0,84,0,33,0,165,0,0,0,103,0,0,0,188,0,116,0,171,0,0,0,116,0,0,0,0,0,190,0,199,0,19,0,85,0,104,0,248,0,165,0,32,0,132,0,230,0,126,0,45,0,16,0,44,0,147,0,0,0,150,0,187,0,0,0,155,0,97,0,238,0,54,0,24,0,53,0,30,0,136,0,64,0,226,0,7,0,89,0,0,0,76,0,96,0,6,0,73,0,161,0,66,0,0,0,129,0,182,0,0,0,144,0,169,0,52,0,135,0,62,0,50,0,159,0,17,0,133,0,127,0,234,0,223,0,6,0,128,0,178,0,12,0,10,0,191,0,0,0,162,0,175,0,190,0,122,0,0,0,36,0,222,0,0,0,164,0,220,0,221,0,11,0,0,0,219,0,169,0,234,0,178,0,0,0,18,0,183,0,31,0,103,0,41,0,220,0,0,0,89,0,134,0,0,0,0,0,0,0,0,0,0,0,0,0,91,0,0,0,120,0,221,0,0,0,228,0,50,0,0,0,227,0,0,0,130,0,0,0,38,0,26,0,163,0,87,0,237,0,0,0,188,0,106,0,233,0,115,0,150,0,47,0,0,0,23,0,0,0,204,0,99,0,184,0,0,0,129,0,195,0,23,0,0,0,0,0,20,0,246,0,170,0,0,0,0,0,66,0,101,0,177,0,38,0,221,0,104,0,66,0,0,0,4,0,25,0,226,0,152,0,123,0,40,0,228,0,0,0,116,0,199,0,24,0,0,0,1,0,0,0,0,0,0,0,53,0,57,0,47,0,0,0,118,0,4,0,0,0,104,0,230,0,9,0,0,0,193,0,115,0,0,0,143,0,0,0,166,0,144,0,135,0,68,0,161,0,0,0,206,0,113,0,6,0,165,0,0,0,212,0,189,0,147,0,94,0,7,0,0,0,21,0,81,0,0,0,168,0,122,0,251,0,0,0,84,0,102,0,0,0,172,0,0,0,122,0,128,0,108,0,228,0,0,0,24,0,93,0,41,0,152,0,89,0,160,0,222,0,196,0,205,0,195,0,117,0,81,0,50,0,0,0,174,0,91,0,219,0,184,0,0,0,33,0,196,0,0,0,0,0,170,0,0,0,105,0,68,0,68,0,132,0,212,0,0,0,80,0,203,0,64,0,199,0,0,0,2,0,77,0,0,0,241,0,239,0,0,0,62,0,128,0,67,0,175,0,95,0,109,0,209,0,8,0,180,0,35,0,0,0,131,0,44,0,89,0,174,0,52,0,98,0,0,0,244,0,244,0,180,0,158,0,152,0,235,0,105,0,0,0,0,0,29,0,0,0,96,0,108,0,112,0,102,0,57,0,197,0,0,0,245,0,48,0,115,0,163,0,103,0,43,0,78,0,74,0,149,0,0,0,79,0,93,0,182,0,84,0,24,0,185,0,28,0,116,0,0,0,0,0,249,0,112,0,224,0,0,0,112,0,144,0,156,0,217,0,0,0,226,0,150,0,25,0,216,0,177,0,112,0,0,0,113,0,32,0,0,0,86,0,54,0,240,0,87,0,58,0,101,0,91,0,68,0,118,0,217,0,51,0,0,0,48,0,49,0,168,0,74,0,121,0,0,0,0,0,63,0,209,0,0,0,200,0,128,0,183,0,134,0,200,0,166,0,247,0,221,0,0,0,105,0,123,0,36,0,226,0,115,0,0,0,87,0,0,0,235,0,139,0,29,0,181,0,185,0,0,0,194,0,217,0,164,0,187,0,246,0,216,0,223,0,163,0,15,0,232,0,129,0,0,0,109,0,0,0,85,0,148,0,83,0,177,0,128,0,8,0,60,0,107,0,156,0,38,0,70,0,56,0,96,0,162,0,91,0,160,0,84,0,176,0,0,0,118,0,56,0,210,0,53,0,252,0,128,0,143,0,129,0,155,0,200,0,193,0,0,0,53,0,103,0,173,0,132,0,0,0,60,0,0,0,156,0,0,0,148,0,78,0,65,0,0,0,5,0,252,0,121,0,146,0,198,0,8,0,244,0,6,0,91,0,0,0,211,0,0,0,252,0,243,0,139,0,115,0,37,0,196,0,111,0,0,0,180,0,101,0,183,0,0,0,198,0,0,0,0,0,0,0,0,0,84,0,43,0,0,0,0,0,110,0,163,0,252,0,154,0,0,0,62,0,242,0,181,0,142,0,86,0,163,0,102,0,0,0,220,0,253,0,152,0,196,0,130,0,4,0,150,0,226,0,125,0,33,0,135,0,102,0,153,0,229,0,0,0,198,0,251,0,76,0,0,0,36,0,120,0,70,0,103,0,89,0,0,0,92,0,57,0,0,0,80,0,75,0,117,0,85,0,165,0,153,0,116,0,0,0,0,0,0,0,170,0,148,0,0,0,243,0,117,0,219,0);
signal scenario_full  : scenario_type := (0,0,139,31,77,31,2,31,86,31,11,31,201,31,92,31,164,31,164,30,164,29,118,31,118,30,16,31,8,31,10,31,191,31,36,31,42,31,32,31,32,30,25,31,238,31,202,31,8,31,8,30,208,31,72,31,33,31,85,31,34,31,34,30,131,31,131,30,12,31,155,31,5,31,41,31,108,31,104,31,4,31,114,31,205,31,248,31,248,30,248,29,249,31,87,31,87,30,131,31,131,30,129,31,34,31,34,30,25,31,25,30,94,31,194,31,99,31,186,31,160,31,145,31,219,31,226,31,33,31,33,30,33,29,227,31,63,31,63,30,221,31,221,30,32,31,46,31,215,31,181,31,181,30,181,29,96,31,170,31,203,31,246,31,138,31,34,31,123,31,44,31,44,30,44,29,44,28,44,27,28,31,40,31,199,31,47,31,91,31,91,30,8,31,228,31,228,30,135,31,203,31,55,31,197,31,81,31,81,30,175,31,59,31,232,31,96,31,135,31,135,30,241,31,49,31,49,30,64,31,197,31,210,31,63,31,146,31,146,30,250,31,254,31,149,31,92,31,111,31,61,31,148,31,68,31,10,31,79,31,147,31,120,31,158,31,219,31,208,31,10,31,44,31,44,30,184,31,184,30,173,31,228,31,9,31,158,31,252,31,164,31,44,31,55,31,238,31,33,31,107,31,199,31,199,30,134,31,117,31,15,31,246,31,2,31,2,30,57,31,233,31,233,30,80,31,18,31,34,31,83,31,83,30,105,31,105,30,101,31,229,31,229,30,122,31,32,31,32,30,58,31,36,31,36,30,224,31,224,30,93,31,93,30,93,29,95,31,210,31,250,31,133,31,174,31,174,30,174,29,210,31,118,31,167,31,167,30,65,31,173,31,140,31,62,31,94,31,17,31,148,31,148,30,148,29,214,31,189,31,209,31,209,30,18,31,55,31,229,31,142,31,9,31,216,31,228,31,46,31,93,31,171,31,124,31,65,31,164,31,164,30,199,31,238,31,238,30,63,31,179,31,179,30,25,31,60,31,60,30,185,31,18,31,57,31,52,31,237,31,49,31,102,31,102,30,116,31,28,31,28,30,28,29,252,31,139,31,68,31,194,31,173,31,88,31,88,30,61,31,68,31,204,31,23,31,23,30,21,31,228,31,231,31,119,31,121,31,38,31,78,31,101,31,188,31,67,31,74,31,131,31,243,31,231,31,106,31,106,30,106,29,238,31,122,31,2,31,198,31,234,31,86,31,254,31,122,31,229,31,229,30,52,31,36,31,36,30,36,29,36,28,73,31,109,31,43,31,218,31,249,31,197,31,132,31,74,31,32,31,163,31,202,31,40,31,189,31,66,31,145,31,198,31,244,31,244,30,247,31,68,31,68,30,68,29,68,28,250,31,250,30,250,29,99,31,98,31,81,31,84,31,33,31,165,31,165,30,103,31,103,30,188,31,116,31,171,31,171,30,116,31,116,30,116,29,190,31,199,31,19,31,85,31,104,31,248,31,165,31,32,31,132,31,230,31,126,31,45,31,16,31,44,31,147,31,147,30,150,31,187,31,187,30,155,31,97,31,238,31,54,31,24,31,53,31,30,31,136,31,64,31,226,31,7,31,89,31,89,30,76,31,96,31,6,31,73,31,161,31,66,31,66,30,129,31,182,31,182,30,144,31,169,31,52,31,135,31,62,31,50,31,159,31,17,31,133,31,127,31,234,31,223,31,6,31,128,31,178,31,12,31,10,31,191,31,191,30,162,31,175,31,190,31,122,31,122,30,36,31,222,31,222,30,164,31,220,31,221,31,11,31,11,30,219,31,169,31,234,31,178,31,178,30,18,31,183,31,31,31,103,31,41,31,220,31,220,30,89,31,134,31,134,30,134,29,134,28,134,27,134,26,134,25,91,31,91,30,120,31,221,31,221,30,228,31,50,31,50,30,227,31,227,30,130,31,130,30,38,31,26,31,163,31,87,31,237,31,237,30,188,31,106,31,233,31,115,31,150,31,47,31,47,30,23,31,23,30,204,31,99,31,184,31,184,30,129,31,195,31,23,31,23,30,23,29,20,31,246,31,170,31,170,30,170,29,66,31,101,31,177,31,38,31,221,31,104,31,66,31,66,30,4,31,25,31,226,31,152,31,123,31,40,31,228,31,228,30,116,31,199,31,24,31,24,30,1,31,1,30,1,29,1,28,53,31,57,31,47,31,47,30,118,31,4,31,4,30,104,31,230,31,9,31,9,30,193,31,115,31,115,30,143,31,143,30,166,31,144,31,135,31,68,31,161,31,161,30,206,31,113,31,6,31,165,31,165,30,212,31,189,31,147,31,94,31,7,31,7,30,21,31,81,31,81,30,168,31,122,31,251,31,251,30,84,31,102,31,102,30,172,31,172,30,122,31,128,31,108,31,228,31,228,30,24,31,93,31,41,31,152,31,89,31,160,31,222,31,196,31,205,31,195,31,117,31,81,31,50,31,50,30,174,31,91,31,219,31,184,31,184,30,33,31,196,31,196,30,196,29,170,31,170,30,105,31,68,31,68,31,132,31,212,31,212,30,80,31,203,31,64,31,199,31,199,30,2,31,77,31,77,30,241,31,239,31,239,30,62,31,128,31,67,31,175,31,95,31,109,31,209,31,8,31,180,31,35,31,35,30,131,31,44,31,89,31,174,31,52,31,98,31,98,30,244,31,244,31,180,31,158,31,152,31,235,31,105,31,105,30,105,29,29,31,29,30,96,31,108,31,112,31,102,31,57,31,197,31,197,30,245,31,48,31,115,31,163,31,103,31,43,31,78,31,74,31,149,31,149,30,79,31,93,31,182,31,84,31,24,31,185,31,28,31,116,31,116,30,116,29,249,31,112,31,224,31,224,30,112,31,144,31,156,31,217,31,217,30,226,31,150,31,25,31,216,31,177,31,112,31,112,30,113,31,32,31,32,30,86,31,54,31,240,31,87,31,58,31,101,31,91,31,68,31,118,31,217,31,51,31,51,30,48,31,49,31,168,31,74,31,121,31,121,30,121,29,63,31,209,31,209,30,200,31,128,31,183,31,134,31,200,31,166,31,247,31,221,31,221,30,105,31,123,31,36,31,226,31,115,31,115,30,87,31,87,30,235,31,139,31,29,31,181,31,185,31,185,30,194,31,217,31,164,31,187,31,246,31,216,31,223,31,163,31,15,31,232,31,129,31,129,30,109,31,109,30,85,31,148,31,83,31,177,31,128,31,8,31,60,31,107,31,156,31,38,31,70,31,56,31,96,31,162,31,91,31,160,31,84,31,176,31,176,30,118,31,56,31,210,31,53,31,252,31,128,31,143,31,129,31,155,31,200,31,193,31,193,30,53,31,103,31,173,31,132,31,132,30,60,31,60,30,156,31,156,30,148,31,78,31,65,31,65,30,5,31,252,31,121,31,146,31,198,31,8,31,244,31,6,31,91,31,91,30,211,31,211,30,252,31,243,31,139,31,115,31,37,31,196,31,111,31,111,30,180,31,101,31,183,31,183,30,198,31,198,30,198,29,198,28,198,27,84,31,43,31,43,30,43,29,110,31,163,31,252,31,154,31,154,30,62,31,242,31,181,31,142,31,86,31,163,31,102,31,102,30,220,31,253,31,152,31,196,31,130,31,4,31,150,31,226,31,125,31,33,31,135,31,102,31,153,31,229,31,229,30,198,31,251,31,76,31,76,30,36,31,120,31,70,31,103,31,89,31,89,30,92,31,57,31,57,30,80,31,75,31,117,31,85,31,165,31,153,31,116,31,116,30,116,29,116,28,170,31,148,31,148,30,243,31,117,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
