-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_122 is
end project_tb_122;

architecture project_tb_arch_122 of project_tb_122 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 167;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,19,0,192,0,176,0,151,0,0,0,0,0,33,0,0,0,41,0,200,0,0,0,115,0,212,0,196,0,6,0,172,0,104,0,73,0,224,0,218,0,185,0,156,0,154,0,71,0,169,0,29,0,143,0,99,0,0,0,227,0,0,0,60,0,167,0,59,0,26,0,95,0,0,0,89,0,196,0,208,0,15,0,171,0,10,0,154,0,0,0,48,0,51,0,35,0,203,0,104,0,82,0,146,0,0,0,169,0,216,0,141,0,53,0,45,0,69,0,246,0,0,0,0,0,68,0,55,0,0,0,241,0,159,0,136,0,93,0,135,0,0,0,111,0,111,0,225,0,142,0,127,0,42,0,128,0,0,0,14,0,122,0,54,0,101,0,31,0,0,0,217,0,234,0,114,0,114,0,106,0,172,0,140,0,53,0,0,0,170,0,33,0,101,0,66,0,92,0,161,0,111,0,95,0,188,0,0,0,155,0,151,0,185,0,0,0,135,0,77,0,226,0,0,0,242,0,113,0,203,0,182,0,1,0,155,0,0,0,22,0,158,0,0,0,222,0,56,0,212,0,79,0,171,0,52,0,30,0,0,0,0,0,0,0,85,0,184,0,76,0,171,0,222,0,108,0,165,0,190,0,137,0,157,0,72,0,172,0,72,0,92,0,182,0,219,0,0,0,17,0,169,0,0,0,223,0,24,0,188,0,0,0,189,0,0,0,0,0,138,0,0,0,53,0,122,0,49,0,0,0,7,0);
signal scenario_full  : scenario_type := (0,0,19,31,192,31,176,31,151,31,151,30,151,29,33,31,33,30,41,31,200,31,200,30,115,31,212,31,196,31,6,31,172,31,104,31,73,31,224,31,218,31,185,31,156,31,154,31,71,31,169,31,29,31,143,31,99,31,99,30,227,31,227,30,60,31,167,31,59,31,26,31,95,31,95,30,89,31,196,31,208,31,15,31,171,31,10,31,154,31,154,30,48,31,51,31,35,31,203,31,104,31,82,31,146,31,146,30,169,31,216,31,141,31,53,31,45,31,69,31,246,31,246,30,246,29,68,31,55,31,55,30,241,31,159,31,136,31,93,31,135,31,135,30,111,31,111,31,225,31,142,31,127,31,42,31,128,31,128,30,14,31,122,31,54,31,101,31,31,31,31,30,217,31,234,31,114,31,114,31,106,31,172,31,140,31,53,31,53,30,170,31,33,31,101,31,66,31,92,31,161,31,111,31,95,31,188,31,188,30,155,31,151,31,185,31,185,30,135,31,77,31,226,31,226,30,242,31,113,31,203,31,182,31,1,31,155,31,155,30,22,31,158,31,158,30,222,31,56,31,212,31,79,31,171,31,52,31,30,31,30,30,30,29,30,28,85,31,184,31,76,31,171,31,222,31,108,31,165,31,190,31,137,31,157,31,72,31,172,31,72,31,92,31,182,31,219,31,219,30,17,31,169,31,169,30,223,31,24,31,188,31,188,30,189,31,189,30,189,29,138,31,138,30,53,31,122,31,49,31,49,30,7,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
