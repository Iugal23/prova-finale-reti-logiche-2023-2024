-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_9 is
end project_tb_9;

architecture project_tb_arch_9 of project_tb_9 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 783;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (25,0,39,0,200,0,226,0,228,0,0,0,213,0,8,0,0,0,125,0,3,0,193,0,247,0,11,0,69,0,0,0,27,0,205,0,246,0,10,0,50,0,33,0,186,0,0,0,244,0,79,0,121,0,0,0,239,0,51,0,0,0,123,0,0,0,179,0,101,0,190,0,204,0,0,0,182,0,91,0,73,0,68,0,70,0,73,0,107,0,57,0,0,0,0,0,0,0,0,0,0,0,91,0,132,0,19,0,0,0,37,0,140,0,17,0,130,0,0,0,177,0,82,0,224,0,4,0,0,0,201,0,40,0,40,0,233,0,27,0,41,0,99,0,15,0,218,0,228,0,0,0,219,0,134,0,182,0,63,0,147,0,73,0,31,0,0,0,161,0,113,0,131,0,84,0,27,0,107,0,211,0,250,0,0,0,0,0,159,0,121,0,0,0,3,0,211,0,0,0,110,0,0,0,156,0,0,0,77,0,86,0,242,0,0,0,138,0,55,0,4,0,163,0,103,0,143,0,177,0,29,0,71,0,117,0,36,0,88,0,0,0,65,0,255,0,27,0,84,0,5,0,0,0,39,0,157,0,35,0,203,0,5,0,144,0,254,0,112,0,237,0,102,0,10,0,0,0,48,0,124,0,222,0,250,0,0,0,204,0,176,0,212,0,251,0,66,0,197,0,211,0,202,0,0,0,253,0,43,0,0,0,194,0,87,0,98,0,163,0,13,0,0,0,147,0,3,0,0,0,230,0,0,0,134,0,0,0,0,0,164,0,230,0,158,0,91,0,0,0,63,0,127,0,88,0,149,0,30,0,0,0,135,0,78,0,0,0,139,0,0,0,162,0,88,0,251,0,236,0,31,0,218,0,112,0,255,0,186,0,29,0,125,0,194,0,139,0,205,0,110,0,62,0,121,0,212,0,221,0,0,0,0,0,132,0,65,0,94,0,52,0,0,0,117,0,154,0,0,0,212,0,69,0,186,0,81,0,0,0,169,0,22,0,47,0,0,0,0,0,164,0,157,0,199,0,180,0,0,0,85,0,14,0,156,0,3,0,134,0,74,0,0,0,73,0,170,0,23,0,87,0,44,0,25,0,199,0,125,0,195,0,66,0,88,0,17,0,158,0,133,0,197,0,92,0,182,0,141,0,82,0,138,0,226,0,163,0,105,0,152,0,215,0,131,0,0,0,66,0,157,0,123,0,110,0,216,0,155,0,5,0,0,0,43,0,36,0,234,0,151,0,139,0,0,0,161,0,185,0,33,0,171,0,0,0,57,0,44,0,252,0,190,0,56,0,6,0,107,0,15,0,14,0,169,0,229,0,129,0,0,0,12,0,0,0,129,0,185,0,158,0,109,0,235,0,87,0,73,0,0,0,2,0,0,0,192,0,108,0,71,0,63,0,185,0,0,0,236,0,0,0,143,0,150,0,251,0,22,0,0,0,87,0,87,0,135,0,132,0,0,0,230,0,128,0,84,0,81,0,235,0,206,0,51,0,87,0,0,0,227,0,0,0,154,0,0,0,113,0,161,0,0,0,177,0,65,0,0,0,109,0,0,0,130,0,44,0,246,0,0,0,221,0,10,0,188,0,0,0,38,0,75,0,64,0,185,0,0,0,18,0,7,0,175,0,168,0,237,0,184,0,82,0,230,0,229,0,234,0,205,0,122,0,33,0,161,0,137,0,12,0,37,0,185,0,197,0,26,0,0,0,60,0,158,0,251,0,109,0,52,0,178,0,0,0,232,0,51,0,0,0,145,0,31,0,194,0,213,0,204,0,76,0,66,0,0,0,174,0,0,0,1,0,170,0,108,0,0,0,196,0,199,0,28,0,155,0,56,0,0,0,201,0,80,0,0,0,87,0,189,0,118,0,237,0,0,0,56,0,0,0,85,0,164,0,30,0,113,0,198,0,0,0,104,0,0,0,172,0,0,0,97,0,223,0,116,0,0,0,154,0,237,0,244,0,235,0,197,0,215,0,28,0,185,0,99,0,0,0,0,0,89,0,252,0,51,0,181,0,151,0,87,0,0,0,36,0,97,0,247,0,0,0,188,0,165,0,140,0,165,0,0,0,0,0,164,0,76,0,255,0,113,0,116,0,0,0,98,0,130,0,0,0,112,0,56,0,78,0,251,0,0,0,0,0,174,0,212,0,161,0,127,0,28,0,250,0,85,0,0,0,59,0,196,0,1,0,54,0,106,0,139,0,179,0,85,0,148,0,0,0,0,0,102,0,32,0,238,0,91,0,193,0,0,0,0,0,231,0,0,0,232,0,71,0,6,0,158,0,0,0,123,0,194,0,136,0,101,0,132,0,160,0,252,0,1,0,0,0,36,0,208,0,0,0,150,0,90,0,85,0,220,0,97,0,249,0,104,0,103,0,0,0,11,0,198,0,184,0,0,0,212,0,36,0,201,0,19,0,58,0,142,0,0,0,152,0,217,0,24,0,253,0,21,0,45,0,106,0,218,0,200,0,28,0,76,0,163,0,221,0,164,0,49,0,56,0,216,0,191,0,14,0,18,0,117,0,171,0,237,0,103,0,88,0,72,0,0,0,148,0,12,0,0,0,110,0,21,0,217,0,57,0,159,0,0,0,111,0,248,0,125,0,1,0,102,0,73,0,0,0,227,0,33,0,59,0,58,0,0,0,7,0,0,0,147,0,116,0,57,0,29,0,36,0,0,0,78,0,137,0,65,0,179,0,153,0,102,0,91,0,0,0,152,0,76,0,254,0,153,0,0,0,4,0,81,0,18,0,186,0,71,0,92,0,3,0,33,0,228,0,194,0,0,0,192,0,249,0,112,0,59,0,26,0,39,0,241,0,0,0,0,0,32,0,8,0,5,0,0,0,236,0,47,0,237,0,199,0,0,0,0,0,242,0,136,0,217,0,114,0,0,0,166,0,0,0,2,0,39,0,0,0,80,0,83,0,199,0,69,0,146,0,86,0,16,0,255,0,0,0,116,0,19,0,183,0,0,0,149,0,175,0,146,0,0,0,73,0,91,0,123,0,71,0,77,0,7,0,245,0,0,0,0,0,0,0,0,0,149,0,235,0,35,0,118,0,0,0,250,0,94,0,190,0,38,0,245,0,185,0,213,0,129,0,25,0,98,0,114,0,42,0,13,0,249,0,0,0,157,0,195,0,254,0,50,0,18,0,254,0,0,0,87,0,58,0,135,0,169,0,202,0,45,0,97,0,164,0,213,0,0,0,144,0,217,0,29,0,174,0,48,0,14,0,209,0,0,0,241,0,173,0,0,0,124,0,99,0,253,0,10,0,33,0,250,0,109,0,187,0,220,0,153,0,30,0,113,0,144,0,73,0,0,0,137,0,128,0,177,0,238,0,185,0,223,0,5,0,35,0,38,0,148,0,120,0,162,0,32,0,184,0,0,0,150,0,0,0,73,0,81,0,5,0,254,0,149,0,32,0,162,0,185,0,211,0,97,0,218,0,162,0,90,0,40,0,62,0,11,0,64,0,76,0,28,0,43,0,123,0,170,0,217,0);
signal scenario_full  : scenario_type := (25,31,39,31,200,31,226,31,228,31,228,30,213,31,8,31,8,30,125,31,3,31,193,31,247,31,11,31,69,31,69,30,27,31,205,31,246,31,10,31,50,31,33,31,186,31,186,30,244,31,79,31,121,31,121,30,239,31,51,31,51,30,123,31,123,30,179,31,101,31,190,31,204,31,204,30,182,31,91,31,73,31,68,31,70,31,73,31,107,31,57,31,57,30,57,29,57,28,57,27,57,26,91,31,132,31,19,31,19,30,37,31,140,31,17,31,130,31,130,30,177,31,82,31,224,31,4,31,4,30,201,31,40,31,40,31,233,31,27,31,41,31,99,31,15,31,218,31,228,31,228,30,219,31,134,31,182,31,63,31,147,31,73,31,31,31,31,30,161,31,113,31,131,31,84,31,27,31,107,31,211,31,250,31,250,30,250,29,159,31,121,31,121,30,3,31,211,31,211,30,110,31,110,30,156,31,156,30,77,31,86,31,242,31,242,30,138,31,55,31,4,31,163,31,103,31,143,31,177,31,29,31,71,31,117,31,36,31,88,31,88,30,65,31,255,31,27,31,84,31,5,31,5,30,39,31,157,31,35,31,203,31,5,31,144,31,254,31,112,31,237,31,102,31,10,31,10,30,48,31,124,31,222,31,250,31,250,30,204,31,176,31,212,31,251,31,66,31,197,31,211,31,202,31,202,30,253,31,43,31,43,30,194,31,87,31,98,31,163,31,13,31,13,30,147,31,3,31,3,30,230,31,230,30,134,31,134,30,134,29,164,31,230,31,158,31,91,31,91,30,63,31,127,31,88,31,149,31,30,31,30,30,135,31,78,31,78,30,139,31,139,30,162,31,88,31,251,31,236,31,31,31,218,31,112,31,255,31,186,31,29,31,125,31,194,31,139,31,205,31,110,31,62,31,121,31,212,31,221,31,221,30,221,29,132,31,65,31,94,31,52,31,52,30,117,31,154,31,154,30,212,31,69,31,186,31,81,31,81,30,169,31,22,31,47,31,47,30,47,29,164,31,157,31,199,31,180,31,180,30,85,31,14,31,156,31,3,31,134,31,74,31,74,30,73,31,170,31,23,31,87,31,44,31,25,31,199,31,125,31,195,31,66,31,88,31,17,31,158,31,133,31,197,31,92,31,182,31,141,31,82,31,138,31,226,31,163,31,105,31,152,31,215,31,131,31,131,30,66,31,157,31,123,31,110,31,216,31,155,31,5,31,5,30,43,31,36,31,234,31,151,31,139,31,139,30,161,31,185,31,33,31,171,31,171,30,57,31,44,31,252,31,190,31,56,31,6,31,107,31,15,31,14,31,169,31,229,31,129,31,129,30,12,31,12,30,129,31,185,31,158,31,109,31,235,31,87,31,73,31,73,30,2,31,2,30,192,31,108,31,71,31,63,31,185,31,185,30,236,31,236,30,143,31,150,31,251,31,22,31,22,30,87,31,87,31,135,31,132,31,132,30,230,31,128,31,84,31,81,31,235,31,206,31,51,31,87,31,87,30,227,31,227,30,154,31,154,30,113,31,161,31,161,30,177,31,65,31,65,30,109,31,109,30,130,31,44,31,246,31,246,30,221,31,10,31,188,31,188,30,38,31,75,31,64,31,185,31,185,30,18,31,7,31,175,31,168,31,237,31,184,31,82,31,230,31,229,31,234,31,205,31,122,31,33,31,161,31,137,31,12,31,37,31,185,31,197,31,26,31,26,30,60,31,158,31,251,31,109,31,52,31,178,31,178,30,232,31,51,31,51,30,145,31,31,31,194,31,213,31,204,31,76,31,66,31,66,30,174,31,174,30,1,31,170,31,108,31,108,30,196,31,199,31,28,31,155,31,56,31,56,30,201,31,80,31,80,30,87,31,189,31,118,31,237,31,237,30,56,31,56,30,85,31,164,31,30,31,113,31,198,31,198,30,104,31,104,30,172,31,172,30,97,31,223,31,116,31,116,30,154,31,237,31,244,31,235,31,197,31,215,31,28,31,185,31,99,31,99,30,99,29,89,31,252,31,51,31,181,31,151,31,87,31,87,30,36,31,97,31,247,31,247,30,188,31,165,31,140,31,165,31,165,30,165,29,164,31,76,31,255,31,113,31,116,31,116,30,98,31,130,31,130,30,112,31,56,31,78,31,251,31,251,30,251,29,174,31,212,31,161,31,127,31,28,31,250,31,85,31,85,30,59,31,196,31,1,31,54,31,106,31,139,31,179,31,85,31,148,31,148,30,148,29,102,31,32,31,238,31,91,31,193,31,193,30,193,29,231,31,231,30,232,31,71,31,6,31,158,31,158,30,123,31,194,31,136,31,101,31,132,31,160,31,252,31,1,31,1,30,36,31,208,31,208,30,150,31,90,31,85,31,220,31,97,31,249,31,104,31,103,31,103,30,11,31,198,31,184,31,184,30,212,31,36,31,201,31,19,31,58,31,142,31,142,30,152,31,217,31,24,31,253,31,21,31,45,31,106,31,218,31,200,31,28,31,76,31,163,31,221,31,164,31,49,31,56,31,216,31,191,31,14,31,18,31,117,31,171,31,237,31,103,31,88,31,72,31,72,30,148,31,12,31,12,30,110,31,21,31,217,31,57,31,159,31,159,30,111,31,248,31,125,31,1,31,102,31,73,31,73,30,227,31,33,31,59,31,58,31,58,30,7,31,7,30,147,31,116,31,57,31,29,31,36,31,36,30,78,31,137,31,65,31,179,31,153,31,102,31,91,31,91,30,152,31,76,31,254,31,153,31,153,30,4,31,81,31,18,31,186,31,71,31,92,31,3,31,33,31,228,31,194,31,194,30,192,31,249,31,112,31,59,31,26,31,39,31,241,31,241,30,241,29,32,31,8,31,5,31,5,30,236,31,47,31,237,31,199,31,199,30,199,29,242,31,136,31,217,31,114,31,114,30,166,31,166,30,2,31,39,31,39,30,80,31,83,31,199,31,69,31,146,31,86,31,16,31,255,31,255,30,116,31,19,31,183,31,183,30,149,31,175,31,146,31,146,30,73,31,91,31,123,31,71,31,77,31,7,31,245,31,245,30,245,29,245,28,245,27,149,31,235,31,35,31,118,31,118,30,250,31,94,31,190,31,38,31,245,31,185,31,213,31,129,31,25,31,98,31,114,31,42,31,13,31,249,31,249,30,157,31,195,31,254,31,50,31,18,31,254,31,254,30,87,31,58,31,135,31,169,31,202,31,45,31,97,31,164,31,213,31,213,30,144,31,217,31,29,31,174,31,48,31,14,31,209,31,209,30,241,31,173,31,173,30,124,31,99,31,253,31,10,31,33,31,250,31,109,31,187,31,220,31,153,31,30,31,113,31,144,31,73,31,73,30,137,31,128,31,177,31,238,31,185,31,223,31,5,31,35,31,38,31,148,31,120,31,162,31,32,31,184,31,184,30,150,31,150,30,73,31,81,31,5,31,254,31,149,31,32,31,162,31,185,31,211,31,97,31,218,31,162,31,90,31,40,31,62,31,11,31,64,31,76,31,28,31,43,31,123,31,170,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
