-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 828;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,186,0,22,0,0,0,163,0,57,0,14,0,0,0,141,0,238,0,93,0,55,0,178,0,0,0,0,0,86,0,236,0,161,0,48,0,12,0,97,0,210,0,0,0,40,0,218,0,77,0,41,0,83,0,100,0,0,0,27,0,3,0,196,0,207,0,134,0,158,0,45,0,153,0,30,0,201,0,243,0,137,0,173,0,112,0,0,0,208,0,198,0,93,0,63,0,12,0,142,0,0,0,44,0,135,0,80,0,231,0,0,0,110,0,75,0,12,0,29,0,0,0,82,0,13,0,0,0,0,0,180,0,226,0,245,0,179,0,51,0,43,0,24,0,223,0,168,0,1,0,249,0,126,0,188,0,0,0,222,0,3,0,219,0,130,0,36,0,64,0,4,0,45,0,250,0,48,0,127,0,84,0,0,0,204,0,43,0,138,0,109,0,181,0,58,0,131,0,190,0,104,0,229,0,62,0,197,0,20,0,0,0,24,0,80,0,119,0,0,0,0,0,220,0,161,0,105,0,29,0,77,0,0,0,32,0,0,0,228,0,207,0,225,0,0,0,230,0,161,0,0,0,172,0,154,0,153,0,145,0,0,0,68,0,158,0,219,0,0,0,59,0,154,0,179,0,141,0,62,0,0,0,0,0,0,0,0,0,0,0,250,0,7,0,3,0,216,0,0,0,164,0,42,0,191,0,92,0,0,0,170,0,135,0,133,0,13,0,73,0,57,0,0,0,124,0,52,0,0,0,0,0,59,0,0,0,3,0,123,0,99,0,0,0,0,0,0,0,68,0,69,0,233,0,137,0,59,0,143,0,103,0,223,0,107,0,143,0,0,0,0,0,134,0,31,0,61,0,20,0,68,0,222,0,140,0,115,0,191,0,157,0,162,0,0,0,241,0,16,0,0,0,247,0,117,0,73,0,23,0,163,0,27,0,185,0,0,0,4,0,253,0,250,0,0,0,73,0,124,0,250,0,97,0,141,0,176,0,175,0,241,0,86,0,0,0,0,0,0,0,67,0,3,0,42,0,217,0,252,0,180,0,0,0,223,0,245,0,35,0,231,0,0,0,222,0,132,0,214,0,255,0,201,0,70,0,225,0,153,0,45,0,100,0,208,0,0,0,0,0,172,0,64,0,149,0,49,0,205,0,26,0,201,0,0,0,143,0,86,0,95,0,0,0,228,0,79,0,0,0,242,0,103,0,89,0,0,0,214,0,0,0,0,0,93,0,1,0,50,0,8,0,52,0,23,0,107,0,121,0,176,0,29,0,0,0,156,0,0,0,141,0,177,0,203,0,208,0,113,0,214,0,254,0,24,0,0,0,28,0,167,0,217,0,191,0,0,0,255,0,0,0,9,0,0,0,251,0,244,0,78,0,187,0,51,0,192,0,61,0,110,0,171,0,82,0,131,0,98,0,63,0,105,0,57,0,72,0,234,0,227,0,112,0,73,0,220,0,1,0,242,0,11,0,181,0,220,0,178,0,149,0,128,0,163,0,182,0,43,0,186,0,10,0,124,0,61,0,201,0,85,0,15,0,48,0,192,0,250,0,192,0,242,0,0,0,55,0,226,0,0,0,144,0,80,0,175,0,51,0,48,0,176,0,205,0,28,0,195,0,176,0,37,0,222,0,174,0,235,0,118,0,139,0,155,0,0,0,142,0,212,0,121,0,28,0,153,0,165,0,161,0,200,0,20,0,185,0,244,0,244,0,97,0,143,0,164,0,115,0,17,0,110,0,236,0,236,0,197,0,5,0,138,0,111,0,0,0,147,0,165,0,181,0,235,0,87,0,0,0,15,0,130,0,0,0,0,0,0,0,182,0,19,0,154,0,227,0,19,0,71,0,42,0,0,0,32,0,238,0,0,0,255,0,213,0,175,0,6,0,0,0,161,0,93,0,82,0,162,0,0,0,216,0,127,0,32,0,226,0,72,0,243,0,13,0,65,0,89,0,221,0,233,0,55,0,0,0,105,0,20,0,39,0,210,0,122,0,35,0,3,0,164,0,0,0,171,0,126,0,26,0,32,0,0,0,209,0,0,0,0,0,167,0,57,0,119,0,144,0,185,0,236,0,112,0,14,0,90,0,0,0,50,0,35,0,12,0,47,0,0,0,139,0,192,0,65,0,20,0,66,0,0,0,107,0,0,0,0,0,114,0,85,0,174,0,47,0,0,0,22,0,250,0,29,0,39,0,103,0,53,0,68,0,142,0,220,0,140,0,137,0,18,0,205,0,247,0,41,0,162,0,157,0,0,0,61,0,243,0,0,0,177,0,45,0,217,0,56,0,206,0,0,0,234,0,177,0,157,0,13,0,0,0,58,0,0,0,0,0,32,0,30,0,39,0,156,0,4,0,69,0,231,0,242,0,62,0,48,0,100,0,0,0,241,0,0,0,93,0,229,0,85,0,81,0,187,0,153,0,240,0,114,0,242,0,0,0,249,0,107,0,6,0,178,0,0,0,0,0,102,0,0,0,221,0,0,0,211,0,70,0,65,0,232,0,0,0,96,0,41,0,195,0,64,0,131,0,253,0,84,0,0,0,210,0,187,0,209,0,26,0,7,0,196,0,39,0,89,0,243,0,75,0,24,0,112,0,238,0,254,0,19,0,7,0,241,0,211,0,118,0,92,0,0,0,59,0,0,0,0,0,133,0,161,0,0,0,0,0,188,0,153,0,66,0,173,0,108,0,0,0,24,0,220,0,173,0,252,0,198,0,0,0,0,0,178,0,155,0,0,0,255,0,162,0,0,0,0,0,0,0,134,0,153,0,248,0,59,0,216,0,222,0,54,0,143,0,226,0,237,0,0,0,0,0,26,0,127,0,99,0,66,0,145,0,79,0,0,0,133,0,130,0,94,0,241,0,217,0,138,0,221,0,45,0,32,0,53,0,204,0,152,0,100,0,0,0,137,0,179,0,116,0,39,0,88,0,155,0,80,0,192,0,13,0,0,0,0,0,127,0,101,0,6,0,39,0,13,0,201,0,101,0,0,0,229,0,73,0,0,0,55,0,0,0,83,0,1,0,0,0,115,0,0,0,65,0,5,0,150,0,224,0,116,0,61,0,0,0,35,0,184,0,90,0,200,0,47,0,237,0,63,0,207,0,20,0,0,0,0,0,173,0,49,0,56,0,144,0,23,0,51,0,2,0,236,0,0,0,251,0,202,0,141,0,33,0,60,0,140,0,12,0,154,0,0,0,0,0,151,0,96,0,133,0,9,0,104,0,0,0,112,0,49,0,137,0,42,0,0,0,102,0,150,0,215,0,123,0,0,0,0,0,129,0,25,0,207,0,42,0,239,0,0,0,201,0,132,0,0,0,135,0,247,0,0,0,0,0,62,0,0,0,97,0,68,0,137,0,243,0,0,0,0,0,199,0,230,0,28,0,94,0,191,0,0,0,193,0,63,0,162,0,0,0,0,0,96,0,222,0,178,0,220,0,120,0,15,0,233,0,50,0,186,0,78,0,243,0,242,0,0,0,161,0,114,0,133,0,140,0,229,0,203,0,160,0,231,0,197,0,166,0,144,0,0,0,220,0,22,0,177,0,170,0,250,0,178,0,95,0,76,0,115,0,52,0,208,0,1,0,0,0,88,0,170,0,116,0,0,0,31,0,67,0,7,0,111,0,16,0,229,0,6,0,0,0,0,0,0,0,63,0,0,0,95,0,80,0,109,0,0,0,0,0,86,0,252,0,0,0,42,0);
signal scenario_full  : scenario_type := (0,0,186,31,22,31,22,30,163,31,57,31,14,31,14,30,141,31,238,31,93,31,55,31,178,31,178,30,178,29,86,31,236,31,161,31,48,31,12,31,97,31,210,31,210,30,40,31,218,31,77,31,41,31,83,31,100,31,100,30,27,31,3,31,196,31,207,31,134,31,158,31,45,31,153,31,30,31,201,31,243,31,137,31,173,31,112,31,112,30,208,31,198,31,93,31,63,31,12,31,142,31,142,30,44,31,135,31,80,31,231,31,231,30,110,31,75,31,12,31,29,31,29,30,82,31,13,31,13,30,13,29,180,31,226,31,245,31,179,31,51,31,43,31,24,31,223,31,168,31,1,31,249,31,126,31,188,31,188,30,222,31,3,31,219,31,130,31,36,31,64,31,4,31,45,31,250,31,48,31,127,31,84,31,84,30,204,31,43,31,138,31,109,31,181,31,58,31,131,31,190,31,104,31,229,31,62,31,197,31,20,31,20,30,24,31,80,31,119,31,119,30,119,29,220,31,161,31,105,31,29,31,77,31,77,30,32,31,32,30,228,31,207,31,225,31,225,30,230,31,161,31,161,30,172,31,154,31,153,31,145,31,145,30,68,31,158,31,219,31,219,30,59,31,154,31,179,31,141,31,62,31,62,30,62,29,62,28,62,27,62,26,250,31,7,31,3,31,216,31,216,30,164,31,42,31,191,31,92,31,92,30,170,31,135,31,133,31,13,31,73,31,57,31,57,30,124,31,52,31,52,30,52,29,59,31,59,30,3,31,123,31,99,31,99,30,99,29,99,28,68,31,69,31,233,31,137,31,59,31,143,31,103,31,223,31,107,31,143,31,143,30,143,29,134,31,31,31,61,31,20,31,68,31,222,31,140,31,115,31,191,31,157,31,162,31,162,30,241,31,16,31,16,30,247,31,117,31,73,31,23,31,163,31,27,31,185,31,185,30,4,31,253,31,250,31,250,30,73,31,124,31,250,31,97,31,141,31,176,31,175,31,241,31,86,31,86,30,86,29,86,28,67,31,3,31,42,31,217,31,252,31,180,31,180,30,223,31,245,31,35,31,231,31,231,30,222,31,132,31,214,31,255,31,201,31,70,31,225,31,153,31,45,31,100,31,208,31,208,30,208,29,172,31,64,31,149,31,49,31,205,31,26,31,201,31,201,30,143,31,86,31,95,31,95,30,228,31,79,31,79,30,242,31,103,31,89,31,89,30,214,31,214,30,214,29,93,31,1,31,50,31,8,31,52,31,23,31,107,31,121,31,176,31,29,31,29,30,156,31,156,30,141,31,177,31,203,31,208,31,113,31,214,31,254,31,24,31,24,30,28,31,167,31,217,31,191,31,191,30,255,31,255,30,9,31,9,30,251,31,244,31,78,31,187,31,51,31,192,31,61,31,110,31,171,31,82,31,131,31,98,31,63,31,105,31,57,31,72,31,234,31,227,31,112,31,73,31,220,31,1,31,242,31,11,31,181,31,220,31,178,31,149,31,128,31,163,31,182,31,43,31,186,31,10,31,124,31,61,31,201,31,85,31,15,31,48,31,192,31,250,31,192,31,242,31,242,30,55,31,226,31,226,30,144,31,80,31,175,31,51,31,48,31,176,31,205,31,28,31,195,31,176,31,37,31,222,31,174,31,235,31,118,31,139,31,155,31,155,30,142,31,212,31,121,31,28,31,153,31,165,31,161,31,200,31,20,31,185,31,244,31,244,31,97,31,143,31,164,31,115,31,17,31,110,31,236,31,236,31,197,31,5,31,138,31,111,31,111,30,147,31,165,31,181,31,235,31,87,31,87,30,15,31,130,31,130,30,130,29,130,28,182,31,19,31,154,31,227,31,19,31,71,31,42,31,42,30,32,31,238,31,238,30,255,31,213,31,175,31,6,31,6,30,161,31,93,31,82,31,162,31,162,30,216,31,127,31,32,31,226,31,72,31,243,31,13,31,65,31,89,31,221,31,233,31,55,31,55,30,105,31,20,31,39,31,210,31,122,31,35,31,3,31,164,31,164,30,171,31,126,31,26,31,32,31,32,30,209,31,209,30,209,29,167,31,57,31,119,31,144,31,185,31,236,31,112,31,14,31,90,31,90,30,50,31,35,31,12,31,47,31,47,30,139,31,192,31,65,31,20,31,66,31,66,30,107,31,107,30,107,29,114,31,85,31,174,31,47,31,47,30,22,31,250,31,29,31,39,31,103,31,53,31,68,31,142,31,220,31,140,31,137,31,18,31,205,31,247,31,41,31,162,31,157,31,157,30,61,31,243,31,243,30,177,31,45,31,217,31,56,31,206,31,206,30,234,31,177,31,157,31,13,31,13,30,58,31,58,30,58,29,32,31,30,31,39,31,156,31,4,31,69,31,231,31,242,31,62,31,48,31,100,31,100,30,241,31,241,30,93,31,229,31,85,31,81,31,187,31,153,31,240,31,114,31,242,31,242,30,249,31,107,31,6,31,178,31,178,30,178,29,102,31,102,30,221,31,221,30,211,31,70,31,65,31,232,31,232,30,96,31,41,31,195,31,64,31,131,31,253,31,84,31,84,30,210,31,187,31,209,31,26,31,7,31,196,31,39,31,89,31,243,31,75,31,24,31,112,31,238,31,254,31,19,31,7,31,241,31,211,31,118,31,92,31,92,30,59,31,59,30,59,29,133,31,161,31,161,30,161,29,188,31,153,31,66,31,173,31,108,31,108,30,24,31,220,31,173,31,252,31,198,31,198,30,198,29,178,31,155,31,155,30,255,31,162,31,162,30,162,29,162,28,134,31,153,31,248,31,59,31,216,31,222,31,54,31,143,31,226,31,237,31,237,30,237,29,26,31,127,31,99,31,66,31,145,31,79,31,79,30,133,31,130,31,94,31,241,31,217,31,138,31,221,31,45,31,32,31,53,31,204,31,152,31,100,31,100,30,137,31,179,31,116,31,39,31,88,31,155,31,80,31,192,31,13,31,13,30,13,29,127,31,101,31,6,31,39,31,13,31,201,31,101,31,101,30,229,31,73,31,73,30,55,31,55,30,83,31,1,31,1,30,115,31,115,30,65,31,5,31,150,31,224,31,116,31,61,31,61,30,35,31,184,31,90,31,200,31,47,31,237,31,63,31,207,31,20,31,20,30,20,29,173,31,49,31,56,31,144,31,23,31,51,31,2,31,236,31,236,30,251,31,202,31,141,31,33,31,60,31,140,31,12,31,154,31,154,30,154,29,151,31,96,31,133,31,9,31,104,31,104,30,112,31,49,31,137,31,42,31,42,30,102,31,150,31,215,31,123,31,123,30,123,29,129,31,25,31,207,31,42,31,239,31,239,30,201,31,132,31,132,30,135,31,247,31,247,30,247,29,62,31,62,30,97,31,68,31,137,31,243,31,243,30,243,29,199,31,230,31,28,31,94,31,191,31,191,30,193,31,63,31,162,31,162,30,162,29,96,31,222,31,178,31,220,31,120,31,15,31,233,31,50,31,186,31,78,31,243,31,242,31,242,30,161,31,114,31,133,31,140,31,229,31,203,31,160,31,231,31,197,31,166,31,144,31,144,30,220,31,22,31,177,31,170,31,250,31,178,31,95,31,76,31,115,31,52,31,208,31,1,31,1,30,88,31,170,31,116,31,116,30,31,31,67,31,7,31,111,31,16,31,229,31,6,31,6,30,6,29,6,28,63,31,63,30,95,31,80,31,109,31,109,30,109,29,86,31,252,31,252,30,42,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
