-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_463 is
end project_tb_463;

architecture project_tb_arch_463 of project_tb_463 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 996;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (98,0,0,0,0,0,136,0,0,0,97,0,192,0,140,0,153,0,210,0,36,0,153,0,222,0,50,0,130,0,251,0,225,0,253,0,162,0,0,0,213,0,239,0,247,0,253,0,176,0,144,0,52,0,148,0,195,0,161,0,248,0,90,0,120,0,36,0,219,0,220,0,227,0,118,0,0,0,178,0,176,0,30,0,238,0,160,0,30,0,93,0,81,0,167,0,169,0,0,0,251,0,133,0,63,0,67,0,155,0,219,0,250,0,248,0,0,0,0,0,142,0,204,0,103,0,221,0,34,0,11,0,60,0,101,0,55,0,226,0,156,0,7,0,137,0,118,0,179,0,0,0,201,0,184,0,213,0,98,0,127,0,0,0,4,0,61,0,133,0,0,0,93,0,216,0,190,0,219,0,154,0,48,0,0,0,160,0,244,0,212,0,213,0,217,0,113,0,229,0,105,0,0,0,0,0,37,0,158,0,243,0,144,0,199,0,240,0,18,0,212,0,237,0,15,0,209,0,41,0,128,0,222,0,82,0,107,0,232,0,178,0,188,0,83,0,177,0,0,0,184,0,0,0,86,0,212,0,53,0,0,0,243,0,255,0,0,0,201,0,0,0,0,0,0,0,95,0,123,0,226,0,234,0,50,0,0,0,21,0,92,0,199,0,21,0,20,0,133,0,0,0,28,0,173,0,97,0,0,0,140,0,206,0,158,0,169,0,180,0,137,0,74,0,219,0,187,0,0,0,83,0,250,0,86,0,2,0,124,0,0,0,18,0,207,0,135,0,0,0,141,0,79,0,174,0,0,0,167,0,19,0,47,0,148,0,0,0,236,0,0,0,10,0,74,0,46,0,147,0,103,0,186,0,63,0,3,0,173,0,249,0,0,0,50,0,27,0,189,0,112,0,169,0,0,0,0,0,125,0,216,0,121,0,239,0,0,0,21,0,0,0,17,0,223,0,197,0,0,0,238,0,192,0,109,0,227,0,91,0,212,0,135,0,58,0,0,0,125,0,158,0,204,0,182,0,221,0,57,0,136,0,23,0,97,0,0,0,242,0,0,0,61,0,102,0,84,0,0,0,38,0,210,0,170,0,21,0,0,0,0,0,0,0,240,0,22,0,0,0,94,0,84,0,96,0,0,0,0,0,82,0,0,0,10,0,0,0,41,0,40,0,58,0,138,0,107,0,0,0,253,0,50,0,170,0,96,0,0,0,112,0,26,0,0,0,0,0,0,0,50,0,243,0,58,0,0,0,250,0,91,0,53,0,151,0,119,0,185,0,0,0,38,0,49,0,0,0,34,0,49,0,0,0,0,0,228,0,28,0,68,0,187,0,155,0,176,0,0,0,0,0,68,0,37,0,231,0,206,0,212,0,58,0,240,0,180,0,28,0,0,0,169,0,0,0,31,0,222,0,221,0,181,0,221,0,0,0,195,0,158,0,0,0,15,0,89,0,52,0,0,0,205,0,0,0,213,0,170,0,0,0,92,0,79,0,0,0,138,0,0,0,35,0,244,0,165,0,199,0,198,0,232,0,95,0,74,0,45,0,67,0,125,0,0,0,235,0,0,0,239,0,98,0,238,0,106,0,160,0,73,0,98,0,30,0,116,0,233,0,246,0,99,0,175,0,124,0,115,0,230,0,54,0,213,0,181,0,14,0,17,0,225,0,45,0,239,0,255,0,42,0,0,0,135,0,0,0,161,0,99,0,69,0,0,0,55,0,145,0,160,0,222,0,3,0,63,0,197,0,247,0,183,0,53,0,14,0,124,0,0,0,66,0,75,0,0,0,9,0,106,0,116,0,0,0,100,0,190,0,0,0,185,0,0,0,0,0,78,0,71,0,140,0,0,0,162,0,229,0,0,0,104,0,0,0,129,0,95,0,192,0,139,0,164,0,241,0,230,0,252,0,29,0,73,0,144,0,58,0,0,0,206,0,0,0,59,0,0,0,36,0,93,0,128,0,54,0,38,0,0,0,165,0,232,0,40,0,209,0,154,0,87,0,0,0,137,0,0,0,87,0,229,0,85,0,177,0,105,0,14,0,215,0,191,0,219,0,0,0,37,0,0,0,0,0,137,0,18,0,0,0,229,0,58,0,0,0,253,0,0,0,117,0,126,0,26,0,185,0,161,0,111,0,87,0,168,0,0,0,142,0,210,0,0,0,252,0,106,0,0,0,0,0,30,0,43,0,4,0,0,0,88,0,0,0,145,0,44,0,152,0,81,0,0,0,40,0,34,0,45,0,0,0,98,0,0,0,157,0,59,0,116,0,0,0,84,0,155,0,0,0,171,0,226,0,0,0,225,0,238,0,139,0,33,0,78,0,176,0,39,0,140,0,162,0,101,0,253,0,74,0,16,0,143,0,230,0,55,0,130,0,0,0,0,0,168,0,130,0,203,0,92,0,0,0,0,0,9,0,247,0,0,0,0,0,0,0,237,0,50,0,53,0,168,0,96,0,10,0,0,0,85,0,51,0,0,0,0,0,206,0,247,0,251,0,253,0,215,0,151,0,227,0,51,0,0,0,0,0,237,0,238,0,88,0,79,0,121,0,61,0,216,0,171,0,0,0,0,0,133,0,71,0,242,0,0,0,19,0,113,0,20,0,125,0,251,0,233,0,0,0,217,0,245,0,181,0,173,0,215,0,0,0,0,0,0,0,4,0,149,0,0,0,0,0,35,0,210,0,0,0,157,0,159,0,251,0,42,0,61,0,226,0,0,0,69,0,19,0,186,0,204,0,0,0,202,0,248,0,80,0,188,0,210,0,54,0,0,0,177,0,231,0,20,0,190,0,166,0,193,0,69,0,230,0,78,0,115,0,137,0,219,0,169,0,0,0,225,0,0,0,113,0,65,0,196,0,0,0,0,0,208,0,0,0,181,0,198,0,2,0,190,0,0,0,0,0,194,0,1,0,184,0,0,0,208,0,254,0,5,0,135,0,58,0,98,0,238,0,0,0,24,0,19,0,90,0,135,0,198,0,135,0,75,0,182,0,39,0,37,0,0,0,13,0,203,0,48,0,228,0,34,0,183,0,250,0,0,0,173,0,58,0,155,0,54,0,55,0,46,0,107,0,15,0,113,0,71,0,21,0,0,0,69,0,0,0,5,0,79,0,3,0,28,0,213,0,0,0,0,0,207,0,0,0,160,0,0,0,141,0,27,0,18,0,77,0,69,0,213,0,89,0,212,0,0,0,8,0,120,0,0,0,129,0,49,0,0,0,0,0,0,0,0,0,158,0,144,0,215,0,0,0,91,0,229,0,182,0,26,0,0,0,67,0,6,0,0,0,202,0,166,0,169,0,0,0,0,0,229,0,1,0,0,0,0,0,0,0,1,0,218,0,161,0,29,0,21,0,0,0,193,0,10,0,187,0,240,0,251,0,59,0,0,0,204,0,46,0,126,0,0,0,148,0,118,0,190,0,0,0,209,0,0,0,0,0,255,0,188,0,0,0,91,0,0,0,81,0,57,0,18,0,250,0,206,0,189,0,115,0,119,0,59,0,229,0,221,0,161,0,0,0,247,0,106,0,70,0,145,0,247,0,175,0,60,0,111,0,218,0,101,0,99,0,79,0,204,0,0,0,26,0,14,0,195,0,3,0,99,0,244,0,0,0,22,0,180,0,184,0,200,0,239,0,139,0,13,0,167,0,0,0,20,0,0,0,23,0,245,0,176,0,141,0,188,0,112,0,69,0,235,0,175,0,254,0,171,0,209,0,108,0,112,0,0,0,64,0,28,0,179,0,252,0,87,0,3,0,173,0,67,0,13,0,224,0,0,0,122,0,0,0,228,0,189,0,106,0,100,0,16,0,0,0,54,0,254,0,249,0,75,0,189,0,0,0,171,0,0,0,108,0,236,0,0,0,77,0,53,0,107,0,59,0,226,0,182,0,0,0,213,0,0,0,179,0,218,0,71,0,126,0,250,0,85,0,30,0,188,0,165,0,89,0,143,0,136,0,203,0,0,0,7,0,220,0,77,0,64,0,236,0,249,0,0,0,131,0,172,0,33,0,0,0,161,0,37,0,246,0,116,0,11,0,230,0,181,0,194,0,0,0,211,0,131,0,237,0,0,0,61,0,0,0,0,0,242,0,165,0,28,0,121,0,77,0,26,0,117,0,5,0,9,0,184,0,0,0,230,0,0,0,123,0,189,0,73,0,148,0,181,0,86,0,228,0,194,0,122,0,67,0,238,0,0,0,227,0,0,0,246,0,0,0,64,0,25,0,247,0,185,0,154,0,0,0,142,0,6,0,151,0,167,0,0,0,206,0,0,0,76,0,85,0,251,0,22,0,63,0,176,0,32,0,17,0,32,0,0,0,200,0,167,0,42,0,68,0,0,0,5,0,101,0,204,0,0,0,114,0,10,0,234,0,0,0,84,0,0,0,0,0,193,0,242,0,191,0,172,0,211,0,0,0,70,0,10,0,0,0,229,0,0,0,60,0,48,0,0,0);
signal scenario_full  : scenario_type := (98,31,98,30,98,29,136,31,136,30,97,31,192,31,140,31,153,31,210,31,36,31,153,31,222,31,50,31,130,31,251,31,225,31,253,31,162,31,162,30,213,31,239,31,247,31,253,31,176,31,144,31,52,31,148,31,195,31,161,31,248,31,90,31,120,31,36,31,219,31,220,31,227,31,118,31,118,30,178,31,176,31,30,31,238,31,160,31,30,31,93,31,81,31,167,31,169,31,169,30,251,31,133,31,63,31,67,31,155,31,219,31,250,31,248,31,248,30,248,29,142,31,204,31,103,31,221,31,34,31,11,31,60,31,101,31,55,31,226,31,156,31,7,31,137,31,118,31,179,31,179,30,201,31,184,31,213,31,98,31,127,31,127,30,4,31,61,31,133,31,133,30,93,31,216,31,190,31,219,31,154,31,48,31,48,30,160,31,244,31,212,31,213,31,217,31,113,31,229,31,105,31,105,30,105,29,37,31,158,31,243,31,144,31,199,31,240,31,18,31,212,31,237,31,15,31,209,31,41,31,128,31,222,31,82,31,107,31,232,31,178,31,188,31,83,31,177,31,177,30,184,31,184,30,86,31,212,31,53,31,53,30,243,31,255,31,255,30,201,31,201,30,201,29,201,28,95,31,123,31,226,31,234,31,50,31,50,30,21,31,92,31,199,31,21,31,20,31,133,31,133,30,28,31,173,31,97,31,97,30,140,31,206,31,158,31,169,31,180,31,137,31,74,31,219,31,187,31,187,30,83,31,250,31,86,31,2,31,124,31,124,30,18,31,207,31,135,31,135,30,141,31,79,31,174,31,174,30,167,31,19,31,47,31,148,31,148,30,236,31,236,30,10,31,74,31,46,31,147,31,103,31,186,31,63,31,3,31,173,31,249,31,249,30,50,31,27,31,189,31,112,31,169,31,169,30,169,29,125,31,216,31,121,31,239,31,239,30,21,31,21,30,17,31,223,31,197,31,197,30,238,31,192,31,109,31,227,31,91,31,212,31,135,31,58,31,58,30,125,31,158,31,204,31,182,31,221,31,57,31,136,31,23,31,97,31,97,30,242,31,242,30,61,31,102,31,84,31,84,30,38,31,210,31,170,31,21,31,21,30,21,29,21,28,240,31,22,31,22,30,94,31,84,31,96,31,96,30,96,29,82,31,82,30,10,31,10,30,41,31,40,31,58,31,138,31,107,31,107,30,253,31,50,31,170,31,96,31,96,30,112,31,26,31,26,30,26,29,26,28,50,31,243,31,58,31,58,30,250,31,91,31,53,31,151,31,119,31,185,31,185,30,38,31,49,31,49,30,34,31,49,31,49,30,49,29,228,31,28,31,68,31,187,31,155,31,176,31,176,30,176,29,68,31,37,31,231,31,206,31,212,31,58,31,240,31,180,31,28,31,28,30,169,31,169,30,31,31,222,31,221,31,181,31,221,31,221,30,195,31,158,31,158,30,15,31,89,31,52,31,52,30,205,31,205,30,213,31,170,31,170,30,92,31,79,31,79,30,138,31,138,30,35,31,244,31,165,31,199,31,198,31,232,31,95,31,74,31,45,31,67,31,125,31,125,30,235,31,235,30,239,31,98,31,238,31,106,31,160,31,73,31,98,31,30,31,116,31,233,31,246,31,99,31,175,31,124,31,115,31,230,31,54,31,213,31,181,31,14,31,17,31,225,31,45,31,239,31,255,31,42,31,42,30,135,31,135,30,161,31,99,31,69,31,69,30,55,31,145,31,160,31,222,31,3,31,63,31,197,31,247,31,183,31,53,31,14,31,124,31,124,30,66,31,75,31,75,30,9,31,106,31,116,31,116,30,100,31,190,31,190,30,185,31,185,30,185,29,78,31,71,31,140,31,140,30,162,31,229,31,229,30,104,31,104,30,129,31,95,31,192,31,139,31,164,31,241,31,230,31,252,31,29,31,73,31,144,31,58,31,58,30,206,31,206,30,59,31,59,30,36,31,93,31,128,31,54,31,38,31,38,30,165,31,232,31,40,31,209,31,154,31,87,31,87,30,137,31,137,30,87,31,229,31,85,31,177,31,105,31,14,31,215,31,191,31,219,31,219,30,37,31,37,30,37,29,137,31,18,31,18,30,229,31,58,31,58,30,253,31,253,30,117,31,126,31,26,31,185,31,161,31,111,31,87,31,168,31,168,30,142,31,210,31,210,30,252,31,106,31,106,30,106,29,30,31,43,31,4,31,4,30,88,31,88,30,145,31,44,31,152,31,81,31,81,30,40,31,34,31,45,31,45,30,98,31,98,30,157,31,59,31,116,31,116,30,84,31,155,31,155,30,171,31,226,31,226,30,225,31,238,31,139,31,33,31,78,31,176,31,39,31,140,31,162,31,101,31,253,31,74,31,16,31,143,31,230,31,55,31,130,31,130,30,130,29,168,31,130,31,203,31,92,31,92,30,92,29,9,31,247,31,247,30,247,29,247,28,237,31,50,31,53,31,168,31,96,31,10,31,10,30,85,31,51,31,51,30,51,29,206,31,247,31,251,31,253,31,215,31,151,31,227,31,51,31,51,30,51,29,237,31,238,31,88,31,79,31,121,31,61,31,216,31,171,31,171,30,171,29,133,31,71,31,242,31,242,30,19,31,113,31,20,31,125,31,251,31,233,31,233,30,217,31,245,31,181,31,173,31,215,31,215,30,215,29,215,28,4,31,149,31,149,30,149,29,35,31,210,31,210,30,157,31,159,31,251,31,42,31,61,31,226,31,226,30,69,31,19,31,186,31,204,31,204,30,202,31,248,31,80,31,188,31,210,31,54,31,54,30,177,31,231,31,20,31,190,31,166,31,193,31,69,31,230,31,78,31,115,31,137,31,219,31,169,31,169,30,225,31,225,30,113,31,65,31,196,31,196,30,196,29,208,31,208,30,181,31,198,31,2,31,190,31,190,30,190,29,194,31,1,31,184,31,184,30,208,31,254,31,5,31,135,31,58,31,98,31,238,31,238,30,24,31,19,31,90,31,135,31,198,31,135,31,75,31,182,31,39,31,37,31,37,30,13,31,203,31,48,31,228,31,34,31,183,31,250,31,250,30,173,31,58,31,155,31,54,31,55,31,46,31,107,31,15,31,113,31,71,31,21,31,21,30,69,31,69,30,5,31,79,31,3,31,28,31,213,31,213,30,213,29,207,31,207,30,160,31,160,30,141,31,27,31,18,31,77,31,69,31,213,31,89,31,212,31,212,30,8,31,120,31,120,30,129,31,49,31,49,30,49,29,49,28,49,27,158,31,144,31,215,31,215,30,91,31,229,31,182,31,26,31,26,30,67,31,6,31,6,30,202,31,166,31,169,31,169,30,169,29,229,31,1,31,1,30,1,29,1,28,1,31,218,31,161,31,29,31,21,31,21,30,193,31,10,31,187,31,240,31,251,31,59,31,59,30,204,31,46,31,126,31,126,30,148,31,118,31,190,31,190,30,209,31,209,30,209,29,255,31,188,31,188,30,91,31,91,30,81,31,57,31,18,31,250,31,206,31,189,31,115,31,119,31,59,31,229,31,221,31,161,31,161,30,247,31,106,31,70,31,145,31,247,31,175,31,60,31,111,31,218,31,101,31,99,31,79,31,204,31,204,30,26,31,14,31,195,31,3,31,99,31,244,31,244,30,22,31,180,31,184,31,200,31,239,31,139,31,13,31,167,31,167,30,20,31,20,30,23,31,245,31,176,31,141,31,188,31,112,31,69,31,235,31,175,31,254,31,171,31,209,31,108,31,112,31,112,30,64,31,28,31,179,31,252,31,87,31,3,31,173,31,67,31,13,31,224,31,224,30,122,31,122,30,228,31,189,31,106,31,100,31,16,31,16,30,54,31,254,31,249,31,75,31,189,31,189,30,171,31,171,30,108,31,236,31,236,30,77,31,53,31,107,31,59,31,226,31,182,31,182,30,213,31,213,30,179,31,218,31,71,31,126,31,250,31,85,31,30,31,188,31,165,31,89,31,143,31,136,31,203,31,203,30,7,31,220,31,77,31,64,31,236,31,249,31,249,30,131,31,172,31,33,31,33,30,161,31,37,31,246,31,116,31,11,31,230,31,181,31,194,31,194,30,211,31,131,31,237,31,237,30,61,31,61,30,61,29,242,31,165,31,28,31,121,31,77,31,26,31,117,31,5,31,9,31,184,31,184,30,230,31,230,30,123,31,189,31,73,31,148,31,181,31,86,31,228,31,194,31,122,31,67,31,238,31,238,30,227,31,227,30,246,31,246,30,64,31,25,31,247,31,185,31,154,31,154,30,142,31,6,31,151,31,167,31,167,30,206,31,206,30,76,31,85,31,251,31,22,31,63,31,176,31,32,31,17,31,32,31,32,30,200,31,167,31,42,31,68,31,68,30,5,31,101,31,204,31,204,30,114,31,10,31,234,31,234,30,84,31,84,30,84,29,193,31,242,31,191,31,172,31,211,31,211,30,70,31,10,31,10,30,229,31,229,30,60,31,48,31,48,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
