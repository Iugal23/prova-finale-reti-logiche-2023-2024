-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_633 is
end project_tb_633;

architecture project_tb_arch_633 of project_tb_633 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 179;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (85,0,0,0,254,0,3,0,24,0,134,0,114,0,84,0,96,0,129,0,82,0,101,0,0,0,218,0,0,0,123,0,180,0,216,0,0,0,64,0,224,0,0,0,0,0,234,0,0,0,0,0,0,0,0,0,192,0,21,0,232,0,0,0,0,0,30,0,202,0,106,0,67,0,112,0,156,0,178,0,7,0,0,0,200,0,123,0,247,0,162,0,205,0,166,0,0,0,219,0,189,0,237,0,135,0,134,0,0,0,246,0,0,0,73,0,5,0,62,0,192,0,60,0,243,0,101,0,83,0,0,0,153,0,116,0,0,0,138,0,0,0,206,0,61,0,0,0,79,0,0,0,112,0,91,0,91,0,182,0,116,0,0,0,161,0,237,0,143,0,208,0,29,0,96,0,212,0,35,0,82,0,0,0,115,0,142,0,0,0,51,0,24,0,235,0,39,0,141,0,186,0,116,0,58,0,145,0,79,0,215,0,232,0,84,0,0,0,0,0,63,0,5,0,0,0,100,0,0,0,228,0,0,0,0,0,162,0,0,0,0,0,235,0,110,0,56,0,146,0,28,0,0,0,226,0,233,0,47,0,155,0,233,0,0,0,71,0,208,0,166,0,137,0,59,0,34,0,55,0,143,0,232,0,137,0,0,0,129,0,182,0,209,0,242,0,77,0,0,0,14,0,0,0,130,0,32,0,228,0,75,0,236,0,130,0,245,0,240,0,250,0,219,0,35,0,195,0,242,0,238,0,70,0,121,0,189,0,37,0,191,0,106,0,0,0,86,0,213,0,88,0,240,0,0,0,148,0);
signal scenario_full  : scenario_type := (85,31,85,30,254,31,3,31,24,31,134,31,114,31,84,31,96,31,129,31,82,31,101,31,101,30,218,31,218,30,123,31,180,31,216,31,216,30,64,31,224,31,224,30,224,29,234,31,234,30,234,29,234,28,234,27,192,31,21,31,232,31,232,30,232,29,30,31,202,31,106,31,67,31,112,31,156,31,178,31,7,31,7,30,200,31,123,31,247,31,162,31,205,31,166,31,166,30,219,31,189,31,237,31,135,31,134,31,134,30,246,31,246,30,73,31,5,31,62,31,192,31,60,31,243,31,101,31,83,31,83,30,153,31,116,31,116,30,138,31,138,30,206,31,61,31,61,30,79,31,79,30,112,31,91,31,91,31,182,31,116,31,116,30,161,31,237,31,143,31,208,31,29,31,96,31,212,31,35,31,82,31,82,30,115,31,142,31,142,30,51,31,24,31,235,31,39,31,141,31,186,31,116,31,58,31,145,31,79,31,215,31,232,31,84,31,84,30,84,29,63,31,5,31,5,30,100,31,100,30,228,31,228,30,228,29,162,31,162,30,162,29,235,31,110,31,56,31,146,31,28,31,28,30,226,31,233,31,47,31,155,31,233,31,233,30,71,31,208,31,166,31,137,31,59,31,34,31,55,31,143,31,232,31,137,31,137,30,129,31,182,31,209,31,242,31,77,31,77,30,14,31,14,30,130,31,32,31,228,31,75,31,236,31,130,31,245,31,240,31,250,31,219,31,35,31,195,31,242,31,238,31,70,31,121,31,189,31,37,31,191,31,106,31,106,30,86,31,213,31,88,31,240,31,240,30,148,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
