-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 258;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (173,0,151,0,101,0,91,0,2,0,0,0,41,0,124,0,129,0,0,0,0,0,0,0,42,0,0,0,201,0,113,0,111,0,124,0,195,0,82,0,247,0,142,0,200,0,72,0,153,0,238,0,0,0,138,0,73,0,167,0,197,0,29,0,199,0,0,0,245,0,149,0,68,0,0,0,41,0,31,0,103,0,48,0,70,0,26,0,150,0,186,0,250,0,26,0,0,0,0,0,2,0,145,0,0,0,184,0,0,0,178,0,78,0,217,0,76,0,84,0,67,0,209,0,218,0,182,0,0,0,57,0,1,0,0,0,207,0,70,0,39,0,188,0,241,0,0,0,204,0,157,0,0,0,94,0,140,0,209,0,163,0,128,0,215,0,45,0,175,0,9,0,0,0,46,0,50,0,8,0,233,0,0,0,206,0,0,0,200,0,0,0,0,0,34,0,64,0,165,0,173,0,37,0,0,0,11,0,113,0,231,0,126,0,215,0,138,0,55,0,0,0,57,0,0,0,118,0,38,0,0,0,0,0,0,0,176,0,144,0,59,0,248,0,24,0,11,0,129,0,61,0,0,0,205,0,17,0,102,0,158,0,0,0,106,0,173,0,56,0,0,0,5,0,124,0,236,0,152,0,0,0,202,0,106,0,0,0,0,0,0,0,80,0,47,0,34,0,64,0,78,0,238,0,58,0,146,0,19,0,178,0,5,0,0,0,0,0,0,0,231,0,101,0,74,0,21,0,26,0,112,0,34,0,112,0,52,0,44,0,246,0,155,0,120,0,86,0,237,0,14,0,76,0,122,0,0,0,37,0,143,0,155,0,0,0,105,0,120,0,177,0,91,0,149,0,57,0,168,0,0,0,0,0,51,0,83,0,123,0,0,0,0,0,0,0,40,0,21,0,138,0,154,0,151,0,2,0,113,0,18,0,199,0,124,0,0,0,110,0,0,0,0,0,36,0,111,0,198,0,0,0,239,0,0,0,137,0,169,0,46,0,154,0,170,0,0,0,89,0,1,0,0,0,157,0,98,0,127,0,222,0,94,0,200,0,0,0,236,0,57,0,117,0,229,0,170,0,0,0,115,0,7,0,0,0,127,0,190,0,128,0,167,0,154,0,36,0,110,0,228,0,73,0,28,0,128,0,155,0,16,0,0,0,179,0);
signal scenario_full  : scenario_type := (173,31,151,31,101,31,91,31,2,31,2,30,41,31,124,31,129,31,129,30,129,29,129,28,42,31,42,30,201,31,113,31,111,31,124,31,195,31,82,31,247,31,142,31,200,31,72,31,153,31,238,31,238,30,138,31,73,31,167,31,197,31,29,31,199,31,199,30,245,31,149,31,68,31,68,30,41,31,31,31,103,31,48,31,70,31,26,31,150,31,186,31,250,31,26,31,26,30,26,29,2,31,145,31,145,30,184,31,184,30,178,31,78,31,217,31,76,31,84,31,67,31,209,31,218,31,182,31,182,30,57,31,1,31,1,30,207,31,70,31,39,31,188,31,241,31,241,30,204,31,157,31,157,30,94,31,140,31,209,31,163,31,128,31,215,31,45,31,175,31,9,31,9,30,46,31,50,31,8,31,233,31,233,30,206,31,206,30,200,31,200,30,200,29,34,31,64,31,165,31,173,31,37,31,37,30,11,31,113,31,231,31,126,31,215,31,138,31,55,31,55,30,57,31,57,30,118,31,38,31,38,30,38,29,38,28,176,31,144,31,59,31,248,31,24,31,11,31,129,31,61,31,61,30,205,31,17,31,102,31,158,31,158,30,106,31,173,31,56,31,56,30,5,31,124,31,236,31,152,31,152,30,202,31,106,31,106,30,106,29,106,28,80,31,47,31,34,31,64,31,78,31,238,31,58,31,146,31,19,31,178,31,5,31,5,30,5,29,5,28,231,31,101,31,74,31,21,31,26,31,112,31,34,31,112,31,52,31,44,31,246,31,155,31,120,31,86,31,237,31,14,31,76,31,122,31,122,30,37,31,143,31,155,31,155,30,105,31,120,31,177,31,91,31,149,31,57,31,168,31,168,30,168,29,51,31,83,31,123,31,123,30,123,29,123,28,40,31,21,31,138,31,154,31,151,31,2,31,113,31,18,31,199,31,124,31,124,30,110,31,110,30,110,29,36,31,111,31,198,31,198,30,239,31,239,30,137,31,169,31,46,31,154,31,170,31,170,30,89,31,1,31,1,30,157,31,98,31,127,31,222,31,94,31,200,31,200,30,236,31,57,31,117,31,229,31,170,31,170,30,115,31,7,31,7,30,127,31,190,31,128,31,167,31,154,31,36,31,110,31,228,31,73,31,28,31,128,31,155,31,16,31,16,30,179,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
