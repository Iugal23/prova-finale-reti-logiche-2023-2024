-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_274 is
end project_tb_274;

architecture project_tb_arch_274 of project_tb_274 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 338;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (63,0,201,0,240,0,203,0,175,0,0,0,181,0,193,0,223,0,12,0,212,0,24,0,250,0,106,0,162,0,0,0,23,0,78,0,32,0,212,0,60,0,19,0,0,0,239,0,153,0,9,0,73,0,42,0,140,0,0,0,109,0,154,0,101,0,134,0,136,0,12,0,250,0,91,0,0,0,105,0,0,0,202,0,238,0,138,0,0,0,8,0,90,0,208,0,0,0,157,0,0,0,0,0,0,0,0,0,164,0,90,0,129,0,0,0,32,0,236,0,80,0,91,0,0,0,0,0,230,0,199,0,110,0,38,0,106,0,0,0,0,0,137,0,216,0,49,0,136,0,253,0,240,0,0,0,84,0,117,0,0,0,53,0,75,0,127,0,67,0,105,0,110,0,0,0,70,0,56,0,112,0,83,0,79,0,192,0,39,0,243,0,0,0,0,0,101,0,205,0,214,0,43,0,190,0,139,0,237,0,0,0,23,0,176,0,0,0,0,0,114,0,114,0,213,0,120,0,0,0,72,0,0,0,0,0,75,0,108,0,53,0,184,0,5,0,83,0,0,0,168,0,79,0,0,0,167,0,128,0,217,0,0,0,135,0,0,0,142,0,110,0,214,0,0,0,178,0,30,0,92,0,163,0,0,0,107,0,66,0,49,0,0,0,64,0,20,0,6,0,238,0,230,0,82,0,0,0,157,0,135,0,125,0,134,0,188,0,42,0,209,0,60,0,20,0,223,0,139,0,0,0,0,0,1,0,0,0,72,0,63,0,140,0,230,0,0,0,199,0,86,0,204,0,118,0,175,0,84,0,93,0,95,0,167,0,0,0,152,0,0,0,227,0,157,0,153,0,248,0,64,0,236,0,0,0,78,0,31,0,18,0,0,0,58,0,45,0,0,0,0,0,0,0,241,0,60,0,59,0,175,0,105,0,198,0,30,0,146,0,32,0,160,0,175,0,222,0,187,0,199,0,215,0,154,0,206,0,0,0,5,0,217,0,217,0,27,0,58,0,32,0,189,0,9,0,254,0,203,0,149,0,120,0,63,0,72,0,0,0,65,0,4,0,150,0,167,0,174,0,0,0,131,0,207,0,0,0,0,0,60,0,0,0,185,0,104,0,0,0,104,0,68,0,78,0,0,0,22,0,40,0,172,0,152,0,67,0,140,0,187,0,54,0,233,0,235,0,126,0,26,0,32,0,156,0,125,0,34,0,135,0,0,0,244,0,0,0,187,0,100,0,228,0,188,0,49,0,83,0,131,0,69,0,0,0,90,0,79,0,174,0,0,0,0,0,24,0,250,0,75,0,250,0,230,0,0,0,81,0,182,0,30,0,0,0,180,0,3,0,202,0,0,0,0,0,189,0,2,0,0,0,9,0,191,0,18,0,133,0,0,0,36,0,247,0,125,0,0,0,129,0,219,0,0,0,112,0,98,0,98,0,149,0,0,0,101,0,87,0,0,0,0,0,85,0,201,0,118,0,183,0,0,0,0,0,0,0,0,0,159,0,156,0,0,0);
signal scenario_full  : scenario_type := (63,31,201,31,240,31,203,31,175,31,175,30,181,31,193,31,223,31,12,31,212,31,24,31,250,31,106,31,162,31,162,30,23,31,78,31,32,31,212,31,60,31,19,31,19,30,239,31,153,31,9,31,73,31,42,31,140,31,140,30,109,31,154,31,101,31,134,31,136,31,12,31,250,31,91,31,91,30,105,31,105,30,202,31,238,31,138,31,138,30,8,31,90,31,208,31,208,30,157,31,157,30,157,29,157,28,157,27,164,31,90,31,129,31,129,30,32,31,236,31,80,31,91,31,91,30,91,29,230,31,199,31,110,31,38,31,106,31,106,30,106,29,137,31,216,31,49,31,136,31,253,31,240,31,240,30,84,31,117,31,117,30,53,31,75,31,127,31,67,31,105,31,110,31,110,30,70,31,56,31,112,31,83,31,79,31,192,31,39,31,243,31,243,30,243,29,101,31,205,31,214,31,43,31,190,31,139,31,237,31,237,30,23,31,176,31,176,30,176,29,114,31,114,31,213,31,120,31,120,30,72,31,72,30,72,29,75,31,108,31,53,31,184,31,5,31,83,31,83,30,168,31,79,31,79,30,167,31,128,31,217,31,217,30,135,31,135,30,142,31,110,31,214,31,214,30,178,31,30,31,92,31,163,31,163,30,107,31,66,31,49,31,49,30,64,31,20,31,6,31,238,31,230,31,82,31,82,30,157,31,135,31,125,31,134,31,188,31,42,31,209,31,60,31,20,31,223,31,139,31,139,30,139,29,1,31,1,30,72,31,63,31,140,31,230,31,230,30,199,31,86,31,204,31,118,31,175,31,84,31,93,31,95,31,167,31,167,30,152,31,152,30,227,31,157,31,153,31,248,31,64,31,236,31,236,30,78,31,31,31,18,31,18,30,58,31,45,31,45,30,45,29,45,28,241,31,60,31,59,31,175,31,105,31,198,31,30,31,146,31,32,31,160,31,175,31,222,31,187,31,199,31,215,31,154,31,206,31,206,30,5,31,217,31,217,31,27,31,58,31,32,31,189,31,9,31,254,31,203,31,149,31,120,31,63,31,72,31,72,30,65,31,4,31,150,31,167,31,174,31,174,30,131,31,207,31,207,30,207,29,60,31,60,30,185,31,104,31,104,30,104,31,68,31,78,31,78,30,22,31,40,31,172,31,152,31,67,31,140,31,187,31,54,31,233,31,235,31,126,31,26,31,32,31,156,31,125,31,34,31,135,31,135,30,244,31,244,30,187,31,100,31,228,31,188,31,49,31,83,31,131,31,69,31,69,30,90,31,79,31,174,31,174,30,174,29,24,31,250,31,75,31,250,31,230,31,230,30,81,31,182,31,30,31,30,30,180,31,3,31,202,31,202,30,202,29,189,31,2,31,2,30,9,31,191,31,18,31,133,31,133,30,36,31,247,31,125,31,125,30,129,31,219,31,219,30,112,31,98,31,98,31,149,31,149,30,101,31,87,31,87,30,87,29,85,31,201,31,118,31,183,31,183,30,183,29,183,28,183,27,159,31,156,31,156,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
