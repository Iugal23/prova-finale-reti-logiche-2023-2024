-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_26 is
end project_tb_26;

architecture project_tb_arch_26 of project_tb_26 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 907;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,250,0,139,0,187,0,124,0,159,0,96,0,27,0,93,0,111,0,214,0,135,0,13,0,203,0,248,0,199,0,48,0,234,0,36,0,190,0,176,0,40,0,242,0,0,0,28,0,34,0,0,0,107,0,73,0,239,0,0,0,0,0,140,0,206,0,122,0,56,0,0,0,250,0,205,0,0,0,189,0,185,0,92,0,85,0,190,0,56,0,42,0,54,0,63,0,140,0,138,0,105,0,35,0,178,0,0,0,54,0,215,0,12,0,245,0,26,0,0,0,0,0,185,0,0,0,49,0,22,0,56,0,0,0,132,0,159,0,186,0,233,0,238,0,232,0,107,0,117,0,152,0,156,0,143,0,221,0,3,0,247,0,114,0,153,0,0,0,9,0,102,0,111,0,190,0,136,0,234,0,65,0,98,0,216,0,0,0,114,0,176,0,51,0,0,0,211,0,193,0,0,0,238,0,4,0,21,0,0,0,166,0,106,0,175,0,128,0,42,0,80,0,22,0,0,0,81,0,226,0,150,0,110,0,0,0,47,0,177,0,0,0,194,0,140,0,182,0,169,0,136,0,78,0,0,0,28,0,4,0,159,0,165,0,115,0,110,0,0,0,190,0,121,0,0,0,152,0,61,0,0,0,214,0,57,0,15,0,0,0,1,0,145,0,83,0,0,0,245,0,0,0,0,0,52,0,154,0,0,0,230,0,185,0,132,0,0,0,0,0,225,0,162,0,124,0,110,0,10,0,27,0,0,0,60,0,11,0,227,0,90,0,147,0,222,0,137,0,107,0,240,0,80,0,193,0,56,0,0,0,0,0,0,0,165,0,0,0,41,0,115,0,24,0,156,0,155,0,197,0,146,0,209,0,42,0,234,0,87,0,74,0,241,0,0,0,180,0,0,0,28,0,136,0,0,0,46,0,248,0,58,0,130,0,226,0,22,0,20,0,0,0,243,0,0,0,43,0,170,0,142,0,198,0,74,0,56,0,67,0,132,0,151,0,229,0,30,0,206,0,204,0,167,0,0,0,13,0,20,0,199,0,73,0,101,0,103,0,7,0,102,0,178,0,255,0,132,0,136,0,235,0,217,0,128,0,71,0,65,0,39,0,168,0,0,0,90,0,13,0,79,0,0,0,187,0,0,0,20,0,67,0,52,0,129,0,191,0,150,0,23,0,11,0,92,0,34,0,0,0,195,0,246,0,121,0,93,0,197,0,35,0,239,0,51,0,0,0,0,0,14,0,152,0,0,0,0,0,88,0,185,0,43,0,0,0,114,0,15,0,162,0,97,0,126,0,227,0,121,0,0,0,33,0,255,0,220,0,212,0,124,0,79,0,38,0,238,0,131,0,182,0,0,0,85,0,32,0,191,0,195,0,181,0,246,0,155,0,0,0,107,0,82,0,29,0,173,0,0,0,190,0,177,0,14,0,26,0,0,0,0,0,64,0,0,0,0,0,116,0,118,0,2,0,0,0,229,0,100,0,121,0,89,0,104,0,188,0,151,0,217,0,40,0,0,0,174,0,76,0,7,0,189,0,25,0,0,0,0,0,120,0,118,0,210,0,0,0,2,0,0,0,250,0,193,0,0,0,0,0,213,0,100,0,226,0,130,0,7,0,4,0,66,0,108,0,22,0,5,0,133,0,0,0,221,0,4,0,150,0,231,0,0,0,183,0,88,0,238,0,183,0,167,0,141,0,0,0,106,0,211,0,0,0,5,0,190,0,111,0,0,0,0,0,0,0,80,0,239,0,85,0,217,0,0,0,231,0,231,0,123,0,0,0,180,0,59,0,5,0,209,0,52,0,15,0,194,0,0,0,0,0,125,0,64,0,9,0,153,0,116,0,74,0,143,0,0,0,0,0,0,0,61,0,0,0,56,0,0,0,88,0,134,0,0,0,53,0,0,0,0,0,0,0,4,0,100,0,225,0,124,0,223,0,0,0,150,0,0,0,22,0,238,0,95,0,149,0,243,0,130,0,195,0,243,0,107,0,239,0,198,0,124,0,79,0,66,0,166,0,0,0,254,0,220,0,97,0,160,0,120,0,88,0,145,0,0,0,238,0,0,0,114,0,216,0,186,0,59,0,88,0,125,0,0,0,140,0,0,0,182,0,64,0,61,0,117,0,216,0,26,0,0,0,114,0,225,0,0,0,40,0,0,0,90,0,254,0,205,0,0,0,117,0,0,0,0,0,139,0,0,0,192,0,0,0,70,0,228,0,165,0,0,0,191,0,0,0,119,0,0,0,201,0,131,0,106,0,53,0,75,0,39,0,0,0,90,0,0,0,157,0,228,0,146,0,191,0,79,0,230,0,191,0,140,0,239,0,23,0,69,0,38,0,37,0,132,0,119,0,139,0,189,0,27,0,145,0,165,0,111,0,242,0,28,0,18,0,178,0,86,0,77,0,123,0,119,0,36,0,86,0,151,0,245,0,56,0,155,0,121,0,208,0,188,0,0,0,128,0,151,0,228,0,131,0,242,0,162,0,0,0,168,0,195,0,150,0,179,0,86,0,233,0,208,0,167,0,17,0,188,0,230,0,233,0,226,0,66,0,233,0,78,0,145,0,93,0,0,0,91,0,99,0,168,0,98,0,0,0,51,0,40,0,95,0,133,0,137,0,0,0,66,0,217,0,141,0,232,0,126,0,208,0,185,0,38,0,92,0,6,0,150,0,251,0,119,0,75,0,0,0,72,0,207,0,194,0,134,0,85,0,197,0,149,0,0,0,0,0,83,0,39,0,0,0,73,0,138,0,57,0,1,0,209,0,0,0,0,0,44,0,136,0,253,0,33,0,213,0,43,0,0,0,140,0,0,0,125,0,206,0,246,0,0,0,20,0,0,0,39,0,81,0,168,0,180,0,36,0,179,0,24,0,215,0,83,0,0,0,0,0,209,0,0,0,212,0,155,0,0,0,88,0,115,0,188,0,38,0,0,0,213,0,166,0,135,0,147,0,171,0,43,0,42,0,159,0,47,0,74,0,199,0,171,0,0,0,117,0,66,0,48,0,10,0,16,0,59,0,235,0,0,0,254,0,154,0,43,0,196,0,57,0,0,0,64,0,205,0,126,0,5,0,241,0,208,0,215,0,121,0,202,0,21,0,0,0,106,0,191,0,8,0,82,0,82,0,100,0,0,0,169,0,158,0,0,0,86,0,137,0,197,0,65,0,52,0,145,0,36,0,193,0,2,0,7,0,167,0,79,0,180,0,7,0,72,0,232,0,42,0,5,0,206,0,140,0,99,0,221,0,190,0,244,0,111,0,0,0,162,0,137,0,255,0,155,0,40,0,0,0,116,0,158,0,0,0,212,0,231,0,165,0,233,0,74,0,240,0,207,0,0,0,205,0,96,0,209,0,105,0,174,0,114,0,200,0,8,0,148,0,226,0,40,0,149,0,75,0,74,0,135,0,58,0,244,0,95,0,245,0,167,0,224,0,0,0,37,0,50,0,136,0,138,0,0,0,158,0,160,0,0,0,111,0,197,0,30,0,68,0,129,0,195,0,163,0,119,0,235,0,205,0,246,0,0,0,187,0,106,0,19,0,172,0,0,0,73,0,219,0,153,0,122,0,252,0,209,0,128,0,230,0,97,0,39,0,0,0,165,0,144,0,0,0,0,0,143,0,214,0,0,0,165,0,116,0,77,0,51,0,37,0,29,0,88,0,0,0,112,0,61,0,234,0,71,0,178,0,100,0,0,0,211,0,151,0,169,0,0,0,12,0,83,0,93,0,144,0,55,0,10,0,186,0,187,0,0,0,57,0,214,0,235,0,93,0,78,0,213,0,93,0,255,0,26,0,74,0,104,0,199,0,132,0,110,0,77,0,0,0,143,0,155,0,48,0,0,0,131,0,248,0,216,0,46,0,0,0,57,0,184,0,210,0,223,0,49,0,0,0,80,0,24,0,32,0,140,0,83,0,0,0,0,0,234,0,19,0,115,0,184,0,92,0,61,0,146,0,8,0,104,0,132,0,38,0,242,0,214,0,28,0,132,0,29,0,130,0,103,0,32,0,0,0,241,0,126,0,102,0,121,0,54,0,110,0,28,0,129,0);
signal scenario_full  : scenario_type := (219,31,250,31,139,31,187,31,124,31,159,31,96,31,27,31,93,31,111,31,214,31,135,31,13,31,203,31,248,31,199,31,48,31,234,31,36,31,190,31,176,31,40,31,242,31,242,30,28,31,34,31,34,30,107,31,73,31,239,31,239,30,239,29,140,31,206,31,122,31,56,31,56,30,250,31,205,31,205,30,189,31,185,31,92,31,85,31,190,31,56,31,42,31,54,31,63,31,140,31,138,31,105,31,35,31,178,31,178,30,54,31,215,31,12,31,245,31,26,31,26,30,26,29,185,31,185,30,49,31,22,31,56,31,56,30,132,31,159,31,186,31,233,31,238,31,232,31,107,31,117,31,152,31,156,31,143,31,221,31,3,31,247,31,114,31,153,31,153,30,9,31,102,31,111,31,190,31,136,31,234,31,65,31,98,31,216,31,216,30,114,31,176,31,51,31,51,30,211,31,193,31,193,30,238,31,4,31,21,31,21,30,166,31,106,31,175,31,128,31,42,31,80,31,22,31,22,30,81,31,226,31,150,31,110,31,110,30,47,31,177,31,177,30,194,31,140,31,182,31,169,31,136,31,78,31,78,30,28,31,4,31,159,31,165,31,115,31,110,31,110,30,190,31,121,31,121,30,152,31,61,31,61,30,214,31,57,31,15,31,15,30,1,31,145,31,83,31,83,30,245,31,245,30,245,29,52,31,154,31,154,30,230,31,185,31,132,31,132,30,132,29,225,31,162,31,124,31,110,31,10,31,27,31,27,30,60,31,11,31,227,31,90,31,147,31,222,31,137,31,107,31,240,31,80,31,193,31,56,31,56,30,56,29,56,28,165,31,165,30,41,31,115,31,24,31,156,31,155,31,197,31,146,31,209,31,42,31,234,31,87,31,74,31,241,31,241,30,180,31,180,30,28,31,136,31,136,30,46,31,248,31,58,31,130,31,226,31,22,31,20,31,20,30,243,31,243,30,43,31,170,31,142,31,198,31,74,31,56,31,67,31,132,31,151,31,229,31,30,31,206,31,204,31,167,31,167,30,13,31,20,31,199,31,73,31,101,31,103,31,7,31,102,31,178,31,255,31,132,31,136,31,235,31,217,31,128,31,71,31,65,31,39,31,168,31,168,30,90,31,13,31,79,31,79,30,187,31,187,30,20,31,67,31,52,31,129,31,191,31,150,31,23,31,11,31,92,31,34,31,34,30,195,31,246,31,121,31,93,31,197,31,35,31,239,31,51,31,51,30,51,29,14,31,152,31,152,30,152,29,88,31,185,31,43,31,43,30,114,31,15,31,162,31,97,31,126,31,227,31,121,31,121,30,33,31,255,31,220,31,212,31,124,31,79,31,38,31,238,31,131,31,182,31,182,30,85,31,32,31,191,31,195,31,181,31,246,31,155,31,155,30,107,31,82,31,29,31,173,31,173,30,190,31,177,31,14,31,26,31,26,30,26,29,64,31,64,30,64,29,116,31,118,31,2,31,2,30,229,31,100,31,121,31,89,31,104,31,188,31,151,31,217,31,40,31,40,30,174,31,76,31,7,31,189,31,25,31,25,30,25,29,120,31,118,31,210,31,210,30,2,31,2,30,250,31,193,31,193,30,193,29,213,31,100,31,226,31,130,31,7,31,4,31,66,31,108,31,22,31,5,31,133,31,133,30,221,31,4,31,150,31,231,31,231,30,183,31,88,31,238,31,183,31,167,31,141,31,141,30,106,31,211,31,211,30,5,31,190,31,111,31,111,30,111,29,111,28,80,31,239,31,85,31,217,31,217,30,231,31,231,31,123,31,123,30,180,31,59,31,5,31,209,31,52,31,15,31,194,31,194,30,194,29,125,31,64,31,9,31,153,31,116,31,74,31,143,31,143,30,143,29,143,28,61,31,61,30,56,31,56,30,88,31,134,31,134,30,53,31,53,30,53,29,53,28,4,31,100,31,225,31,124,31,223,31,223,30,150,31,150,30,22,31,238,31,95,31,149,31,243,31,130,31,195,31,243,31,107,31,239,31,198,31,124,31,79,31,66,31,166,31,166,30,254,31,220,31,97,31,160,31,120,31,88,31,145,31,145,30,238,31,238,30,114,31,216,31,186,31,59,31,88,31,125,31,125,30,140,31,140,30,182,31,64,31,61,31,117,31,216,31,26,31,26,30,114,31,225,31,225,30,40,31,40,30,90,31,254,31,205,31,205,30,117,31,117,30,117,29,139,31,139,30,192,31,192,30,70,31,228,31,165,31,165,30,191,31,191,30,119,31,119,30,201,31,131,31,106,31,53,31,75,31,39,31,39,30,90,31,90,30,157,31,228,31,146,31,191,31,79,31,230,31,191,31,140,31,239,31,23,31,69,31,38,31,37,31,132,31,119,31,139,31,189,31,27,31,145,31,165,31,111,31,242,31,28,31,18,31,178,31,86,31,77,31,123,31,119,31,36,31,86,31,151,31,245,31,56,31,155,31,121,31,208,31,188,31,188,30,128,31,151,31,228,31,131,31,242,31,162,31,162,30,168,31,195,31,150,31,179,31,86,31,233,31,208,31,167,31,17,31,188,31,230,31,233,31,226,31,66,31,233,31,78,31,145,31,93,31,93,30,91,31,99,31,168,31,98,31,98,30,51,31,40,31,95,31,133,31,137,31,137,30,66,31,217,31,141,31,232,31,126,31,208,31,185,31,38,31,92,31,6,31,150,31,251,31,119,31,75,31,75,30,72,31,207,31,194,31,134,31,85,31,197,31,149,31,149,30,149,29,83,31,39,31,39,30,73,31,138,31,57,31,1,31,209,31,209,30,209,29,44,31,136,31,253,31,33,31,213,31,43,31,43,30,140,31,140,30,125,31,206,31,246,31,246,30,20,31,20,30,39,31,81,31,168,31,180,31,36,31,179,31,24,31,215,31,83,31,83,30,83,29,209,31,209,30,212,31,155,31,155,30,88,31,115,31,188,31,38,31,38,30,213,31,166,31,135,31,147,31,171,31,43,31,42,31,159,31,47,31,74,31,199,31,171,31,171,30,117,31,66,31,48,31,10,31,16,31,59,31,235,31,235,30,254,31,154,31,43,31,196,31,57,31,57,30,64,31,205,31,126,31,5,31,241,31,208,31,215,31,121,31,202,31,21,31,21,30,106,31,191,31,8,31,82,31,82,31,100,31,100,30,169,31,158,31,158,30,86,31,137,31,197,31,65,31,52,31,145,31,36,31,193,31,2,31,7,31,167,31,79,31,180,31,7,31,72,31,232,31,42,31,5,31,206,31,140,31,99,31,221,31,190,31,244,31,111,31,111,30,162,31,137,31,255,31,155,31,40,31,40,30,116,31,158,31,158,30,212,31,231,31,165,31,233,31,74,31,240,31,207,31,207,30,205,31,96,31,209,31,105,31,174,31,114,31,200,31,8,31,148,31,226,31,40,31,149,31,75,31,74,31,135,31,58,31,244,31,95,31,245,31,167,31,224,31,224,30,37,31,50,31,136,31,138,31,138,30,158,31,160,31,160,30,111,31,197,31,30,31,68,31,129,31,195,31,163,31,119,31,235,31,205,31,246,31,246,30,187,31,106,31,19,31,172,31,172,30,73,31,219,31,153,31,122,31,252,31,209,31,128,31,230,31,97,31,39,31,39,30,165,31,144,31,144,30,144,29,143,31,214,31,214,30,165,31,116,31,77,31,51,31,37,31,29,31,88,31,88,30,112,31,61,31,234,31,71,31,178,31,100,31,100,30,211,31,151,31,169,31,169,30,12,31,83,31,93,31,144,31,55,31,10,31,186,31,187,31,187,30,57,31,214,31,235,31,93,31,78,31,213,31,93,31,255,31,26,31,74,31,104,31,199,31,132,31,110,31,77,31,77,30,143,31,155,31,48,31,48,30,131,31,248,31,216,31,46,31,46,30,57,31,184,31,210,31,223,31,49,31,49,30,80,31,24,31,32,31,140,31,83,31,83,30,83,29,234,31,19,31,115,31,184,31,92,31,61,31,146,31,8,31,104,31,132,31,38,31,242,31,214,31,28,31,132,31,29,31,130,31,103,31,32,31,32,30,241,31,126,31,102,31,121,31,54,31,110,31,28,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
