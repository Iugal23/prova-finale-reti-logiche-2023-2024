-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_757 is
end project_tb_757;

architecture project_tb_arch_757 of project_tb_757 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 760;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,66,0,194,0,122,0,81,0,98,0,132,0,96,0,10,0,155,0,180,0,182,0,165,0,51,0,36,0,33,0,0,0,255,0,0,0,179,0,0,0,201,0,94,0,226,0,90,0,72,0,179,0,124,0,130,0,71,0,0,0,35,0,21,0,42,0,113,0,142,0,197,0,20,0,0,0,0,0,89,0,145,0,133,0,78,0,54,0,165,0,116,0,0,0,210,0,210,0,27,0,157,0,226,0,250,0,0,0,0,0,0,0,97,0,95,0,6,0,236,0,229,0,159,0,0,0,16,0,114,0,215,0,101,0,244,0,234,0,84,0,20,0,54,0,119,0,179,0,250,0,165,0,188,0,3,0,108,0,0,0,220,0,128,0,191,0,30,0,250,0,73,0,117,0,65,0,59,0,234,0,51,0,88,0,223,0,32,0,144,0,56,0,32,0,168,0,0,0,16,0,0,0,0,0,238,0,198,0,12,0,163,0,0,0,230,0,234,0,188,0,55,0,148,0,46,0,4,0,146,0,69,0,93,0,215,0,99,0,241,0,158,0,0,0,133,0,146,0,14,0,118,0,218,0,13,0,92,0,167,0,82,0,193,0,0,0,0,0,193,0,230,0,186,0,0,0,68,0,88,0,85,0,0,0,65,0,107,0,0,0,33,0,143,0,222,0,84,0,142,0,0,0,129,0,131,0,149,0,209,0,85,0,254,0,211,0,34,0,171,0,68,0,123,0,13,0,62,0,6,0,0,0,228,0,0,0,117,0,181,0,0,0,19,0,124,0,0,0,0,0,137,0,131,0,0,0,0,0,93,0,170,0,27,0,0,0,0,0,9,0,42,0,132,0,198,0,213,0,91,0,11,0,198,0,176,0,151,0,147,0,0,0,143,0,239,0,150,0,45,0,165,0,124,0,236,0,0,0,0,0,14,0,0,0,221,0,210,0,221,0,202,0,224,0,187,0,61,0,99,0,0,0,125,0,72,0,0,0,200,0,83,0,0,0,230,0,200,0,0,0,47,0,34,0,77,0,145,0,251,0,22,0,79,0,235,0,85,0,76,0,242,0,0,0,253,0,176,0,152,0,133,0,155,0,209,0,74,0,232,0,0,0,0,0,0,0,0,0,222,0,65,0,147,0,241,0,141,0,205,0,122,0,170,0,185,0,0,0,27,0,120,0,139,0,145,0,139,0,191,0,0,0,0,0,125,0,60,0,0,0,246,0,92,0,233,0,215,0,115,0,230,0,164,0,57,0,0,0,42,0,38,0,160,0,56,0,0,0,44,0,144,0,171,0,0,0,157,0,23,0,188,0,0,0,0,0,179,0,134,0,230,0,108,0,203,0,22,0,60,0,166,0,31,0,3,0,190,0,0,0,28,0,204,0,65,0,76,0,170,0,239,0,179,0,170,0,111,0,182,0,252,0,247,0,30,0,176,0,188,0,0,0,101,0,0,0,209,0,196,0,217,0,132,0,0,0,176,0,180,0,0,0,0,0,0,0,200,0,174,0,16,0,23,0,0,0,33,0,111,0,224,0,161,0,26,0,12,0,0,0,186,0,238,0,63,0,20,0,85,0,164,0,215,0,21,0,78,0,96,0,0,0,122,0,113,0,31,0,146,0,111,0,150,0,89,0,0,0,37,0,114,0,223,0,242,0,0,0,0,0,172,0,203,0,0,0,237,0,0,0,148,0,137,0,221,0,117,0,254,0,0,0,77,0,157,0,211,0,0,0,194,0,139,0,65,0,172,0,0,0,55,0,131,0,63,0,115,0,245,0,228,0,155,0,66,0,70,0,0,0,0,0,0,0,0,0,0,0,136,0,63,0,171,0,20,0,109,0,252,0,0,0,238,0,145,0,0,0,185,0,134,0,188,0,127,0,0,0,30,0,150,0,141,0,52,0,31,0,63,0,0,0,42,0,141,0,153,0,0,0,245,0,21,0,217,0,69,0,203,0,35,0,246,0,134,0,0,0,101,0,218,0,0,0,0,0,0,0,148,0,236,0,239,0,33,0,0,0,140,0,0,0,66,0,202,0,19,0,99,0,29,0,112,0,176,0,22,0,239,0,247,0,0,0,132,0,183,0,118,0,102,0,206,0,222,0,3,0,168,0,6,0,204,0,7,0,68,0,0,0,135,0,174,0,226,0,0,0,254,0,133,0,239,0,80,0,194,0,0,0,186,0,0,0,119,0,107,0,196,0,0,0,110,0,95,0,69,0,0,0,0,0,166,0,171,0,52,0,205,0,247,0,0,0,114,0,209,0,226,0,17,0,147,0,0,0,21,0,0,0,212,0,209,0,0,0,180,0,0,0,0,0,39,0,195,0,0,0,131,0,107,0,221,0,77,0,75,0,0,0,56,0,0,0,127,0,75,0,71,0,201,0,43,0,0,0,0,0,117,0,0,0,0,0,172,0,167,0,199,0,155,0,145,0,0,0,232,0,13,0,12,0,159,0,0,0,190,0,130,0,83,0,0,0,0,0,101,0,203,0,34,0,249,0,229,0,127,0,0,0,167,0,39,0,62,0,141,0,6,0,0,0,12,0,163,0,128,0,35,0,135,0,194,0,112,0,0,0,0,0,140,0,139,0,0,0,178,0,210,0,0,0,0,0,162,0,148,0,24,0,207,0,86,0,110,0,175,0,54,0,231,0,47,0,114,0,141,0,236,0,49,0,61,0,83,0,104,0,143,0,88,0,184,0,0,0,118,0,226,0,251,0,93,0,35,0,0,0,119,0,115,0,0,0,34,0,75,0,0,0,0,0,50,0,128,0,120,0,38,0,184,0,147,0,116,0,107,0,118,0,59,0,36,0,248,0,214,0,0,0,0,0,62,0,102,0,154,0,100,0,0,0,169,0,3,0,28,0,87,0,32,0,237,0,0,0,0,0,92,0,44,0,195,0,0,0,0,0,0,0,187,0,96,0,187,0,0,0,0,0,149,0,140,0,0,0,99,0,60,0,193,0,111,0,120,0,29,0,142,0,235,0,37,0,12,0,62,0,187,0,0,0,223,0,251,0,223,0,0,0,218,0,0,0,67,0,0,0,53,0,46,0,134,0,15,0,118,0,193,0,62,0,0,0,0,0,108,0,55,0,0,0,106,0,54,0,0,0,137,0,200,0,192,0,203,0,129,0,123,0,25,0,5,0,189,0,116,0,251,0,21,0,0,0,109,0,247,0,121,0,7,0,117,0,94,0,98,0,0,0,29,0,53,0,97,0,232,0,246,0,210,0,232,0,164,0,59,0,239,0,29,0,97,0,155,0,113,0,215,0,169,0,182,0,175,0,230,0,228,0,23,0,0,0,76,0,251,0,0,0,0,0,0,0,7,0,0,0,0,0,0,0,232,0,209,0,0,0,98,0,0,0,0,0,240,0,111,0,165,0,30,0,99,0,228,0,59,0);
signal scenario_full  : scenario_type := (0,0,66,31,194,31,122,31,81,31,98,31,132,31,96,31,10,31,155,31,180,31,182,31,165,31,51,31,36,31,33,31,33,30,255,31,255,30,179,31,179,30,201,31,94,31,226,31,90,31,72,31,179,31,124,31,130,31,71,31,71,30,35,31,21,31,42,31,113,31,142,31,197,31,20,31,20,30,20,29,89,31,145,31,133,31,78,31,54,31,165,31,116,31,116,30,210,31,210,31,27,31,157,31,226,31,250,31,250,30,250,29,250,28,97,31,95,31,6,31,236,31,229,31,159,31,159,30,16,31,114,31,215,31,101,31,244,31,234,31,84,31,20,31,54,31,119,31,179,31,250,31,165,31,188,31,3,31,108,31,108,30,220,31,128,31,191,31,30,31,250,31,73,31,117,31,65,31,59,31,234,31,51,31,88,31,223,31,32,31,144,31,56,31,32,31,168,31,168,30,16,31,16,30,16,29,238,31,198,31,12,31,163,31,163,30,230,31,234,31,188,31,55,31,148,31,46,31,4,31,146,31,69,31,93,31,215,31,99,31,241,31,158,31,158,30,133,31,146,31,14,31,118,31,218,31,13,31,92,31,167,31,82,31,193,31,193,30,193,29,193,31,230,31,186,31,186,30,68,31,88,31,85,31,85,30,65,31,107,31,107,30,33,31,143,31,222,31,84,31,142,31,142,30,129,31,131,31,149,31,209,31,85,31,254,31,211,31,34,31,171,31,68,31,123,31,13,31,62,31,6,31,6,30,228,31,228,30,117,31,181,31,181,30,19,31,124,31,124,30,124,29,137,31,131,31,131,30,131,29,93,31,170,31,27,31,27,30,27,29,9,31,42,31,132,31,198,31,213,31,91,31,11,31,198,31,176,31,151,31,147,31,147,30,143,31,239,31,150,31,45,31,165,31,124,31,236,31,236,30,236,29,14,31,14,30,221,31,210,31,221,31,202,31,224,31,187,31,61,31,99,31,99,30,125,31,72,31,72,30,200,31,83,31,83,30,230,31,200,31,200,30,47,31,34,31,77,31,145,31,251,31,22,31,79,31,235,31,85,31,76,31,242,31,242,30,253,31,176,31,152,31,133,31,155,31,209,31,74,31,232,31,232,30,232,29,232,28,232,27,222,31,65,31,147,31,241,31,141,31,205,31,122,31,170,31,185,31,185,30,27,31,120,31,139,31,145,31,139,31,191,31,191,30,191,29,125,31,60,31,60,30,246,31,92,31,233,31,215,31,115,31,230,31,164,31,57,31,57,30,42,31,38,31,160,31,56,31,56,30,44,31,144,31,171,31,171,30,157,31,23,31,188,31,188,30,188,29,179,31,134,31,230,31,108,31,203,31,22,31,60,31,166,31,31,31,3,31,190,31,190,30,28,31,204,31,65,31,76,31,170,31,239,31,179,31,170,31,111,31,182,31,252,31,247,31,30,31,176,31,188,31,188,30,101,31,101,30,209,31,196,31,217,31,132,31,132,30,176,31,180,31,180,30,180,29,180,28,200,31,174,31,16,31,23,31,23,30,33,31,111,31,224,31,161,31,26,31,12,31,12,30,186,31,238,31,63,31,20,31,85,31,164,31,215,31,21,31,78,31,96,31,96,30,122,31,113,31,31,31,146,31,111,31,150,31,89,31,89,30,37,31,114,31,223,31,242,31,242,30,242,29,172,31,203,31,203,30,237,31,237,30,148,31,137,31,221,31,117,31,254,31,254,30,77,31,157,31,211,31,211,30,194,31,139,31,65,31,172,31,172,30,55,31,131,31,63,31,115,31,245,31,228,31,155,31,66,31,70,31,70,30,70,29,70,28,70,27,70,26,136,31,63,31,171,31,20,31,109,31,252,31,252,30,238,31,145,31,145,30,185,31,134,31,188,31,127,31,127,30,30,31,150,31,141,31,52,31,31,31,63,31,63,30,42,31,141,31,153,31,153,30,245,31,21,31,217,31,69,31,203,31,35,31,246,31,134,31,134,30,101,31,218,31,218,30,218,29,218,28,148,31,236,31,239,31,33,31,33,30,140,31,140,30,66,31,202,31,19,31,99,31,29,31,112,31,176,31,22,31,239,31,247,31,247,30,132,31,183,31,118,31,102,31,206,31,222,31,3,31,168,31,6,31,204,31,7,31,68,31,68,30,135,31,174,31,226,31,226,30,254,31,133,31,239,31,80,31,194,31,194,30,186,31,186,30,119,31,107,31,196,31,196,30,110,31,95,31,69,31,69,30,69,29,166,31,171,31,52,31,205,31,247,31,247,30,114,31,209,31,226,31,17,31,147,31,147,30,21,31,21,30,212,31,209,31,209,30,180,31,180,30,180,29,39,31,195,31,195,30,131,31,107,31,221,31,77,31,75,31,75,30,56,31,56,30,127,31,75,31,71,31,201,31,43,31,43,30,43,29,117,31,117,30,117,29,172,31,167,31,199,31,155,31,145,31,145,30,232,31,13,31,12,31,159,31,159,30,190,31,130,31,83,31,83,30,83,29,101,31,203,31,34,31,249,31,229,31,127,31,127,30,167,31,39,31,62,31,141,31,6,31,6,30,12,31,163,31,128,31,35,31,135,31,194,31,112,31,112,30,112,29,140,31,139,31,139,30,178,31,210,31,210,30,210,29,162,31,148,31,24,31,207,31,86,31,110,31,175,31,54,31,231,31,47,31,114,31,141,31,236,31,49,31,61,31,83,31,104,31,143,31,88,31,184,31,184,30,118,31,226,31,251,31,93,31,35,31,35,30,119,31,115,31,115,30,34,31,75,31,75,30,75,29,50,31,128,31,120,31,38,31,184,31,147,31,116,31,107,31,118,31,59,31,36,31,248,31,214,31,214,30,214,29,62,31,102,31,154,31,100,31,100,30,169,31,3,31,28,31,87,31,32,31,237,31,237,30,237,29,92,31,44,31,195,31,195,30,195,29,195,28,187,31,96,31,187,31,187,30,187,29,149,31,140,31,140,30,99,31,60,31,193,31,111,31,120,31,29,31,142,31,235,31,37,31,12,31,62,31,187,31,187,30,223,31,251,31,223,31,223,30,218,31,218,30,67,31,67,30,53,31,46,31,134,31,15,31,118,31,193,31,62,31,62,30,62,29,108,31,55,31,55,30,106,31,54,31,54,30,137,31,200,31,192,31,203,31,129,31,123,31,25,31,5,31,189,31,116,31,251,31,21,31,21,30,109,31,247,31,121,31,7,31,117,31,94,31,98,31,98,30,29,31,53,31,97,31,232,31,246,31,210,31,232,31,164,31,59,31,239,31,29,31,97,31,155,31,113,31,215,31,169,31,182,31,175,31,230,31,228,31,23,31,23,30,76,31,251,31,251,30,251,29,251,28,7,31,7,30,7,29,7,28,232,31,209,31,209,30,98,31,98,30,98,29,240,31,111,31,165,31,30,31,99,31,228,31,59,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
