-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_850 is
end project_tb_850;

architecture project_tb_arch_850 of project_tb_850 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 962;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (171,0,78,0,141,0,255,0,214,0,191,0,191,0,137,0,8,0,193,0,71,0,0,0,0,0,163,0,130,0,135,0,193,0,169,0,70,0,17,0,96,0,96,0,0,0,210,0,225,0,202,0,0,0,233,0,10,0,119,0,110,0,0,0,63,0,0,0,0,0,121,0,66,0,210,0,74,0,194,0,202,0,0,0,177,0,97,0,17,0,58,0,250,0,127,0,0,0,165,0,0,0,159,0,124,0,169,0,0,0,125,0,227,0,118,0,3,0,0,0,135,0,53,0,186,0,0,0,253,0,121,0,237,0,145,0,184,0,176,0,238,0,0,0,172,0,198,0,0,0,0,0,177,0,65,0,182,0,54,0,113,0,148,0,49,0,53,0,0,0,37,0,196,0,217,0,0,0,191,0,166,0,0,0,81,0,0,0,0,0,254,0,6,0,131,0,31,0,111,0,231,0,140,0,22,0,175,0,7,0,78,0,109,0,237,0,0,0,150,0,0,0,0,0,132,0,23,0,0,0,216,0,31,0,90,0,0,0,121,0,153,0,85,0,185,0,79,0,94,0,109,0,96,0,28,0,164,0,217,0,0,0,250,0,160,0,120,0,43,0,0,0,178,0,125,0,127,0,0,0,125,0,140,0,252,0,182,0,149,0,18,0,252,0,98,0,244,0,50,0,0,0,132,0,146,0,65,0,0,0,120,0,75,0,222,0,128,0,134,0,255,0,154,0,239,0,127,0,149,0,55,0,99,0,100,0,82,0,239,0,220,0,0,0,179,0,221,0,84,0,223,0,71,0,223,0,253,0,158,0,113,0,134,0,0,0,63,0,161,0,223,0,44,0,21,0,58,0,42,0,189,0,71,0,183,0,113,0,242,0,0,0,0,0,47,0,133,0,215,0,127,0,0,0,0,0,0,0,69,0,168,0,4,0,122,0,138,0,0,0,22,0,0,0,189,0,0,0,13,0,112,0,126,0,178,0,130,0,248,0,172,0,65,0,175,0,87,0,148,0,109,0,23,0,103,0,0,0,76,0,173,0,231,0,47,0,176,0,93,0,84,0,227,0,186,0,82,0,73,0,0,0,137,0,205,0,0,0,59,0,178,0,243,0,0,0,121,0,18,0,5,0,255,0,0,0,0,0,3,0,0,0,136,0,0,0,9,0,10,0,146,0,226,0,59,0,234,0,82,0,129,0,125,0,88,0,82,0,126,0,6,0,247,0,0,0,152,0,246,0,0,0,184,0,61,0,124,0,8,0,0,0,164,0,0,0,0,0,41,0,200,0,149,0,0,0,216,0,254,0,0,0,226,0,214,0,149,0,0,0,0,0,206,0,64,0,39,0,125,0,117,0,98,0,12,0,0,0,0,0,144,0,143,0,35,0,129,0,99,0,34,0,195,0,83,0,0,0,124,0,40,0,122,0,114,0,0,0,251,0,192,0,131,0,197,0,91,0,112,0,3,0,137,0,63,0,33,0,2,0,0,0,224,0,113,0,0,0,143,0,28,0,0,0,7,0,239,0,132,0,0,0,0,0,23,0,146,0,177,0,131,0,101,0,0,0,0,0,53,0,65,0,0,0,182,0,0,0,190,0,0,0,61,0,239,0,0,0,96,0,0,0,64,0,226,0,0,0,95,0,158,0,101,0,151,0,0,0,105,0,140,0,0,0,61,0,74,0,0,0,0,0,254,0,243,0,0,0,33,0,33,0,0,0,0,0,12,0,141,0,0,0,190,0,230,0,0,0,123,0,214,0,174,0,83,0,129,0,94,0,218,0,74,0,24,0,21,0,253,0,228,0,0,0,90,0,0,0,182,0,42,0,8,0,0,0,220,0,185,0,222,0,242,0,5,0,110,0,110,0,34,0,0,0,19,0,150,0,227,0,202,0,62,0,116,0,7,0,96,0,17,0,177,0,95,0,0,0,205,0,255,0,41,0,95,0,67,0,1,0,34,0,187,0,234,0,228,0,43,0,131,0,92,0,0,0,203,0,0,0,251,0,90,0,125,0,61,0,0,0,15,0,124,0,86,0,232,0,250,0,181,0,140,0,157,0,0,0,87,0,244,0,39,0,66,0,36,0,140,0,204,0,199,0,0,0,81,0,255,0,96,0,0,0,61,0,70,0,207,0,173,0,205,0,0,0,137,0,232,0,193,0,0,0,10,0,0,0,93,0,0,0,247,0,64,0,177,0,254,0,76,0,97,0,41,0,20,0,65,0,110,0,243,0,170,0,168,0,28,0,34,0,0,0,4,0,0,0,26,0,180,0,105,0,45,0,233,0,97,0,0,0,172,0,173,0,0,0,154,0,184,0,67,0,0,0,183,0,204,0,0,0,0,0,48,0,166,0,0,0,63,0,0,0,229,0,190,0,38,0,126,0,152,0,146,0,53,0,63,0,208,0,135,0,35,0,112,0,0,0,243,0,0,0,101,0,78,0,60,0,69,0,161,0,189,0,134,0,0,0,229,0,55,0,13,0,228,0,0,0,178,0,192,0,116,0,46,0,118,0,72,0,244,0,0,0,0,0,2,0,219,0,225,0,0,0,0,0,42,0,22,0,66,0,23,0,0,0,0,0,235,0,184,0,55,0,93,0,94,0,133,0,0,0,102,0,152,0,104,0,89,0,179,0,227,0,1,0,58,0,172,0,14,0,0,0,183,0,0,0,240,0,70,0,35,0,130,0,0,0,186,0,36,0,96,0,63,0,146,0,109,0,190,0,94,0,242,0,0,0,54,0,67,0,163,0,233,0,119,0,206,0,0,0,184,0,27,0,0,0,62,0,131,0,10,0,112,0,21,0,124,0,100,0,57,0,0,0,242,0,252,0,177,0,213,0,252,0,47,0,0,0,0,0,71,0,207,0,241,0,155,0,228,0,24,0,0,0,0,0,172,0,46,0,210,0,40,0,37,0,0,0,209,0,193,0,154,0,0,0,220,0,63,0,141,0,133,0,59,0,174,0,34,0,0,0,0,0,10,0,116,0,117,0,0,0,0,0,80,0,0,0,138,0,5,0,75,0,55,0,26,0,115,0,66,0,0,0,133,0,117,0,134,0,222,0,41,0,72,0,143,0,29,0,0,0,192,0,129,0,142,0,153,0,254,0,152,0,0,0,55,0,102,0,0,0,180,0,3,0,0,0,7,0,149,0,183,0,201,0,93,0,38,0,0,0,0,0,0,0,170,0,1,0,0,0,210,0,114,0,219,0,146,0,0,0,0,0,140,0,0,0,211,0,20,0,0,0,79,0,121,0,197,0,106,0,0,0,119,0,0,0,89,0,183,0,9,0,69,0,94,0,69,0,147,0,84,0,0,0,175,0,163,0,89,0,30,0,0,0,140,0,116,0,55,0,78,0,0,0,0,0,0,0,200,0,0,0,0,0,0,0,102,0,0,0,0,0,53,0,124,0,54,0,0,0,0,0,93,0,173,0,8,0,179,0,111,0,0,0,0,0,210,0,56,0,0,0,12,0,104,0,8,0,25,0,0,0,119,0,248,0,186,0,102,0,40,0,213,0,200,0,219,0,243,0,0,0,102,0,172,0,0,0,32,0,192,0,0,0,195,0,199,0,147,0,27,0,175,0,18,0,75,0,200,0,157,0,0,0,81,0,147,0,0,0,147,0,51,0,0,0,0,0,80,0,97,0,73,0,0,0,179,0,138,0,0,0,15,0,22,0,76,0,0,0,146,0,0,0,113,0,145,0,224,0,253,0,46,0,216,0,211,0,0,0,42,0,196,0,218,0,226,0,169,0,180,0,0,0,221,0,6,0,126,0,190,0,0,0,251,0,116,0,0,0,185,0,198,0,3,0,0,0,158,0,0,0,174,0,77,0,157,0,201,0,146,0,0,0,106,0,235,0,150,0,93,0,140,0,190,0,62,0,104,0,60,0,115,0,0,0,148,0,0,0,186,0,123,0,124,0,196,0,18,0,216,0,153,0,11,0,23,0,0,0,198,0,49,0,64,0,110,0,119,0,49,0,94,0,0,0,92,0,135,0,239,0,0,0,154,0,0,0,196,0,63,0,147,0,96,0,232,0,0,0,191,0,234,0,193,0,155,0,72,0,0,0,27,0,213,0,40,0,74,0,203,0,11,0,213,0,0,0,164,0,253,0,0,0,110,0,23,0,111,0,125,0,151,0,0,0,254,0,18,0,155,0,134,0,109,0,73,0,28,0,0,0,0,0,159,0,84,0,0,0,0,0,168,0,160,0,60,0,0,0,115,0,120,0,0,0,214,0,154,0,22,0,76,0,40,0,172,0,6,0,196,0,67,0,219,0,171,0,52,0,101,0,97,0,11,0,0,0);
signal scenario_full  : scenario_type := (171,31,78,31,141,31,255,31,214,31,191,31,191,31,137,31,8,31,193,31,71,31,71,30,71,29,163,31,130,31,135,31,193,31,169,31,70,31,17,31,96,31,96,31,96,30,210,31,225,31,202,31,202,30,233,31,10,31,119,31,110,31,110,30,63,31,63,30,63,29,121,31,66,31,210,31,74,31,194,31,202,31,202,30,177,31,97,31,17,31,58,31,250,31,127,31,127,30,165,31,165,30,159,31,124,31,169,31,169,30,125,31,227,31,118,31,3,31,3,30,135,31,53,31,186,31,186,30,253,31,121,31,237,31,145,31,184,31,176,31,238,31,238,30,172,31,198,31,198,30,198,29,177,31,65,31,182,31,54,31,113,31,148,31,49,31,53,31,53,30,37,31,196,31,217,31,217,30,191,31,166,31,166,30,81,31,81,30,81,29,254,31,6,31,131,31,31,31,111,31,231,31,140,31,22,31,175,31,7,31,78,31,109,31,237,31,237,30,150,31,150,30,150,29,132,31,23,31,23,30,216,31,31,31,90,31,90,30,121,31,153,31,85,31,185,31,79,31,94,31,109,31,96,31,28,31,164,31,217,31,217,30,250,31,160,31,120,31,43,31,43,30,178,31,125,31,127,31,127,30,125,31,140,31,252,31,182,31,149,31,18,31,252,31,98,31,244,31,50,31,50,30,132,31,146,31,65,31,65,30,120,31,75,31,222,31,128,31,134,31,255,31,154,31,239,31,127,31,149,31,55,31,99,31,100,31,82,31,239,31,220,31,220,30,179,31,221,31,84,31,223,31,71,31,223,31,253,31,158,31,113,31,134,31,134,30,63,31,161,31,223,31,44,31,21,31,58,31,42,31,189,31,71,31,183,31,113,31,242,31,242,30,242,29,47,31,133,31,215,31,127,31,127,30,127,29,127,28,69,31,168,31,4,31,122,31,138,31,138,30,22,31,22,30,189,31,189,30,13,31,112,31,126,31,178,31,130,31,248,31,172,31,65,31,175,31,87,31,148,31,109,31,23,31,103,31,103,30,76,31,173,31,231,31,47,31,176,31,93,31,84,31,227,31,186,31,82,31,73,31,73,30,137,31,205,31,205,30,59,31,178,31,243,31,243,30,121,31,18,31,5,31,255,31,255,30,255,29,3,31,3,30,136,31,136,30,9,31,10,31,146,31,226,31,59,31,234,31,82,31,129,31,125,31,88,31,82,31,126,31,6,31,247,31,247,30,152,31,246,31,246,30,184,31,61,31,124,31,8,31,8,30,164,31,164,30,164,29,41,31,200,31,149,31,149,30,216,31,254,31,254,30,226,31,214,31,149,31,149,30,149,29,206,31,64,31,39,31,125,31,117,31,98,31,12,31,12,30,12,29,144,31,143,31,35,31,129,31,99,31,34,31,195,31,83,31,83,30,124,31,40,31,122,31,114,31,114,30,251,31,192,31,131,31,197,31,91,31,112,31,3,31,137,31,63,31,33,31,2,31,2,30,224,31,113,31,113,30,143,31,28,31,28,30,7,31,239,31,132,31,132,30,132,29,23,31,146,31,177,31,131,31,101,31,101,30,101,29,53,31,65,31,65,30,182,31,182,30,190,31,190,30,61,31,239,31,239,30,96,31,96,30,64,31,226,31,226,30,95,31,158,31,101,31,151,31,151,30,105,31,140,31,140,30,61,31,74,31,74,30,74,29,254,31,243,31,243,30,33,31,33,31,33,30,33,29,12,31,141,31,141,30,190,31,230,31,230,30,123,31,214,31,174,31,83,31,129,31,94,31,218,31,74,31,24,31,21,31,253,31,228,31,228,30,90,31,90,30,182,31,42,31,8,31,8,30,220,31,185,31,222,31,242,31,5,31,110,31,110,31,34,31,34,30,19,31,150,31,227,31,202,31,62,31,116,31,7,31,96,31,17,31,177,31,95,31,95,30,205,31,255,31,41,31,95,31,67,31,1,31,34,31,187,31,234,31,228,31,43,31,131,31,92,31,92,30,203,31,203,30,251,31,90,31,125,31,61,31,61,30,15,31,124,31,86,31,232,31,250,31,181,31,140,31,157,31,157,30,87,31,244,31,39,31,66,31,36,31,140,31,204,31,199,31,199,30,81,31,255,31,96,31,96,30,61,31,70,31,207,31,173,31,205,31,205,30,137,31,232,31,193,31,193,30,10,31,10,30,93,31,93,30,247,31,64,31,177,31,254,31,76,31,97,31,41,31,20,31,65,31,110,31,243,31,170,31,168,31,28,31,34,31,34,30,4,31,4,30,26,31,180,31,105,31,45,31,233,31,97,31,97,30,172,31,173,31,173,30,154,31,184,31,67,31,67,30,183,31,204,31,204,30,204,29,48,31,166,31,166,30,63,31,63,30,229,31,190,31,38,31,126,31,152,31,146,31,53,31,63,31,208,31,135,31,35,31,112,31,112,30,243,31,243,30,101,31,78,31,60,31,69,31,161,31,189,31,134,31,134,30,229,31,55,31,13,31,228,31,228,30,178,31,192,31,116,31,46,31,118,31,72,31,244,31,244,30,244,29,2,31,219,31,225,31,225,30,225,29,42,31,22,31,66,31,23,31,23,30,23,29,235,31,184,31,55,31,93,31,94,31,133,31,133,30,102,31,152,31,104,31,89,31,179,31,227,31,1,31,58,31,172,31,14,31,14,30,183,31,183,30,240,31,70,31,35,31,130,31,130,30,186,31,36,31,96,31,63,31,146,31,109,31,190,31,94,31,242,31,242,30,54,31,67,31,163,31,233,31,119,31,206,31,206,30,184,31,27,31,27,30,62,31,131,31,10,31,112,31,21,31,124,31,100,31,57,31,57,30,242,31,252,31,177,31,213,31,252,31,47,31,47,30,47,29,71,31,207,31,241,31,155,31,228,31,24,31,24,30,24,29,172,31,46,31,210,31,40,31,37,31,37,30,209,31,193,31,154,31,154,30,220,31,63,31,141,31,133,31,59,31,174,31,34,31,34,30,34,29,10,31,116,31,117,31,117,30,117,29,80,31,80,30,138,31,5,31,75,31,55,31,26,31,115,31,66,31,66,30,133,31,117,31,134,31,222,31,41,31,72,31,143,31,29,31,29,30,192,31,129,31,142,31,153,31,254,31,152,31,152,30,55,31,102,31,102,30,180,31,3,31,3,30,7,31,149,31,183,31,201,31,93,31,38,31,38,30,38,29,38,28,170,31,1,31,1,30,210,31,114,31,219,31,146,31,146,30,146,29,140,31,140,30,211,31,20,31,20,30,79,31,121,31,197,31,106,31,106,30,119,31,119,30,89,31,183,31,9,31,69,31,94,31,69,31,147,31,84,31,84,30,175,31,163,31,89,31,30,31,30,30,140,31,116,31,55,31,78,31,78,30,78,29,78,28,200,31,200,30,200,29,200,28,102,31,102,30,102,29,53,31,124,31,54,31,54,30,54,29,93,31,173,31,8,31,179,31,111,31,111,30,111,29,210,31,56,31,56,30,12,31,104,31,8,31,25,31,25,30,119,31,248,31,186,31,102,31,40,31,213,31,200,31,219,31,243,31,243,30,102,31,172,31,172,30,32,31,192,31,192,30,195,31,199,31,147,31,27,31,175,31,18,31,75,31,200,31,157,31,157,30,81,31,147,31,147,30,147,31,51,31,51,30,51,29,80,31,97,31,73,31,73,30,179,31,138,31,138,30,15,31,22,31,76,31,76,30,146,31,146,30,113,31,145,31,224,31,253,31,46,31,216,31,211,31,211,30,42,31,196,31,218,31,226,31,169,31,180,31,180,30,221,31,6,31,126,31,190,31,190,30,251,31,116,31,116,30,185,31,198,31,3,31,3,30,158,31,158,30,174,31,77,31,157,31,201,31,146,31,146,30,106,31,235,31,150,31,93,31,140,31,190,31,62,31,104,31,60,31,115,31,115,30,148,31,148,30,186,31,123,31,124,31,196,31,18,31,216,31,153,31,11,31,23,31,23,30,198,31,49,31,64,31,110,31,119,31,49,31,94,31,94,30,92,31,135,31,239,31,239,30,154,31,154,30,196,31,63,31,147,31,96,31,232,31,232,30,191,31,234,31,193,31,155,31,72,31,72,30,27,31,213,31,40,31,74,31,203,31,11,31,213,31,213,30,164,31,253,31,253,30,110,31,23,31,111,31,125,31,151,31,151,30,254,31,18,31,155,31,134,31,109,31,73,31,28,31,28,30,28,29,159,31,84,31,84,30,84,29,168,31,160,31,60,31,60,30,115,31,120,31,120,30,214,31,154,31,22,31,76,31,40,31,172,31,6,31,196,31,67,31,219,31,171,31,52,31,101,31,97,31,11,31,11,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
