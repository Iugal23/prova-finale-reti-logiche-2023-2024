-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_191 is
end project_tb_191;

architecture project_tb_arch_191 of project_tb_191 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 825;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,77,0,163,0,123,0,128,0,253,0,108,0,255,0,123,0,0,0,210,0,202,0,63,0,57,0,194,0,149,0,47,0,234,0,255,0,113,0,222,0,46,0,226,0,97,0,53,0,0,0,196,0,19,0,0,0,0,0,251,0,72,0,117,0,110,0,158,0,0,0,0,0,232,0,152,0,10,0,17,0,86,0,153,0,146,0,122,0,203,0,115,0,251,0,159,0,151,0,254,0,184,0,0,0,53,0,225,0,87,0,195,0,4,0,148,0,98,0,218,0,103,0,255,0,0,0,44,0,0,0,0,0,42,0,84,0,0,0,151,0,72,0,232,0,207,0,0,0,140,0,38,0,0,0,0,0,0,0,169,0,87,0,175,0,243,0,0,0,131,0,104,0,41,0,82,0,137,0,108,0,42,0,192,0,0,0,166,0,212,0,195,0,94,0,129,0,0,0,27,0,71,0,0,0,0,0,96,0,154,0,179,0,230,0,0,0,146,0,159,0,23,0,71,0,0,0,77,0,112,0,158,0,46,0,72,0,234,0,107,0,0,0,36,0,36,0,48,0,0,0,226,0,170,0,199,0,179,0,229,0,0,0,127,0,117,0,52,0,142,0,0,0,197,0,132,0,221,0,214,0,159,0,163,0,74,0,176,0,63,0,16,0,39,0,202,0,55,0,210,0,140,0,125,0,89,0,250,0,88,0,0,0,205,0,84,0,64,0,231,0,165,0,0,0,0,0,40,0,234,0,114,0,0,0,246,0,219,0,150,0,51,0,0,0,0,0,177,0,160,0,245,0,124,0,165,0,200,0,144,0,113,0,136,0,0,0,100,0,21,0,0,0,243,0,221,0,0,0,0,0,134,0,233,0,0,0,140,0,96,0,0,0,174,0,203,0,186,0,160,0,158,0,66,0,225,0,43,0,0,0,176,0,42,0,103,0,135,0,0,0,90,0,228,0,141,0,45,0,204,0,0,0,155,0,196,0,0,0,213,0,37,0,0,0,33,0,62,0,157,0,245,0,123,0,1,0,59,0,11,0,226,0,50,0,83,0,0,0,35,0,148,0,147,0,0,0,155,0,155,0,197,0,38,0,55,0,0,0,153,0,87,0,184,0,0,0,52,0,128,0,104,0,164,0,191,0,224,0,253,0,18,0,56,0,125,0,0,0,153,0,213,0,249,0,0,0,163,0,232,0,89,0,227,0,227,0,0,0,0,0,83,0,166,0,16,0,132,0,25,0,109,0,63,0,222,0,0,0,250,0,0,0,26,0,141,0,28,0,0,0,43,0,0,0,36,0,212,0,0,0,179,0,99,0,50,0,151,0,50,0,192,0,154,0,136,0,76,0,74,0,181,0,91,0,0,0,237,0,249,0,0,0,183,0,22,0,252,0,0,0,0,0,50,0,116,0,151,0,134,0,163,0,187,0,70,0,193,0,0,0,50,0,174,0,39,0,192,0,18,0,218,0,129,0,78,0,0,0,0,0,0,0,78,0,89,0,222,0,68,0,110,0,6,0,209,0,153,0,220,0,87,0,199,0,80,0,85,0,118,0,0,0,241,0,0,0,0,0,71,0,0,0,48,0,57,0,0,0,0,0,105,0,199,0,210,0,209,0,101,0,0,0,159,0,146,0,72,0,0,0,211,0,56,0,113,0,0,0,0,0,161,0,49,0,162,0,76,0,8,0,32,0,147,0,184,0,0,0,255,0,209,0,216,0,225,0,0,0,234,0,0,0,171,0,0,0,78,0,156,0,34,0,0,0,14,0,0,0,227,0,250,0,142,0,191,0,100,0,52,0,0,0,84,0,140,0,129,0,0,0,48,0,111,0,92,0,100,0,186,0,243,0,236,0,95,0,197,0,0,0,213,0,223,0,0,0,21,0,93,0,214,0,83,0,0,0,208,0,196,0,0,0,64,0,11,0,127,0,116,0,61,0,201,0,240,0,121,0,167,0,231,0,72,0,76,0,0,0,154,0,136,0,9,0,196,0,205,0,122,0,48,0,171,0,231,0,99,0,233,0,216,0,0,0,0,0,51,0,0,0,0,0,217,0,0,0,192,0,180,0,85,0,251,0,54,0,230,0,105,0,70,0,63,0,48,0,105,0,160,0,196,0,75,0,0,0,232,0,236,0,111,0,101,0,206,0,22,0,21,0,24,0,35,0,109,0,153,0,0,0,75,0,48,0,53,0,86,0,0,0,109,0,0,0,176,0,221,0,2,0,32,0,98,0,146,0,74,0,11,0,60,0,193,0,254,0,2,0,55,0,104,0,0,0,0,0,89,0,36,0,0,0,124,0,11,0,33,0,142,0,177,0,0,0,133,0,157,0,126,0,58,0,209,0,22,0,214,0,0,0,57,0,207,0,203,0,80,0,140,0,110,0,0,0,154,0,0,0,242,0,90,0,233,0,0,0,81,0,47,0,139,0,235,0,0,0,233,0,4,0,239,0,51,0,70,0,70,0,196,0,0,0,0,0,232,0,144,0,53,0,254,0,0,0,35,0,0,0,0,0,90,0,72,0,219,0,19,0,101,0,107,0,124,0,0,0,0,0,104,0,13,0,122,0,52,0,46,0,160,0,65,0,0,0,221,0,229,0,0,0,77,0,22,0,219,0,94,0,0,0,147,0,242,0,252,0,192,0,192,0,33,0,178,0,130,0,201,0,0,0,202,0,30,0,143,0,141,0,61,0,177,0,88,0,238,0,69,0,137,0,63,0,159,0,124,0,25,0,59,0,0,0,67,0,37,0,43,0,163,0,232,0,232,0,180,0,37,0,91,0,0,0,137,0,29,0,175,0,90,0,191,0,94,0,189,0,5,0,190,0,0,0,123,0,126,0,0,0,252,0,95,0,225,0,0,0,19,0,140,0,0,0,128,0,195,0,52,0,83,0,3,0,222,0,251,0,230,0,191,0,250,0,0,0,234,0,251,0,0,0,165,0,49,0,152,0,66,0,0,0,232,0,132,0,39,0,0,0,64,0,84,0,76,0,108,0,163,0,71,0,75,0,120,0,13,0,46,0,141,0,101,0,100,0,0,0,142,0,10,0,187,0,0,0,0,0,87,0,196,0,49,0,22,0,0,0,0,0,52,0,61,0,0,0,143,0,75,0,93,0,49,0,138,0,49,0,51,0,156,0,196,0,82,0,0,0,20,0,0,0,50,0,245,0,79,0,41,0,123,0,0,0,235,0,201,0,71,0,222,0,207,0,105,0,174,0,81,0,143,0,0,0,82,0,191,0,241,0,171,0,10,0,0,0,103,0,0,0,0,0,255,0,0,0,0,0,142,0,232,0,229,0,33,0,232,0,0,0,108,0,157,0,1,0,59,0,129,0,0,0,0,0,78,0,181,0,159,0,188,0,26,0,81,0,221,0,0,0,160,0,0,0,231,0,175,0,0,0,205,0,233,0,5,0,117,0,147,0,37,0,40,0,0,0,90,0,201,0,50,0,173,0,47,0,0,0,52,0,0,0,135,0,228,0,189,0,0,0,0,0,76,0,0,0,209,0,0,0,175,0,124,0,190,0,4,0,128,0,131,0,0,0,73,0,146,0,108,0,17,0,0,0,158,0,197,0,90,0,0,0,0,0,163,0,4,0,125,0,60,0,96,0,230,0,227,0,212,0,145,0,58,0,19,0,230,0,19,0,209,0,20,0,0,0,219,0,48,0,0,0,103,0,154,0,44,0,0,0);
signal scenario_full  : scenario_type := (134,31,77,31,163,31,123,31,128,31,253,31,108,31,255,31,123,31,123,30,210,31,202,31,63,31,57,31,194,31,149,31,47,31,234,31,255,31,113,31,222,31,46,31,226,31,97,31,53,31,53,30,196,31,19,31,19,30,19,29,251,31,72,31,117,31,110,31,158,31,158,30,158,29,232,31,152,31,10,31,17,31,86,31,153,31,146,31,122,31,203,31,115,31,251,31,159,31,151,31,254,31,184,31,184,30,53,31,225,31,87,31,195,31,4,31,148,31,98,31,218,31,103,31,255,31,255,30,44,31,44,30,44,29,42,31,84,31,84,30,151,31,72,31,232,31,207,31,207,30,140,31,38,31,38,30,38,29,38,28,169,31,87,31,175,31,243,31,243,30,131,31,104,31,41,31,82,31,137,31,108,31,42,31,192,31,192,30,166,31,212,31,195,31,94,31,129,31,129,30,27,31,71,31,71,30,71,29,96,31,154,31,179,31,230,31,230,30,146,31,159,31,23,31,71,31,71,30,77,31,112,31,158,31,46,31,72,31,234,31,107,31,107,30,36,31,36,31,48,31,48,30,226,31,170,31,199,31,179,31,229,31,229,30,127,31,117,31,52,31,142,31,142,30,197,31,132,31,221,31,214,31,159,31,163,31,74,31,176,31,63,31,16,31,39,31,202,31,55,31,210,31,140,31,125,31,89,31,250,31,88,31,88,30,205,31,84,31,64,31,231,31,165,31,165,30,165,29,40,31,234,31,114,31,114,30,246,31,219,31,150,31,51,31,51,30,51,29,177,31,160,31,245,31,124,31,165,31,200,31,144,31,113,31,136,31,136,30,100,31,21,31,21,30,243,31,221,31,221,30,221,29,134,31,233,31,233,30,140,31,96,31,96,30,174,31,203,31,186,31,160,31,158,31,66,31,225,31,43,31,43,30,176,31,42,31,103,31,135,31,135,30,90,31,228,31,141,31,45,31,204,31,204,30,155,31,196,31,196,30,213,31,37,31,37,30,33,31,62,31,157,31,245,31,123,31,1,31,59,31,11,31,226,31,50,31,83,31,83,30,35,31,148,31,147,31,147,30,155,31,155,31,197,31,38,31,55,31,55,30,153,31,87,31,184,31,184,30,52,31,128,31,104,31,164,31,191,31,224,31,253,31,18,31,56,31,125,31,125,30,153,31,213,31,249,31,249,30,163,31,232,31,89,31,227,31,227,31,227,30,227,29,83,31,166,31,16,31,132,31,25,31,109,31,63,31,222,31,222,30,250,31,250,30,26,31,141,31,28,31,28,30,43,31,43,30,36,31,212,31,212,30,179,31,99,31,50,31,151,31,50,31,192,31,154,31,136,31,76,31,74,31,181,31,91,31,91,30,237,31,249,31,249,30,183,31,22,31,252,31,252,30,252,29,50,31,116,31,151,31,134,31,163,31,187,31,70,31,193,31,193,30,50,31,174,31,39,31,192,31,18,31,218,31,129,31,78,31,78,30,78,29,78,28,78,31,89,31,222,31,68,31,110,31,6,31,209,31,153,31,220,31,87,31,199,31,80,31,85,31,118,31,118,30,241,31,241,30,241,29,71,31,71,30,48,31,57,31,57,30,57,29,105,31,199,31,210,31,209,31,101,31,101,30,159,31,146,31,72,31,72,30,211,31,56,31,113,31,113,30,113,29,161,31,49,31,162,31,76,31,8,31,32,31,147,31,184,31,184,30,255,31,209,31,216,31,225,31,225,30,234,31,234,30,171,31,171,30,78,31,156,31,34,31,34,30,14,31,14,30,227,31,250,31,142,31,191,31,100,31,52,31,52,30,84,31,140,31,129,31,129,30,48,31,111,31,92,31,100,31,186,31,243,31,236,31,95,31,197,31,197,30,213,31,223,31,223,30,21,31,93,31,214,31,83,31,83,30,208,31,196,31,196,30,64,31,11,31,127,31,116,31,61,31,201,31,240,31,121,31,167,31,231,31,72,31,76,31,76,30,154,31,136,31,9,31,196,31,205,31,122,31,48,31,171,31,231,31,99,31,233,31,216,31,216,30,216,29,51,31,51,30,51,29,217,31,217,30,192,31,180,31,85,31,251,31,54,31,230,31,105,31,70,31,63,31,48,31,105,31,160,31,196,31,75,31,75,30,232,31,236,31,111,31,101,31,206,31,22,31,21,31,24,31,35,31,109,31,153,31,153,30,75,31,48,31,53,31,86,31,86,30,109,31,109,30,176,31,221,31,2,31,32,31,98,31,146,31,74,31,11,31,60,31,193,31,254,31,2,31,55,31,104,31,104,30,104,29,89,31,36,31,36,30,124,31,11,31,33,31,142,31,177,31,177,30,133,31,157,31,126,31,58,31,209,31,22,31,214,31,214,30,57,31,207,31,203,31,80,31,140,31,110,31,110,30,154,31,154,30,242,31,90,31,233,31,233,30,81,31,47,31,139,31,235,31,235,30,233,31,4,31,239,31,51,31,70,31,70,31,196,31,196,30,196,29,232,31,144,31,53,31,254,31,254,30,35,31,35,30,35,29,90,31,72,31,219,31,19,31,101,31,107,31,124,31,124,30,124,29,104,31,13,31,122,31,52,31,46,31,160,31,65,31,65,30,221,31,229,31,229,30,77,31,22,31,219,31,94,31,94,30,147,31,242,31,252,31,192,31,192,31,33,31,178,31,130,31,201,31,201,30,202,31,30,31,143,31,141,31,61,31,177,31,88,31,238,31,69,31,137,31,63,31,159,31,124,31,25,31,59,31,59,30,67,31,37,31,43,31,163,31,232,31,232,31,180,31,37,31,91,31,91,30,137,31,29,31,175,31,90,31,191,31,94,31,189,31,5,31,190,31,190,30,123,31,126,31,126,30,252,31,95,31,225,31,225,30,19,31,140,31,140,30,128,31,195,31,52,31,83,31,3,31,222,31,251,31,230,31,191,31,250,31,250,30,234,31,251,31,251,30,165,31,49,31,152,31,66,31,66,30,232,31,132,31,39,31,39,30,64,31,84,31,76,31,108,31,163,31,71,31,75,31,120,31,13,31,46,31,141,31,101,31,100,31,100,30,142,31,10,31,187,31,187,30,187,29,87,31,196,31,49,31,22,31,22,30,22,29,52,31,61,31,61,30,143,31,75,31,93,31,49,31,138,31,49,31,51,31,156,31,196,31,82,31,82,30,20,31,20,30,50,31,245,31,79,31,41,31,123,31,123,30,235,31,201,31,71,31,222,31,207,31,105,31,174,31,81,31,143,31,143,30,82,31,191,31,241,31,171,31,10,31,10,30,103,31,103,30,103,29,255,31,255,30,255,29,142,31,232,31,229,31,33,31,232,31,232,30,108,31,157,31,1,31,59,31,129,31,129,30,129,29,78,31,181,31,159,31,188,31,26,31,81,31,221,31,221,30,160,31,160,30,231,31,175,31,175,30,205,31,233,31,5,31,117,31,147,31,37,31,40,31,40,30,90,31,201,31,50,31,173,31,47,31,47,30,52,31,52,30,135,31,228,31,189,31,189,30,189,29,76,31,76,30,209,31,209,30,175,31,124,31,190,31,4,31,128,31,131,31,131,30,73,31,146,31,108,31,17,31,17,30,158,31,197,31,90,31,90,30,90,29,163,31,4,31,125,31,60,31,96,31,230,31,227,31,212,31,145,31,58,31,19,31,230,31,19,31,209,31,20,31,20,30,219,31,48,31,48,30,103,31,154,31,44,31,44,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
