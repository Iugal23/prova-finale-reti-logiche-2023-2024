-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1006;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (183,0,21,0,123,0,195,0,2,0,162,0,148,0,78,0,33,0,102,0,140,0,0,0,0,0,0,0,117,0,106,0,0,0,133,0,0,0,180,0,120,0,111,0,71,0,0,0,156,0,0,0,154,0,36,0,0,0,60,0,189,0,139,0,0,0,223,0,0,0,56,0,0,0,106,0,96,0,101,0,108,0,17,0,81,0,78,0,0,0,0,0,58,0,0,0,82,0,15,0,0,0,119,0,166,0,82,0,37,0,118,0,24,0,175,0,166,0,151,0,142,0,122,0,156,0,247,0,248,0,111,0,0,0,203,0,0,0,106,0,237,0,0,0,0,0,169,0,0,0,167,0,75,0,91,0,222,0,0,0,205,0,138,0,0,0,96,0,0,0,0,0,170,0,98,0,59,0,68,0,38,0,166,0,172,0,26,0,33,0,138,0,173,0,0,0,50,0,181,0,36,0,0,0,185,0,125,0,0,0,185,0,74,0,0,0,0,0,100,0,34,0,72,0,255,0,5,0,192,0,153,0,61,0,201,0,0,0,127,0,7,0,46,0,32,0,159,0,183,0,210,0,203,0,15,0,0,0,0,0,223,0,178,0,180,0,99,0,129,0,104,0,0,0,147,0,196,0,170,0,169,0,212,0,182,0,133,0,27,0,175,0,0,0,146,0,175,0,234,0,184,0,113,0,194,0,159,0,66,0,173,0,63,0,239,0,78,0,0,0,0,0,0,0,155,0,129,0,0,0,36,0,88,0,247,0,197,0,0,0,15,0,88,0,0,0,153,0,30,0,193,0,0,0,112,0,197,0,108,0,0,0,47,0,20,0,0,0,0,0,118,0,0,0,234,0,144,0,69,0,98,0,0,0,0,0,0,0,198,0,164,0,32,0,0,0,118,0,184,0,71,0,109,0,207,0,0,0,58,0,0,0,0,0,94,0,214,0,104,0,21,0,52,0,210,0,0,0,0,0,147,0,214,0,23,0,49,0,144,0,74,0,241,0,115,0,101,0,178,0,206,0,198,0,244,0,97,0,0,0,72,0,0,0,209,0,253,0,205,0,231,0,207,0,0,0,125,0,60,0,0,0,163,0,26,0,160,0,156,0,33,0,26,0,155,0,99,0,32,0,0,0,28,0,80,0,235,0,0,0,42,0,121,0,11,0,189,0,220,0,34,0,171,0,109,0,0,0,61,0,231,0,230,0,66,0,11,0,35,0,44,0,66,0,192,0,253,0,0,0,4,0,172,0,192,0,0,0,133,0,0,0,200,0,0,0,252,0,0,0,58,0,188,0,0,0,0,0,225,0,197,0,210,0,0,0,55,0,191,0,132,0,242,0,0,0,0,0,0,0,0,0,69,0,0,0,0,0,100,0,0,0,16,0,0,0,153,0,0,0,234,0,211,0,91,0,133,0,98,0,121,0,180,0,0,0,249,0,0,0,170,0,0,0,168,0,239,0,74,0,244,0,29,0,223,0,79,0,143,0,0,0,212,0,88,0,163,0,0,0,213,0,225,0,0,0,25,0,95,0,51,0,96,0,43,0,76,0,0,0,236,0,224,0,169,0,178,0,29,0,229,0,217,0,0,0,0,0,0,0,160,0,165,0,27,0,71,0,196,0,66,0,125,0,34,0,180,0,29,0,38,0,137,0,31,0,95,0,55,0,220,0,111,0,101,0,192,0,145,0,0,0,0,0,231,0,0,0,99,0,0,0,164,0,224,0,0,0,72,0,0,0,208,0,208,0,152,0,93,0,204,0,14,0,28,0,0,0,102,0,177,0,45,0,160,0,38,0,185,0,22,0,172,0,222,0,161,0,3,0,2,0,49,0,46,0,159,0,197,0,100,0,197,0,68,0,130,0,0,0,206,0,251,0,0,0,86,0,0,0,109,0,225,0,206,0,223,0,12,0,244,0,44,0,97,0,9,0,200,0,68,0,87,0,182,0,182,0,170,0,87,0,0,0,135,0,42,0,240,0,14,0,47,0,92,0,148,0,0,0,0,0,208,0,91,0,0,0,118,0,217,0,169,0,187,0,154,0,238,0,69,0,0,0,114,0,4,0,196,0,0,0,0,0,229,0,0,0,17,0,205,0,235,0,167,0,154,0,18,0,0,0,20,0,98,0,0,0,137,0,103,0,171,0,210,0,0,0,234,0,54,0,0,0,0,0,33,0,0,0,93,0,143,0,111,0,83,0,116,0,97,0,139,0,101,0,108,0,0,0,140,0,209,0,31,0,109,0,100,0,210,0,230,0,192,0,172,0,82,0,57,0,29,0,27,0,235,0,218,0,92,0,177,0,108,0,32,0,125,0,73,0,112,0,0,0,0,0,0,0,68,0,191,0,0,0,129,0,0,0,147,0,217,0,0,0,12,0,241,0,208,0,191,0,212,0,84,0,0,0,0,0,9,0,184,0,80,0,61,0,148,0,56,0,14,0,116,0,36,0,29,0,152,0,84,0,0,0,243,0,0,0,122,0,37,0,240,0,184,0,28,0,227,0,220,0,121,0,0,0,178,0,46,0,122,0,0,0,90,0,223,0,35,0,137,0,0,0,79,0,93,0,251,0,176,0,71,0,175,0,34,0,73,0,235,0,51,0,41,0,92,0,136,0,107,0,109,0,187,0,252,0,169,0,0,0,162,0,134,0,136,0,67,0,0,0,59,0,133,0,123,0,102,0,157,0,230,0,0,0,69,0,63,0,182,0,0,0,228,0,38,0,0,0,124,0,0,0,161,0,194,0,25,0,8,0,195,0,104,0,25,0,0,0,203,0,208,0,179,0,210,0,22,0,0,0,0,0,244,0,23,0,40,0,92,0,58,0,204,0,111,0,160,0,196,0,0,0,0,0,82,0,145,0,0,0,170,0,7,0,231,0,85,0,0,0,0,0,0,0,13,0,215,0,122,0,61,0,190,0,133,0,20,0,245,0,121,0,166,0,242,0,142,0,232,0,0,0,36,0,0,0,4,0,226,0,0,0,0,0,0,0,145,0,0,0,154,0,12,0,95,0,214,0,128,0,0,0,144,0,68,0,251,0,135,0,0,0,0,0,30,0,0,0,21,0,242,0,255,0,0,0,152,0,136,0,66,0,0,0,0,0,236,0,25,0,50,0,39,0,66,0,67,0,214,0,0,0,160,0,176,0,41,0,26,0,116,0,0,0,169,0,235,0,204,0,158,0,255,0,0,0,0,0,66,0,0,0,207,0,0,0,76,0,75,0,127,0,79,0,113,0,7,0,208,0,69,0,147,0,113,0,123,0,29,0,168,0,224,0,195,0,0,0,179,0,0,0,181,0,218,0,181,0,85,0,140,0,70,0,244,0,5,0,245,0,222,0,1,0,99,0,247,0,245,0,166,0,10,0,139,0,0,0,0,0,42,0,249,0,210,0,145,0,142,0,243,0,228,0,0,0,49,0,0,0,53,0,99,0,89,0,146,0,199,0,242,0,0,0,178,0,187,0,0,0,0,0,0,0,63,0,154,0,31,0,207,0,168,0,35,0,202,0,90,0,0,0,157,0,14,0,140,0,83,0,176,0,193,0,203,0,33,0,243,0,71,0,5,0,2,0,79,0,0,0,113,0,137,0,43,0,198,0,209,0,0,0,229,0,6,0,58,0,98,0,89,0,203,0,113,0,37,0,0,0,69,0,155,0,20,0,43,0,124,0,0,0,205,0,253,0,209,0,184,0,79,0,124,0,143,0,85,0,0,0,99,0,57,0,56,0,183,0,200,0,0,0,184,0,142,0,122,0,243,0,124,0,250,0,138,0,0,0,0,0,9,0,0,0,0,0,0,0,49,0,176,0,0,0,0,0,205,0,98,0,124,0,213,0,0,0,38,0,104,0,194,0,0,0,126,0,194,0,220,0,139,0,172,0,3,0,245,0,169,0,20,0,155,0,32,0,0,0,172,0,0,0,105,0,128,0,55,0,123,0,109,0,0,0,244,0,202,0,25,0,150,0,53,0,99,0,46,0,180,0,146,0,0,0,25,0,109,0,37,0,85,0,123,0,0,0,41,0,230,0,164,0,102,0,105,0,216,0,161,0,234,0,77,0,229,0,123,0,0,0,127,0,228,0,0,0,208,0,146,0,11,0,167,0,0,0,0,0,39,0,153,0,179,0,231,0,52,0,1,0,219,0,170,0,0,0,35,0,149,0,13,0,196,0,110,0,36,0,221,0,66,0,187,0,40,0,192,0,88,0,9,0,0,0,116,0,0,0,0,0,34,0,120,0,239,0,20,0,0,0,108,0,52,0,0,0,131,0,200,0,123,0,96,0,195,0,106,0,24,0,0,0,181,0,0,0,79,0,142,0,196,0,0,0,89,0,0,0,170,0,181,0,118,0,221,0,0,0,107,0,222,0,97,0,150,0,198,0,253,0,179,0,234,0,113,0,4,0,250,0,218,0,255,0,166,0,192,0,25,0,101,0,149,0,170,0,133,0,202,0,64,0,216,0,0,0,192,0,118,0,0,0,153,0,110,0,2,0,0,0,134,0,5,0,140,0);
signal scenario_full  : scenario_type := (183,31,21,31,123,31,195,31,2,31,162,31,148,31,78,31,33,31,102,31,140,31,140,30,140,29,140,28,117,31,106,31,106,30,133,31,133,30,180,31,120,31,111,31,71,31,71,30,156,31,156,30,154,31,36,31,36,30,60,31,189,31,139,31,139,30,223,31,223,30,56,31,56,30,106,31,96,31,101,31,108,31,17,31,81,31,78,31,78,30,78,29,58,31,58,30,82,31,15,31,15,30,119,31,166,31,82,31,37,31,118,31,24,31,175,31,166,31,151,31,142,31,122,31,156,31,247,31,248,31,111,31,111,30,203,31,203,30,106,31,237,31,237,30,237,29,169,31,169,30,167,31,75,31,91,31,222,31,222,30,205,31,138,31,138,30,96,31,96,30,96,29,170,31,98,31,59,31,68,31,38,31,166,31,172,31,26,31,33,31,138,31,173,31,173,30,50,31,181,31,36,31,36,30,185,31,125,31,125,30,185,31,74,31,74,30,74,29,100,31,34,31,72,31,255,31,5,31,192,31,153,31,61,31,201,31,201,30,127,31,7,31,46,31,32,31,159,31,183,31,210,31,203,31,15,31,15,30,15,29,223,31,178,31,180,31,99,31,129,31,104,31,104,30,147,31,196,31,170,31,169,31,212,31,182,31,133,31,27,31,175,31,175,30,146,31,175,31,234,31,184,31,113,31,194,31,159,31,66,31,173,31,63,31,239,31,78,31,78,30,78,29,78,28,155,31,129,31,129,30,36,31,88,31,247,31,197,31,197,30,15,31,88,31,88,30,153,31,30,31,193,31,193,30,112,31,197,31,108,31,108,30,47,31,20,31,20,30,20,29,118,31,118,30,234,31,144,31,69,31,98,31,98,30,98,29,98,28,198,31,164,31,32,31,32,30,118,31,184,31,71,31,109,31,207,31,207,30,58,31,58,30,58,29,94,31,214,31,104,31,21,31,52,31,210,31,210,30,210,29,147,31,214,31,23,31,49,31,144,31,74,31,241,31,115,31,101,31,178,31,206,31,198,31,244,31,97,31,97,30,72,31,72,30,209,31,253,31,205,31,231,31,207,31,207,30,125,31,60,31,60,30,163,31,26,31,160,31,156,31,33,31,26,31,155,31,99,31,32,31,32,30,28,31,80,31,235,31,235,30,42,31,121,31,11,31,189,31,220,31,34,31,171,31,109,31,109,30,61,31,231,31,230,31,66,31,11,31,35,31,44,31,66,31,192,31,253,31,253,30,4,31,172,31,192,31,192,30,133,31,133,30,200,31,200,30,252,31,252,30,58,31,188,31,188,30,188,29,225,31,197,31,210,31,210,30,55,31,191,31,132,31,242,31,242,30,242,29,242,28,242,27,69,31,69,30,69,29,100,31,100,30,16,31,16,30,153,31,153,30,234,31,211,31,91,31,133,31,98,31,121,31,180,31,180,30,249,31,249,30,170,31,170,30,168,31,239,31,74,31,244,31,29,31,223,31,79,31,143,31,143,30,212,31,88,31,163,31,163,30,213,31,225,31,225,30,25,31,95,31,51,31,96,31,43,31,76,31,76,30,236,31,224,31,169,31,178,31,29,31,229,31,217,31,217,30,217,29,217,28,160,31,165,31,27,31,71,31,196,31,66,31,125,31,34,31,180,31,29,31,38,31,137,31,31,31,95,31,55,31,220,31,111,31,101,31,192,31,145,31,145,30,145,29,231,31,231,30,99,31,99,30,164,31,224,31,224,30,72,31,72,30,208,31,208,31,152,31,93,31,204,31,14,31,28,31,28,30,102,31,177,31,45,31,160,31,38,31,185,31,22,31,172,31,222,31,161,31,3,31,2,31,49,31,46,31,159,31,197,31,100,31,197,31,68,31,130,31,130,30,206,31,251,31,251,30,86,31,86,30,109,31,225,31,206,31,223,31,12,31,244,31,44,31,97,31,9,31,200,31,68,31,87,31,182,31,182,31,170,31,87,31,87,30,135,31,42,31,240,31,14,31,47,31,92,31,148,31,148,30,148,29,208,31,91,31,91,30,118,31,217,31,169,31,187,31,154,31,238,31,69,31,69,30,114,31,4,31,196,31,196,30,196,29,229,31,229,30,17,31,205,31,235,31,167,31,154,31,18,31,18,30,20,31,98,31,98,30,137,31,103,31,171,31,210,31,210,30,234,31,54,31,54,30,54,29,33,31,33,30,93,31,143,31,111,31,83,31,116,31,97,31,139,31,101,31,108,31,108,30,140,31,209,31,31,31,109,31,100,31,210,31,230,31,192,31,172,31,82,31,57,31,29,31,27,31,235,31,218,31,92,31,177,31,108,31,32,31,125,31,73,31,112,31,112,30,112,29,112,28,68,31,191,31,191,30,129,31,129,30,147,31,217,31,217,30,12,31,241,31,208,31,191,31,212,31,84,31,84,30,84,29,9,31,184,31,80,31,61,31,148,31,56,31,14,31,116,31,36,31,29,31,152,31,84,31,84,30,243,31,243,30,122,31,37,31,240,31,184,31,28,31,227,31,220,31,121,31,121,30,178,31,46,31,122,31,122,30,90,31,223,31,35,31,137,31,137,30,79,31,93,31,251,31,176,31,71,31,175,31,34,31,73,31,235,31,51,31,41,31,92,31,136,31,107,31,109,31,187,31,252,31,169,31,169,30,162,31,134,31,136,31,67,31,67,30,59,31,133,31,123,31,102,31,157,31,230,31,230,30,69,31,63,31,182,31,182,30,228,31,38,31,38,30,124,31,124,30,161,31,194,31,25,31,8,31,195,31,104,31,25,31,25,30,203,31,208,31,179,31,210,31,22,31,22,30,22,29,244,31,23,31,40,31,92,31,58,31,204,31,111,31,160,31,196,31,196,30,196,29,82,31,145,31,145,30,170,31,7,31,231,31,85,31,85,30,85,29,85,28,13,31,215,31,122,31,61,31,190,31,133,31,20,31,245,31,121,31,166,31,242,31,142,31,232,31,232,30,36,31,36,30,4,31,226,31,226,30,226,29,226,28,145,31,145,30,154,31,12,31,95,31,214,31,128,31,128,30,144,31,68,31,251,31,135,31,135,30,135,29,30,31,30,30,21,31,242,31,255,31,255,30,152,31,136,31,66,31,66,30,66,29,236,31,25,31,50,31,39,31,66,31,67,31,214,31,214,30,160,31,176,31,41,31,26,31,116,31,116,30,169,31,235,31,204,31,158,31,255,31,255,30,255,29,66,31,66,30,207,31,207,30,76,31,75,31,127,31,79,31,113,31,7,31,208,31,69,31,147,31,113,31,123,31,29,31,168,31,224,31,195,31,195,30,179,31,179,30,181,31,218,31,181,31,85,31,140,31,70,31,244,31,5,31,245,31,222,31,1,31,99,31,247,31,245,31,166,31,10,31,139,31,139,30,139,29,42,31,249,31,210,31,145,31,142,31,243,31,228,31,228,30,49,31,49,30,53,31,99,31,89,31,146,31,199,31,242,31,242,30,178,31,187,31,187,30,187,29,187,28,63,31,154,31,31,31,207,31,168,31,35,31,202,31,90,31,90,30,157,31,14,31,140,31,83,31,176,31,193,31,203,31,33,31,243,31,71,31,5,31,2,31,79,31,79,30,113,31,137,31,43,31,198,31,209,31,209,30,229,31,6,31,58,31,98,31,89,31,203,31,113,31,37,31,37,30,69,31,155,31,20,31,43,31,124,31,124,30,205,31,253,31,209,31,184,31,79,31,124,31,143,31,85,31,85,30,99,31,57,31,56,31,183,31,200,31,200,30,184,31,142,31,122,31,243,31,124,31,250,31,138,31,138,30,138,29,9,31,9,30,9,29,9,28,49,31,176,31,176,30,176,29,205,31,98,31,124,31,213,31,213,30,38,31,104,31,194,31,194,30,126,31,194,31,220,31,139,31,172,31,3,31,245,31,169,31,20,31,155,31,32,31,32,30,172,31,172,30,105,31,128,31,55,31,123,31,109,31,109,30,244,31,202,31,25,31,150,31,53,31,99,31,46,31,180,31,146,31,146,30,25,31,109,31,37,31,85,31,123,31,123,30,41,31,230,31,164,31,102,31,105,31,216,31,161,31,234,31,77,31,229,31,123,31,123,30,127,31,228,31,228,30,208,31,146,31,11,31,167,31,167,30,167,29,39,31,153,31,179,31,231,31,52,31,1,31,219,31,170,31,170,30,35,31,149,31,13,31,196,31,110,31,36,31,221,31,66,31,187,31,40,31,192,31,88,31,9,31,9,30,116,31,116,30,116,29,34,31,120,31,239,31,20,31,20,30,108,31,52,31,52,30,131,31,200,31,123,31,96,31,195,31,106,31,24,31,24,30,181,31,181,30,79,31,142,31,196,31,196,30,89,31,89,30,170,31,181,31,118,31,221,31,221,30,107,31,222,31,97,31,150,31,198,31,253,31,179,31,234,31,113,31,4,31,250,31,218,31,255,31,166,31,192,31,25,31,101,31,149,31,170,31,133,31,202,31,64,31,216,31,216,30,192,31,118,31,118,30,153,31,110,31,2,31,2,30,134,31,5,31,140,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
