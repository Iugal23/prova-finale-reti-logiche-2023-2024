-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_39 is
end project_tb_39;

architecture project_tb_arch_39 of project_tb_39 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 754;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (94,0,63,0,124,0,0,0,92,0,46,0,0,0,33,0,72,0,31,0,138,0,153,0,237,0,215,0,152,0,153,0,6,0,122,0,13,0,28,0,24,0,135,0,32,0,195,0,0,0,178,0,155,0,251,0,197,0,221,0,17,0,48,0,0,0,189,0,248,0,115,0,193,0,151,0,215,0,26,0,32,0,227,0,143,0,216,0,131,0,125,0,229,0,172,0,23,0,0,0,19,0,13,0,249,0,90,0,215,0,108,0,195,0,125,0,40,0,191,0,180,0,237,0,0,0,180,0,239,0,33,0,177,0,105,0,208,0,206,0,0,0,196,0,0,0,226,0,96,0,17,0,82,0,35,0,151,0,6,0,255,0,125,0,13,0,14,0,89,0,37,0,247,0,0,0,0,0,0,0,215,0,133,0,149,0,0,0,0,0,194,0,96,0,89,0,209,0,127,0,238,0,45,0,211,0,97,0,0,0,87,0,237,0,159,0,7,0,0,0,73,0,193,0,222,0,20,0,41,0,28,0,7,0,189,0,50,0,96,0,199,0,95,0,98,0,196,0,0,0,162,0,4,0,0,0,28,0,139,0,104,0,195,0,0,0,48,0,175,0,8,0,0,0,0,0,211,0,0,0,61,0,191,0,26,0,0,0,2,0,228,0,110,0,62,0,0,0,110,0,225,0,52,0,22,0,44,0,174,0,103,0,92,0,100,0,164,0,87,0,213,0,187,0,143,0,167,0,170,0,159,0,131,0,242,0,0,0,225,0,229,0,245,0,55,0,126,0,227,0,55,0,0,0,166,0,0,0,0,0,37,0,198,0,36,0,65,0,185,0,184,0,69,0,37,0,236,0,7,0,0,0,86,0,31,0,170,0,0,0,16,0,246,0,34,0,124,0,112,0,45,0,85,0,87,0,143,0,102,0,99,0,174,0,0,0,150,0,254,0,0,0,0,0,225,0,28,0,0,0,51,0,0,0,134,0,0,0,0,0,100,0,248,0,252,0,201,0,171,0,136,0,0,0,177,0,0,0,55,0,51,0,25,0,248,0,121,0,75,0,62,0,38,0,133,0,234,0,0,0,221,0,101,0,0,0,23,0,198,0,182,0,153,0,0,0,164,0,51,0,95,0,246,0,0,0,0,0,132,0,0,0,163,0,193,0,50,0,194,0,65,0,72,0,122,0,227,0,25,0,141,0,0,0,131,0,221,0,170,0,0,0,194,0,141,0,188,0,0,0,132,0,177,0,110,0,245,0,188,0,132,0,9,0,73,0,80,0,83,0,64,0,144,0,65,0,0,0,116,0,149,0,54,0,206,0,26,0,0,0,0,0,155,0,189,0,212,0,64,0,11,0,181,0,16,0,0,0,0,0,144,0,0,0,92,0,133,0,24,0,154,0,163,0,254,0,48,0,12,0,56,0,4,0,158,0,103,0,180,0,0,0,163,0,0,0,105,0,121,0,248,0,155,0,131,0,167,0,0,0,161,0,38,0,207,0,224,0,0,0,0,0,62,0,0,0,36,0,0,0,252,0,0,0,234,0,123,0,222,0,12,0,125,0,189,0,238,0,139,0,245,0,0,0,169,0,44,0,245,0,210,0,0,0,0,0,0,0,89,0,84,0,177,0,7,0,159,0,0,0,183,0,203,0,18,0,28,0,64,0,88,0,71,0,15,0,249,0,193,0,122,0,0,0,142,0,114,0,122,0,94,0,247,0,219,0,176,0,111,0,157,0,202,0,0,0,36,0,212,0,190,0,165,0,2,0,177,0,0,0,191,0,63,0,18,0,104,0,0,0,176,0,84,0,110,0,140,0,193,0,161,0,50,0,176,0,0,0,151,0,174,0,25,0,0,0,0,0,114,0,168,0,118,0,218,0,77,0,75,0,64,0,85,0,103,0,96,0,12,0,232,0,0,0,0,0,19,0,18,0,143,0,219,0,48,0,0,0,50,0,0,0,20,0,254,0,77,0,87,0,19,0,151,0,185,0,247,0,0,0,42,0,197,0,0,0,44,0,230,0,50,0,247,0,93,0,22,0,247,0,229,0,0,0,0,0,148,0,44,0,51,0,0,0,46,0,79,0,0,0,0,0,177,0,0,0,221,0,41,0,0,0,0,0,115,0,2,0,0,0,22,0,0,0,0,0,65,0,9,0,191,0,117,0,81,0,156,0,242,0,0,0,0,0,0,0,112,0,31,0,0,0,161,0,6,0,38,0,160,0,165,0,127,0,164,0,240,0,214,0,162,0,66,0,106,0,43,0,121,0,19,0,77,0,182,0,67,0,127,0,0,0,167,0,237,0,154,0,180,0,94,0,57,0,0,0,137,0,32,0,97,0,0,0,195,0,66,0,66,0,76,0,127,0,233,0,0,0,205,0,0,0,175,0,232,0,153,0,165,0,0,0,216,0,110,0,254,0,130,0,102,0,0,0,67,0,0,0,104,0,86,0,61,0,87,0,0,0,19,0,143,0,118,0,158,0,159,0,0,0,220,0,61,0,121,0,120,0,25,0,157,0,147,0,80,0,13,0,0,0,102,0,129,0,112,0,87,0,130,0,43,0,108,0,137,0,41,0,88,0,113,0,73,0,0,0,110,0,27,0,45,0,0,0,0,0,0,0,3,0,115,0,0,0,146,0,129,0,153,0,152,0,0,0,228,0,244,0,0,0,132,0,0,0,225,0,0,0,71,0,21,0,32,0,30,0,149,0,109,0,6,0,59,0,13,0,77,0,249,0,48,0,49,0,0,0,85,0,0,0,116,0,231,0,144,0,248,0,56,0,171,0,9,0,104,0,238,0,22,0,83,0,200,0,250,0,44,0,200,0,0,0,71,0,183,0,57,0,180,0,58,0,238,0,0,0,102,0,0,0,16,0,139,0,46,0,158,0,107,0,214,0,84,0,151,0,238,0,149,0,22,0,228,0,0,0,127,0,0,0,144,0,231,0,73,0,0,0,165,0,53,0,89,0,55,0,116,0,60,0,75,0,179,0,248,0,0,0,93,0,104,0,144,0,114,0,45,0,145,0,206,0,0,0,0,0,0,0,229,0,33,0,250,0,237,0,32,0,170,0,168,0,233,0,203,0,139,0,148,0,14,0,2,0,0,0,132,0,198,0,187,0,14,0,164,0,0,0,67,0,241,0,167,0,0,0,132,0,88,0,0,0,33,0,180,0,118,0,52,0,242,0,121,0,82,0,195,0,231,0,150,0,215,0,94,0,117,0,0,0,8,0,252,0,0,0,201,0,207,0,201,0,0,0,224,0,0,0,238,0,18,0,63,0,188,0,71,0,0,0,206,0,58,0,0,0,24,0,141,0,39,0,16,0,0,0,78,0,219,0,33,0,101,0,191,0,23,0,81,0,12,0,134,0,211,0,66,0);
signal scenario_full  : scenario_type := (94,31,63,31,124,31,124,30,92,31,46,31,46,30,33,31,72,31,31,31,138,31,153,31,237,31,215,31,152,31,153,31,6,31,122,31,13,31,28,31,24,31,135,31,32,31,195,31,195,30,178,31,155,31,251,31,197,31,221,31,17,31,48,31,48,30,189,31,248,31,115,31,193,31,151,31,215,31,26,31,32,31,227,31,143,31,216,31,131,31,125,31,229,31,172,31,23,31,23,30,19,31,13,31,249,31,90,31,215,31,108,31,195,31,125,31,40,31,191,31,180,31,237,31,237,30,180,31,239,31,33,31,177,31,105,31,208,31,206,31,206,30,196,31,196,30,226,31,96,31,17,31,82,31,35,31,151,31,6,31,255,31,125,31,13,31,14,31,89,31,37,31,247,31,247,30,247,29,247,28,215,31,133,31,149,31,149,30,149,29,194,31,96,31,89,31,209,31,127,31,238,31,45,31,211,31,97,31,97,30,87,31,237,31,159,31,7,31,7,30,73,31,193,31,222,31,20,31,41,31,28,31,7,31,189,31,50,31,96,31,199,31,95,31,98,31,196,31,196,30,162,31,4,31,4,30,28,31,139,31,104,31,195,31,195,30,48,31,175,31,8,31,8,30,8,29,211,31,211,30,61,31,191,31,26,31,26,30,2,31,228,31,110,31,62,31,62,30,110,31,225,31,52,31,22,31,44,31,174,31,103,31,92,31,100,31,164,31,87,31,213,31,187,31,143,31,167,31,170,31,159,31,131,31,242,31,242,30,225,31,229,31,245,31,55,31,126,31,227,31,55,31,55,30,166,31,166,30,166,29,37,31,198,31,36,31,65,31,185,31,184,31,69,31,37,31,236,31,7,31,7,30,86,31,31,31,170,31,170,30,16,31,246,31,34,31,124,31,112,31,45,31,85,31,87,31,143,31,102,31,99,31,174,31,174,30,150,31,254,31,254,30,254,29,225,31,28,31,28,30,51,31,51,30,134,31,134,30,134,29,100,31,248,31,252,31,201,31,171,31,136,31,136,30,177,31,177,30,55,31,51,31,25,31,248,31,121,31,75,31,62,31,38,31,133,31,234,31,234,30,221,31,101,31,101,30,23,31,198,31,182,31,153,31,153,30,164,31,51,31,95,31,246,31,246,30,246,29,132,31,132,30,163,31,193,31,50,31,194,31,65,31,72,31,122,31,227,31,25,31,141,31,141,30,131,31,221,31,170,31,170,30,194,31,141,31,188,31,188,30,132,31,177,31,110,31,245,31,188,31,132,31,9,31,73,31,80,31,83,31,64,31,144,31,65,31,65,30,116,31,149,31,54,31,206,31,26,31,26,30,26,29,155,31,189,31,212,31,64,31,11,31,181,31,16,31,16,30,16,29,144,31,144,30,92,31,133,31,24,31,154,31,163,31,254,31,48,31,12,31,56,31,4,31,158,31,103,31,180,31,180,30,163,31,163,30,105,31,121,31,248,31,155,31,131,31,167,31,167,30,161,31,38,31,207,31,224,31,224,30,224,29,62,31,62,30,36,31,36,30,252,31,252,30,234,31,123,31,222,31,12,31,125,31,189,31,238,31,139,31,245,31,245,30,169,31,44,31,245,31,210,31,210,30,210,29,210,28,89,31,84,31,177,31,7,31,159,31,159,30,183,31,203,31,18,31,28,31,64,31,88,31,71,31,15,31,249,31,193,31,122,31,122,30,142,31,114,31,122,31,94,31,247,31,219,31,176,31,111,31,157,31,202,31,202,30,36,31,212,31,190,31,165,31,2,31,177,31,177,30,191,31,63,31,18,31,104,31,104,30,176,31,84,31,110,31,140,31,193,31,161,31,50,31,176,31,176,30,151,31,174,31,25,31,25,30,25,29,114,31,168,31,118,31,218,31,77,31,75,31,64,31,85,31,103,31,96,31,12,31,232,31,232,30,232,29,19,31,18,31,143,31,219,31,48,31,48,30,50,31,50,30,20,31,254,31,77,31,87,31,19,31,151,31,185,31,247,31,247,30,42,31,197,31,197,30,44,31,230,31,50,31,247,31,93,31,22,31,247,31,229,31,229,30,229,29,148,31,44,31,51,31,51,30,46,31,79,31,79,30,79,29,177,31,177,30,221,31,41,31,41,30,41,29,115,31,2,31,2,30,22,31,22,30,22,29,65,31,9,31,191,31,117,31,81,31,156,31,242,31,242,30,242,29,242,28,112,31,31,31,31,30,161,31,6,31,38,31,160,31,165,31,127,31,164,31,240,31,214,31,162,31,66,31,106,31,43,31,121,31,19,31,77,31,182,31,67,31,127,31,127,30,167,31,237,31,154,31,180,31,94,31,57,31,57,30,137,31,32,31,97,31,97,30,195,31,66,31,66,31,76,31,127,31,233,31,233,30,205,31,205,30,175,31,232,31,153,31,165,31,165,30,216,31,110,31,254,31,130,31,102,31,102,30,67,31,67,30,104,31,86,31,61,31,87,31,87,30,19,31,143,31,118,31,158,31,159,31,159,30,220,31,61,31,121,31,120,31,25,31,157,31,147,31,80,31,13,31,13,30,102,31,129,31,112,31,87,31,130,31,43,31,108,31,137,31,41,31,88,31,113,31,73,31,73,30,110,31,27,31,45,31,45,30,45,29,45,28,3,31,115,31,115,30,146,31,129,31,153,31,152,31,152,30,228,31,244,31,244,30,132,31,132,30,225,31,225,30,71,31,21,31,32,31,30,31,149,31,109,31,6,31,59,31,13,31,77,31,249,31,48,31,49,31,49,30,85,31,85,30,116,31,231,31,144,31,248,31,56,31,171,31,9,31,104,31,238,31,22,31,83,31,200,31,250,31,44,31,200,31,200,30,71,31,183,31,57,31,180,31,58,31,238,31,238,30,102,31,102,30,16,31,139,31,46,31,158,31,107,31,214,31,84,31,151,31,238,31,149,31,22,31,228,31,228,30,127,31,127,30,144,31,231,31,73,31,73,30,165,31,53,31,89,31,55,31,116,31,60,31,75,31,179,31,248,31,248,30,93,31,104,31,144,31,114,31,45,31,145,31,206,31,206,30,206,29,206,28,229,31,33,31,250,31,237,31,32,31,170,31,168,31,233,31,203,31,139,31,148,31,14,31,2,31,2,30,132,31,198,31,187,31,14,31,164,31,164,30,67,31,241,31,167,31,167,30,132,31,88,31,88,30,33,31,180,31,118,31,52,31,242,31,121,31,82,31,195,31,231,31,150,31,215,31,94,31,117,31,117,30,8,31,252,31,252,30,201,31,207,31,201,31,201,30,224,31,224,30,238,31,18,31,63,31,188,31,71,31,71,30,206,31,58,31,58,30,24,31,141,31,39,31,16,31,16,30,78,31,219,31,33,31,101,31,191,31,23,31,81,31,12,31,134,31,211,31,66,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
