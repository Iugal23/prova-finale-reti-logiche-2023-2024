-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_970 is
end project_tb_970;

architecture project_tb_arch_970 of project_tb_970 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 901;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (103,0,0,0,198,0,209,0,3,0,85,0,145,0,204,0,60,0,115,0,113,0,26,0,130,0,105,0,59,0,193,0,215,0,162,0,0,0,0,0,176,0,34,0,84,0,233,0,0,0,83,0,149,0,45,0,104,0,88,0,0,0,149,0,0,0,38,0,5,0,21,0,0,0,34,0,182,0,95,0,180,0,116,0,0,0,221,0,209,0,0,0,115,0,28,0,102,0,69,0,79,0,0,0,90,0,0,0,175,0,28,0,124,0,0,0,6,0,245,0,2,0,14,0,48,0,184,0,0,0,160,0,228,0,69,0,7,0,78,0,231,0,77,0,76,0,0,0,76,0,143,0,147,0,79,0,0,0,0,0,9,0,108,0,155,0,85,0,41,0,87,0,0,0,8,0,229,0,0,0,51,0,0,0,151,0,151,0,0,0,1,0,0,0,157,0,165,0,0,0,0,0,0,0,0,0,32,0,0,0,0,0,146,0,141,0,108,0,17,0,220,0,218,0,216,0,71,0,199,0,0,0,197,0,125,0,0,0,36,0,64,0,188,0,95,0,154,0,194,0,226,0,238,0,233,0,254,0,169,0,0,0,242,0,201,0,238,0,87,0,188,0,142,0,19,0,107,0,99,0,75,0,44,0,40,0,85,0,220,0,141,0,108,0,246,0,110,0,95,0,0,0,194,0,246,0,29,0,183,0,49,0,152,0,0,0,0,0,227,0,0,0,8,0,67,0,0,0,208,0,0,0,0,0,10,0,27,0,147,0,0,0,142,0,238,0,114,0,248,0,232,0,161,0,108,0,68,0,202,0,0,0,0,0,161,0,48,0,0,0,0,0,181,0,145,0,101,0,82,0,139,0,56,0,0,0,0,0,133,0,230,0,23,0,0,0,0,0,0,0,12,0,190,0,221,0,118,0,255,0,190,0,84,0,101,0,215,0,0,0,110,0,33,0,213,0,149,0,0,0,198,0,8,0,0,0,239,0,89,0,115,0,219,0,229,0,117,0,10,0,180,0,191,0,116,0,86,0,203,0,250,0,196,0,214,0,237,0,36,0,0,0,253,0,98,0,80,0,96,0,175,0,247,0,0,0,0,0,149,0,99,0,22,0,233,0,71,0,86,0,0,0,85,0,92,0,0,0,223,0,95,0,0,0,71,0,0,0,254,0,143,0,103,0,0,0,149,0,74,0,191,0,178,0,63,0,23,0,9,0,71,0,187,0,201,0,65,0,149,0,0,0,5,0,223,0,0,0,195,0,1,0,0,0,77,0,252,0,130,0,8,0,154,0,224,0,129,0,95,0,125,0,14,0,109,0,59,0,248,0,0,0,83,0,46,0,0,0,21,0,35,0,0,0,160,0,147,0,0,0,134,0,34,0,0,0,142,0,157,0,135,0,72,0,0,0,157,0,209,0,71,0,70,0,42,0,118,0,47,0,0,0,37,0,56,0,47,0,0,0,118,0,158,0,158,0,29,0,20,0,187,0,118,0,71,0,159,0,228,0,109,0,0,0,55,0,166,0,143,0,4,0,211,0,0,0,134,0,13,0,0,0,214,0,127,0,69,0,139,0,0,0,180,0,138,0,150,0,0,0,61,0,206,0,39,0,184,0,221,0,51,0,127,0,193,0,30,0,32,0,0,0,240,0,71,0,0,0,233,0,52,0,179,0,100,0,83,0,166,0,42,0,0,0,0,0,37,0,0,0,52,0,0,0,162,0,42,0,217,0,0,0,211,0,18,0,173,0,0,0,200,0,54,0,48,0,78,0,145,0,0,0,0,0,220,0,180,0,246,0,16,0,235,0,144,0,75,0,0,0,0,0,243,0,0,0,228,0,113,0,55,0,74,0,65,0,73,0,242,0,189,0,251,0,77,0,64,0,131,0,0,0,99,0,149,0,240,0,179,0,207,0,114,0,69,0,250,0,82,0,223,0,34,0,0,0,231,0,139,0,99,0,67,0,0,0,199,0,0,0,108,0,22,0,239,0,81,0,159,0,0,0,214,0,0,0,202,0,0,0,162,0,176,0,5,0,0,0,192,0,140,0,0,0,60,0,78,0,178,0,12,0,255,0,0,0,0,0,133,0,0,0,152,0,229,0,50,0,147,0,211,0,0,0,244,0,91,0,234,0,0,0,150,0,0,0,51,0,43,0,34,0,124,0,0,0,0,0,115,0,0,0,0,0,146,0,168,0,195,0,66,0,74,0,5,0,0,0,67,0,204,0,113,0,43,0,0,0,214,0,18,0,0,0,0,0,200,0,83,0,135,0,17,0,9,0,115,0,122,0,133,0,80,0,19,0,78,0,190,0,168,0,163,0,60,0,155,0,87,0,127,0,123,0,189,0,132,0,35,0,35,0,184,0,207,0,235,0,39,0,155,0,215,0,115,0,98,0,191,0,0,0,243,0,224,0,0,0,221,0,162,0,38,0,196,0,197,0,251,0,242,0,0,0,112,0,7,0,61,0,108,0,68,0,110,0,31,0,0,0,0,0,0,0,88,0,0,0,66,0,186,0,69,0,155,0,0,0,18,0,136,0,66,0,160,0,0,0,148,0,122,0,173,0,158,0,212,0,31,0,156,0,41,0,144,0,0,0,0,0,202,0,58,0,56,0,0,0,0,0,63,0,188,0,162,0,0,0,0,0,198,0,68,0,0,0,194,0,35,0,0,0,250,0,247,0,201,0,151,0,0,0,21,0,0,0,103,0,0,0,108,0,77,0,251,0,66,0,10,0,105,0,0,0,0,0,248,0,98,0,0,0,209,0,54,0,42,0,143,0,62,0,109,0,87,0,0,0,0,0,174,0,36,0,61,0,43,0,211,0,87,0,0,0,216,0,7,0,55,0,105,0,0,0,234,0,0,0,0,0,200,0,237,0,232,0,154,0,192,0,65,0,72,0,222,0,254,0,0,0,0,0,39,0,89,0,130,0,0,0,131,0,189,0,137,0,47,0,126,0,138,0,58,0,92,0,170,0,0,0,0,0,55,0,126,0,176,0,150,0,105,0,236,0,0,0,0,0,253,0,162,0,0,0,193,0,109,0,0,0,125,0,123,0,170,0,0,0,92,0,24,0,249,0,0,0,0,0,75,0,135,0,142,0,0,0,79,0,0,0,127,0,205,0,112,0,9,0,26,0,96,0,118,0,140,0,0,0,0,0,185,0,24,0,12,0,214,0,0,0,0,0,0,0,94,0,0,0,204,0,0,0,36,0,54,0,76,0,122,0,30,0,193,0,87,0,0,0,226,0,218,0,45,0,201,0,194,0,187,0,123,0,238,0,0,0,221,0,168,0,130,0,74,0,98,0,37,0,165,0,209,0,0,0,54,0,0,0,81,0,213,0,29,0,220,0,117,0,8,0,0,0,240,0,35,0,0,0,171,0,0,0,53,0,137,0,0,0,146,0,25,0,1,0,241,0,27,0,13,0,111,0,167,0,0,0,192,0,12,0,74,0,37,0,0,0,102,0,85,0,72,0,46,0,23,0,0,0,128,0,43,0,112,0,219,0,130,0,106,0,0,0,0,0,176,0,217,0,40,0,23,0,85,0,31,0,6,0,126,0,206,0,0,0,194,0,61,0,191,0,0,0,0,0,89,0,0,0,225,0,79,0,157,0,62,0,12,0,96,0,0,0,87,0,67,0,2,0,156,0,29,0,24,0,30,0,159,0,228,0,193,0,80,0,142,0,225,0,0,0,168,0,181,0,125,0,220,0,171,0,172,0,130,0,29,0,237,0,62,0,67,0,73,0,0,0,113,0,91,0,0,0,116,0,81,0,241,0,180,0,99,0,59,0,102,0,62,0,39,0,66,0,219,0,247,0,200,0,216,0,143,0,110,0,174,0,103,0,201,0,173,0,6,0,18,0,0,0,221,0,2,0,95,0,124,0,158,0,0,0,154,0,255,0,125,0,42,0,0,0,172,0,204,0,0,0,0,0,165,0,28,0,217,0,0,0,0,0,0,0,213,0,78,0,32,0,224,0,0,0,96,0,14,0,128,0,140,0,69,0,127,0,0,0,173,0,5,0,125,0,139,0);
signal scenario_full  : scenario_type := (103,31,103,30,198,31,209,31,3,31,85,31,145,31,204,31,60,31,115,31,113,31,26,31,130,31,105,31,59,31,193,31,215,31,162,31,162,30,162,29,176,31,34,31,84,31,233,31,233,30,83,31,149,31,45,31,104,31,88,31,88,30,149,31,149,30,38,31,5,31,21,31,21,30,34,31,182,31,95,31,180,31,116,31,116,30,221,31,209,31,209,30,115,31,28,31,102,31,69,31,79,31,79,30,90,31,90,30,175,31,28,31,124,31,124,30,6,31,245,31,2,31,14,31,48,31,184,31,184,30,160,31,228,31,69,31,7,31,78,31,231,31,77,31,76,31,76,30,76,31,143,31,147,31,79,31,79,30,79,29,9,31,108,31,155,31,85,31,41,31,87,31,87,30,8,31,229,31,229,30,51,31,51,30,151,31,151,31,151,30,1,31,1,30,157,31,165,31,165,30,165,29,165,28,165,27,32,31,32,30,32,29,146,31,141,31,108,31,17,31,220,31,218,31,216,31,71,31,199,31,199,30,197,31,125,31,125,30,36,31,64,31,188,31,95,31,154,31,194,31,226,31,238,31,233,31,254,31,169,31,169,30,242,31,201,31,238,31,87,31,188,31,142,31,19,31,107,31,99,31,75,31,44,31,40,31,85,31,220,31,141,31,108,31,246,31,110,31,95,31,95,30,194,31,246,31,29,31,183,31,49,31,152,31,152,30,152,29,227,31,227,30,8,31,67,31,67,30,208,31,208,30,208,29,10,31,27,31,147,31,147,30,142,31,238,31,114,31,248,31,232,31,161,31,108,31,68,31,202,31,202,30,202,29,161,31,48,31,48,30,48,29,181,31,145,31,101,31,82,31,139,31,56,31,56,30,56,29,133,31,230,31,23,31,23,30,23,29,23,28,12,31,190,31,221,31,118,31,255,31,190,31,84,31,101,31,215,31,215,30,110,31,33,31,213,31,149,31,149,30,198,31,8,31,8,30,239,31,89,31,115,31,219,31,229,31,117,31,10,31,180,31,191,31,116,31,86,31,203,31,250,31,196,31,214,31,237,31,36,31,36,30,253,31,98,31,80,31,96,31,175,31,247,31,247,30,247,29,149,31,99,31,22,31,233,31,71,31,86,31,86,30,85,31,92,31,92,30,223,31,95,31,95,30,71,31,71,30,254,31,143,31,103,31,103,30,149,31,74,31,191,31,178,31,63,31,23,31,9,31,71,31,187,31,201,31,65,31,149,31,149,30,5,31,223,31,223,30,195,31,1,31,1,30,77,31,252,31,130,31,8,31,154,31,224,31,129,31,95,31,125,31,14,31,109,31,59,31,248,31,248,30,83,31,46,31,46,30,21,31,35,31,35,30,160,31,147,31,147,30,134,31,34,31,34,30,142,31,157,31,135,31,72,31,72,30,157,31,209,31,71,31,70,31,42,31,118,31,47,31,47,30,37,31,56,31,47,31,47,30,118,31,158,31,158,31,29,31,20,31,187,31,118,31,71,31,159,31,228,31,109,31,109,30,55,31,166,31,143,31,4,31,211,31,211,30,134,31,13,31,13,30,214,31,127,31,69,31,139,31,139,30,180,31,138,31,150,31,150,30,61,31,206,31,39,31,184,31,221,31,51,31,127,31,193,31,30,31,32,31,32,30,240,31,71,31,71,30,233,31,52,31,179,31,100,31,83,31,166,31,42,31,42,30,42,29,37,31,37,30,52,31,52,30,162,31,42,31,217,31,217,30,211,31,18,31,173,31,173,30,200,31,54,31,48,31,78,31,145,31,145,30,145,29,220,31,180,31,246,31,16,31,235,31,144,31,75,31,75,30,75,29,243,31,243,30,228,31,113,31,55,31,74,31,65,31,73,31,242,31,189,31,251,31,77,31,64,31,131,31,131,30,99,31,149,31,240,31,179,31,207,31,114,31,69,31,250,31,82,31,223,31,34,31,34,30,231,31,139,31,99,31,67,31,67,30,199,31,199,30,108,31,22,31,239,31,81,31,159,31,159,30,214,31,214,30,202,31,202,30,162,31,176,31,5,31,5,30,192,31,140,31,140,30,60,31,78,31,178,31,12,31,255,31,255,30,255,29,133,31,133,30,152,31,229,31,50,31,147,31,211,31,211,30,244,31,91,31,234,31,234,30,150,31,150,30,51,31,43,31,34,31,124,31,124,30,124,29,115,31,115,30,115,29,146,31,168,31,195,31,66,31,74,31,5,31,5,30,67,31,204,31,113,31,43,31,43,30,214,31,18,31,18,30,18,29,200,31,83,31,135,31,17,31,9,31,115,31,122,31,133,31,80,31,19,31,78,31,190,31,168,31,163,31,60,31,155,31,87,31,127,31,123,31,189,31,132,31,35,31,35,31,184,31,207,31,235,31,39,31,155,31,215,31,115,31,98,31,191,31,191,30,243,31,224,31,224,30,221,31,162,31,38,31,196,31,197,31,251,31,242,31,242,30,112,31,7,31,61,31,108,31,68,31,110,31,31,31,31,30,31,29,31,28,88,31,88,30,66,31,186,31,69,31,155,31,155,30,18,31,136,31,66,31,160,31,160,30,148,31,122,31,173,31,158,31,212,31,31,31,156,31,41,31,144,31,144,30,144,29,202,31,58,31,56,31,56,30,56,29,63,31,188,31,162,31,162,30,162,29,198,31,68,31,68,30,194,31,35,31,35,30,250,31,247,31,201,31,151,31,151,30,21,31,21,30,103,31,103,30,108,31,77,31,251,31,66,31,10,31,105,31,105,30,105,29,248,31,98,31,98,30,209,31,54,31,42,31,143,31,62,31,109,31,87,31,87,30,87,29,174,31,36,31,61,31,43,31,211,31,87,31,87,30,216,31,7,31,55,31,105,31,105,30,234,31,234,30,234,29,200,31,237,31,232,31,154,31,192,31,65,31,72,31,222,31,254,31,254,30,254,29,39,31,89,31,130,31,130,30,131,31,189,31,137,31,47,31,126,31,138,31,58,31,92,31,170,31,170,30,170,29,55,31,126,31,176,31,150,31,105,31,236,31,236,30,236,29,253,31,162,31,162,30,193,31,109,31,109,30,125,31,123,31,170,31,170,30,92,31,24,31,249,31,249,30,249,29,75,31,135,31,142,31,142,30,79,31,79,30,127,31,205,31,112,31,9,31,26,31,96,31,118,31,140,31,140,30,140,29,185,31,24,31,12,31,214,31,214,30,214,29,214,28,94,31,94,30,204,31,204,30,36,31,54,31,76,31,122,31,30,31,193,31,87,31,87,30,226,31,218,31,45,31,201,31,194,31,187,31,123,31,238,31,238,30,221,31,168,31,130,31,74,31,98,31,37,31,165,31,209,31,209,30,54,31,54,30,81,31,213,31,29,31,220,31,117,31,8,31,8,30,240,31,35,31,35,30,171,31,171,30,53,31,137,31,137,30,146,31,25,31,1,31,241,31,27,31,13,31,111,31,167,31,167,30,192,31,12,31,74,31,37,31,37,30,102,31,85,31,72,31,46,31,23,31,23,30,128,31,43,31,112,31,219,31,130,31,106,31,106,30,106,29,176,31,217,31,40,31,23,31,85,31,31,31,6,31,126,31,206,31,206,30,194,31,61,31,191,31,191,30,191,29,89,31,89,30,225,31,79,31,157,31,62,31,12,31,96,31,96,30,87,31,67,31,2,31,156,31,29,31,24,31,30,31,159,31,228,31,193,31,80,31,142,31,225,31,225,30,168,31,181,31,125,31,220,31,171,31,172,31,130,31,29,31,237,31,62,31,67,31,73,31,73,30,113,31,91,31,91,30,116,31,81,31,241,31,180,31,99,31,59,31,102,31,62,31,39,31,66,31,219,31,247,31,200,31,216,31,143,31,110,31,174,31,103,31,201,31,173,31,6,31,18,31,18,30,221,31,2,31,95,31,124,31,158,31,158,30,154,31,255,31,125,31,42,31,42,30,172,31,204,31,204,30,204,29,165,31,28,31,217,31,217,30,217,29,217,28,213,31,78,31,32,31,224,31,224,30,96,31,14,31,128,31,140,31,69,31,127,31,127,30,173,31,5,31,125,31,139,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
