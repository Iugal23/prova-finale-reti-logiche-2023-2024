-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 823;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,0,0,0,0,16,0,10,0,210,0,133,0,29,0,145,0,236,0,226,0,8,0,252,0,3,0,128,0,246,0,3,0,0,0,45,0,196,0,14,0,144,0,52,0,228,0,153,0,125,0,86,0,151,0,0,0,3,0,0,0,224,0,187,0,71,0,230,0,190,0,0,0,0,0,166,0,226,0,0,0,0,0,0,0,142,0,227,0,0,0,113,0,185,0,0,0,0,0,59,0,169,0,19,0,0,0,201,0,225,0,160,0,180,0,0,0,25,0,89,0,165,0,208,0,82,0,114,0,36,0,245,0,52,0,161,0,116,0,141,0,196,0,0,0,5,0,0,0,221,0,0,0,209,0,81,0,0,0,0,0,23,0,37,0,4,0,39,0,226,0,106,0,0,0,231,0,106,0,22,0,209,0,251,0,0,0,15,0,0,0,30,0,5,0,0,0,74,0,0,0,15,0,202,0,162,0,0,0,81,0,232,0,87,0,0,0,7,0,165,0,247,0,209,0,238,0,81,0,0,0,27,0,201,0,48,0,5,0,132,0,6,0,38,0,154,0,119,0,211,0,22,0,145,0,179,0,204,0,0,0,0,0,0,0,30,0,30,0,0,0,144,0,0,0,117,0,0,0,0,0,92,0,81,0,0,0,181,0,0,0,79,0,13,0,20,0,187,0,7,0,219,0,221,0,71,0,236,0,0,0,208,0,62,0,226,0,57,0,0,0,20,0,0,0,218,0,84,0,0,0,0,0,176,0,170,0,254,0,212,0,192,0,132,0,251,0,125,0,159,0,104,0,17,0,194,0,70,0,210,0,244,0,153,0,34,0,206,0,4,0,241,0,12,0,167,0,226,0,228,0,245,0,90,0,167,0,200,0,0,0,10,0,203,0,195,0,36,0,0,0,223,0,218,0,62,0,177,0,222,0,187,0,223,0,0,0,231,0,164,0,83,0,0,0,248,0,180,0,11,0,0,0,70,0,190,0,214,0,40,0,0,0,0,0,190,0,166,0,95,0,99,0,142,0,117,0,0,0,0,0,142,0,123,0,0,0,0,0,0,0,194,0,71,0,86,0,131,0,0,0,0,0,98,0,90,0,14,0,95,0,218,0,5,0,6,0,249,0,0,0,157,0,61,0,162,0,56,0,0,0,30,0,0,0,223,0,230,0,41,0,103,0,83,0,61,0,109,0,131,0,106,0,0,0,96,0,19,0,139,0,113,0,142,0,26,0,218,0,226,0,201,0,110,0,96,0,142,0,188,0,0,0,4,0,0,0,252,0,58,0,0,0,0,0,73,0,184,0,111,0,0,0,116,0,166,0,0,0,0,0,0,0,75,0,248,0,195,0,131,0,166,0,155,0,129,0,0,0,202,0,155,0,2,0,72,0,0,0,165,0,4,0,240,0,0,0,0,0,0,0,253,0,1,0,0,0,248,0,121,0,250,0,70,0,50,0,217,0,196,0,0,0,204,0,0,0,0,0,122,0,126,0,83,0,115,0,47,0,110,0,10,0,31,0,19,0,164,0,139,0,53,0,63,0,68,0,126,0,0,0,188,0,229,0,96,0,0,0,0,0,120,0,130,0,232,0,0,0,238,0,205,0,23,0,175,0,102,0,191,0,0,0,210,0,221,0,216,0,218,0,115,0,35,0,249,0,208,0,76,0,52,0,250,0,0,0,87,0,99,0,82,0,42,0,131,0,198,0,210,0,0,0,27,0,192,0,55,0,120,0,9,0,46,0,0,0,67,0,143,0,62,0,114,0,237,0,188,0,154,0,250,0,248,0,0,0,101,0,79,0,145,0,0,0,0,0,94,0,103,0,148,0,126,0,237,0,92,0,32,0,108,0,74,0,68,0,255,0,84,0,146,0,57,0,127,0,63,0,29,0,0,0,175,0,231,0,205,0,45,0,28,0,207,0,55,0,0,0,7,0,166,0,3,0,107,0,220,0,0,0,60,0,149,0,44,0,135,0,208,0,238,0,81,0,0,0,0,0,129,0,240,0,118,0,187,0,143,0,29,0,171,0,116,0,53,0,143,0,163,0,143,0,99,0,168,0,155,0,0,0,0,0,0,0,0,0,123,0,120,0,144,0,207,0,0,0,85,0,0,0,134,0,40,0,226,0,204,0,246,0,30,0,0,0,0,0,94,0,163,0,208,0,21,0,17,0,238,0,8,0,0,0,187,0,107,0,0,0,189,0,157,0,24,0,175,0,213,0,0,0,34,0,112,0,64,0,249,0,0,0,41,0,237,0,151,0,89,0,164,0,55,0,247,0,141,0,89,0,0,0,125,0,148,0,45,0,225,0,217,0,122,0,88,0,104,0,56,0,0,0,251,0,0,0,170,0,250,0,77,0,0,0,0,0,210,0,242,0,0,0,0,0,241,0,0,0,0,0,195,0,197,0,93,0,0,0,246,0,0,0,153,0,0,0,91,0,232,0,236,0,170,0,188,0,0,0,59,0,63,0,226,0,148,0,141,0,228,0,111,0,170,0,44,0,8,0,225,0,202,0,229,0,0,0,0,0,90,0,184,0,207,0,141,0,0,0,238,0,239,0,197,0,112,0,238,0,92,0,60,0,20,0,138,0,32,0,20,0,115,0,120,0,38,0,211,0,233,0,113,0,187,0,193,0,0,0,183,0,0,0,44,0,39,0,107,0,25,0,49,0,0,0,0,0,0,0,146,0,247,0,191,0,191,0,135,0,0,0,188,0,237,0,121,0,206,0,0,0,0,0,217,0,28,0,240,0,222,0,76,0,0,0,168,0,170,0,84,0,114,0,88,0,1,0,209,0,0,0,0,0,137,0,0,0,198,0,208,0,166,0,167,0,0,0,248,0,249,0,138,0,128,0,0,0,40,0,144,0,130,0,200,0,0,0,0,0,137,0,102,0,27,0,182,0,120,0,224,0,0,0,218,0,89,0,77,0,83,0,20,0,181,0,246,0,19,0,123,0,17,0,112,0,28,0,148,0,19,0,145,0,223,0,185,0,183,0,103,0,172,0,68,0,203,0,224,0,68,0,89,0,152,0,250,0,248,0,251,0,117,0,194,0,222,0,0,0,0,0,0,0,0,0,0,0,0,0,193,0,190,0,8,0,0,0,154,0,15,0,155,0,184,0,0,0,0,0,42,0,233,0,107,0,122,0,42,0,216,0,202,0,90,0,82,0,79,0,182,0,11,0,0,0,76,0,0,0,26,0,0,0,88,0,0,0,0,0,0,0,0,0,48,0,148,0,0,0,39,0,0,0,97,0,35,0,26,0,0,0,0,0,6,0,170,0,4,0,0,0,0,0,0,0,194,0,96,0,31,0,0,0,215,0,0,0,184,0,175,0,218,0,39,0,165,0,0,0,230,0,172,0,22,0,34,0,75,0,72,0,98,0,132,0,0,0,12,0,0,0,0,0,12,0,117,0,0,0,187,0,171,0,0,0,158,0,197,0,176,0,254,0,233,0,30,0,0,0,60,0,88,0,2,0,107,0,6,0,64,0,34,0,1,0,12,0,19,0,0,0,38,0,0,0,166,0,0,0,0,0,119,0,153,0,119,0,158,0,135,0,0,0,152,0,231,0,169,0,38,0,169,0,0,0,122,0,19,0,162,0,0,0,200,0,22,0,255,0,36,0,138,0,88,0,0,0,0,0,206,0,46,0,55,0,206,0,73,0,218,0,86,0,195,0,247,0);
signal scenario_full  : scenario_type := (56,31,56,30,56,29,16,31,10,31,210,31,133,31,29,31,145,31,236,31,226,31,8,31,252,31,3,31,128,31,246,31,3,31,3,30,45,31,196,31,14,31,144,31,52,31,228,31,153,31,125,31,86,31,151,31,151,30,3,31,3,30,224,31,187,31,71,31,230,31,190,31,190,30,190,29,166,31,226,31,226,30,226,29,226,28,142,31,227,31,227,30,113,31,185,31,185,30,185,29,59,31,169,31,19,31,19,30,201,31,225,31,160,31,180,31,180,30,25,31,89,31,165,31,208,31,82,31,114,31,36,31,245,31,52,31,161,31,116,31,141,31,196,31,196,30,5,31,5,30,221,31,221,30,209,31,81,31,81,30,81,29,23,31,37,31,4,31,39,31,226,31,106,31,106,30,231,31,106,31,22,31,209,31,251,31,251,30,15,31,15,30,30,31,5,31,5,30,74,31,74,30,15,31,202,31,162,31,162,30,81,31,232,31,87,31,87,30,7,31,165,31,247,31,209,31,238,31,81,31,81,30,27,31,201,31,48,31,5,31,132,31,6,31,38,31,154,31,119,31,211,31,22,31,145,31,179,31,204,31,204,30,204,29,204,28,30,31,30,31,30,30,144,31,144,30,117,31,117,30,117,29,92,31,81,31,81,30,181,31,181,30,79,31,13,31,20,31,187,31,7,31,219,31,221,31,71,31,236,31,236,30,208,31,62,31,226,31,57,31,57,30,20,31,20,30,218,31,84,31,84,30,84,29,176,31,170,31,254,31,212,31,192,31,132,31,251,31,125,31,159,31,104,31,17,31,194,31,70,31,210,31,244,31,153,31,34,31,206,31,4,31,241,31,12,31,167,31,226,31,228,31,245,31,90,31,167,31,200,31,200,30,10,31,203,31,195,31,36,31,36,30,223,31,218,31,62,31,177,31,222,31,187,31,223,31,223,30,231,31,164,31,83,31,83,30,248,31,180,31,11,31,11,30,70,31,190,31,214,31,40,31,40,30,40,29,190,31,166,31,95,31,99,31,142,31,117,31,117,30,117,29,142,31,123,31,123,30,123,29,123,28,194,31,71,31,86,31,131,31,131,30,131,29,98,31,90,31,14,31,95,31,218,31,5,31,6,31,249,31,249,30,157,31,61,31,162,31,56,31,56,30,30,31,30,30,223,31,230,31,41,31,103,31,83,31,61,31,109,31,131,31,106,31,106,30,96,31,19,31,139,31,113,31,142,31,26,31,218,31,226,31,201,31,110,31,96,31,142,31,188,31,188,30,4,31,4,30,252,31,58,31,58,30,58,29,73,31,184,31,111,31,111,30,116,31,166,31,166,30,166,29,166,28,75,31,248,31,195,31,131,31,166,31,155,31,129,31,129,30,202,31,155,31,2,31,72,31,72,30,165,31,4,31,240,31,240,30,240,29,240,28,253,31,1,31,1,30,248,31,121,31,250,31,70,31,50,31,217,31,196,31,196,30,204,31,204,30,204,29,122,31,126,31,83,31,115,31,47,31,110,31,10,31,31,31,19,31,164,31,139,31,53,31,63,31,68,31,126,31,126,30,188,31,229,31,96,31,96,30,96,29,120,31,130,31,232,31,232,30,238,31,205,31,23,31,175,31,102,31,191,31,191,30,210,31,221,31,216,31,218,31,115,31,35,31,249,31,208,31,76,31,52,31,250,31,250,30,87,31,99,31,82,31,42,31,131,31,198,31,210,31,210,30,27,31,192,31,55,31,120,31,9,31,46,31,46,30,67,31,143,31,62,31,114,31,237,31,188,31,154,31,250,31,248,31,248,30,101,31,79,31,145,31,145,30,145,29,94,31,103,31,148,31,126,31,237,31,92,31,32,31,108,31,74,31,68,31,255,31,84,31,146,31,57,31,127,31,63,31,29,31,29,30,175,31,231,31,205,31,45,31,28,31,207,31,55,31,55,30,7,31,166,31,3,31,107,31,220,31,220,30,60,31,149,31,44,31,135,31,208,31,238,31,81,31,81,30,81,29,129,31,240,31,118,31,187,31,143,31,29,31,171,31,116,31,53,31,143,31,163,31,143,31,99,31,168,31,155,31,155,30,155,29,155,28,155,27,123,31,120,31,144,31,207,31,207,30,85,31,85,30,134,31,40,31,226,31,204,31,246,31,30,31,30,30,30,29,94,31,163,31,208,31,21,31,17,31,238,31,8,31,8,30,187,31,107,31,107,30,189,31,157,31,24,31,175,31,213,31,213,30,34,31,112,31,64,31,249,31,249,30,41,31,237,31,151,31,89,31,164,31,55,31,247,31,141,31,89,31,89,30,125,31,148,31,45,31,225,31,217,31,122,31,88,31,104,31,56,31,56,30,251,31,251,30,170,31,250,31,77,31,77,30,77,29,210,31,242,31,242,30,242,29,241,31,241,30,241,29,195,31,197,31,93,31,93,30,246,31,246,30,153,31,153,30,91,31,232,31,236,31,170,31,188,31,188,30,59,31,63,31,226,31,148,31,141,31,228,31,111,31,170,31,44,31,8,31,225,31,202,31,229,31,229,30,229,29,90,31,184,31,207,31,141,31,141,30,238,31,239,31,197,31,112,31,238,31,92,31,60,31,20,31,138,31,32,31,20,31,115,31,120,31,38,31,211,31,233,31,113,31,187,31,193,31,193,30,183,31,183,30,44,31,39,31,107,31,25,31,49,31,49,30,49,29,49,28,146,31,247,31,191,31,191,31,135,31,135,30,188,31,237,31,121,31,206,31,206,30,206,29,217,31,28,31,240,31,222,31,76,31,76,30,168,31,170,31,84,31,114,31,88,31,1,31,209,31,209,30,209,29,137,31,137,30,198,31,208,31,166,31,167,31,167,30,248,31,249,31,138,31,128,31,128,30,40,31,144,31,130,31,200,31,200,30,200,29,137,31,102,31,27,31,182,31,120,31,224,31,224,30,218,31,89,31,77,31,83,31,20,31,181,31,246,31,19,31,123,31,17,31,112,31,28,31,148,31,19,31,145,31,223,31,185,31,183,31,103,31,172,31,68,31,203,31,224,31,68,31,89,31,152,31,250,31,248,31,251,31,117,31,194,31,222,31,222,30,222,29,222,28,222,27,222,26,222,25,193,31,190,31,8,31,8,30,154,31,15,31,155,31,184,31,184,30,184,29,42,31,233,31,107,31,122,31,42,31,216,31,202,31,90,31,82,31,79,31,182,31,11,31,11,30,76,31,76,30,26,31,26,30,88,31,88,30,88,29,88,28,88,27,48,31,148,31,148,30,39,31,39,30,97,31,35,31,26,31,26,30,26,29,6,31,170,31,4,31,4,30,4,29,4,28,194,31,96,31,31,31,31,30,215,31,215,30,184,31,175,31,218,31,39,31,165,31,165,30,230,31,172,31,22,31,34,31,75,31,72,31,98,31,132,31,132,30,12,31,12,30,12,29,12,31,117,31,117,30,187,31,171,31,171,30,158,31,197,31,176,31,254,31,233,31,30,31,30,30,60,31,88,31,2,31,107,31,6,31,64,31,34,31,1,31,12,31,19,31,19,30,38,31,38,30,166,31,166,30,166,29,119,31,153,31,119,31,158,31,135,31,135,30,152,31,231,31,169,31,38,31,169,31,169,30,122,31,19,31,162,31,162,30,200,31,22,31,255,31,36,31,138,31,88,31,88,30,88,29,206,31,46,31,55,31,206,31,73,31,218,31,86,31,195,31,247,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
