-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_445 is
end project_tb_445;

architecture project_tb_arch_445 of project_tb_445 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 875;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (184,0,0,0,197,0,175,0,179,0,0,0,141,0,123,0,162,0,239,0,0,0,200,0,156,0,0,0,0,0,216,0,59,0,139,0,0,0,1,0,219,0,0,0,73,0,20,0,0,0,135,0,92,0,122,0,0,0,107,0,0,0,17,0,84,0,0,0,23,0,207,0,48,0,62,0,0,0,0,0,0,0,249,0,115,0,0,0,219,0,0,0,157,0,166,0,227,0,164,0,243,0,0,0,47,0,171,0,0,0,90,0,4,0,71,0,102,0,134,0,53,0,230,0,147,0,93,0,122,0,138,0,0,0,147,0,82,0,229,0,164,0,171,0,0,0,0,0,223,0,65,0,0,0,114,0,154,0,152,0,91,0,222,0,249,0,150,0,250,0,99,0,0,0,226,0,9,0,146,0,64,0,169,0,0,0,115,0,0,0,235,0,81,0,240,0,0,0,161,0,43,0,184,0,243,0,25,0,215,0,229,0,94,0,0,0,0,0,0,0,225,0,223,0,0,0,167,0,230,0,18,0,45,0,0,0,165,0,138,0,230,0,194,0,98,0,27,0,0,0,223,0,137,0,210,0,147,0,46,0,196,0,12,0,110,0,121,0,217,0,157,0,71,0,0,0,172,0,64,0,0,0,171,0,195,0,34,0,216,0,217,0,0,0,0,0,14,0,174,0,116,0,187,0,224,0,24,0,0,0,54,0,0,0,175,0,24,0,157,0,136,0,99,0,91,0,0,0,183,0,234,0,70,0,0,0,15,0,174,0,189,0,0,0,167,0,0,0,17,0,134,0,158,0,0,0,119,0,104,0,164,0,150,0,149,0,137,0,70,0,151,0,34,0,0,0,195,0,117,0,110,0,73,0,0,0,0,0,0,0,168,0,160,0,0,0,154,0,241,0,0,0,69,0,95,0,0,0,242,0,222,0,202,0,71,0,163,0,103,0,14,0,57,0,44,0,97,0,98,0,251,0,132,0,235,0,83,0,195,0,0,0,240,0,88,0,16,0,185,0,176,0,235,0,224,0,0,0,224,0,61,0,228,0,77,0,0,0,24,0,156,0,104,0,0,0,71,0,30,0,147,0,140,0,75,0,200,0,192,0,0,0,0,0,213,0,0,0,10,0,206,0,102,0,69,0,133,0,68,0,153,0,115,0,66,0,0,0,92,0,223,0,210,0,124,0,94,0,213,0,199,0,92,0,233,0,45,0,56,0,131,0,159,0,187,0,9,0,97,0,5,0,30,0,0,0,222,0,157,0,32,0,197,0,254,0,206,0,0,0,34,0,70,0,116,0,169,0,162,0,212,0,138,0,217,0,14,0,106,0,199,0,102,0,162,0,115,0,125,0,103,0,117,0,220,0,131,0,95,0,89,0,28,0,244,0,0,0,0,0,240,0,124,0,235,0,102,0,144,0,218,0,48,0,0,0,172,0,0,0,151,0,207,0,44,0,50,0,62,0,157,0,39,0,96,0,214,0,52,0,0,0,1,0,247,0,97,0,0,0,20,0,175,0,0,0,6,0,0,0,230,0,166,0,0,0,86,0,87,0,56,0,163,0,164,0,59,0,226,0,16,0,20,0,97,0,161,0,39,0,185,0,69,0,133,0,186,0,0,0,0,0,75,0,31,0,167,0,177,0,212,0,243,0,223,0,64,0,137,0,233,0,65,0,0,0,9,0,210,0,190,0,182,0,247,0,175,0,107,0,46,0,191,0,209,0,19,0,105,0,66,0,41,0,34,0,234,0,79,0,88,0,193,0,7,0,232,0,0,0,125,0,14,0,0,0,0,0,0,0,213,0,227,0,0,0,60,0,0,0,68,0,206,0,36,0,162,0,147,0,42,0,226,0,244,0,0,0,13,0,0,0,0,0,211,0,100,0,14,0,0,0,0,0,19,0,6,0,180,0,84,0,0,0,113,0,38,0,32,0,123,0,84,0,31,0,0,0,168,0,148,0,135,0,103,0,187,0,145,0,224,0,190,0,200,0,193,0,42,0,12,0,0,0,48,0,214,0,181,0,163,0,161,0,10,0,158,0,88,0,44,0,113,0,0,0,0,0,193,0,28,0,21,0,22,0,225,0,166,0,191,0,58,0,0,0,175,0,0,0,0,0,0,0,176,0,165,0,0,0,89,0,0,0,104,0,245,0,134,0,74,0,0,0,251,0,226,0,0,0,0,0,190,0,85,0,0,0,152,0,217,0,0,0,254,0,0,0,157,0,139,0,36,0,0,0,255,0,143,0,0,0,28,0,168,0,160,0,225,0,11,0,0,0,99,0,0,0,96,0,111,0,219,0,200,0,150,0,53,0,151,0,201,0,93,0,0,0,38,0,0,0,135,0,155,0,0,0,234,0,118,0,210,0,18,0,31,0,121,0,246,0,211,0,43,0,29,0,16,0,165,0,0,0,0,0,132,0,86,0,52,0,176,0,0,0,45,0,126,0,0,0,0,0,18,0,0,0,201,0,82,0,157,0,0,0,0,0,214,0,235,0,185,0,0,0,52,0,0,0,2,0,64,0,129,0,209,0,50,0,145,0,107,0,126,0,228,0,147,0,109,0,231,0,145,0,0,0,58,0,70,0,30,0,31,0,0,0,0,0,27,0,0,0,82,0,203,0,0,0,137,0,102,0,91,0,118,0,100,0,18,0,185,0,241,0,17,0,139,0,140,0,92,0,252,0,55,0,0,0,155,0,225,0,173,0,170,0,158,0,227,0,187,0,0,0,227,0,98,0,47,0,110,0,105,0,192,0,107,0,0,0,154,0,250,0,0,0,0,0,0,0,61,0,32,0,0,0,137,0,149,0,12,0,216,0,169,0,192,0,80,0,91,0,14,0,195,0,40,0,210,0,7,0,170,0,59,0,0,0,196,0,45,0,239,0,216,0,164,0,207,0,133,0,153,0,173,0,17,0,176,0,120,0,0,0,48,0,219,0,0,0,219,0,18,0,157,0,194,0,0,0,4,0,83,0,5,0,204,0,0,0,122,0,249,0,180,0,96,0,182,0,54,0,0,0,0,0,156,0,0,0,204,0,150,0,0,0,0,0,68,0,165,0,49,0,25,0,0,0,65,0,0,0,217,0,217,0,37,0,106,0,67,0,44,0,162,0,25,0,114,0,103,0,25,0,229,0,17,0,154,0,0,0,0,0,69,0,0,0,248,0,44,0,0,0,0,0,0,0,0,0,45,0,204,0,50,0,2,0,0,0,0,0,231,0,179,0,87,0,63,0,0,0,73,0,0,0,34,0,0,0,82,0,59,0,0,0,0,0,26,0,143,0,124,0,0,0,0,0,121,0,116,0,0,0,39,0,119,0,3,0,59,0,101,0,74,0,0,0,164,0,60,0,93,0,186,0,53,0,0,0,0,0,63,0,52,0,189,0,40,0,122,0,231,0,70,0,111,0,135,0,197,0,211,0,245,0,0,0,247,0,0,0,0,0,197,0,0,0,117,0,0,0,0,0,143,0,100,0,75,0,0,0,165,0,83,0,35,0,0,0,222,0,224,0,0,0,4,0,244,0,30,0,0,0,194,0,139,0,253,0,0,0,225,0,206,0,0,0,0,0,0,0,126,0,152,0,169,0,206,0,94,0,50,0,168,0,0,0,247,0,171,0,159,0,61,0,38,0,160,0,67,0,0,0,0,0,137,0,28,0,34,0,0,0,4,0,202,0,116,0,204,0,218,0,144,0,255,0,130,0,123,0,194,0,0,0,4,0,65,0,0,0,0,0,102,0,37,0,240,0,136,0,27,0,1,0,0,0,101,0,67,0,209,0,189,0,37,0,225,0,8,0,29,0,0,0,49,0,124,0,203,0,84,0,37,0,0,0,0,0,49,0,38,0,229,0,21,0,4,0,241,0,237,0,0,0,171,0,0,0,25,0,44,0,197,0,183,0,210,0,76,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (184,31,184,30,197,31,175,31,179,31,179,30,141,31,123,31,162,31,239,31,239,30,200,31,156,31,156,30,156,29,216,31,59,31,139,31,139,30,1,31,219,31,219,30,73,31,20,31,20,30,135,31,92,31,122,31,122,30,107,31,107,30,17,31,84,31,84,30,23,31,207,31,48,31,62,31,62,30,62,29,62,28,249,31,115,31,115,30,219,31,219,30,157,31,166,31,227,31,164,31,243,31,243,30,47,31,171,31,171,30,90,31,4,31,71,31,102,31,134,31,53,31,230,31,147,31,93,31,122,31,138,31,138,30,147,31,82,31,229,31,164,31,171,31,171,30,171,29,223,31,65,31,65,30,114,31,154,31,152,31,91,31,222,31,249,31,150,31,250,31,99,31,99,30,226,31,9,31,146,31,64,31,169,31,169,30,115,31,115,30,235,31,81,31,240,31,240,30,161,31,43,31,184,31,243,31,25,31,215,31,229,31,94,31,94,30,94,29,94,28,225,31,223,31,223,30,167,31,230,31,18,31,45,31,45,30,165,31,138,31,230,31,194,31,98,31,27,31,27,30,223,31,137,31,210,31,147,31,46,31,196,31,12,31,110,31,121,31,217,31,157,31,71,31,71,30,172,31,64,31,64,30,171,31,195,31,34,31,216,31,217,31,217,30,217,29,14,31,174,31,116,31,187,31,224,31,24,31,24,30,54,31,54,30,175,31,24,31,157,31,136,31,99,31,91,31,91,30,183,31,234,31,70,31,70,30,15,31,174,31,189,31,189,30,167,31,167,30,17,31,134,31,158,31,158,30,119,31,104,31,164,31,150,31,149,31,137,31,70,31,151,31,34,31,34,30,195,31,117,31,110,31,73,31,73,30,73,29,73,28,168,31,160,31,160,30,154,31,241,31,241,30,69,31,95,31,95,30,242,31,222,31,202,31,71,31,163,31,103,31,14,31,57,31,44,31,97,31,98,31,251,31,132,31,235,31,83,31,195,31,195,30,240,31,88,31,16,31,185,31,176,31,235,31,224,31,224,30,224,31,61,31,228,31,77,31,77,30,24,31,156,31,104,31,104,30,71,31,30,31,147,31,140,31,75,31,200,31,192,31,192,30,192,29,213,31,213,30,10,31,206,31,102,31,69,31,133,31,68,31,153,31,115,31,66,31,66,30,92,31,223,31,210,31,124,31,94,31,213,31,199,31,92,31,233,31,45,31,56,31,131,31,159,31,187,31,9,31,97,31,5,31,30,31,30,30,222,31,157,31,32,31,197,31,254,31,206,31,206,30,34,31,70,31,116,31,169,31,162,31,212,31,138,31,217,31,14,31,106,31,199,31,102,31,162,31,115,31,125,31,103,31,117,31,220,31,131,31,95,31,89,31,28,31,244,31,244,30,244,29,240,31,124,31,235,31,102,31,144,31,218,31,48,31,48,30,172,31,172,30,151,31,207,31,44,31,50,31,62,31,157,31,39,31,96,31,214,31,52,31,52,30,1,31,247,31,97,31,97,30,20,31,175,31,175,30,6,31,6,30,230,31,166,31,166,30,86,31,87,31,56,31,163,31,164,31,59,31,226,31,16,31,20,31,97,31,161,31,39,31,185,31,69,31,133,31,186,31,186,30,186,29,75,31,31,31,167,31,177,31,212,31,243,31,223,31,64,31,137,31,233,31,65,31,65,30,9,31,210,31,190,31,182,31,247,31,175,31,107,31,46,31,191,31,209,31,19,31,105,31,66,31,41,31,34,31,234,31,79,31,88,31,193,31,7,31,232,31,232,30,125,31,14,31,14,30,14,29,14,28,213,31,227,31,227,30,60,31,60,30,68,31,206,31,36,31,162,31,147,31,42,31,226,31,244,31,244,30,13,31,13,30,13,29,211,31,100,31,14,31,14,30,14,29,19,31,6,31,180,31,84,31,84,30,113,31,38,31,32,31,123,31,84,31,31,31,31,30,168,31,148,31,135,31,103,31,187,31,145,31,224,31,190,31,200,31,193,31,42,31,12,31,12,30,48,31,214,31,181,31,163,31,161,31,10,31,158,31,88,31,44,31,113,31,113,30,113,29,193,31,28,31,21,31,22,31,225,31,166,31,191,31,58,31,58,30,175,31,175,30,175,29,175,28,176,31,165,31,165,30,89,31,89,30,104,31,245,31,134,31,74,31,74,30,251,31,226,31,226,30,226,29,190,31,85,31,85,30,152,31,217,31,217,30,254,31,254,30,157,31,139,31,36,31,36,30,255,31,143,31,143,30,28,31,168,31,160,31,225,31,11,31,11,30,99,31,99,30,96,31,111,31,219,31,200,31,150,31,53,31,151,31,201,31,93,31,93,30,38,31,38,30,135,31,155,31,155,30,234,31,118,31,210,31,18,31,31,31,121,31,246,31,211,31,43,31,29,31,16,31,165,31,165,30,165,29,132,31,86,31,52,31,176,31,176,30,45,31,126,31,126,30,126,29,18,31,18,30,201,31,82,31,157,31,157,30,157,29,214,31,235,31,185,31,185,30,52,31,52,30,2,31,64,31,129,31,209,31,50,31,145,31,107,31,126,31,228,31,147,31,109,31,231,31,145,31,145,30,58,31,70,31,30,31,31,31,31,30,31,29,27,31,27,30,82,31,203,31,203,30,137,31,102,31,91,31,118,31,100,31,18,31,185,31,241,31,17,31,139,31,140,31,92,31,252,31,55,31,55,30,155,31,225,31,173,31,170,31,158,31,227,31,187,31,187,30,227,31,98,31,47,31,110,31,105,31,192,31,107,31,107,30,154,31,250,31,250,30,250,29,250,28,61,31,32,31,32,30,137,31,149,31,12,31,216,31,169,31,192,31,80,31,91,31,14,31,195,31,40,31,210,31,7,31,170,31,59,31,59,30,196,31,45,31,239,31,216,31,164,31,207,31,133,31,153,31,173,31,17,31,176,31,120,31,120,30,48,31,219,31,219,30,219,31,18,31,157,31,194,31,194,30,4,31,83,31,5,31,204,31,204,30,122,31,249,31,180,31,96,31,182,31,54,31,54,30,54,29,156,31,156,30,204,31,150,31,150,30,150,29,68,31,165,31,49,31,25,31,25,30,65,31,65,30,217,31,217,31,37,31,106,31,67,31,44,31,162,31,25,31,114,31,103,31,25,31,229,31,17,31,154,31,154,30,154,29,69,31,69,30,248,31,44,31,44,30,44,29,44,28,44,27,45,31,204,31,50,31,2,31,2,30,2,29,231,31,179,31,87,31,63,31,63,30,73,31,73,30,34,31,34,30,82,31,59,31,59,30,59,29,26,31,143,31,124,31,124,30,124,29,121,31,116,31,116,30,39,31,119,31,3,31,59,31,101,31,74,31,74,30,164,31,60,31,93,31,186,31,53,31,53,30,53,29,63,31,52,31,189,31,40,31,122,31,231,31,70,31,111,31,135,31,197,31,211,31,245,31,245,30,247,31,247,30,247,29,197,31,197,30,117,31,117,30,117,29,143,31,100,31,75,31,75,30,165,31,83,31,35,31,35,30,222,31,224,31,224,30,4,31,244,31,30,31,30,30,194,31,139,31,253,31,253,30,225,31,206,31,206,30,206,29,206,28,126,31,152,31,169,31,206,31,94,31,50,31,168,31,168,30,247,31,171,31,159,31,61,31,38,31,160,31,67,31,67,30,67,29,137,31,28,31,34,31,34,30,4,31,202,31,116,31,204,31,218,31,144,31,255,31,130,31,123,31,194,31,194,30,4,31,65,31,65,30,65,29,102,31,37,31,240,31,136,31,27,31,1,31,1,30,101,31,67,31,209,31,189,31,37,31,225,31,8,31,29,31,29,30,49,31,124,31,203,31,84,31,37,31,37,30,37,29,49,31,38,31,229,31,21,31,4,31,241,31,237,31,237,30,171,31,171,30,25,31,44,31,197,31,183,31,210,31,76,31,76,30,76,29,76,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
