-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 242;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,0,0,237,0,133,0,244,0,79,0,93,0,178,0,106,0,0,0,38,0,195,0,73,0,246,0,197,0,10,0,100,0,0,0,253,0,0,0,0,0,183,0,0,0,19,0,132,0,130,0,101,0,49,0,118,0,74,0,44,0,225,0,202,0,148,0,162,0,168,0,38,0,0,0,215,0,110,0,15,0,0,0,165,0,0,0,195,0,155,0,189,0,226,0,129,0,55,0,13,0,0,0,0,0,250,0,98,0,0,0,150,0,2,0,92,0,0,0,103,0,89,0,5,0,38,0,0,0,0,0,139,0,81,0,216,0,167,0,0,0,238,0,115,0,0,0,0,0,32,0,185,0,0,0,0,0,0,0,94,0,0,0,0,0,75,0,111,0,98,0,105,0,0,0,124,0,179,0,246,0,116,0,34,0,0,0,0,0,247,0,192,0,0,0,40,0,220,0,73,0,179,0,18,0,149,0,136,0,49,0,117,0,32,0,127,0,0,0,0,0,31,0,22,0,85,0,0,0,12,0,0,0,0,0,161,0,0,0,110,0,82,0,172,0,0,0,59,0,168,0,239,0,225,0,48,0,116,0,155,0,252,0,203,0,150,0,218,0,59,0,196,0,173,0,185,0,189,0,70,0,0,0,179,0,0,0,121,0,24,0,158,0,68,0,249,0,80,0,84,0,194,0,144,0,0,0,232,0,92,0,119,0,177,0,18,0,253,0,163,0,224,0,203,0,220,0,6,0,115,0,0,0,197,0,158,0,171,0,205,0,0,0,0,0,0,0,90,0,16,0,152,0,149,0,55,0,174,0,128,0,234,0,243,0,96,0,29,0,202,0,199,0,251,0,0,0,0,0,129,0,121,0,0,0,39,0,3,0,0,0,94,0,161,0,215,0,205,0,125,0,71,0,227,0,61,0,176,0,0,0,238,0,241,0,206,0,0,0,171,0,26,0,216,0,10,0,18,0,138,0,233,0,13,0,11,0,0,0,142,0,109,0,245,0,67,0,0,0,65,0,0,0,213,0,254,0,139,0,26,0,4,0,0,0,0,0,5,0,18,0,25,0,17,0,221,0,109,0,0,0,194,0);
signal scenario_full  : scenario_type := (219,31,219,30,237,31,133,31,244,31,79,31,93,31,178,31,106,31,106,30,38,31,195,31,73,31,246,31,197,31,10,31,100,31,100,30,253,31,253,30,253,29,183,31,183,30,19,31,132,31,130,31,101,31,49,31,118,31,74,31,44,31,225,31,202,31,148,31,162,31,168,31,38,31,38,30,215,31,110,31,15,31,15,30,165,31,165,30,195,31,155,31,189,31,226,31,129,31,55,31,13,31,13,30,13,29,250,31,98,31,98,30,150,31,2,31,92,31,92,30,103,31,89,31,5,31,38,31,38,30,38,29,139,31,81,31,216,31,167,31,167,30,238,31,115,31,115,30,115,29,32,31,185,31,185,30,185,29,185,28,94,31,94,30,94,29,75,31,111,31,98,31,105,31,105,30,124,31,179,31,246,31,116,31,34,31,34,30,34,29,247,31,192,31,192,30,40,31,220,31,73,31,179,31,18,31,149,31,136,31,49,31,117,31,32,31,127,31,127,30,127,29,31,31,22,31,85,31,85,30,12,31,12,30,12,29,161,31,161,30,110,31,82,31,172,31,172,30,59,31,168,31,239,31,225,31,48,31,116,31,155,31,252,31,203,31,150,31,218,31,59,31,196,31,173,31,185,31,189,31,70,31,70,30,179,31,179,30,121,31,24,31,158,31,68,31,249,31,80,31,84,31,194,31,144,31,144,30,232,31,92,31,119,31,177,31,18,31,253,31,163,31,224,31,203,31,220,31,6,31,115,31,115,30,197,31,158,31,171,31,205,31,205,30,205,29,205,28,90,31,16,31,152,31,149,31,55,31,174,31,128,31,234,31,243,31,96,31,29,31,202,31,199,31,251,31,251,30,251,29,129,31,121,31,121,30,39,31,3,31,3,30,94,31,161,31,215,31,205,31,125,31,71,31,227,31,61,31,176,31,176,30,238,31,241,31,206,31,206,30,171,31,26,31,216,31,10,31,18,31,138,31,233,31,13,31,11,31,11,30,142,31,109,31,245,31,67,31,67,30,65,31,65,30,213,31,254,31,139,31,26,31,4,31,4,30,4,29,5,31,18,31,25,31,17,31,221,31,109,31,109,30,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
