-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 909;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (253,0,254,0,0,0,106,0,0,0,11,0,1,0,65,0,135,0,53,0,238,0,105,0,0,0,217,0,82,0,163,0,123,0,0,0,47,0,188,0,59,0,65,0,119,0,111,0,110,0,87,0,87,0,240,0,72,0,0,0,116,0,91,0,139,0,0,0,169,0,100,0,144,0,0,0,179,0,46,0,180,0,244,0,27,0,36,0,242,0,90,0,216,0,96,0,242,0,0,0,0,0,39,0,0,0,241,0,0,0,71,0,83,0,17,0,24,0,116,0,77,0,59,0,0,0,123,0,0,0,73,0,1,0,185,0,105,0,130,0,48,0,84,0,244,0,0,0,0,0,0,0,80,0,75,0,46,0,93,0,0,0,111,0,88,0,141,0,27,0,137,0,29,0,0,0,96,0,56,0,169,0,0,0,113,0,212,0,87,0,123,0,92,0,0,0,0,0,116,0,0,0,168,0,10,0,0,0,56,0,222,0,187,0,232,0,23,0,127,0,8,0,0,0,142,0,128,0,116,0,173,0,13,0,158,0,21,0,173,0,167,0,147,0,127,0,0,0,103,0,102,0,227,0,242,0,129,0,0,0,118,0,107,0,133,0,25,0,218,0,0,0,75,0,120,0,166,0,75,0,151,0,0,0,46,0,0,0,50,0,11,0,90,0,246,0,228,0,0,0,225,0,0,0,186,0,0,0,118,0,187,0,79,0,189,0,89,0,74,0,204,0,57,0,22,0,255,0,51,0,17,0,0,0,125,0,218,0,236,0,11,0,225,0,0,0,106,0,0,0,67,0,4,0,0,0,0,0,36,0,55,0,0,0,230,0,160,0,169,0,167,0,124,0,54,0,216,0,167,0,220,0,69,0,0,0,173,0,24,0,11,0,34,0,121,0,6,0,222,0,213,0,230,0,127,0,226,0,50,0,249,0,150,0,46,0,148,0,21,0,177,0,204,0,51,0,34,0,215,0,0,0,56,0,114,0,156,0,17,0,58,0,236,0,129,0,0,0,143,0,164,0,162,0,31,0,67,0,131,0,0,0,151,0,76,0,179,0,0,0,0,0,0,0,0,0,168,0,154,0,0,0,60,0,247,0,204,0,0,0,73,0,185,0,167,0,242,0,242,0,107,0,114,0,201,0,112,0,114,0,37,0,0,0,181,0,0,0,26,0,54,0,242,0,114,0,182,0,124,0,0,0,230,0,42,0,64,0,83,0,156,0,119,0,106,0,233,0,0,0,135,0,244,0,133,0,45,0,113,0,11,0,42,0,56,0,17,0,202,0,0,0,96,0,0,0,134,0,153,0,111,0,0,0,43,0,207,0,234,0,0,0,135,0,0,0,0,0,195,0,176,0,143,0,84,0,250,0,0,0,146,0,122,0,203,0,46,0,197,0,81,0,69,0,20,0,0,0,20,0,38,0,4,0,203,0,16,0,120,0,247,0,225,0,182,0,7,0,171,0,146,0,29,0,0,0,135,0,219,0,58,0,136,0,82,0,202,0,228,0,255,0,70,0,6,0,186,0,202,0,34,0,200,0,223,0,69,0,69,0,0,0,32,0,199,0,175,0,132,0,181,0,0,0,55,0,174,0,164,0,155,0,55,0,0,0,0,0,238,0,15,0,234,0,72,0,150,0,0,0,110,0,67,0,234,0,220,0,26,0,0,0,0,0,233,0,40,0,67,0,178,0,0,0,15,0,13,0,153,0,104,0,125,0,231,0,0,0,41,0,217,0,2,0,206,0,10,0,85,0,0,0,181,0,33,0,156,0,186,0,42,0,110,0,189,0,49,0,0,0,197,0,110,0,166,0,75,0,198,0,91,0,27,0,66,0,151,0,123,0,214,0,14,0,229,0,0,0,123,0,0,0,75,0,142,0,148,0,233,0,85,0,0,0,0,0,0,0,34,0,0,0,220,0,192,0,92,0,123,0,167,0,230,0,218,0,0,0,44,0,25,0,60,0,83,0,233,0,142,0,58,0,209,0,91,0,0,0,208,0,94,0,130,0,64,0,190,0,211,0,0,0,0,0,170,0,0,0,255,0,168,0,245,0,79,0,0,0,0,0,14,0,99,0,200,0,45,0,186,0,0,0,68,0,204,0,98,0,217,0,186,0,0,0,195,0,5,0,188,0,226,0,202,0,113,0,0,0,171,0,3,0,17,0,36,0,188,0,23,0,0,0,21,0,180,0,242,0,147,0,0,0,56,0,0,0,182,0,0,0,0,0,0,0,23,0,36,0,150,0,43,0,98,0,78,0,246,0,58,0,228,0,245,0,206,0,119,0,111,0,192,0,0,0,226,0,230,0,45,0,189,0,103,0,9,0,31,0,16,0,0,0,40,0,159,0,0,0,44,0,9,0,124,0,0,0,0,0,0,0,150,0,18,0,36,0,113,0,70,0,226,0,233,0,171,0,0,0,88,0,75,0,0,0,253,0,44,0,204,0,23,0,11,0,0,0,0,0,204,0,253,0,100,0,150,0,92,0,211,0,153,0,0,0,73,0,0,0,68,0,211,0,14,0,131,0,0,0,19,0,91,0,142,0,0,0,26,0,185,0,0,0,240,0,230,0,3,0,254,0,144,0,191,0,208,0,29,0,243,0,0,0,167,0,81,0,174,0,67,0,208,0,0,0,66,0,172,0,248,0,0,0,173,0,140,0,241,0,0,0,48,0,111,0,83,0,63,0,95,0,119,0,36,0,0,0,0,0,0,0,0,0,113,0,183,0,60,0,109,0,38,0,216,0,116,0,92,0,122,0,102,0,248,0,136,0,103,0,148,0,59,0,0,0,10,0,41,0,148,0,89,0,38,0,156,0,0,0,56,0,229,0,74,0,0,0,212,0,0,0,35,0,236,0,247,0,0,0,41,0,82,0,0,0,155,0,126,0,67,0,107,0,0,0,36,0,217,0,85,0,78,0,251,0,0,0,116,0,251,0,187,0,0,0,179,0,90,0,88,0,160,0,0,0,234,0,123,0,250,0,46,0,209,0,0,0,252,0,239,0,48,0,204,0,199,0,53,0,126,0,5,0,87,0,6,0,126,0,101,0,161,0,197,0,135,0,89,0,120,0,70,0,91,0,204,0,100,0,0,0,0,0,103,0,123,0,84,0,0,0,51,0,0,0,231,0,0,0,215,0,158,0,177,0,0,0,206,0,141,0,64,0,0,0,187,0,110,0,0,0,41,0,234,0,202,0,197,0,223,0,83,0,141,0,36,0,68,0,10,0,121,0,151,0,40,0,0,0,95,0,156,0,212,0,42,0,37,0,113,0,0,0,30,0,0,0,165,0,78,0,146,0,0,0,0,0,0,0,140,0,203,0,0,0,224,0,119,0,2,0,49,0,121,0,35,0,61,0,179,0,0,0,147,0,148,0,240,0,58,0,147,0,61,0,184,0,205,0,84,0,211,0,0,0,0,0,200,0,11,0,94,0,140,0,12,0,24,0,0,0,12,0,254,0,141,0,191,0,29,0,145,0,69,0,166,0,114,0,175,0,223,0,112,0,91,0,127,0,0,0,0,0,152,0,0,0,19,0,200,0,25,0,110,0,58,0,37,0,99,0,0,0,162,0,115,0,100,0,0,0,120,0,240,0,156,0,214,0,165,0,0,0,146,0,166,0,148,0,66,0,168,0,0,0,86,0,21,0,24,0,140,0,0,0,68,0,209,0,112,0,22,0,142,0,152,0,17,0,0,0,102,0,0,0,138,0,176,0,204,0,162,0,186,0,151,0,150,0,112,0,0,0,117,0,0,0,3,0,0,0,115,0,0,0,168,0,145,0,202,0,9,0,249,0,54,0,229,0,118,0,148,0,192,0,154,0,244,0,123,0,0,0,0,0,0,0,0,0,208,0,0,0,59,0,60,0,112,0,215,0,121,0,0,0,0,0,246,0,175,0,125,0,96,0,65,0,70,0,149,0,141,0,56,0,0,0,0,0,175,0,33,0,227,0,32,0,154,0,140,0,136,0,245,0,14,0,235,0,57,0,98,0,69,0,6,0,119,0,21,0,29,0,191,0,167,0,167,0,233,0,66,0,0,0,0,0,27,0,245,0,97,0,73,0,0,0,79,0);
signal scenario_full  : scenario_type := (253,31,254,31,254,30,106,31,106,30,11,31,1,31,65,31,135,31,53,31,238,31,105,31,105,30,217,31,82,31,163,31,123,31,123,30,47,31,188,31,59,31,65,31,119,31,111,31,110,31,87,31,87,31,240,31,72,31,72,30,116,31,91,31,139,31,139,30,169,31,100,31,144,31,144,30,179,31,46,31,180,31,244,31,27,31,36,31,242,31,90,31,216,31,96,31,242,31,242,30,242,29,39,31,39,30,241,31,241,30,71,31,83,31,17,31,24,31,116,31,77,31,59,31,59,30,123,31,123,30,73,31,1,31,185,31,105,31,130,31,48,31,84,31,244,31,244,30,244,29,244,28,80,31,75,31,46,31,93,31,93,30,111,31,88,31,141,31,27,31,137,31,29,31,29,30,96,31,56,31,169,31,169,30,113,31,212,31,87,31,123,31,92,31,92,30,92,29,116,31,116,30,168,31,10,31,10,30,56,31,222,31,187,31,232,31,23,31,127,31,8,31,8,30,142,31,128,31,116,31,173,31,13,31,158,31,21,31,173,31,167,31,147,31,127,31,127,30,103,31,102,31,227,31,242,31,129,31,129,30,118,31,107,31,133,31,25,31,218,31,218,30,75,31,120,31,166,31,75,31,151,31,151,30,46,31,46,30,50,31,11,31,90,31,246,31,228,31,228,30,225,31,225,30,186,31,186,30,118,31,187,31,79,31,189,31,89,31,74,31,204,31,57,31,22,31,255,31,51,31,17,31,17,30,125,31,218,31,236,31,11,31,225,31,225,30,106,31,106,30,67,31,4,31,4,30,4,29,36,31,55,31,55,30,230,31,160,31,169,31,167,31,124,31,54,31,216,31,167,31,220,31,69,31,69,30,173,31,24,31,11,31,34,31,121,31,6,31,222,31,213,31,230,31,127,31,226,31,50,31,249,31,150,31,46,31,148,31,21,31,177,31,204,31,51,31,34,31,215,31,215,30,56,31,114,31,156,31,17,31,58,31,236,31,129,31,129,30,143,31,164,31,162,31,31,31,67,31,131,31,131,30,151,31,76,31,179,31,179,30,179,29,179,28,179,27,168,31,154,31,154,30,60,31,247,31,204,31,204,30,73,31,185,31,167,31,242,31,242,31,107,31,114,31,201,31,112,31,114,31,37,31,37,30,181,31,181,30,26,31,54,31,242,31,114,31,182,31,124,31,124,30,230,31,42,31,64,31,83,31,156,31,119,31,106,31,233,31,233,30,135,31,244,31,133,31,45,31,113,31,11,31,42,31,56,31,17,31,202,31,202,30,96,31,96,30,134,31,153,31,111,31,111,30,43,31,207,31,234,31,234,30,135,31,135,30,135,29,195,31,176,31,143,31,84,31,250,31,250,30,146,31,122,31,203,31,46,31,197,31,81,31,69,31,20,31,20,30,20,31,38,31,4,31,203,31,16,31,120,31,247,31,225,31,182,31,7,31,171,31,146,31,29,31,29,30,135,31,219,31,58,31,136,31,82,31,202,31,228,31,255,31,70,31,6,31,186,31,202,31,34,31,200,31,223,31,69,31,69,31,69,30,32,31,199,31,175,31,132,31,181,31,181,30,55,31,174,31,164,31,155,31,55,31,55,30,55,29,238,31,15,31,234,31,72,31,150,31,150,30,110,31,67,31,234,31,220,31,26,31,26,30,26,29,233,31,40,31,67,31,178,31,178,30,15,31,13,31,153,31,104,31,125,31,231,31,231,30,41,31,217,31,2,31,206,31,10,31,85,31,85,30,181,31,33,31,156,31,186,31,42,31,110,31,189,31,49,31,49,30,197,31,110,31,166,31,75,31,198,31,91,31,27,31,66,31,151,31,123,31,214,31,14,31,229,31,229,30,123,31,123,30,75,31,142,31,148,31,233,31,85,31,85,30,85,29,85,28,34,31,34,30,220,31,192,31,92,31,123,31,167,31,230,31,218,31,218,30,44,31,25,31,60,31,83,31,233,31,142,31,58,31,209,31,91,31,91,30,208,31,94,31,130,31,64,31,190,31,211,31,211,30,211,29,170,31,170,30,255,31,168,31,245,31,79,31,79,30,79,29,14,31,99,31,200,31,45,31,186,31,186,30,68,31,204,31,98,31,217,31,186,31,186,30,195,31,5,31,188,31,226,31,202,31,113,31,113,30,171,31,3,31,17,31,36,31,188,31,23,31,23,30,21,31,180,31,242,31,147,31,147,30,56,31,56,30,182,31,182,30,182,29,182,28,23,31,36,31,150,31,43,31,98,31,78,31,246,31,58,31,228,31,245,31,206,31,119,31,111,31,192,31,192,30,226,31,230,31,45,31,189,31,103,31,9,31,31,31,16,31,16,30,40,31,159,31,159,30,44,31,9,31,124,31,124,30,124,29,124,28,150,31,18,31,36,31,113,31,70,31,226,31,233,31,171,31,171,30,88,31,75,31,75,30,253,31,44,31,204,31,23,31,11,31,11,30,11,29,204,31,253,31,100,31,150,31,92,31,211,31,153,31,153,30,73,31,73,30,68,31,211,31,14,31,131,31,131,30,19,31,91,31,142,31,142,30,26,31,185,31,185,30,240,31,230,31,3,31,254,31,144,31,191,31,208,31,29,31,243,31,243,30,167,31,81,31,174,31,67,31,208,31,208,30,66,31,172,31,248,31,248,30,173,31,140,31,241,31,241,30,48,31,111,31,83,31,63,31,95,31,119,31,36,31,36,30,36,29,36,28,36,27,113,31,183,31,60,31,109,31,38,31,216,31,116,31,92,31,122,31,102,31,248,31,136,31,103,31,148,31,59,31,59,30,10,31,41,31,148,31,89,31,38,31,156,31,156,30,56,31,229,31,74,31,74,30,212,31,212,30,35,31,236,31,247,31,247,30,41,31,82,31,82,30,155,31,126,31,67,31,107,31,107,30,36,31,217,31,85,31,78,31,251,31,251,30,116,31,251,31,187,31,187,30,179,31,90,31,88,31,160,31,160,30,234,31,123,31,250,31,46,31,209,31,209,30,252,31,239,31,48,31,204,31,199,31,53,31,126,31,5,31,87,31,6,31,126,31,101,31,161,31,197,31,135,31,89,31,120,31,70,31,91,31,204,31,100,31,100,30,100,29,103,31,123,31,84,31,84,30,51,31,51,30,231,31,231,30,215,31,158,31,177,31,177,30,206,31,141,31,64,31,64,30,187,31,110,31,110,30,41,31,234,31,202,31,197,31,223,31,83,31,141,31,36,31,68,31,10,31,121,31,151,31,40,31,40,30,95,31,156,31,212,31,42,31,37,31,113,31,113,30,30,31,30,30,165,31,78,31,146,31,146,30,146,29,146,28,140,31,203,31,203,30,224,31,119,31,2,31,49,31,121,31,35,31,61,31,179,31,179,30,147,31,148,31,240,31,58,31,147,31,61,31,184,31,205,31,84,31,211,31,211,30,211,29,200,31,11,31,94,31,140,31,12,31,24,31,24,30,12,31,254,31,141,31,191,31,29,31,145,31,69,31,166,31,114,31,175,31,223,31,112,31,91,31,127,31,127,30,127,29,152,31,152,30,19,31,200,31,25,31,110,31,58,31,37,31,99,31,99,30,162,31,115,31,100,31,100,30,120,31,240,31,156,31,214,31,165,31,165,30,146,31,166,31,148,31,66,31,168,31,168,30,86,31,21,31,24,31,140,31,140,30,68,31,209,31,112,31,22,31,142,31,152,31,17,31,17,30,102,31,102,30,138,31,176,31,204,31,162,31,186,31,151,31,150,31,112,31,112,30,117,31,117,30,3,31,3,30,115,31,115,30,168,31,145,31,202,31,9,31,249,31,54,31,229,31,118,31,148,31,192,31,154,31,244,31,123,31,123,30,123,29,123,28,123,27,208,31,208,30,59,31,60,31,112,31,215,31,121,31,121,30,121,29,246,31,175,31,125,31,96,31,65,31,70,31,149,31,141,31,56,31,56,30,56,29,175,31,33,31,227,31,32,31,154,31,140,31,136,31,245,31,14,31,235,31,57,31,98,31,69,31,6,31,119,31,21,31,29,31,191,31,167,31,167,31,233,31,66,31,66,30,66,29,27,31,245,31,97,31,73,31,73,30,79,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
