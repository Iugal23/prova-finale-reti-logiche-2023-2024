-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 290;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,150,0,51,0,99,0,0,0,0,0,1,0,23,0,0,0,78,0,0,0,40,0,8,0,181,0,149,0,24,0,69,0,56,0,243,0,236,0,212,0,0,0,201,0,23,0,20,0,197,0,136,0,228,0,180,0,0,0,251,0,0,0,183,0,172,0,0,0,0,0,155,0,141,0,214,0,99,0,71,0,18,0,0,0,0,0,67,0,240,0,48,0,210,0,0,0,222,0,215,0,111,0,62,0,222,0,24,0,0,0,114,0,171,0,145,0,68,0,233,0,76,0,3,0,143,0,101,0,66,0,40,0,37,0,98,0,154,0,22,0,76,0,39,0,13,0,0,0,229,0,11,0,74,0,158,0,88,0,43,0,0,0,191,0,227,0,252,0,138,0,188,0,34,0,140,0,0,0,0,0,43,0,207,0,110,0,188,0,161,0,0,0,52,0,12,0,65,0,116,0,141,0,94,0,168,0,142,0,0,0,0,0,0,0,158,0,31,0,127,0,134,0,164,0,179,0,0,0,207,0,62,0,186,0,39,0,164,0,63,0,0,0,132,0,199,0,0,0,135,0,85,0,189,0,210,0,162,0,106,0,213,0,21,0,62,0,42,0,19,0,234,0,0,0,0,0,239,0,0,0,248,0,149,0,164,0,0,0,0,0,68,0,96,0,158,0,0,0,52,0,243,0,0,0,0,0,213,0,142,0,235,0,125,0,0,0,165,0,0,0,0,0,95,0,187,0,34,0,160,0,7,0,23,0,146,0,28,0,0,0,32,0,0,0,61,0,110,0,154,0,9,0,158,0,181,0,140,0,0,0,172,0,132,0,0,0,180,0,85,0,0,0,212,0,150,0,9,0,19,0,106,0,0,0,140,0,239,0,66,0,108,0,211,0,189,0,106,0,122,0,40,0,237,0,173,0,0,0,243,0,0,0,0,0,57,0,80,0,106,0,115,0,0,0,217,0,29,0,153,0,0,0,235,0,227,0,183,0,143,0,93,0,0,0,0,0,116,0,94,0,0,0,239,0,0,0,204,0,0,0,72,0,0,0,131,0,75,0,173,0,101,0,51,0,146,0,234,0,214,0,211,0,116,0,248,0,21,0,147,0,185,0,59,0,83,0,74,0,136,0,129,0,211,0,79,0,54,0,99,0,0,0,0,0,138,0,113,0,97,0,20,0,0,0,153,0,26,0,111,0,117,0,202,0,233,0,21,0,158,0,0,0,7,0,28,0,196,0,114,0,133,0,0,0,0,0,31,0,27,0,0,0,187,0,65,0,0,0,0,0,152,0,164,0,72,0,104,0);
signal scenario_full  : scenario_type := (7,31,150,31,51,31,99,31,99,30,99,29,1,31,23,31,23,30,78,31,78,30,40,31,8,31,181,31,149,31,24,31,69,31,56,31,243,31,236,31,212,31,212,30,201,31,23,31,20,31,197,31,136,31,228,31,180,31,180,30,251,31,251,30,183,31,172,31,172,30,172,29,155,31,141,31,214,31,99,31,71,31,18,31,18,30,18,29,67,31,240,31,48,31,210,31,210,30,222,31,215,31,111,31,62,31,222,31,24,31,24,30,114,31,171,31,145,31,68,31,233,31,76,31,3,31,143,31,101,31,66,31,40,31,37,31,98,31,154,31,22,31,76,31,39,31,13,31,13,30,229,31,11,31,74,31,158,31,88,31,43,31,43,30,191,31,227,31,252,31,138,31,188,31,34,31,140,31,140,30,140,29,43,31,207,31,110,31,188,31,161,31,161,30,52,31,12,31,65,31,116,31,141,31,94,31,168,31,142,31,142,30,142,29,142,28,158,31,31,31,127,31,134,31,164,31,179,31,179,30,207,31,62,31,186,31,39,31,164,31,63,31,63,30,132,31,199,31,199,30,135,31,85,31,189,31,210,31,162,31,106,31,213,31,21,31,62,31,42,31,19,31,234,31,234,30,234,29,239,31,239,30,248,31,149,31,164,31,164,30,164,29,68,31,96,31,158,31,158,30,52,31,243,31,243,30,243,29,213,31,142,31,235,31,125,31,125,30,165,31,165,30,165,29,95,31,187,31,34,31,160,31,7,31,23,31,146,31,28,31,28,30,32,31,32,30,61,31,110,31,154,31,9,31,158,31,181,31,140,31,140,30,172,31,132,31,132,30,180,31,85,31,85,30,212,31,150,31,9,31,19,31,106,31,106,30,140,31,239,31,66,31,108,31,211,31,189,31,106,31,122,31,40,31,237,31,173,31,173,30,243,31,243,30,243,29,57,31,80,31,106,31,115,31,115,30,217,31,29,31,153,31,153,30,235,31,227,31,183,31,143,31,93,31,93,30,93,29,116,31,94,31,94,30,239,31,239,30,204,31,204,30,72,31,72,30,131,31,75,31,173,31,101,31,51,31,146,31,234,31,214,31,211,31,116,31,248,31,21,31,147,31,185,31,59,31,83,31,74,31,136,31,129,31,211,31,79,31,54,31,99,31,99,30,99,29,138,31,113,31,97,31,20,31,20,30,153,31,26,31,111,31,117,31,202,31,233,31,21,31,158,31,158,30,7,31,28,31,196,31,114,31,133,31,133,30,133,29,31,31,27,31,27,30,187,31,65,31,65,30,65,29,152,31,164,31,72,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
