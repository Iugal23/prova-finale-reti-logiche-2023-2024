-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_276 is
end project_tb_276;

architecture project_tb_arch_276 of project_tb_276 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 738;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (26,0,0,0,11,0,171,0,204,0,40,0,59,0,50,0,190,0,77,0,0,0,0,0,220,0,65,0,147,0,162,0,104,0,72,0,15,0,86,0,125,0,174,0,0,0,5,0,124,0,142,0,162,0,0,0,241,0,173,0,13,0,122,0,135,0,183,0,41,0,120,0,35,0,32,0,251,0,36,0,0,0,19,0,219,0,0,0,131,0,185,0,228,0,97,0,70,0,214,0,95,0,0,0,111,0,0,0,206,0,0,0,236,0,40,0,134,0,40,0,0,0,242,0,0,0,106,0,249,0,131,0,118,0,10,0,219,0,0,0,157,0,86,0,227,0,4,0,174,0,0,0,110,0,101,0,127,0,213,0,252,0,89,0,144,0,111,0,241,0,0,0,67,0,207,0,0,0,121,0,91,0,228,0,0,0,253,0,19,0,125,0,73,0,19,0,156,0,180,0,125,0,55,0,161,0,240,0,188,0,68,0,5,0,253,0,49,0,3,0,0,0,0,0,0,0,46,0,140,0,0,0,129,0,148,0,89,0,0,0,158,0,60,0,18,0,214,0,213,0,254,0,224,0,151,0,18,0,113,0,188,0,17,0,117,0,105,0,0,0,103,0,208,0,37,0,152,0,21,0,177,0,99,0,197,0,0,0,34,0,115,0,0,0,193,0,167,0,0,0,0,0,232,0,161,0,45,0,33,0,39,0,99,0,218,0,12,0,245,0,51,0,215,0,143,0,95,0,0,0,47,0,109,0,0,0,99,0,155,0,0,0,80,0,225,0,161,0,105,0,78,0,53,0,54,0,62,0,0,0,165,0,237,0,0,0,55,0,206,0,177,0,1,0,237,0,121,0,57,0,80,0,0,0,85,0,34,0,249,0,8,0,36,0,0,0,115,0,98,0,158,0,251,0,42,0,134,0,240,0,143,0,75,0,98,0,0,0,212,0,203,0,79,0,61,0,0,0,143,0,38,0,0,0,128,0,67,0,54,0,81,0,0,0,253,0,58,0,90,0,59,0,0,0,23,0,114,0,0,0,203,0,0,0,0,0,0,0,122,0,28,0,59,0,80,0,129,0,0,0,121,0,150,0,56,0,0,0,77,0,182,0,251,0,29,0,0,0,4,0,148,0,221,0,0,0,37,0,248,0,234,0,208,0,223,0,171,0,0,0,0,0,104,0,84,0,20,0,0,0,0,0,15,0,242,0,0,0,30,0,199,0,46,0,251,0,232,0,73,0,20,0,0,0,158,0,240,0,149,0,248,0,119,0,157,0,101,0,0,0,148,0,230,0,149,0,46,0,13,0,208,0,76,0,244,0,240,0,91,0,0,0,80,0,106,0,224,0,52,0,100,0,191,0,251,0,71,0,140,0,143,0,159,0,11,0,212,0,160,0,153,0,152,0,0,0,0,0,127,0,30,0,160,0,252,0,0,0,236,0,0,0,0,0,165,0,152,0,124,0,1,0,248,0,248,0,14,0,0,0,45,0,0,0,104,0,200,0,230,0,250,0,14,0,44,0,191,0,93,0,108,0,0,0,100,0,18,0,123,0,244,0,138,0,130,0,70,0,93,0,188,0,112,0,119,0,201,0,12,0,0,0,0,0,187,0,71,0,67,0,169,0,99,0,98,0,119,0,170,0,61,0,33,0,91,0,171,0,186,0,7,0,201,0,246,0,5,0,58,0,0,0,0,0,29,0,146,0,2,0,38,0,41,0,151,0,104,0,0,0,134,0,0,0,221,0,0,0,205,0,111,0,238,0,0,0,187,0,0,0,28,0,0,0,13,0,0,0,131,0,58,0,235,0,0,0,42,0,0,0,157,0,0,0,32,0,0,0,4,0,214,0,208,0,251,0,120,0,154,0,0,0,0,0,159,0,48,0,67,0,187,0,81,0,53,0,57,0,117,0,44,0,231,0,0,0,166,0,0,0,0,0,114,0,244,0,242,0,7,0,160,0,0,0,179,0,195,0,150,0,20,0,0,0,136,0,180,0,186,0,199,0,74,0,111,0,74,0,218,0,0,0,197,0,43,0,238,0,0,0,144,0,153,0,0,0,105,0,0,0,0,0,237,0,129,0,190,0,20,0,85,0,236,0,218,0,0,0,44,0,0,0,80,0,219,0,238,0,47,0,137,0,156,0,215,0,153,0,0,0,27,0,218,0,78,0,134,0,29,0,231,0,0,0,237,0,67,0,47,0,205,0,153,0,186,0,5,0,252,0,217,0,49,0,146,0,221,0,167,0,148,0,252,0,95,0,235,0,240,0,0,0,166,0,190,0,201,0,23,0,217,0,0,0,227,0,202,0,105,0,15,0,90,0,129,0,245,0,1,0,69,0,0,0,96,0,0,0,0,0,3,0,252,0,198,0,85,0,0,0,113,0,38,0,223,0,32,0,219,0,0,0,18,0,0,0,103,0,201,0,35,0,35,0,76,0,149,0,139,0,207,0,193,0,144,0,0,0,0,0,92,0,94,0,211,0,197,0,47,0,0,0,236,0,102,0,206,0,8,0,34,0,163,0,0,0,45,0,61,0,51,0,251,0,0,0,0,0,245,0,137,0,225,0,149,0,107,0,238,0,41,0,203,0,141,0,67,0,73,0,52,0,67,0,72,0,0,0,4,0,60,0,106,0,60,0,46,0,138,0,29,0,82,0,0,0,251,0,138,0,209,0,152,0,138,0,156,0,0,0,178,0,169,0,0,0,203,0,237,0,0,0,109,0,234,0,0,0,81,0,26,0,235,0,61,0,246,0,155,0,171,0,94,0,0,0,0,0,29,0,19,0,247,0,210,0,0,0,234,0,0,0,155,0,160,0,126,0,181,0,0,0,149,0,182,0,0,0,0,0,6,0,76,0,39,0,49,0,110,0,0,0,2,0,120,0,0,0,0,0,66,0,183,0,148,0,248,0,0,0,0,0,249,0,48,0,44,0,24,0,193,0,202,0,73,0,198,0,180,0,60,0,191,0,75,0,77,0,213,0,180,0,206,0,2,0,203,0,246,0,85,0,0,0,228,0,101,0,136,0,84,0,248,0,0,0,6,0,130,0,188,0,252,0,0,0,66,0,0,0,132,0,94,0,55,0,198,0,52,0,138,0,0,0,131,0,141,0,141,0,0,0,119,0,0,0,187,0,28,0,244,0,74,0,55,0,208,0,178,0,0,0,223,0,46,0,196,0,0,0,124,0,139,0,5,0,13,0,0,0,226,0,149,0,64,0,78,0,66,0,12,0,0,0,0,0,245,0,7,0,47,0,80,0,220,0,38,0,0,0,184,0,171,0,124,0,169,0,190,0,0,0,0,0,40,0);
signal scenario_full  : scenario_type := (26,31,26,30,11,31,171,31,204,31,40,31,59,31,50,31,190,31,77,31,77,30,77,29,220,31,65,31,147,31,162,31,104,31,72,31,15,31,86,31,125,31,174,31,174,30,5,31,124,31,142,31,162,31,162,30,241,31,173,31,13,31,122,31,135,31,183,31,41,31,120,31,35,31,32,31,251,31,36,31,36,30,19,31,219,31,219,30,131,31,185,31,228,31,97,31,70,31,214,31,95,31,95,30,111,31,111,30,206,31,206,30,236,31,40,31,134,31,40,31,40,30,242,31,242,30,106,31,249,31,131,31,118,31,10,31,219,31,219,30,157,31,86,31,227,31,4,31,174,31,174,30,110,31,101,31,127,31,213,31,252,31,89,31,144,31,111,31,241,31,241,30,67,31,207,31,207,30,121,31,91,31,228,31,228,30,253,31,19,31,125,31,73,31,19,31,156,31,180,31,125,31,55,31,161,31,240,31,188,31,68,31,5,31,253,31,49,31,3,31,3,30,3,29,3,28,46,31,140,31,140,30,129,31,148,31,89,31,89,30,158,31,60,31,18,31,214,31,213,31,254,31,224,31,151,31,18,31,113,31,188,31,17,31,117,31,105,31,105,30,103,31,208,31,37,31,152,31,21,31,177,31,99,31,197,31,197,30,34,31,115,31,115,30,193,31,167,31,167,30,167,29,232,31,161,31,45,31,33,31,39,31,99,31,218,31,12,31,245,31,51,31,215,31,143,31,95,31,95,30,47,31,109,31,109,30,99,31,155,31,155,30,80,31,225,31,161,31,105,31,78,31,53,31,54,31,62,31,62,30,165,31,237,31,237,30,55,31,206,31,177,31,1,31,237,31,121,31,57,31,80,31,80,30,85,31,34,31,249,31,8,31,36,31,36,30,115,31,98,31,158,31,251,31,42,31,134,31,240,31,143,31,75,31,98,31,98,30,212,31,203,31,79,31,61,31,61,30,143,31,38,31,38,30,128,31,67,31,54,31,81,31,81,30,253,31,58,31,90,31,59,31,59,30,23,31,114,31,114,30,203,31,203,30,203,29,203,28,122,31,28,31,59,31,80,31,129,31,129,30,121,31,150,31,56,31,56,30,77,31,182,31,251,31,29,31,29,30,4,31,148,31,221,31,221,30,37,31,248,31,234,31,208,31,223,31,171,31,171,30,171,29,104,31,84,31,20,31,20,30,20,29,15,31,242,31,242,30,30,31,199,31,46,31,251,31,232,31,73,31,20,31,20,30,158,31,240,31,149,31,248,31,119,31,157,31,101,31,101,30,148,31,230,31,149,31,46,31,13,31,208,31,76,31,244,31,240,31,91,31,91,30,80,31,106,31,224,31,52,31,100,31,191,31,251,31,71,31,140,31,143,31,159,31,11,31,212,31,160,31,153,31,152,31,152,30,152,29,127,31,30,31,160,31,252,31,252,30,236,31,236,30,236,29,165,31,152,31,124,31,1,31,248,31,248,31,14,31,14,30,45,31,45,30,104,31,200,31,230,31,250,31,14,31,44,31,191,31,93,31,108,31,108,30,100,31,18,31,123,31,244,31,138,31,130,31,70,31,93,31,188,31,112,31,119,31,201,31,12,31,12,30,12,29,187,31,71,31,67,31,169,31,99,31,98,31,119,31,170,31,61,31,33,31,91,31,171,31,186,31,7,31,201,31,246,31,5,31,58,31,58,30,58,29,29,31,146,31,2,31,38,31,41,31,151,31,104,31,104,30,134,31,134,30,221,31,221,30,205,31,111,31,238,31,238,30,187,31,187,30,28,31,28,30,13,31,13,30,131,31,58,31,235,31,235,30,42,31,42,30,157,31,157,30,32,31,32,30,4,31,214,31,208,31,251,31,120,31,154,31,154,30,154,29,159,31,48,31,67,31,187,31,81,31,53,31,57,31,117,31,44,31,231,31,231,30,166,31,166,30,166,29,114,31,244,31,242,31,7,31,160,31,160,30,179,31,195,31,150,31,20,31,20,30,136,31,180,31,186,31,199,31,74,31,111,31,74,31,218,31,218,30,197,31,43,31,238,31,238,30,144,31,153,31,153,30,105,31,105,30,105,29,237,31,129,31,190,31,20,31,85,31,236,31,218,31,218,30,44,31,44,30,80,31,219,31,238,31,47,31,137,31,156,31,215,31,153,31,153,30,27,31,218,31,78,31,134,31,29,31,231,31,231,30,237,31,67,31,47,31,205,31,153,31,186,31,5,31,252,31,217,31,49,31,146,31,221,31,167,31,148,31,252,31,95,31,235,31,240,31,240,30,166,31,190,31,201,31,23,31,217,31,217,30,227,31,202,31,105,31,15,31,90,31,129,31,245,31,1,31,69,31,69,30,96,31,96,30,96,29,3,31,252,31,198,31,85,31,85,30,113,31,38,31,223,31,32,31,219,31,219,30,18,31,18,30,103,31,201,31,35,31,35,31,76,31,149,31,139,31,207,31,193,31,144,31,144,30,144,29,92,31,94,31,211,31,197,31,47,31,47,30,236,31,102,31,206,31,8,31,34,31,163,31,163,30,45,31,61,31,51,31,251,31,251,30,251,29,245,31,137,31,225,31,149,31,107,31,238,31,41,31,203,31,141,31,67,31,73,31,52,31,67,31,72,31,72,30,4,31,60,31,106,31,60,31,46,31,138,31,29,31,82,31,82,30,251,31,138,31,209,31,152,31,138,31,156,31,156,30,178,31,169,31,169,30,203,31,237,31,237,30,109,31,234,31,234,30,81,31,26,31,235,31,61,31,246,31,155,31,171,31,94,31,94,30,94,29,29,31,19,31,247,31,210,31,210,30,234,31,234,30,155,31,160,31,126,31,181,31,181,30,149,31,182,31,182,30,182,29,6,31,76,31,39,31,49,31,110,31,110,30,2,31,120,31,120,30,120,29,66,31,183,31,148,31,248,31,248,30,248,29,249,31,48,31,44,31,24,31,193,31,202,31,73,31,198,31,180,31,60,31,191,31,75,31,77,31,213,31,180,31,206,31,2,31,203,31,246,31,85,31,85,30,228,31,101,31,136,31,84,31,248,31,248,30,6,31,130,31,188,31,252,31,252,30,66,31,66,30,132,31,94,31,55,31,198,31,52,31,138,31,138,30,131,31,141,31,141,31,141,30,119,31,119,30,187,31,28,31,244,31,74,31,55,31,208,31,178,31,178,30,223,31,46,31,196,31,196,30,124,31,139,31,5,31,13,31,13,30,226,31,149,31,64,31,78,31,66,31,12,31,12,30,12,29,245,31,7,31,47,31,80,31,220,31,38,31,38,30,184,31,171,31,124,31,169,31,190,31,190,30,190,29,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
