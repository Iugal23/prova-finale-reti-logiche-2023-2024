-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 783;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,215,0,0,0,0,0,83,0,216,0,10,0,126,0,160,0,104,0,91,0,71,0,98,0,0,0,222,0,0,0,102,0,233,0,72,0,225,0,0,0,42,0,30,0,207,0,12,0,202,0,163,0,185,0,171,0,47,0,27,0,159,0,0,0,0,0,131,0,25,0,77,0,108,0,36,0,41,0,0,0,53,0,233,0,55,0,86,0,62,0,0,0,174,0,33,0,87,0,159,0,26,0,94,0,180,0,116,0,0,0,44,0,172,0,99,0,0,0,157,0,204,0,99,0,80,0,120,0,184,0,214,0,205,0,0,0,158,0,0,0,147,0,115,0,207,0,146,0,157,0,0,0,6,0,193,0,122,0,72,0,243,0,179,0,235,0,245,0,133,0,51,0,158,0,0,0,39,0,7,0,143,0,0,0,0,0,0,0,114,0,0,0,0,0,0,0,0,0,7,0,248,0,144,0,0,0,248,0,234,0,202,0,139,0,0,0,57,0,190,0,246,0,165,0,233,0,0,0,56,0,0,0,136,0,0,0,80,0,60,0,107,0,76,0,217,0,160,0,126,0,119,0,211,0,38,0,255,0,183,0,0,0,0,0,250,0,138,0,117,0,218,0,39,0,206,0,152,0,16,0,60,0,235,0,25,0,131,0,0,0,25,0,166,0,0,0,94,0,184,0,16,0,128,0,244,0,0,0,0,0,39,0,53,0,18,0,74,0,28,0,217,0,93,0,50,0,218,0,6,0,174,0,36,0,119,0,147,0,0,0,56,0,68,0,247,0,155,0,209,0,76,0,208,0,212,0,0,0,93,0,136,0,0,0,0,0,48,0,251,0,0,0,120,0,116,0,5,0,0,0,239,0,0,0,183,0,204,0,1,0,118,0,0,0,0,0,0,0,24,0,78,0,28,0,90,0,126,0,70,0,0,0,221,0,236,0,190,0,74,0,68,0,0,0,221,0,128,0,86,0,0,0,58,0,125,0,187,0,0,0,145,0,0,0,135,0,40,0,0,0,219,0,255,0,116,0,131,0,0,0,98,0,0,0,17,0,16,0,4,0,235,0,0,0,0,0,0,0,139,0,0,0,35,0,222,0,60,0,11,0,0,0,0,0,23,0,135,0,249,0,63,0,0,0,0,0,74,0,0,0,101,0,0,0,0,0,230,0,51,0,231,0,7,0,0,0,0,0,18,0,27,0,0,0,105,0,0,0,144,0,249,0,211,0,0,0,89,0,212,0,162,0,173,0,242,0,156,0,15,0,156,0,0,0,217,0,0,0,169,0,168,0,235,0,0,0,47,0,85,0,242,0,72,0,207,0,145,0,77,0,156,0,148,0,136,0,121,0,160,0,0,0,198,0,148,0,214,0,139,0,0,0,0,0,116,0,62,0,42,0,182,0,106,0,0,0,0,0,0,0,154,0,40,0,0,0,100,0,213,0,170,0,66,0,153,0,165,0,65,0,25,0,103,0,142,0,173,0,148,0,105,0,233,0,255,0,158,0,76,0,120,0,46,0,205,0,253,0,2,0,0,0,116,0,249,0,115,0,0,0,32,0,17,0,227,0,0,0,170,0,233,0,96,0,200,0,88,0,140,0,169,0,90,0,14,0,250,0,168,0,158,0,26,0,32,0,0,0,234,0,183,0,159,0,0,0,0,0,0,0,0,0,0,0,0,0,189,0,114,0,147,0,34,0,134,0,12,0,231,0,220,0,201,0,29,0,38,0,84,0,21,0,206,0,56,0,210,0,129,0,218,0,156,0,16,0,130,0,14,0,17,0,210,0,89,0,145,0,0,0,79,0,0,0,72,0,6,0,137,0,158,0,28,0,241,0,213,0,53,0,67,0,139,0,31,0,112,0,155,0,0,0,0,0,168,0,136,0,0,0,7,0,78,0,0,0,95,0,230,0,143,0,228,0,107,0,0,0,26,0,41,0,0,0,23,0,133,0,246,0,18,0,202,0,182,0,235,0,85,0,160,0,65,0,0,0,139,0,108,0,101,0,0,0,202,0,185,0,234,0,14,0,0,0,74,0,75,0,0,0,99,0,153,0,198,0,165,0,1,0,109,0,230,0,182,0,135,0,69,0,215,0,244,0,170,0,190,0,89,0,21,0,33,0,0,0,164,0,155,0,74,0,170,0,0,0,168,0,53,0,0,0,244,0,13,0,50,0,68,0,140,0,0,0,95,0,95,0,159,0,126,0,233,0,0,0,4,0,203,0,136,0,88,0,44,0,154,0,133,0,230,0,186,0,0,0,42,0,141,0,0,0,96,0,29,0,2,0,0,0,166,0,0,0,0,0,0,0,0,0,28,0,0,0,22,0,229,0,101,0,158,0,63,0,89,0,89,0,189,0,157,0,237,0,235,0,13,0,26,0,0,0,186,0,8,0,163,0,81,0,100,0,30,0,144,0,0,0,56,0,102,0,208,0,225,0,28,0,83,0,0,0,116,0,88,0,106,0,77,0,235,0,73,0,245,0,2,0,153,0,219,0,165,0,76,0,245,0,0,0,143,0,42,0,0,0,101,0,172,0,254,0,115,0,0,0,103,0,216,0,78,0,35,0,245,0,0,0,127,0,0,0,40,0,102,0,168,0,244,0,72,0,111,0,0,0,179,0,207,0,0,0,159,0,0,0,0,0,238,0,180,0,57,0,146,0,191,0,172,0,115,0,8,0,64,0,0,0,18,0,212,0,1,0,72,0,85,0,226,0,0,0,0,0,245,0,129,0,112,0,4,0,31,0,108,0,84,0,131,0,247,0,223,0,84,0,187,0,215,0,105,0,156,0,152,0,179,0,0,0,35,0,90,0,159,0,0,0,19,0,208,0,184,0,201,0,236,0,0,0,249,0,0,0,215,0,0,0,132,0,34,0,228,0,173,0,0,0,0,0,160,0,135,0,162,0,41,0,0,0,0,0,219,0,73,0,0,0,235,0,54,0,166,0,164,0,135,0,0,0,100,0,162,0,209,0,0,0,203,0,26,0,163,0,0,0,6,0,78,0,178,0,154,0,0,0,246,0,163,0,218,0,162,0,94,0,0,0,141,0,91,0,143,0,38,0,155,0,113,0,23,0,0,0,110,0,46,0,156,0,22,0,0,0,8,0,146,0,0,0,123,0,0,0,221,0,0,0,0,0,197,0,42,0,168,0,0,0,156,0,7,0,104,0,8,0,83,0,224,0,0,0,41,0,72,0,177,0,0,0,69,0,120,0,232,0,155,0,0,0,49,0,0,0,109,0,173,0,236,0,0,0,7,0,181,0,114,0,74,0,207,0,244,0,134,0,107,0,206,0,87,0,97,0,242,0,30,0,212,0,192,0,223,0,183,0,0,0,0,0,165,0,0,0,0,0,101,0,0,0,99,0,0,0,85,0,0,0,142,0,139,0,79,0,248,0,255,0,0,0,0,0,89,0,0,0,102,0,62,0,154,0,114,0,0,0,0,0,252,0,38,0,55,0,92,0,0,0,146,0,76,0,158,0,174,0,0,0,14,0,0,0,112,0);
signal scenario_full  : scenario_type := (0,0,215,31,215,30,215,29,83,31,216,31,10,31,126,31,160,31,104,31,91,31,71,31,98,31,98,30,222,31,222,30,102,31,233,31,72,31,225,31,225,30,42,31,30,31,207,31,12,31,202,31,163,31,185,31,171,31,47,31,27,31,159,31,159,30,159,29,131,31,25,31,77,31,108,31,36,31,41,31,41,30,53,31,233,31,55,31,86,31,62,31,62,30,174,31,33,31,87,31,159,31,26,31,94,31,180,31,116,31,116,30,44,31,172,31,99,31,99,30,157,31,204,31,99,31,80,31,120,31,184,31,214,31,205,31,205,30,158,31,158,30,147,31,115,31,207,31,146,31,157,31,157,30,6,31,193,31,122,31,72,31,243,31,179,31,235,31,245,31,133,31,51,31,158,31,158,30,39,31,7,31,143,31,143,30,143,29,143,28,114,31,114,30,114,29,114,28,114,27,7,31,248,31,144,31,144,30,248,31,234,31,202,31,139,31,139,30,57,31,190,31,246,31,165,31,233,31,233,30,56,31,56,30,136,31,136,30,80,31,60,31,107,31,76,31,217,31,160,31,126,31,119,31,211,31,38,31,255,31,183,31,183,30,183,29,250,31,138,31,117,31,218,31,39,31,206,31,152,31,16,31,60,31,235,31,25,31,131,31,131,30,25,31,166,31,166,30,94,31,184,31,16,31,128,31,244,31,244,30,244,29,39,31,53,31,18,31,74,31,28,31,217,31,93,31,50,31,218,31,6,31,174,31,36,31,119,31,147,31,147,30,56,31,68,31,247,31,155,31,209,31,76,31,208,31,212,31,212,30,93,31,136,31,136,30,136,29,48,31,251,31,251,30,120,31,116,31,5,31,5,30,239,31,239,30,183,31,204,31,1,31,118,31,118,30,118,29,118,28,24,31,78,31,28,31,90,31,126,31,70,31,70,30,221,31,236,31,190,31,74,31,68,31,68,30,221,31,128,31,86,31,86,30,58,31,125,31,187,31,187,30,145,31,145,30,135,31,40,31,40,30,219,31,255,31,116,31,131,31,131,30,98,31,98,30,17,31,16,31,4,31,235,31,235,30,235,29,235,28,139,31,139,30,35,31,222,31,60,31,11,31,11,30,11,29,23,31,135,31,249,31,63,31,63,30,63,29,74,31,74,30,101,31,101,30,101,29,230,31,51,31,231,31,7,31,7,30,7,29,18,31,27,31,27,30,105,31,105,30,144,31,249,31,211,31,211,30,89,31,212,31,162,31,173,31,242,31,156,31,15,31,156,31,156,30,217,31,217,30,169,31,168,31,235,31,235,30,47,31,85,31,242,31,72,31,207,31,145,31,77,31,156,31,148,31,136,31,121,31,160,31,160,30,198,31,148,31,214,31,139,31,139,30,139,29,116,31,62,31,42,31,182,31,106,31,106,30,106,29,106,28,154,31,40,31,40,30,100,31,213,31,170,31,66,31,153,31,165,31,65,31,25,31,103,31,142,31,173,31,148,31,105,31,233,31,255,31,158,31,76,31,120,31,46,31,205,31,253,31,2,31,2,30,116,31,249,31,115,31,115,30,32,31,17,31,227,31,227,30,170,31,233,31,96,31,200,31,88,31,140,31,169,31,90,31,14,31,250,31,168,31,158,31,26,31,32,31,32,30,234,31,183,31,159,31,159,30,159,29,159,28,159,27,159,26,159,25,189,31,114,31,147,31,34,31,134,31,12,31,231,31,220,31,201,31,29,31,38,31,84,31,21,31,206,31,56,31,210,31,129,31,218,31,156,31,16,31,130,31,14,31,17,31,210,31,89,31,145,31,145,30,79,31,79,30,72,31,6,31,137,31,158,31,28,31,241,31,213,31,53,31,67,31,139,31,31,31,112,31,155,31,155,30,155,29,168,31,136,31,136,30,7,31,78,31,78,30,95,31,230,31,143,31,228,31,107,31,107,30,26,31,41,31,41,30,23,31,133,31,246,31,18,31,202,31,182,31,235,31,85,31,160,31,65,31,65,30,139,31,108,31,101,31,101,30,202,31,185,31,234,31,14,31,14,30,74,31,75,31,75,30,99,31,153,31,198,31,165,31,1,31,109,31,230,31,182,31,135,31,69,31,215,31,244,31,170,31,190,31,89,31,21,31,33,31,33,30,164,31,155,31,74,31,170,31,170,30,168,31,53,31,53,30,244,31,13,31,50,31,68,31,140,31,140,30,95,31,95,31,159,31,126,31,233,31,233,30,4,31,203,31,136,31,88,31,44,31,154,31,133,31,230,31,186,31,186,30,42,31,141,31,141,30,96,31,29,31,2,31,2,30,166,31,166,30,166,29,166,28,166,27,28,31,28,30,22,31,229,31,101,31,158,31,63,31,89,31,89,31,189,31,157,31,237,31,235,31,13,31,26,31,26,30,186,31,8,31,163,31,81,31,100,31,30,31,144,31,144,30,56,31,102,31,208,31,225,31,28,31,83,31,83,30,116,31,88,31,106,31,77,31,235,31,73,31,245,31,2,31,153,31,219,31,165,31,76,31,245,31,245,30,143,31,42,31,42,30,101,31,172,31,254,31,115,31,115,30,103,31,216,31,78,31,35,31,245,31,245,30,127,31,127,30,40,31,102,31,168,31,244,31,72,31,111,31,111,30,179,31,207,31,207,30,159,31,159,30,159,29,238,31,180,31,57,31,146,31,191,31,172,31,115,31,8,31,64,31,64,30,18,31,212,31,1,31,72,31,85,31,226,31,226,30,226,29,245,31,129,31,112,31,4,31,31,31,108,31,84,31,131,31,247,31,223,31,84,31,187,31,215,31,105,31,156,31,152,31,179,31,179,30,35,31,90,31,159,31,159,30,19,31,208,31,184,31,201,31,236,31,236,30,249,31,249,30,215,31,215,30,132,31,34,31,228,31,173,31,173,30,173,29,160,31,135,31,162,31,41,31,41,30,41,29,219,31,73,31,73,30,235,31,54,31,166,31,164,31,135,31,135,30,100,31,162,31,209,31,209,30,203,31,26,31,163,31,163,30,6,31,78,31,178,31,154,31,154,30,246,31,163,31,218,31,162,31,94,31,94,30,141,31,91,31,143,31,38,31,155,31,113,31,23,31,23,30,110,31,46,31,156,31,22,31,22,30,8,31,146,31,146,30,123,31,123,30,221,31,221,30,221,29,197,31,42,31,168,31,168,30,156,31,7,31,104,31,8,31,83,31,224,31,224,30,41,31,72,31,177,31,177,30,69,31,120,31,232,31,155,31,155,30,49,31,49,30,109,31,173,31,236,31,236,30,7,31,181,31,114,31,74,31,207,31,244,31,134,31,107,31,206,31,87,31,97,31,242,31,30,31,212,31,192,31,223,31,183,31,183,30,183,29,165,31,165,30,165,29,101,31,101,30,99,31,99,30,85,31,85,30,142,31,139,31,79,31,248,31,255,31,255,30,255,29,89,31,89,30,102,31,62,31,154,31,114,31,114,30,114,29,252,31,38,31,55,31,92,31,92,30,146,31,76,31,158,31,174,31,174,30,14,31,14,30,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
