-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 875;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (72,0,38,0,0,0,206,0,160,0,56,0,0,0,9,0,255,0,174,0,0,0,147,0,121,0,50,0,203,0,106,0,200,0,0,0,0,0,42,0,180,0,59,0,27,0,55,0,125,0,30,0,0,0,0,0,3,0,55,0,71,0,0,0,192,0,0,0,200,0,145,0,0,0,62,0,130,0,240,0,74,0,169,0,202,0,212,0,37,0,178,0,162,0,120,0,71,0,116,0,47,0,0,0,0,0,217,0,113,0,207,0,175,0,214,0,17,0,49,0,27,0,139,0,184,0,137,0,31,0,0,0,218,0,109,0,0,0,176,0,114,0,199,0,165,0,70,0,135,0,67,0,177,0,228,0,0,0,180,0,252,0,170,0,0,0,27,0,21,0,0,0,178,0,11,0,238,0,83,0,142,0,103,0,47,0,167,0,159,0,113,0,0,0,101,0,251,0,226,0,0,0,0,0,28,0,74,0,196,0,25,0,219,0,10,0,123,0,149,0,0,0,130,0,25,0,103,0,198,0,89,0,2,0,56,0,221,0,196,0,72,0,241,0,241,0,0,0,63,0,218,0,0,0,85,0,0,0,36,0,188,0,154,0,0,0,134,0,116,0,93,0,188,0,178,0,62,0,249,0,97,0,0,0,0,0,47,0,143,0,0,0,30,0,178,0,65,0,0,0,66,0,37,0,192,0,46,0,35,0,109,0,123,0,87,0,238,0,22,0,139,0,97,0,0,0,110,0,0,0,101,0,199,0,183,0,0,0,237,0,245,0,206,0,129,0,161,0,0,0,187,0,0,0,7,0,111,0,136,0,28,0,162,0,35,0,218,0,73,0,0,0,0,0,214,0,49,0,32,0,251,0,136,0,0,0,234,0,214,0,226,0,175,0,0,0,169,0,95,0,134,0,233,0,69,0,176,0,46,0,67,0,64,0,139,0,221,0,145,0,0,0,19,0,7,0,244,0,14,0,47,0,82,0,128,0,99,0,245,0,163,0,0,0,239,0,96,0,215,0,0,0,233,0,0,0,0,0,0,0,37,0,0,0,0,0,58,0,160,0,73,0,28,0,0,0,0,0,0,0,60,0,103,0,127,0,47,0,33,0,37,0,0,0,123,0,74,0,0,0,0,0,2,0,0,0,0,0,210,0,112,0,125,0,129,0,206,0,78,0,82,0,224,0,81,0,0,0,110,0,162,0,171,0,0,0,161,0,63,0,55,0,0,0,242,0,0,0,221,0,181,0,155,0,0,0,254,0,223,0,110,0,70,0,144,0,10,0,133,0,124,0,207,0,8,0,22,0,0,0,15,0,200,0,157,0,252,0,0,0,62,0,49,0,109,0,238,0,189,0,0,0,46,0,73,0,129,0,228,0,0,0,0,0,0,0,0,0,23,0,165,0,173,0,12,0,107,0,41,0,87,0,177,0,56,0,7,0,47,0,131,0,0,0,91,0,201,0,163,0,242,0,134,0,0,0,182,0,181,0,27,0,220,0,161,0,0,0,195,0,70,0,237,0,211,0,0,0,0,0,203,0,77,0,63,0,218,0,64,0,211,0,131,0,187,0,0,0,142,0,231,0,198,0,95,0,39,0,76,0,0,0,230,0,50,0,187,0,115,0,0,0,175,0,154,0,0,0,12,0,77,0,0,0,89,0,47,0,0,0,0,0,66,0,28,0,81,0,213,0,0,0,0,0,8,0,65,0,127,0,172,0,0,0,138,0,105,0,45,0,0,0,90,0,0,0,98,0,245,0,249,0,53,0,50,0,76,0,18,0,98,0,170,0,0,0,177,0,220,0,51,0,88,0,46,0,141,0,97,0,69,0,68,0,19,0,70,0,6,0,11,0,88,0,15,0,162,0,119,0,1,0,0,0,0,0,236,0,152,0,0,0,111,0,63,0,199,0,250,0,226,0,156,0,0,0,0,0,0,0,200,0,40,0,0,0,206,0,208,0,238,0,5,0,154,0,251,0,221,0,0,0,0,0,172,0,0,0,104,0,141,0,0,0,0,0,0,0,58,0,0,0,42,0,75,0,0,0,51,0,89,0,186,0,141,0,36,0,226,0,72,0,117,0,120,0,206,0,180,0,3,0,46,0,99,0,0,0,145,0,185,0,59,0,137,0,0,0,195,0,45,0,31,0,236,0,146,0,136,0,249,0,161,0,212,0,234,0,247,0,220,0,0,0,11,0,0,0,137,0,0,0,3,0,117,0,0,0,102,0,233,0,224,0,170,0,181,0,0,0,6,0,239,0,42,0,115,0,0,0,50,0,0,0,245,0,146,0,166,0,73,0,182,0,20,0,0,0,0,0,43,0,213,0,109,0,47,0,56,0,55,0,56,0,108,0,32,0,0,0,0,0,0,0,0,0,0,0,45,0,224,0,0,0,241,0,9,0,245,0,96,0,120,0,235,0,0,0,78,0,118,0,40,0,250,0,118,0,51,0,215,0,43,0,0,0,124,0,141,0,246,0,169,0,118,0,25,0,87,0,32,0,139,0,146,0,84,0,132,0,126,0,199,0,215,0,0,0,58,0,14,0,0,0,45,0,0,0,199,0,226,0,168,0,0,0,192,0,21,0,229,0,179,0,88,0,237,0,49,0,196,0,222,0,60,0,211,0,0,0,144,0,188,0,0,0,45,0,126,0,76,0,50,0,178,0,32,0,0,0,124,0,133,0,174,0,0,0,138,0,0,0,168,0,0,0,246,0,100,0,185,0,0,0,186,0,166,0,157,0,221,0,189,0,133,0,54,0,0,0,153,0,114,0,0,0,192,0,104,0,178,0,227,0,3,0,172,0,49,0,155,0,60,0,0,0,99,0,135,0,24,0,171,0,0,0,40,0,38,0,0,0,12,0,110,0,34,0,0,0,110,0,103,0,205,0,138,0,200,0,248,0,174,0,234,0,116,0,0,0,132,0,0,0,231,0,52,0,0,0,0,0,182,0,243,0,216,0,10,0,190,0,10,0,25,0,160,0,81,0,96,0,146,0,246,0,0,0,208,0,185,0,192,0,17,0,178,0,118,0,0,0,77,0,0,0,0,0,62,0,0,0,17,0,214,0,41,0,216,0,0,0,8,0,243,0,30,0,0,0,154,0,84,0,124,0,0,0,144,0,85,0,133,0,33,0,64,0,110,0,69,0,82,0,48,0,197,0,235,0,186,0,6,0,20,0,24,0,0,0,254,0,97,0,129,0,78,0,207,0,0,0,177,0,210,0,3,0,165,0,166,0,142,0,129,0,167,0,97,0,0,0,0,0,69,0,0,0,37,0,146,0,95,0,0,0,15,0,168,0,211,0,0,0,145,0,244,0,77,0,130,0,0,0,231,0,255,0,150,0,209,0,203,0,0,0,0,0,123,0,250,0,248,0,213,0,114,0,9,0,1,0,0,0,125,0,142,0,1,0,80,0,0,0,159,0,0,0,141,0,111,0,228,0,196,0,169,0,94,0,103,0,23,0,138,0,0,0,6,0,0,0,238,0,14,0,22,0,133,0,13,0,112,0,169,0,2,0,0,0,225,0,0,0,0,0,117,0,2,0,0,0,0,0,36,0,255,0,0,0,12,0,205,0,190,0,176,0,98,0,0,0,159,0,240,0,134,0,66,0,29,0,193,0,241,0,163,0,148,0,166,0,45,0,86,0,48,0,0,0,21,0,205,0,0,0,10,0,69,0,177,0,150,0,227,0,0,0,7,0,0,0,0,0,207,0,0,0,0,0,5,0,52,0,70,0,0,0,149,0,0,0,75,0,186,0,185,0,24,0,0,0,224,0,0,0,20,0,27,0,45,0,207,0,10,0,202,0,254,0,0,0,51,0,0,0,29,0,73,0,252,0,89,0,89,0,0,0,113,0,0,0,0,0,0,0,0,0,40,0,45,0,157,0,0,0,2,0,13,0,241,0,0,0,57,0,197,0,126,0);
signal scenario_full  : scenario_type := (72,31,38,31,38,30,206,31,160,31,56,31,56,30,9,31,255,31,174,31,174,30,147,31,121,31,50,31,203,31,106,31,200,31,200,30,200,29,42,31,180,31,59,31,27,31,55,31,125,31,30,31,30,30,30,29,3,31,55,31,71,31,71,30,192,31,192,30,200,31,145,31,145,30,62,31,130,31,240,31,74,31,169,31,202,31,212,31,37,31,178,31,162,31,120,31,71,31,116,31,47,31,47,30,47,29,217,31,113,31,207,31,175,31,214,31,17,31,49,31,27,31,139,31,184,31,137,31,31,31,31,30,218,31,109,31,109,30,176,31,114,31,199,31,165,31,70,31,135,31,67,31,177,31,228,31,228,30,180,31,252,31,170,31,170,30,27,31,21,31,21,30,178,31,11,31,238,31,83,31,142,31,103,31,47,31,167,31,159,31,113,31,113,30,101,31,251,31,226,31,226,30,226,29,28,31,74,31,196,31,25,31,219,31,10,31,123,31,149,31,149,30,130,31,25,31,103,31,198,31,89,31,2,31,56,31,221,31,196,31,72,31,241,31,241,31,241,30,63,31,218,31,218,30,85,31,85,30,36,31,188,31,154,31,154,30,134,31,116,31,93,31,188,31,178,31,62,31,249,31,97,31,97,30,97,29,47,31,143,31,143,30,30,31,178,31,65,31,65,30,66,31,37,31,192,31,46,31,35,31,109,31,123,31,87,31,238,31,22,31,139,31,97,31,97,30,110,31,110,30,101,31,199,31,183,31,183,30,237,31,245,31,206,31,129,31,161,31,161,30,187,31,187,30,7,31,111,31,136,31,28,31,162,31,35,31,218,31,73,31,73,30,73,29,214,31,49,31,32,31,251,31,136,31,136,30,234,31,214,31,226,31,175,31,175,30,169,31,95,31,134,31,233,31,69,31,176,31,46,31,67,31,64,31,139,31,221,31,145,31,145,30,19,31,7,31,244,31,14,31,47,31,82,31,128,31,99,31,245,31,163,31,163,30,239,31,96,31,215,31,215,30,233,31,233,30,233,29,233,28,37,31,37,30,37,29,58,31,160,31,73,31,28,31,28,30,28,29,28,28,60,31,103,31,127,31,47,31,33,31,37,31,37,30,123,31,74,31,74,30,74,29,2,31,2,30,2,29,210,31,112,31,125,31,129,31,206,31,78,31,82,31,224,31,81,31,81,30,110,31,162,31,171,31,171,30,161,31,63,31,55,31,55,30,242,31,242,30,221,31,181,31,155,31,155,30,254,31,223,31,110,31,70,31,144,31,10,31,133,31,124,31,207,31,8,31,22,31,22,30,15,31,200,31,157,31,252,31,252,30,62,31,49,31,109,31,238,31,189,31,189,30,46,31,73,31,129,31,228,31,228,30,228,29,228,28,228,27,23,31,165,31,173,31,12,31,107,31,41,31,87,31,177,31,56,31,7,31,47,31,131,31,131,30,91,31,201,31,163,31,242,31,134,31,134,30,182,31,181,31,27,31,220,31,161,31,161,30,195,31,70,31,237,31,211,31,211,30,211,29,203,31,77,31,63,31,218,31,64,31,211,31,131,31,187,31,187,30,142,31,231,31,198,31,95,31,39,31,76,31,76,30,230,31,50,31,187,31,115,31,115,30,175,31,154,31,154,30,12,31,77,31,77,30,89,31,47,31,47,30,47,29,66,31,28,31,81,31,213,31,213,30,213,29,8,31,65,31,127,31,172,31,172,30,138,31,105,31,45,31,45,30,90,31,90,30,98,31,245,31,249,31,53,31,50,31,76,31,18,31,98,31,170,31,170,30,177,31,220,31,51,31,88,31,46,31,141,31,97,31,69,31,68,31,19,31,70,31,6,31,11,31,88,31,15,31,162,31,119,31,1,31,1,30,1,29,236,31,152,31,152,30,111,31,63,31,199,31,250,31,226,31,156,31,156,30,156,29,156,28,200,31,40,31,40,30,206,31,208,31,238,31,5,31,154,31,251,31,221,31,221,30,221,29,172,31,172,30,104,31,141,31,141,30,141,29,141,28,58,31,58,30,42,31,75,31,75,30,51,31,89,31,186,31,141,31,36,31,226,31,72,31,117,31,120,31,206,31,180,31,3,31,46,31,99,31,99,30,145,31,185,31,59,31,137,31,137,30,195,31,45,31,31,31,236,31,146,31,136,31,249,31,161,31,212,31,234,31,247,31,220,31,220,30,11,31,11,30,137,31,137,30,3,31,117,31,117,30,102,31,233,31,224,31,170,31,181,31,181,30,6,31,239,31,42,31,115,31,115,30,50,31,50,30,245,31,146,31,166,31,73,31,182,31,20,31,20,30,20,29,43,31,213,31,109,31,47,31,56,31,55,31,56,31,108,31,32,31,32,30,32,29,32,28,32,27,32,26,45,31,224,31,224,30,241,31,9,31,245,31,96,31,120,31,235,31,235,30,78,31,118,31,40,31,250,31,118,31,51,31,215,31,43,31,43,30,124,31,141,31,246,31,169,31,118,31,25,31,87,31,32,31,139,31,146,31,84,31,132,31,126,31,199,31,215,31,215,30,58,31,14,31,14,30,45,31,45,30,199,31,226,31,168,31,168,30,192,31,21,31,229,31,179,31,88,31,237,31,49,31,196,31,222,31,60,31,211,31,211,30,144,31,188,31,188,30,45,31,126,31,76,31,50,31,178,31,32,31,32,30,124,31,133,31,174,31,174,30,138,31,138,30,168,31,168,30,246,31,100,31,185,31,185,30,186,31,166,31,157,31,221,31,189,31,133,31,54,31,54,30,153,31,114,31,114,30,192,31,104,31,178,31,227,31,3,31,172,31,49,31,155,31,60,31,60,30,99,31,135,31,24,31,171,31,171,30,40,31,38,31,38,30,12,31,110,31,34,31,34,30,110,31,103,31,205,31,138,31,200,31,248,31,174,31,234,31,116,31,116,30,132,31,132,30,231,31,52,31,52,30,52,29,182,31,243,31,216,31,10,31,190,31,10,31,25,31,160,31,81,31,96,31,146,31,246,31,246,30,208,31,185,31,192,31,17,31,178,31,118,31,118,30,77,31,77,30,77,29,62,31,62,30,17,31,214,31,41,31,216,31,216,30,8,31,243,31,30,31,30,30,154,31,84,31,124,31,124,30,144,31,85,31,133,31,33,31,64,31,110,31,69,31,82,31,48,31,197,31,235,31,186,31,6,31,20,31,24,31,24,30,254,31,97,31,129,31,78,31,207,31,207,30,177,31,210,31,3,31,165,31,166,31,142,31,129,31,167,31,97,31,97,30,97,29,69,31,69,30,37,31,146,31,95,31,95,30,15,31,168,31,211,31,211,30,145,31,244,31,77,31,130,31,130,30,231,31,255,31,150,31,209,31,203,31,203,30,203,29,123,31,250,31,248,31,213,31,114,31,9,31,1,31,1,30,125,31,142,31,1,31,80,31,80,30,159,31,159,30,141,31,111,31,228,31,196,31,169,31,94,31,103,31,23,31,138,31,138,30,6,31,6,30,238,31,14,31,22,31,133,31,13,31,112,31,169,31,2,31,2,30,225,31,225,30,225,29,117,31,2,31,2,30,2,29,36,31,255,31,255,30,12,31,205,31,190,31,176,31,98,31,98,30,159,31,240,31,134,31,66,31,29,31,193,31,241,31,163,31,148,31,166,31,45,31,86,31,48,31,48,30,21,31,205,31,205,30,10,31,69,31,177,31,150,31,227,31,227,30,7,31,7,30,7,29,207,31,207,30,207,29,5,31,52,31,70,31,70,30,149,31,149,30,75,31,186,31,185,31,24,31,24,30,224,31,224,30,20,31,27,31,45,31,207,31,10,31,202,31,254,31,254,30,51,31,51,30,29,31,73,31,252,31,89,31,89,31,89,30,113,31,113,30,113,29,113,28,113,27,40,31,45,31,157,31,157,30,2,31,13,31,241,31,241,30,57,31,197,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
