-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_931 is
end project_tb_931;

architecture project_tb_arch_931 of project_tb_931 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 577;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (97,0,0,0,142,0,36,0,0,0,160,0,129,0,87,0,250,0,80,0,4,0,207,0,7,0,203,0,153,0,199,0,117,0,70,0,0,0,90,0,186,0,21,0,185,0,253,0,200,0,161,0,73,0,104,0,49,0,8,0,138,0,0,0,60,0,116,0,163,0,69,0,3,0,164,0,37,0,83,0,0,0,0,0,143,0,0,0,0,0,0,0,169,0,0,0,0,0,120,0,98,0,88,0,13,0,241,0,98,0,131,0,203,0,105,0,217,0,6,0,179,0,193,0,0,0,39,0,0,0,220,0,96,0,44,0,114,0,224,0,102,0,0,0,113,0,176,0,163,0,147,0,222,0,60,0,0,0,152,0,199,0,181,0,49,0,0,0,0,0,108,0,142,0,72,0,0,0,242,0,65,0,74,0,147,0,10,0,192,0,42,0,71,0,0,0,0,0,120,0,132,0,80,0,168,0,0,0,143,0,147,0,54,0,0,0,0,0,155,0,173,0,0,0,35,0,105,0,82,0,118,0,0,0,0,0,54,0,0,0,32,0,62,0,0,0,212,0,0,0,48,0,144,0,167,0,239,0,27,0,0,0,24,0,218,0,0,0,0,0,0,0,0,0,94,0,4,0,29,0,56,0,122,0,25,0,181,0,160,0,183,0,38,0,180,0,27,0,221,0,69,0,196,0,9,0,184,0,178,0,49,0,154,0,163,0,151,0,115,0,115,0,67,0,21,0,0,0,240,0,0,0,201,0,188,0,205,0,153,0,108,0,19,0,0,0,0,0,0,0,125,0,140,0,84,0,139,0,0,0,100,0,13,0,0,0,240,0,69,0,166,0,29,0,144,0,87,0,80,0,11,0,0,0,98,0,11,0,226,0,214,0,170,0,105,0,39,0,65,0,0,0,143,0,211,0,74,0,224,0,0,0,73,0,55,0,2,0,0,0,69,0,173,0,0,0,44,0,73,0,100,0,140,0,0,0,205,0,72,0,217,0,0,0,233,0,54,0,0,0,221,0,0,0,80,0,117,0,169,0,156,0,154,0,174,0,87,0,0,0,207,0,3,0,0,0,0,0,34,0,222,0,199,0,129,0,201,0,180,0,3,0,161,0,43,0,0,0,228,0,16,0,48,0,246,0,242,0,92,0,185,0,75,0,243,0,152,0,13,0,32,0,211,0,112,0,5,0,162,0,222,0,0,0,61,0,0,0,8,0,41,0,159,0,114,0,7,0,53,0,74,0,0,0,237,0,148,0,0,0,0,0,235,0,10,0,0,0,4,0,61,0,62,0,0,0,222,0,0,0,124,0,211,0,83,0,185,0,133,0,0,0,234,0,221,0,0,0,144,0,201,0,44,0,186,0,182,0,178,0,96,0,14,0,253,0,0,0,8,0,22,0,9,0,9,0,0,0,230,0,0,0,147,0,177,0,0,0,245,0,126,0,46,0,52,0,53,0,0,0,239,0,159,0,11,0,0,0,47,0,233,0,55,0,110,0,0,0,97,0,185,0,208,0,10,0,127,0,0,0,0,0,155,0,133,0,204,0,80,0,0,0,152,0,0,0,171,0,57,0,202,0,174,0,79,0,16,0,0,0,92,0,45,0,0,0,20,0,36,0,211,0,85,0,0,0,254,0,52,0,106,0,0,0,194,0,251,0,24,0,61,0,71,0,53,0,219,0,73,0,95,0,0,0,13,0,176,0,0,0,0,0,192,0,61,0,1,0,192,0,53,0,217,0,0,0,173,0,234,0,0,0,64,0,0,0,92,0,119,0,181,0,139,0,7,0,0,0,102,0,0,0,151,0,0,0,176,0,197,0,0,0,228,0,28,0,118,0,96,0,174,0,60,0,0,0,123,0,41,0,215,0,0,0,55,0,195,0,0,0,172,0,198,0,0,0,69,0,0,0,171,0,0,0,7,0,129,0,6,0,102,0,232,0,125,0,0,0,22,0,223,0,242,0,28,0,182,0,0,0,111,0,70,0,248,0,109,0,139,0,151,0,0,0,0,0,164,0,52,0,171,0,13,0,229,0,173,0,182,0,167,0,245,0,40,0,195,0,0,0,75,0,252,0,53,0,76,0,52,0,191,0,222,0,91,0,226,0,141,0,130,0,25,0,0,0,231,0,0,0,0,0,255,0,0,0,245,0,103,0,5,0,0,0,250,0,170,0,135,0,170,0,155,0,0,0,196,0,127,0,114,0,87,0,65,0,30,0,228,0,0,0,116,0,156,0,246,0,215,0,0,0,188,0,217,0,227,0,0,0,150,0,183,0,120,0,6,0,0,0,0,0,8,0,116,0,108,0,10,0,78,0,207,0,144,0,136,0,129,0,21,0,52,0,31,0,52,0,0,0,172,0,0,0,116,0,115,0,221,0,33,0,0,0,0,0,179,0,0,0,49,0,168,0,50,0,22,0,14,0,0,0,121,0,94,0,0,0,30,0,115,0,112,0,0,0,75,0,0,0,58,0,0,0,240,0,201,0,196,0,58,0,0,0,69,0,0,0,148,0,107,0,103,0,106,0,157,0,114,0,115,0,0,0,0,0,0,0,220,0,169,0,203,0,222,0,16,0,92,0,0,0,80,0);
signal scenario_full  : scenario_type := (97,31,97,30,142,31,36,31,36,30,160,31,129,31,87,31,250,31,80,31,4,31,207,31,7,31,203,31,153,31,199,31,117,31,70,31,70,30,90,31,186,31,21,31,185,31,253,31,200,31,161,31,73,31,104,31,49,31,8,31,138,31,138,30,60,31,116,31,163,31,69,31,3,31,164,31,37,31,83,31,83,30,83,29,143,31,143,30,143,29,143,28,169,31,169,30,169,29,120,31,98,31,88,31,13,31,241,31,98,31,131,31,203,31,105,31,217,31,6,31,179,31,193,31,193,30,39,31,39,30,220,31,96,31,44,31,114,31,224,31,102,31,102,30,113,31,176,31,163,31,147,31,222,31,60,31,60,30,152,31,199,31,181,31,49,31,49,30,49,29,108,31,142,31,72,31,72,30,242,31,65,31,74,31,147,31,10,31,192,31,42,31,71,31,71,30,71,29,120,31,132,31,80,31,168,31,168,30,143,31,147,31,54,31,54,30,54,29,155,31,173,31,173,30,35,31,105,31,82,31,118,31,118,30,118,29,54,31,54,30,32,31,62,31,62,30,212,31,212,30,48,31,144,31,167,31,239,31,27,31,27,30,24,31,218,31,218,30,218,29,218,28,218,27,94,31,4,31,29,31,56,31,122,31,25,31,181,31,160,31,183,31,38,31,180,31,27,31,221,31,69,31,196,31,9,31,184,31,178,31,49,31,154,31,163,31,151,31,115,31,115,31,67,31,21,31,21,30,240,31,240,30,201,31,188,31,205,31,153,31,108,31,19,31,19,30,19,29,19,28,125,31,140,31,84,31,139,31,139,30,100,31,13,31,13,30,240,31,69,31,166,31,29,31,144,31,87,31,80,31,11,31,11,30,98,31,11,31,226,31,214,31,170,31,105,31,39,31,65,31,65,30,143,31,211,31,74,31,224,31,224,30,73,31,55,31,2,31,2,30,69,31,173,31,173,30,44,31,73,31,100,31,140,31,140,30,205,31,72,31,217,31,217,30,233,31,54,31,54,30,221,31,221,30,80,31,117,31,169,31,156,31,154,31,174,31,87,31,87,30,207,31,3,31,3,30,3,29,34,31,222,31,199,31,129,31,201,31,180,31,3,31,161,31,43,31,43,30,228,31,16,31,48,31,246,31,242,31,92,31,185,31,75,31,243,31,152,31,13,31,32,31,211,31,112,31,5,31,162,31,222,31,222,30,61,31,61,30,8,31,41,31,159,31,114,31,7,31,53,31,74,31,74,30,237,31,148,31,148,30,148,29,235,31,10,31,10,30,4,31,61,31,62,31,62,30,222,31,222,30,124,31,211,31,83,31,185,31,133,31,133,30,234,31,221,31,221,30,144,31,201,31,44,31,186,31,182,31,178,31,96,31,14,31,253,31,253,30,8,31,22,31,9,31,9,31,9,30,230,31,230,30,147,31,177,31,177,30,245,31,126,31,46,31,52,31,53,31,53,30,239,31,159,31,11,31,11,30,47,31,233,31,55,31,110,31,110,30,97,31,185,31,208,31,10,31,127,31,127,30,127,29,155,31,133,31,204,31,80,31,80,30,152,31,152,30,171,31,57,31,202,31,174,31,79,31,16,31,16,30,92,31,45,31,45,30,20,31,36,31,211,31,85,31,85,30,254,31,52,31,106,31,106,30,194,31,251,31,24,31,61,31,71,31,53,31,219,31,73,31,95,31,95,30,13,31,176,31,176,30,176,29,192,31,61,31,1,31,192,31,53,31,217,31,217,30,173,31,234,31,234,30,64,31,64,30,92,31,119,31,181,31,139,31,7,31,7,30,102,31,102,30,151,31,151,30,176,31,197,31,197,30,228,31,28,31,118,31,96,31,174,31,60,31,60,30,123,31,41,31,215,31,215,30,55,31,195,31,195,30,172,31,198,31,198,30,69,31,69,30,171,31,171,30,7,31,129,31,6,31,102,31,232,31,125,31,125,30,22,31,223,31,242,31,28,31,182,31,182,30,111,31,70,31,248,31,109,31,139,31,151,31,151,30,151,29,164,31,52,31,171,31,13,31,229,31,173,31,182,31,167,31,245,31,40,31,195,31,195,30,75,31,252,31,53,31,76,31,52,31,191,31,222,31,91,31,226,31,141,31,130,31,25,31,25,30,231,31,231,30,231,29,255,31,255,30,245,31,103,31,5,31,5,30,250,31,170,31,135,31,170,31,155,31,155,30,196,31,127,31,114,31,87,31,65,31,30,31,228,31,228,30,116,31,156,31,246,31,215,31,215,30,188,31,217,31,227,31,227,30,150,31,183,31,120,31,6,31,6,30,6,29,8,31,116,31,108,31,10,31,78,31,207,31,144,31,136,31,129,31,21,31,52,31,31,31,52,31,52,30,172,31,172,30,116,31,115,31,221,31,33,31,33,30,33,29,179,31,179,30,49,31,168,31,50,31,22,31,14,31,14,30,121,31,94,31,94,30,30,31,115,31,112,31,112,30,75,31,75,30,58,31,58,30,240,31,201,31,196,31,58,31,58,30,69,31,69,30,148,31,107,31,103,31,106,31,157,31,114,31,115,31,115,30,115,29,115,28,220,31,169,31,203,31,222,31,16,31,92,31,92,30,80,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
