-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 760;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (151,0,12,0,103,0,0,0,0,0,168,0,66,0,61,0,206,0,184,0,242,0,0,0,0,0,134,0,61,0,174,0,27,0,6,0,0,0,60,0,132,0,145,0,45,0,173,0,115,0,7,0,36,0,20,0,42,0,37,0,110,0,103,0,169,0,238,0,0,0,0,0,139,0,181,0,68,0,178,0,198,0,147,0,128,0,170,0,184,0,106,0,64,0,92,0,47,0,29,0,0,0,40,0,194,0,2,0,0,0,18,0,69,0,0,0,100,0,118,0,174,0,148,0,17,0,246,0,112,0,76,0,142,0,235,0,72,0,231,0,201,0,222,0,0,0,224,0,210,0,84,0,43,0,145,0,154,0,112,0,123,0,251,0,0,0,37,0,75,0,230,0,100,0,236,0,96,0,124,0,230,0,148,0,0,0,0,0,231,0,30,0,146,0,0,0,0,0,68,0,0,0,0,0,241,0,214,0,45,0,101,0,165,0,68,0,75,0,198,0,164,0,0,0,0,0,50,0,238,0,242,0,40,0,0,0,52,0,0,0,128,0,26,0,0,0,71,0,0,0,22,0,138,0,0,0,47,0,76,0,48,0,0,0,97,0,226,0,174,0,8,0,47,0,75,0,0,0,0,0,222,0,0,0,207,0,137,0,193,0,135,0,0,0,105,0,53,0,174,0,0,0,0,0,174,0,111,0,195,0,49,0,35,0,108,0,100,0,61,0,213,0,84,0,45,0,162,0,186,0,0,0,11,0,10,0,35,0,18,0,148,0,128,0,205,0,32,0,0,0,183,0,88,0,95,0,85,0,205,0,118,0,0,0,210,0,242,0,13,0,51,0,0,0,38,0,0,0,0,0,0,0,0,0,105,0,76,0,202,0,134,0,14,0,143,0,207,0,161,0,0,0,0,0,69,0,91,0,0,0,195,0,96,0,121,0,166,0,118,0,150,0,3,0,82,0,86,0,209,0,22,0,29,0,109,0,0,0,17,0,44,0,45,0,0,0,14,0,154,0,176,0,116,0,41,0,104,0,135,0,75,0,154,0,0,0,225,0,0,0,0,0,32,0,169,0,235,0,0,0,118,0,251,0,45,0,49,0,131,0,88,0,145,0,0,0,12,0,124,0,188,0,108,0,0,0,0,0,50,0,0,0,0,0,196,0,0,0,131,0,190,0,2,0,195,0,0,0,0,0,116,0,35,0,115,0,43,0,80,0,234,0,0,0,80,0,0,0,156,0,78,0,0,0,233,0,157,0,134,0,0,0,88,0,0,0,189,0,23,0,124,0,27,0,232,0,140,0,104,0,43,0,94,0,0,0,123,0,158,0,90,0,103,0,0,0,216,0,125,0,111,0,168,0,116,0,207,0,84,0,230,0,161,0,41,0,17,0,0,0,145,0,0,0,187,0,88,0,127,0,104,0,0,0,178,0,77,0,179,0,6,0,26,0,31,0,211,0,211,0,206,0,71,0,72,0,237,0,0,0,0,0,0,0,31,0,0,0,67,0,57,0,5,0,53,0,212,0,233,0,253,0,0,0,6,0,0,0,169,0,76,0,83,0,0,0,0,0,23,0,0,0,0,0,0,0,0,0,0,0,197,0,206,0,234,0,43,0,174,0,1,0,58,0,225,0,79,0,149,0,102,0,78,0,138,0,115,0,183,0,0,0,5,0,0,0,227,0,37,0,0,0,0,0,0,0,0,0,80,0,0,0,150,0,41,0,218,0,0,0,3,0,178,0,0,0,115,0,237,0,20,0,130,0,75,0,67,0,124,0,117,0,0,0,16,0,0,0,214,0,12,0,0,0,182,0,241,0,62,0,172,0,26,0,56,0,59,0,128,0,112,0,239,0,131,0,113,0,171,0,0,0,3,0,224,0,56,0,176,0,0,0,194,0,137,0,0,0,21,0,76,0,126,0,39,0,108,0,145,0,161,0,0,0,66,0,144,0,0,0,132,0,86,0,253,0,0,0,0,0,198,0,0,0,0,0,179,0,56,0,172,0,244,0,157,0,209,0,8,0,253,0,220,0,154,0,135,0,132,0,9,0,0,0,37,0,121,0,27,0,169,0,0,0,185,0,111,0,89,0,0,0,169,0,0,0,138,0,86,0,0,0,0,0,16,0,206,0,105,0,158,0,0,0,35,0,71,0,222,0,219,0,83,0,60,0,0,0,244,0,91,0,249,0,59,0,246,0,189,0,0,0,67,0,197,0,147,0,135,0,132,0,0,0,0,0,0,0,170,0,59,0,151,0,167,0,36,0,0,0,189,0,106,0,205,0,167,0,174,0,27,0,193,0,243,0,158,0,21,0,91,0,1,0,0,0,0,0,0,0,0,0,200,0,32,0,114,0,0,0,243,0,34,0,0,0,77,0,76,0,27,0,0,0,26,0,0,0,0,0,66,0,237,0,48,0,0,0,90,0,7,0,139,0,112,0,19,0,245,0,44,0,245,0,127,0,166,0,194,0,33,0,116,0,0,0,238,0,0,0,0,0,0,0,237,0,96,0,172,0,243,0,105,0,157,0,124,0,33,0,219,0,115,0,160,0,192,0,0,0,108,0,228,0,0,0,119,0,161,0,138,0,122,0,230,0,0,0,43,0,85,0,0,0,205,0,180,0,0,0,64,0,0,0,49,0,96,0,75,0,149,0,0,0,5,0,248,0,139,0,0,0,35,0,191,0,0,0,0,0,6,0,136,0,164,0,221,0,144,0,0,0,102,0,166,0,140,0,82,0,149,0,15,0,0,0,82,0,177,0,110,0,126,0,30,0,150,0,0,0,45,0,32,0,171,0,68,0,235,0,210,0,201,0,117,0,220,0,200,0,0,0,205,0,0,0,43,0,141,0,58,0,37,0,0,0,57,0,121,0,103,0,141,0,63,0,96,0,20,0,193,0,206,0,172,0,0,0,123,0,206,0,87,0,142,0,40,0,204,0,65,0,0,0,80,0,230,0,152,0,80,0,26,0,0,0,0,0,170,0,0,0,0,0,42,0,0,0,193,0,166,0,250,0,0,0,147,0,0,0,227,0,102,0,42,0,27,0,118,0,0,0,65,0,196,0,244,0,44,0,93,0,0,0,146,0,63,0,68,0,113,0,89,0,78,0,81,0,16,0,42,0,57,0,190,0,118,0,127,0,180,0,209,0,94,0,55,0,245,0,99,0,167,0,53,0,97,0,98,0,0,0,0,0,75,0,34,0,250,0,0,0,153,0,214,0,114,0,171,0,211,0,75,0,0,0,156,0,203,0,114,0,79,0,118,0,223,0,0,0,82,0,0,0,156,0,62,0,41,0,210,0,128,0,117,0,0,0,120,0,138,0,21,0,80,0,158,0,31,0,0,0,28,0,102,0,0,0,145,0,254,0,18,0,50,0,29,0,160,0,0,0,164,0,99,0,184,0,85,0);
signal scenario_full  : scenario_type := (151,31,12,31,103,31,103,30,103,29,168,31,66,31,61,31,206,31,184,31,242,31,242,30,242,29,134,31,61,31,174,31,27,31,6,31,6,30,60,31,132,31,145,31,45,31,173,31,115,31,7,31,36,31,20,31,42,31,37,31,110,31,103,31,169,31,238,31,238,30,238,29,139,31,181,31,68,31,178,31,198,31,147,31,128,31,170,31,184,31,106,31,64,31,92,31,47,31,29,31,29,30,40,31,194,31,2,31,2,30,18,31,69,31,69,30,100,31,118,31,174,31,148,31,17,31,246,31,112,31,76,31,142,31,235,31,72,31,231,31,201,31,222,31,222,30,224,31,210,31,84,31,43,31,145,31,154,31,112,31,123,31,251,31,251,30,37,31,75,31,230,31,100,31,236,31,96,31,124,31,230,31,148,31,148,30,148,29,231,31,30,31,146,31,146,30,146,29,68,31,68,30,68,29,241,31,214,31,45,31,101,31,165,31,68,31,75,31,198,31,164,31,164,30,164,29,50,31,238,31,242,31,40,31,40,30,52,31,52,30,128,31,26,31,26,30,71,31,71,30,22,31,138,31,138,30,47,31,76,31,48,31,48,30,97,31,226,31,174,31,8,31,47,31,75,31,75,30,75,29,222,31,222,30,207,31,137,31,193,31,135,31,135,30,105,31,53,31,174,31,174,30,174,29,174,31,111,31,195,31,49,31,35,31,108,31,100,31,61,31,213,31,84,31,45,31,162,31,186,31,186,30,11,31,10,31,35,31,18,31,148,31,128,31,205,31,32,31,32,30,183,31,88,31,95,31,85,31,205,31,118,31,118,30,210,31,242,31,13,31,51,31,51,30,38,31,38,30,38,29,38,28,38,27,105,31,76,31,202,31,134,31,14,31,143,31,207,31,161,31,161,30,161,29,69,31,91,31,91,30,195,31,96,31,121,31,166,31,118,31,150,31,3,31,82,31,86,31,209,31,22,31,29,31,109,31,109,30,17,31,44,31,45,31,45,30,14,31,154,31,176,31,116,31,41,31,104,31,135,31,75,31,154,31,154,30,225,31,225,30,225,29,32,31,169,31,235,31,235,30,118,31,251,31,45,31,49,31,131,31,88,31,145,31,145,30,12,31,124,31,188,31,108,31,108,30,108,29,50,31,50,30,50,29,196,31,196,30,131,31,190,31,2,31,195,31,195,30,195,29,116,31,35,31,115,31,43,31,80,31,234,31,234,30,80,31,80,30,156,31,78,31,78,30,233,31,157,31,134,31,134,30,88,31,88,30,189,31,23,31,124,31,27,31,232,31,140,31,104,31,43,31,94,31,94,30,123,31,158,31,90,31,103,31,103,30,216,31,125,31,111,31,168,31,116,31,207,31,84,31,230,31,161,31,41,31,17,31,17,30,145,31,145,30,187,31,88,31,127,31,104,31,104,30,178,31,77,31,179,31,6,31,26,31,31,31,211,31,211,31,206,31,71,31,72,31,237,31,237,30,237,29,237,28,31,31,31,30,67,31,57,31,5,31,53,31,212,31,233,31,253,31,253,30,6,31,6,30,169,31,76,31,83,31,83,30,83,29,23,31,23,30,23,29,23,28,23,27,23,26,197,31,206,31,234,31,43,31,174,31,1,31,58,31,225,31,79,31,149,31,102,31,78,31,138,31,115,31,183,31,183,30,5,31,5,30,227,31,37,31,37,30,37,29,37,28,37,27,80,31,80,30,150,31,41,31,218,31,218,30,3,31,178,31,178,30,115,31,237,31,20,31,130,31,75,31,67,31,124,31,117,31,117,30,16,31,16,30,214,31,12,31,12,30,182,31,241,31,62,31,172,31,26,31,56,31,59,31,128,31,112,31,239,31,131,31,113,31,171,31,171,30,3,31,224,31,56,31,176,31,176,30,194,31,137,31,137,30,21,31,76,31,126,31,39,31,108,31,145,31,161,31,161,30,66,31,144,31,144,30,132,31,86,31,253,31,253,30,253,29,198,31,198,30,198,29,179,31,56,31,172,31,244,31,157,31,209,31,8,31,253,31,220,31,154,31,135,31,132,31,9,31,9,30,37,31,121,31,27,31,169,31,169,30,185,31,111,31,89,31,89,30,169,31,169,30,138,31,86,31,86,30,86,29,16,31,206,31,105,31,158,31,158,30,35,31,71,31,222,31,219,31,83,31,60,31,60,30,244,31,91,31,249,31,59,31,246,31,189,31,189,30,67,31,197,31,147,31,135,31,132,31,132,30,132,29,132,28,170,31,59,31,151,31,167,31,36,31,36,30,189,31,106,31,205,31,167,31,174,31,27,31,193,31,243,31,158,31,21,31,91,31,1,31,1,30,1,29,1,28,1,27,200,31,32,31,114,31,114,30,243,31,34,31,34,30,77,31,76,31,27,31,27,30,26,31,26,30,26,29,66,31,237,31,48,31,48,30,90,31,7,31,139,31,112,31,19,31,245,31,44,31,245,31,127,31,166,31,194,31,33,31,116,31,116,30,238,31,238,30,238,29,238,28,237,31,96,31,172,31,243,31,105,31,157,31,124,31,33,31,219,31,115,31,160,31,192,31,192,30,108,31,228,31,228,30,119,31,161,31,138,31,122,31,230,31,230,30,43,31,85,31,85,30,205,31,180,31,180,30,64,31,64,30,49,31,96,31,75,31,149,31,149,30,5,31,248,31,139,31,139,30,35,31,191,31,191,30,191,29,6,31,136,31,164,31,221,31,144,31,144,30,102,31,166,31,140,31,82,31,149,31,15,31,15,30,82,31,177,31,110,31,126,31,30,31,150,31,150,30,45,31,32,31,171,31,68,31,235,31,210,31,201,31,117,31,220,31,200,31,200,30,205,31,205,30,43,31,141,31,58,31,37,31,37,30,57,31,121,31,103,31,141,31,63,31,96,31,20,31,193,31,206,31,172,31,172,30,123,31,206,31,87,31,142,31,40,31,204,31,65,31,65,30,80,31,230,31,152,31,80,31,26,31,26,30,26,29,170,31,170,30,170,29,42,31,42,30,193,31,166,31,250,31,250,30,147,31,147,30,227,31,102,31,42,31,27,31,118,31,118,30,65,31,196,31,244,31,44,31,93,31,93,30,146,31,63,31,68,31,113,31,89,31,78,31,81,31,16,31,42,31,57,31,190,31,118,31,127,31,180,31,209,31,94,31,55,31,245,31,99,31,167,31,53,31,97,31,98,31,98,30,98,29,75,31,34,31,250,31,250,30,153,31,214,31,114,31,171,31,211,31,75,31,75,30,156,31,203,31,114,31,79,31,118,31,223,31,223,30,82,31,82,30,156,31,62,31,41,31,210,31,128,31,117,31,117,30,120,31,138,31,21,31,80,31,158,31,31,31,31,30,28,31,102,31,102,30,145,31,254,31,18,31,50,31,29,31,160,31,160,30,164,31,99,31,184,31,85,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
