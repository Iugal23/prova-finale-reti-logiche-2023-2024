-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 369;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,127,0,73,0,40,0,164,0,246,0,0,0,59,0,0,0,207,0,193,0,44,0,73,0,117,0,144,0,127,0,0,0,0,0,115,0,43,0,113,0,95,0,38,0,194,0,67,0,18,0,0,0,0,0,115,0,242,0,141,0,157,0,33,0,252,0,158,0,0,0,43,0,0,0,155,0,138,0,220,0,201,0,209,0,160,0,0,0,86,0,0,0,0,0,73,0,145,0,0,0,209,0,163,0,86,0,21,0,0,0,0,0,172,0,0,0,93,0,152,0,172,0,155,0,0,0,106,0,166,0,183,0,106,0,182,0,0,0,0,0,122,0,41,0,192,0,216,0,94,0,218,0,18,0,7,0,201,0,105,0,176,0,145,0,210,0,0,0,243,0,183,0,0,0,234,0,201,0,134,0,94,0,0,0,186,0,38,0,94,0,52,0,141,0,47,0,233,0,151,0,0,0,190,0,156,0,65,0,213,0,216,0,212,0,214,0,168,0,0,0,207,0,52,0,143,0,44,0,44,0,0,0,8,0,222,0,0,0,100,0,179,0,146,0,102,0,104,0,186,0,40,0,131,0,237,0,189,0,0,0,0,0,0,0,0,0,9,0,0,0,69,0,48,0,97,0,100,0,19,0,179,0,16,0,50,0,220,0,220,0,55,0,227,0,23,0,228,0,0,0,0,0,186,0,169,0,22,0,190,0,197,0,0,0,198,0,25,0,0,0,88,0,155,0,113,0,0,0,123,0,21,0,184,0,138,0,162,0,78,0,191,0,0,0,0,0,139,0,80,0,40,0,52,0,155,0,22,0,102,0,180,0,0,0,83,0,164,0,102,0,151,0,226,0,201,0,61,0,0,0,132,0,0,0,20,0,233,0,186,0,0,0,123,0,207,0,34,0,71,0,13,0,210,0,196,0,32,0,218,0,37,0,73,0,117,0,51,0,64,0,189,0,12,0,10,0,218,0,226,0,156,0,248,0,0,0,234,0,214,0,116,0,58,0,55,0,0,0,0,0,164,0,68,0,40,0,141,0,148,0,132,0,0,0,58,0,24,0,0,0,0,0,163,0,186,0,0,0,184,0,139,0,0,0,49,0,164,0,95,0,193,0,175,0,60,0,0,0,130,0,225,0,215,0,14,0,186,0,165,0,172,0,17,0,69,0,0,0,45,0,0,0,36,0,0,0,138,0,11,0,155,0,183,0,72,0,0,0,0,0,53,0,141,0,26,0,218,0,138,0,0,0,31,0,8,0,93,0,10,0,194,0,108,0,205,0,109,0,205,0,0,0,249,0,254,0,108,0,0,0,30,0,0,0,28,0,0,0,13,0,201,0,200,0,0,0,218,0,0,0,66,0,110,0,0,0,35,0,254,0,0,0,189,0,21,0,0,0,251,0,0,0,205,0,33,0,4,0,0,0,0,0,21,0,180,0,199,0,0,0,20,0,189,0,171,0,76,0,127,0,75,0,226,0,235,0,111,0,112,0,0,0,198,0,208,0,159,0,70,0,50,0,231,0,0,0,0,0,16,0,157,0,0,0,0,0,115,0,175,0,70,0,178,0,73,0,146,0,168,0,156,0,0,0,70,0,176,0,20,0,126,0,44,0,36,0,0,0,0,0,160,0,49,0,95,0,33,0,218,0,166,0,0,0,0,0);
signal scenario_full  : scenario_type := (1,31,127,31,73,31,40,31,164,31,246,31,246,30,59,31,59,30,207,31,193,31,44,31,73,31,117,31,144,31,127,31,127,30,127,29,115,31,43,31,113,31,95,31,38,31,194,31,67,31,18,31,18,30,18,29,115,31,242,31,141,31,157,31,33,31,252,31,158,31,158,30,43,31,43,30,155,31,138,31,220,31,201,31,209,31,160,31,160,30,86,31,86,30,86,29,73,31,145,31,145,30,209,31,163,31,86,31,21,31,21,30,21,29,172,31,172,30,93,31,152,31,172,31,155,31,155,30,106,31,166,31,183,31,106,31,182,31,182,30,182,29,122,31,41,31,192,31,216,31,94,31,218,31,18,31,7,31,201,31,105,31,176,31,145,31,210,31,210,30,243,31,183,31,183,30,234,31,201,31,134,31,94,31,94,30,186,31,38,31,94,31,52,31,141,31,47,31,233,31,151,31,151,30,190,31,156,31,65,31,213,31,216,31,212,31,214,31,168,31,168,30,207,31,52,31,143,31,44,31,44,31,44,30,8,31,222,31,222,30,100,31,179,31,146,31,102,31,104,31,186,31,40,31,131,31,237,31,189,31,189,30,189,29,189,28,189,27,9,31,9,30,69,31,48,31,97,31,100,31,19,31,179,31,16,31,50,31,220,31,220,31,55,31,227,31,23,31,228,31,228,30,228,29,186,31,169,31,22,31,190,31,197,31,197,30,198,31,25,31,25,30,88,31,155,31,113,31,113,30,123,31,21,31,184,31,138,31,162,31,78,31,191,31,191,30,191,29,139,31,80,31,40,31,52,31,155,31,22,31,102,31,180,31,180,30,83,31,164,31,102,31,151,31,226,31,201,31,61,31,61,30,132,31,132,30,20,31,233,31,186,31,186,30,123,31,207,31,34,31,71,31,13,31,210,31,196,31,32,31,218,31,37,31,73,31,117,31,51,31,64,31,189,31,12,31,10,31,218,31,226,31,156,31,248,31,248,30,234,31,214,31,116,31,58,31,55,31,55,30,55,29,164,31,68,31,40,31,141,31,148,31,132,31,132,30,58,31,24,31,24,30,24,29,163,31,186,31,186,30,184,31,139,31,139,30,49,31,164,31,95,31,193,31,175,31,60,31,60,30,130,31,225,31,215,31,14,31,186,31,165,31,172,31,17,31,69,31,69,30,45,31,45,30,36,31,36,30,138,31,11,31,155,31,183,31,72,31,72,30,72,29,53,31,141,31,26,31,218,31,138,31,138,30,31,31,8,31,93,31,10,31,194,31,108,31,205,31,109,31,205,31,205,30,249,31,254,31,108,31,108,30,30,31,30,30,28,31,28,30,13,31,201,31,200,31,200,30,218,31,218,30,66,31,110,31,110,30,35,31,254,31,254,30,189,31,21,31,21,30,251,31,251,30,205,31,33,31,4,31,4,30,4,29,21,31,180,31,199,31,199,30,20,31,189,31,171,31,76,31,127,31,75,31,226,31,235,31,111,31,112,31,112,30,198,31,208,31,159,31,70,31,50,31,231,31,231,30,231,29,16,31,157,31,157,30,157,29,115,31,175,31,70,31,178,31,73,31,146,31,168,31,156,31,156,30,70,31,176,31,20,31,126,31,44,31,36,31,36,30,36,29,160,31,49,31,95,31,33,31,218,31,166,31,166,30,166,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
