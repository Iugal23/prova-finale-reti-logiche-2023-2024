-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 662;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (113,0,0,0,211,0,99,0,68,0,161,0,119,0,113,0,41,0,4,0,107,0,120,0,116,0,13,0,27,0,166,0,210,0,0,0,65,0,0,0,193,0,140,0,81,0,225,0,149,0,251,0,0,0,47,0,0,0,95,0,76,0,244,0,6,0,0,0,216,0,95,0,93,0,237,0,218,0,127,0,0,0,89,0,12,0,55,0,93,0,67,0,43,0,77,0,79,0,164,0,12,0,130,0,18,0,155,0,19,0,3,0,120,0,155,0,49,0,164,0,191,0,215,0,0,0,0,0,163,0,205,0,191,0,43,0,190,0,0,0,253,0,205,0,66,0,231,0,215,0,15,0,163,0,161,0,110,0,144,0,0,0,26,0,204,0,30,0,0,0,53,0,104,0,222,0,106,0,105,0,0,0,176,0,147,0,21,0,105,0,83,0,116,0,117,0,237,0,177,0,190,0,136,0,0,0,36,0,109,0,195,0,225,0,50,0,0,0,93,0,7,0,104,0,0,0,173,0,25,0,251,0,0,0,244,0,0,0,117,0,0,0,243,0,0,0,119,0,249,0,31,0,240,0,185,0,0,0,130,0,32,0,0,0,182,0,228,0,0,0,170,0,165,0,67,0,244,0,13,0,99,0,210,0,87,0,112,0,0,0,2,0,167,0,224,0,248,0,144,0,152,0,136,0,11,0,237,0,97,0,150,0,0,0,194,0,0,0,238,0,143,0,244,0,157,0,142,0,136,0,117,0,26,0,34,0,110,0,0,0,113,0,208,0,251,0,6,0,0,0,241,0,87,0,45,0,217,0,164,0,229,0,1,0,0,0,0,0,226,0,164,0,0,0,114,0,0,0,135,0,47,0,90,0,71,0,0,0,144,0,149,0,190,0,230,0,58,0,226,0,197,0,23,0,78,0,0,0,223,0,61,0,40,0,210,0,212,0,196,0,205,0,26,0,166,0,103,0,2,0,218,0,253,0,250,0,0,0,142,0,139,0,0,0,88,0,1,0,238,0,254,0,0,0,149,0,218,0,39,0,183,0,0,0,0,0,0,0,66,0,11,0,0,0,247,0,215,0,35,0,226,0,161,0,30,0,67,0,0,0,0,0,225,0,177,0,167,0,186,0,104,0,248,0,217,0,176,0,0,0,231,0,109,0,111,0,190,0,95,0,164,0,91,0,250,0,129,0,66,0,81,0,0,0,31,0,198,0,0,0,160,0,177,0,99,0,66,0,51,0,22,0,97,0,170,0,235,0,127,0,34,0,157,0,219,0,149,0,248,0,137,0,0,0,172,0,79,0,16,0,246,0,208,0,253,0,173,0,101,0,173,0,241,0,24,0,175,0,128,0,211,0,128,0,221,0,242,0,0,0,208,0,228,0,143,0,25,0,86,0,214,0,198,0,81,0,223,0,231,0,120,0,226,0,157,0,187,0,55,0,150,0,190,0,179,0,41,0,12,0,209,0,0,0,18,0,0,0,3,0,178,0,207,0,123,0,233,0,37,0,42,0,106,0,175,0,14,0,198,0,91,0,139,0,69,0,135,0,131,0,90,0,0,0,148,0,197,0,60,0,115,0,59,0,167,0,93,0,244,0,235,0,201,0,218,0,80,0,116,0,194,0,8,0,89,0,10,0,0,0,129,0,173,0,69,0,18,0,75,0,220,0,133,0,68,0,146,0,60,0,82,0,0,0,197,0,68,0,43,0,45,0,95,0,228,0,65,0,92,0,0,0,223,0,41,0,2,0,238,0,0,0,0,0,0,0,10,0,108,0,13,0,183,0,250,0,171,0,0,0,112,0,0,0,249,0,19,0,86,0,76,0,253,0,0,0,231,0,18,0,183,0,76,0,190,0,0,0,162,0,0,0,20,0,0,0,0,0,231,0,23,0,40,0,157,0,141,0,54,0,72,0,59,0,97,0,150,0,227,0,15,0,0,0,17,0,0,0,141,0,172,0,0,0,44,0,82,0,241,0,133,0,167,0,61,0,143,0,56,0,171,0,76,0,70,0,167,0,238,0,90,0,0,0,183,0,0,0,20,0,177,0,117,0,92,0,64,0,87,0,152,0,91,0,254,0,0,0,243,0,98,0,58,0,132,0,0,0,101,0,73,0,161,0,172,0,128,0,0,0,22,0,142,0,0,0,125,0,64,0,0,0,191,0,214,0,13,0,86,0,0,0,140,0,233,0,217,0,81,0,33,0,29,0,219,0,32,0,91,0,128,0,17,0,233,0,231,0,104,0,0,0,223,0,134,0,236,0,0,0,0,0,199,0,0,0,157,0,0,0,185,0,64,0,198,0,97,0,48,0,77,0,107,0,20,0,5,0,87,0,190,0,37,0,170,0,0,0,201,0,0,0,0,0,47,0,57,0,174,0,37,0,243,0,36,0,85,0,170,0,48,0,248,0,50,0,51,0,215,0,140,0,124,0,151,0,250,0,109,0,138,0,26,0,0,0,187,0,0,0,207,0,48,0,133,0,178,0,0,0,245,0,227,0,215,0,89,0,12,0,222,0,101,0,231,0,84,0,24,0,70,0,254,0,0,0,6,0,0,0,72,0,0,0,22,0,0,0,114,0,0,0,145,0,0,0,151,0,0,0,63,0,223,0,0,0,0,0,138,0,177,0,0,0,134,0,40,0,111,0,169,0,26,0,154,0,49,0,60,0,123,0,241,0,80,0,0,0,0,0,79,0,0,0,30,0,49,0,154,0,19,0,5,0,0,0,152,0,0,0,228,0,0,0,0,0,234,0,168,0,41,0,228,0,0,0,49,0,0,0,64,0,216,0,2,0,195,0,127,0,81,0,143,0,157,0,0,0,177,0,106,0,59,0,0,0,67,0,147,0,33,0,139,0,30,0,33,0,106,0,0,0,6,0,45,0,225,0,153,0,73,0,0,0,0,0,242,0,151,0,139,0,0,0,122,0,222,0,39,0,0,0,130,0,37,0,59,0,253,0,138,0,144,0);
signal scenario_full  : scenario_type := (113,31,113,30,211,31,99,31,68,31,161,31,119,31,113,31,41,31,4,31,107,31,120,31,116,31,13,31,27,31,166,31,210,31,210,30,65,31,65,30,193,31,140,31,81,31,225,31,149,31,251,31,251,30,47,31,47,30,95,31,76,31,244,31,6,31,6,30,216,31,95,31,93,31,237,31,218,31,127,31,127,30,89,31,12,31,55,31,93,31,67,31,43,31,77,31,79,31,164,31,12,31,130,31,18,31,155,31,19,31,3,31,120,31,155,31,49,31,164,31,191,31,215,31,215,30,215,29,163,31,205,31,191,31,43,31,190,31,190,30,253,31,205,31,66,31,231,31,215,31,15,31,163,31,161,31,110,31,144,31,144,30,26,31,204,31,30,31,30,30,53,31,104,31,222,31,106,31,105,31,105,30,176,31,147,31,21,31,105,31,83,31,116,31,117,31,237,31,177,31,190,31,136,31,136,30,36,31,109,31,195,31,225,31,50,31,50,30,93,31,7,31,104,31,104,30,173,31,25,31,251,31,251,30,244,31,244,30,117,31,117,30,243,31,243,30,119,31,249,31,31,31,240,31,185,31,185,30,130,31,32,31,32,30,182,31,228,31,228,30,170,31,165,31,67,31,244,31,13,31,99,31,210,31,87,31,112,31,112,30,2,31,167,31,224,31,248,31,144,31,152,31,136,31,11,31,237,31,97,31,150,31,150,30,194,31,194,30,238,31,143,31,244,31,157,31,142,31,136,31,117,31,26,31,34,31,110,31,110,30,113,31,208,31,251,31,6,31,6,30,241,31,87,31,45,31,217,31,164,31,229,31,1,31,1,30,1,29,226,31,164,31,164,30,114,31,114,30,135,31,47,31,90,31,71,31,71,30,144,31,149,31,190,31,230,31,58,31,226,31,197,31,23,31,78,31,78,30,223,31,61,31,40,31,210,31,212,31,196,31,205,31,26,31,166,31,103,31,2,31,218,31,253,31,250,31,250,30,142,31,139,31,139,30,88,31,1,31,238,31,254,31,254,30,149,31,218,31,39,31,183,31,183,30,183,29,183,28,66,31,11,31,11,30,247,31,215,31,35,31,226,31,161,31,30,31,67,31,67,30,67,29,225,31,177,31,167,31,186,31,104,31,248,31,217,31,176,31,176,30,231,31,109,31,111,31,190,31,95,31,164,31,91,31,250,31,129,31,66,31,81,31,81,30,31,31,198,31,198,30,160,31,177,31,99,31,66,31,51,31,22,31,97,31,170,31,235,31,127,31,34,31,157,31,219,31,149,31,248,31,137,31,137,30,172,31,79,31,16,31,246,31,208,31,253,31,173,31,101,31,173,31,241,31,24,31,175,31,128,31,211,31,128,31,221,31,242,31,242,30,208,31,228,31,143,31,25,31,86,31,214,31,198,31,81,31,223,31,231,31,120,31,226,31,157,31,187,31,55,31,150,31,190,31,179,31,41,31,12,31,209,31,209,30,18,31,18,30,3,31,178,31,207,31,123,31,233,31,37,31,42,31,106,31,175,31,14,31,198,31,91,31,139,31,69,31,135,31,131,31,90,31,90,30,148,31,197,31,60,31,115,31,59,31,167,31,93,31,244,31,235,31,201,31,218,31,80,31,116,31,194,31,8,31,89,31,10,31,10,30,129,31,173,31,69,31,18,31,75,31,220,31,133,31,68,31,146,31,60,31,82,31,82,30,197,31,68,31,43,31,45,31,95,31,228,31,65,31,92,31,92,30,223,31,41,31,2,31,238,31,238,30,238,29,238,28,10,31,108,31,13,31,183,31,250,31,171,31,171,30,112,31,112,30,249,31,19,31,86,31,76,31,253,31,253,30,231,31,18,31,183,31,76,31,190,31,190,30,162,31,162,30,20,31,20,30,20,29,231,31,23,31,40,31,157,31,141,31,54,31,72,31,59,31,97,31,150,31,227,31,15,31,15,30,17,31,17,30,141,31,172,31,172,30,44,31,82,31,241,31,133,31,167,31,61,31,143,31,56,31,171,31,76,31,70,31,167,31,238,31,90,31,90,30,183,31,183,30,20,31,177,31,117,31,92,31,64,31,87,31,152,31,91,31,254,31,254,30,243,31,98,31,58,31,132,31,132,30,101,31,73,31,161,31,172,31,128,31,128,30,22,31,142,31,142,30,125,31,64,31,64,30,191,31,214,31,13,31,86,31,86,30,140,31,233,31,217,31,81,31,33,31,29,31,219,31,32,31,91,31,128,31,17,31,233,31,231,31,104,31,104,30,223,31,134,31,236,31,236,30,236,29,199,31,199,30,157,31,157,30,185,31,64,31,198,31,97,31,48,31,77,31,107,31,20,31,5,31,87,31,190,31,37,31,170,31,170,30,201,31,201,30,201,29,47,31,57,31,174,31,37,31,243,31,36,31,85,31,170,31,48,31,248,31,50,31,51,31,215,31,140,31,124,31,151,31,250,31,109,31,138,31,26,31,26,30,187,31,187,30,207,31,48,31,133,31,178,31,178,30,245,31,227,31,215,31,89,31,12,31,222,31,101,31,231,31,84,31,24,31,70,31,254,31,254,30,6,31,6,30,72,31,72,30,22,31,22,30,114,31,114,30,145,31,145,30,151,31,151,30,63,31,223,31,223,30,223,29,138,31,177,31,177,30,134,31,40,31,111,31,169,31,26,31,154,31,49,31,60,31,123,31,241,31,80,31,80,30,80,29,79,31,79,30,30,31,49,31,154,31,19,31,5,31,5,30,152,31,152,30,228,31,228,30,228,29,234,31,168,31,41,31,228,31,228,30,49,31,49,30,64,31,216,31,2,31,195,31,127,31,81,31,143,31,157,31,157,30,177,31,106,31,59,31,59,30,67,31,147,31,33,31,139,31,30,31,33,31,106,31,106,30,6,31,45,31,225,31,153,31,73,31,73,30,73,29,242,31,151,31,139,31,139,30,122,31,222,31,39,31,39,30,130,31,37,31,59,31,253,31,138,31,144,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
