-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 446;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (251,0,182,0,0,0,157,0,201,0,14,0,119,0,106,0,0,0,109,0,227,0,0,0,105,0,0,0,103,0,0,0,156,0,0,0,238,0,0,0,158,0,0,0,225,0,8,0,189,0,0,0,114,0,54,0,66,0,28,0,0,0,38,0,195,0,0,0,118,0,62,0,189,0,37,0,219,0,158,0,0,0,81,0,97,0,151,0,46,0,46,0,33,0,186,0,0,0,243,0,144,0,0,0,160,0,75,0,143,0,136,0,2,0,0,0,64,0,161,0,124,0,142,0,56,0,250,0,0,0,186,0,0,0,119,0,131,0,0,0,0,0,240,0,0,0,0,0,0,0,174,0,0,0,5,0,0,0,201,0,40,0,11,0,87,0,127,0,142,0,0,0,61,0,158,0,236,0,11,0,4,0,0,0,187,0,174,0,137,0,220,0,39,0,0,0,37,0,225,0,0,0,164,0,15,0,45,0,0,0,225,0,223,0,213,0,161,0,0,0,166,0,37,0,0,0,0,0,176,0,13,0,0,0,26,0,209,0,72,0,52,0,216,0,126,0,216,0,19,0,20,0,65,0,0,0,206,0,151,0,0,0,237,0,0,0,177,0,225,0,192,0,207,0,86,0,54,0,20,0,168,0,241,0,55,0,80,0,176,0,220,0,0,0,187,0,118,0,28,0,168,0,198,0,2,0,0,0,236,0,29,0,201,0,201,0,58,0,10,0,230,0,102,0,205,0,87,0,155,0,218,0,55,0,215,0,197,0,223,0,0,0,30,0,32,0,0,0,243,0,230,0,47,0,0,0,105,0,227,0,29,0,129,0,170,0,220,0,0,0,0,0,46,0,5,0,0,0,155,0,109,0,233,0,118,0,22,0,144,0,195,0,58,0,0,0,183,0,129,0,0,0,13,0,16,0,208,0,113,0,72,0,134,0,248,0,0,0,234,0,107,0,26,0,58,0,63,0,206,0,165,0,228,0,110,0,102,0,166,0,37,0,105,0,36,0,171,0,162,0,218,0,0,0,46,0,14,0,233,0,0,0,0,0,223,0,228,0,4,0,19,0,5,0,107,0,46,0,173,0,0,0,133,0,233,0,6,0,0,0,157,0,24,0,158,0,233,0,59,0,240,0,115,0,0,0,106,0,242,0,163,0,44,0,0,0,101,0,91,0,29,0,206,0,0,0,238,0,233,0,69,0,96,0,174,0,76,0,32,0,241,0,223,0,139,0,216,0,196,0,93,0,0,0,11,0,90,0,5,0,109,0,0,0,202,0,122,0,231,0,230,0,11,0,3,0,206,0,7,0,93,0,0,0,45,0,102,0,101,0,148,0,161,0,142,0,245,0,0,0,160,0,2,0,0,0,146,0,9,0,249,0,145,0,246,0,248,0,30,0,244,0,169,0,0,0,153,0,227,0,0,0,241,0,179,0,0,0,0,0,0,0,0,0,0,0,127,0,66,0,51,0,23,0,169,0,0,0,224,0,1,0,152,0,116,0,0,0,24,0,176,0,231,0,222,0,246,0,194,0,58,0,77,0,103,0,188,0,34,0,3,0,63,0,66,0,234,0,21,0,100,0,0,0,236,0,85,0,80,0,123,0,75,0,0,0,47,0,214,0,192,0,55,0,53,0,247,0,64,0,46,0,153,0,199,0,159,0,201,0,85,0,84,0,244,0,68,0,240,0,89,0,242,0,161,0,232,0,224,0,119,0,0,0,233,0,130,0,181,0,44,0,227,0,0,0,45,0,0,0,217,0,4,0,0,0,191,0,41,0,0,0,46,0,234,0,179,0,106,0,120,0,211,0,63,0,172,0,108,0,211,0,36,0,140,0,38,0,200,0,205,0,0,0,180,0,218,0,159,0,225,0,83,0,162,0,88,0,167,0,1,0,187,0,177,0,172,0,81,0,222,0,197,0,103,0,0,0,201,0,0,0,0,0,136,0,69,0,0,0,253,0,0,0,171,0,0,0,126,0,40,0,0,0,60,0,240,0,178,0,203,0);
signal scenario_full  : scenario_type := (251,31,182,31,182,30,157,31,201,31,14,31,119,31,106,31,106,30,109,31,227,31,227,30,105,31,105,30,103,31,103,30,156,31,156,30,238,31,238,30,158,31,158,30,225,31,8,31,189,31,189,30,114,31,54,31,66,31,28,31,28,30,38,31,195,31,195,30,118,31,62,31,189,31,37,31,219,31,158,31,158,30,81,31,97,31,151,31,46,31,46,31,33,31,186,31,186,30,243,31,144,31,144,30,160,31,75,31,143,31,136,31,2,31,2,30,64,31,161,31,124,31,142,31,56,31,250,31,250,30,186,31,186,30,119,31,131,31,131,30,131,29,240,31,240,30,240,29,240,28,174,31,174,30,5,31,5,30,201,31,40,31,11,31,87,31,127,31,142,31,142,30,61,31,158,31,236,31,11,31,4,31,4,30,187,31,174,31,137,31,220,31,39,31,39,30,37,31,225,31,225,30,164,31,15,31,45,31,45,30,225,31,223,31,213,31,161,31,161,30,166,31,37,31,37,30,37,29,176,31,13,31,13,30,26,31,209,31,72,31,52,31,216,31,126,31,216,31,19,31,20,31,65,31,65,30,206,31,151,31,151,30,237,31,237,30,177,31,225,31,192,31,207,31,86,31,54,31,20,31,168,31,241,31,55,31,80,31,176,31,220,31,220,30,187,31,118,31,28,31,168,31,198,31,2,31,2,30,236,31,29,31,201,31,201,31,58,31,10,31,230,31,102,31,205,31,87,31,155,31,218,31,55,31,215,31,197,31,223,31,223,30,30,31,32,31,32,30,243,31,230,31,47,31,47,30,105,31,227,31,29,31,129,31,170,31,220,31,220,30,220,29,46,31,5,31,5,30,155,31,109,31,233,31,118,31,22,31,144,31,195,31,58,31,58,30,183,31,129,31,129,30,13,31,16,31,208,31,113,31,72,31,134,31,248,31,248,30,234,31,107,31,26,31,58,31,63,31,206,31,165,31,228,31,110,31,102,31,166,31,37,31,105,31,36,31,171,31,162,31,218,31,218,30,46,31,14,31,233,31,233,30,233,29,223,31,228,31,4,31,19,31,5,31,107,31,46,31,173,31,173,30,133,31,233,31,6,31,6,30,157,31,24,31,158,31,233,31,59,31,240,31,115,31,115,30,106,31,242,31,163,31,44,31,44,30,101,31,91,31,29,31,206,31,206,30,238,31,233,31,69,31,96,31,174,31,76,31,32,31,241,31,223,31,139,31,216,31,196,31,93,31,93,30,11,31,90,31,5,31,109,31,109,30,202,31,122,31,231,31,230,31,11,31,3,31,206,31,7,31,93,31,93,30,45,31,102,31,101,31,148,31,161,31,142,31,245,31,245,30,160,31,2,31,2,30,146,31,9,31,249,31,145,31,246,31,248,31,30,31,244,31,169,31,169,30,153,31,227,31,227,30,241,31,179,31,179,30,179,29,179,28,179,27,179,26,127,31,66,31,51,31,23,31,169,31,169,30,224,31,1,31,152,31,116,31,116,30,24,31,176,31,231,31,222,31,246,31,194,31,58,31,77,31,103,31,188,31,34,31,3,31,63,31,66,31,234,31,21,31,100,31,100,30,236,31,85,31,80,31,123,31,75,31,75,30,47,31,214,31,192,31,55,31,53,31,247,31,64,31,46,31,153,31,199,31,159,31,201,31,85,31,84,31,244,31,68,31,240,31,89,31,242,31,161,31,232,31,224,31,119,31,119,30,233,31,130,31,181,31,44,31,227,31,227,30,45,31,45,30,217,31,4,31,4,30,191,31,41,31,41,30,46,31,234,31,179,31,106,31,120,31,211,31,63,31,172,31,108,31,211,31,36,31,140,31,38,31,200,31,205,31,205,30,180,31,218,31,159,31,225,31,83,31,162,31,88,31,167,31,1,31,187,31,177,31,172,31,81,31,222,31,197,31,103,31,103,30,201,31,201,30,201,29,136,31,69,31,69,30,253,31,253,30,171,31,171,30,126,31,40,31,40,30,60,31,240,31,178,31,203,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
