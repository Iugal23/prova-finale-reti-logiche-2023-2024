-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 287;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,50,0,0,0,66,0,43,0,193,0,14,0,112,0,179,0,13,0,169,0,64,0,193,0,234,0,251,0,165,0,181,0,0,0,235,0,224,0,34,0,35,0,0,0,72,0,144,0,6,0,90,0,71,0,0,0,59,0,0,0,42,0,193,0,0,0,210,0,56,0,17,0,0,0,229,0,167,0,84,0,166,0,56,0,158,0,205,0,83,0,126,0,209,0,0,0,84,0,252,0,182,0,0,0,194,0,6,0,118,0,73,0,234,0,0,0,25,0,138,0,0,0,5,0,0,0,215,0,0,0,13,0,67,0,0,0,80,0,0,0,182,0,119,0,0,0,230,0,224,0,0,0,11,0,156,0,84,0,167,0,14,0,189,0,124,0,212,0,248,0,56,0,115,0,122,0,62,0,0,0,199,0,215,0,170,0,165,0,0,0,2,0,77,0,0,0,187,0,188,0,0,0,3,0,0,0,0,0,219,0,125,0,60,0,3,0,93,0,63,0,0,0,0,0,29,0,75,0,151,0,125,0,0,0,84,0,100,0,175,0,0,0,103,0,63,0,137,0,52,0,73,0,16,0,105,0,167,0,0,0,160,0,110,0,252,0,130,0,116,0,159,0,117,0,100,0,0,0,157,0,168,0,2,0,136,0,190,0,212,0,180,0,21,0,177,0,0,0,58,0,0,0,0,0,179,0,7,0,72,0,248,0,246,0,139,0,67,0,129,0,182,0,143,0,28,0,0,0,132,0,179,0,44,0,65,0,82,0,73,0,58,0,96,0,1,0,214,0,0,0,104,0,0,0,88,0,212,0,142,0,166,0,100,0,215,0,33,0,0,0,0,0,134,0,10,0,0,0,40,0,170,0,0,0,126,0,151,0,18,0,171,0,32,0,111,0,113,0,56,0,132,0,132,0,30,0,0,0,170,0,136,0,26,0,0,0,168,0,109,0,133,0,24,0,19,0,183,0,43,0,74,0,22,0,45,0,219,0,232,0,0,0,246,0,0,0,244,0,127,0,34,0,79,0,87,0,0,0,0,0,0,0,234,0,176,0,200,0,10,0,163,0,99,0,51,0,0,0,228,0,44,0,182,0,36,0,245,0,205,0,170,0,174,0,230,0,121,0,189,0,114,0,185,0,165,0,148,0,0,0,0,0,173,0,42,0,201,0,0,0,57,0,108,0,116,0,156,0,83,0,227,0,254,0,0,0,0,0,126,0,114,0,233,0,191,0,0,0,238,0,18,0,107,0,134,0,50,0,250,0,162,0,172,0,38,0,127,0,108,0,236,0);
signal scenario_full  : scenario_type := (133,31,50,31,50,30,66,31,43,31,193,31,14,31,112,31,179,31,13,31,169,31,64,31,193,31,234,31,251,31,165,31,181,31,181,30,235,31,224,31,34,31,35,31,35,30,72,31,144,31,6,31,90,31,71,31,71,30,59,31,59,30,42,31,193,31,193,30,210,31,56,31,17,31,17,30,229,31,167,31,84,31,166,31,56,31,158,31,205,31,83,31,126,31,209,31,209,30,84,31,252,31,182,31,182,30,194,31,6,31,118,31,73,31,234,31,234,30,25,31,138,31,138,30,5,31,5,30,215,31,215,30,13,31,67,31,67,30,80,31,80,30,182,31,119,31,119,30,230,31,224,31,224,30,11,31,156,31,84,31,167,31,14,31,189,31,124,31,212,31,248,31,56,31,115,31,122,31,62,31,62,30,199,31,215,31,170,31,165,31,165,30,2,31,77,31,77,30,187,31,188,31,188,30,3,31,3,30,3,29,219,31,125,31,60,31,3,31,93,31,63,31,63,30,63,29,29,31,75,31,151,31,125,31,125,30,84,31,100,31,175,31,175,30,103,31,63,31,137,31,52,31,73,31,16,31,105,31,167,31,167,30,160,31,110,31,252,31,130,31,116,31,159,31,117,31,100,31,100,30,157,31,168,31,2,31,136,31,190,31,212,31,180,31,21,31,177,31,177,30,58,31,58,30,58,29,179,31,7,31,72,31,248,31,246,31,139,31,67,31,129,31,182,31,143,31,28,31,28,30,132,31,179,31,44,31,65,31,82,31,73,31,58,31,96,31,1,31,214,31,214,30,104,31,104,30,88,31,212,31,142,31,166,31,100,31,215,31,33,31,33,30,33,29,134,31,10,31,10,30,40,31,170,31,170,30,126,31,151,31,18,31,171,31,32,31,111,31,113,31,56,31,132,31,132,31,30,31,30,30,170,31,136,31,26,31,26,30,168,31,109,31,133,31,24,31,19,31,183,31,43,31,74,31,22,31,45,31,219,31,232,31,232,30,246,31,246,30,244,31,127,31,34,31,79,31,87,31,87,30,87,29,87,28,234,31,176,31,200,31,10,31,163,31,99,31,51,31,51,30,228,31,44,31,182,31,36,31,245,31,205,31,170,31,174,31,230,31,121,31,189,31,114,31,185,31,165,31,148,31,148,30,148,29,173,31,42,31,201,31,201,30,57,31,108,31,116,31,156,31,83,31,227,31,254,31,254,30,254,29,126,31,114,31,233,31,191,31,191,30,238,31,18,31,107,31,134,31,50,31,250,31,162,31,172,31,38,31,127,31,108,31,236,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
