-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 648;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (146,0,243,0,26,0,222,0,75,0,51,0,62,0,100,0,0,0,233,0,10,0,113,0,0,0,62,0,12,0,14,0,0,0,35,0,178,0,118,0,255,0,197,0,114,0,112,0,92,0,52,0,0,0,155,0,59,0,183,0,0,0,167,0,0,0,93,0,172,0,0,0,175,0,116,0,149,0,199,0,225,0,173,0,11,0,1,0,221,0,0,0,0,0,163,0,0,0,126,0,143,0,12,0,253,0,0,0,90,0,0,0,70,0,199,0,219,0,0,0,160,0,65,0,172,0,0,0,32,0,0,0,87,0,225,0,175,0,208,0,168,0,196,0,147,0,135,0,0,0,160,0,98,0,188,0,75,0,95,0,229,0,0,0,159,0,100,0,253,0,63,0,172,0,148,0,0,0,183,0,127,0,0,0,0,0,0,0,94,0,0,0,201,0,177,0,212,0,74,0,24,0,107,0,153,0,38,0,5,0,98,0,202,0,49,0,215,0,77,0,48,0,220,0,99,0,249,0,150,0,41,0,235,0,65,0,108,0,70,0,238,0,226,0,40,0,71,0,239,0,90,0,16,0,89,0,11,0,103,0,198,0,0,0,222,0,21,0,186,0,238,0,242,0,0,0,228,0,220,0,75,0,243,0,27,0,69,0,91,0,40,0,0,0,234,0,70,0,164,0,167,0,77,0,0,0,169,0,152,0,231,0,104,0,250,0,204,0,35,0,54,0,208,0,0,0,253,0,66,0,56,0,141,0,149,0,0,0,226,0,0,0,121,0,0,0,203,0,0,0,122,0,194,0,72,0,233,0,102,0,77,0,253,0,35,0,55,0,0,0,102,0,0,0,0,0,77,0,140,0,0,0,41,0,157,0,53,0,90,0,252,0,0,0,0,0,0,0,176,0,0,0,113,0,0,0,0,0,25,0,216,0,34,0,0,0,203,0,57,0,82,0,41,0,246,0,208,0,92,0,161,0,126,0,127,0,131,0,209,0,0,0,144,0,0,0,0,0,46,0,0,0,176,0,78,0,60,0,51,0,100,0,31,0,61,0,4,0,73,0,156,0,5,0,254,0,130,0,243,0,0,0,153,0,0,0,31,0,63,0,109,0,222,0,236,0,0,0,0,0,107,0,183,0,98,0,0,0,141,0,242,0,108,0,98,0,0,0,95,0,0,0,254,0,87,0,24,0,171,0,156,0,234,0,155,0,0,0,0,0,107,0,0,0,242,0,0,0,0,0,123,0,82,0,0,0,222,0,121,0,206,0,0,0,169,0,38,0,6,0,246,0,83,0,142,0,147,0,214,0,1,0,0,0,0,0,121,0,41,0,234,0,0,0,144,0,244,0,0,0,115,0,103,0,222,0,149,0,107,0,94,0,170,0,0,0,0,0,101,0,112,0,218,0,154,0,119,0,236,0,45,0,41,0,19,0,104,0,221,0,224,0,103,0,112,0,46,0,201,0,30,0,203,0,123,0,183,0,0,0,0,0,148,0,14,0,43,0,14,0,0,0,123,0,205,0,58,0,215,0,33,0,98,0,0,0,65,0,0,0,18,0,130,0,0,0,239,0,24,0,61,0,75,0,15,0,243,0,86,0,217,0,91,0,0,0,86,0,102,0,124,0,0,0,35,0,147,0,0,0,204,0,202,0,164,0,231,0,134,0,191,0,72,0,14,0,0,0,245,0,54,0,139,0,0,0,97,0,217,0,94,0,94,0,76,0,236,0,115,0,213,0,158,0,96,0,210,0,94,0,70,0,0,0,203,0,169,0,0,0,170,0,0,0,138,0,215,0,82,0,0,0,186,0,51,0,65,0,185,0,107,0,201,0,157,0,0,0,213,0,140,0,65,0,30,0,38,0,38,0,0,0,164,0,185,0,46,0,105,0,0,0,63,0,0,0,0,0,108,0,231,0,90,0,131,0,112,0,125,0,0,0,252,0,36,0,165,0,0,0,6,0,12,0,104,0,70,0,81,0,41,0,255,0,133,0,236,0,105,0,0,0,239,0,255,0,132,0,160,0,0,0,0,0,64,0,0,0,108,0,114,0,190,0,57,0,225,0,80,0,72,0,172,0,44,0,121,0,25,0,18,0,51,0,171,0,0,0,173,0,229,0,12,0,137,0,0,0,4,0,170,0,4,0,134,0,195,0,118,0,231,0,0,0,39,0,167,0,204,0,107,0,103,0,55,0,170,0,23,0,0,0,0,0,0,0,14,0,11,0,33,0,7,0,92,0,42,0,28,0,132,0,0,0,0,0,132,0,142,0,251,0,0,0,61,0,5,0,80,0,212,0,237,0,86,0,11,0,134,0,46,0,70,0,222,0,184,0,83,0,67,0,214,0,6,0,19,0,0,0,122,0,108,0,114,0,47,0,181,0,0,0,202,0,139,0,173,0,152,0,56,0,215,0,123,0,197,0,179,0,0,0,191,0,117,0,0,0,159,0,106,0,57,0,143,0,174,0,92,0,129,0,249,0,70,0,0,0,0,0,68,0,0,0,33,0,116,0,224,0,22,0,148,0,116,0,97,0,65,0,228,0,0,0,127,0,16,0,205,0,49,0,220,0,5,0,187,0,0,0,21,0,32,0,98,0,209,0,66,0,103,0,0,0,148,0,30,0,91,0,19,0,226,0,168,0,252,0,52,0,48,0,156,0,248,0,152,0,55,0,147,0,200,0,0,0,54,0,145,0,26,0,79,0,176,0,235,0,0,0,0,0,0,0,225,0,99,0,0,0,0,0,188,0,0,0,0,0,196,0,0,0,106,0,126,0,133,0,0,0,195,0,66,0,0,0,178,0,87,0,89,0,0,0,241,0,4,0,219,0,211,0,142,0,98,0,192,0,0,0,0,0,53,0,79,0,0,0,0,0,255,0,136,0,0,0,177,0,51,0,152,0,21,0,21,0);
signal scenario_full  : scenario_type := (146,31,243,31,26,31,222,31,75,31,51,31,62,31,100,31,100,30,233,31,10,31,113,31,113,30,62,31,12,31,14,31,14,30,35,31,178,31,118,31,255,31,197,31,114,31,112,31,92,31,52,31,52,30,155,31,59,31,183,31,183,30,167,31,167,30,93,31,172,31,172,30,175,31,116,31,149,31,199,31,225,31,173,31,11,31,1,31,221,31,221,30,221,29,163,31,163,30,126,31,143,31,12,31,253,31,253,30,90,31,90,30,70,31,199,31,219,31,219,30,160,31,65,31,172,31,172,30,32,31,32,30,87,31,225,31,175,31,208,31,168,31,196,31,147,31,135,31,135,30,160,31,98,31,188,31,75,31,95,31,229,31,229,30,159,31,100,31,253,31,63,31,172,31,148,31,148,30,183,31,127,31,127,30,127,29,127,28,94,31,94,30,201,31,177,31,212,31,74,31,24,31,107,31,153,31,38,31,5,31,98,31,202,31,49,31,215,31,77,31,48,31,220,31,99,31,249,31,150,31,41,31,235,31,65,31,108,31,70,31,238,31,226,31,40,31,71,31,239,31,90,31,16,31,89,31,11,31,103,31,198,31,198,30,222,31,21,31,186,31,238,31,242,31,242,30,228,31,220,31,75,31,243,31,27,31,69,31,91,31,40,31,40,30,234,31,70,31,164,31,167,31,77,31,77,30,169,31,152,31,231,31,104,31,250,31,204,31,35,31,54,31,208,31,208,30,253,31,66,31,56,31,141,31,149,31,149,30,226,31,226,30,121,31,121,30,203,31,203,30,122,31,194,31,72,31,233,31,102,31,77,31,253,31,35,31,55,31,55,30,102,31,102,30,102,29,77,31,140,31,140,30,41,31,157,31,53,31,90,31,252,31,252,30,252,29,252,28,176,31,176,30,113,31,113,30,113,29,25,31,216,31,34,31,34,30,203,31,57,31,82,31,41,31,246,31,208,31,92,31,161,31,126,31,127,31,131,31,209,31,209,30,144,31,144,30,144,29,46,31,46,30,176,31,78,31,60,31,51,31,100,31,31,31,61,31,4,31,73,31,156,31,5,31,254,31,130,31,243,31,243,30,153,31,153,30,31,31,63,31,109,31,222,31,236,31,236,30,236,29,107,31,183,31,98,31,98,30,141,31,242,31,108,31,98,31,98,30,95,31,95,30,254,31,87,31,24,31,171,31,156,31,234,31,155,31,155,30,155,29,107,31,107,30,242,31,242,30,242,29,123,31,82,31,82,30,222,31,121,31,206,31,206,30,169,31,38,31,6,31,246,31,83,31,142,31,147,31,214,31,1,31,1,30,1,29,121,31,41,31,234,31,234,30,144,31,244,31,244,30,115,31,103,31,222,31,149,31,107,31,94,31,170,31,170,30,170,29,101,31,112,31,218,31,154,31,119,31,236,31,45,31,41,31,19,31,104,31,221,31,224,31,103,31,112,31,46,31,201,31,30,31,203,31,123,31,183,31,183,30,183,29,148,31,14,31,43,31,14,31,14,30,123,31,205,31,58,31,215,31,33,31,98,31,98,30,65,31,65,30,18,31,130,31,130,30,239,31,24,31,61,31,75,31,15,31,243,31,86,31,217,31,91,31,91,30,86,31,102,31,124,31,124,30,35,31,147,31,147,30,204,31,202,31,164,31,231,31,134,31,191,31,72,31,14,31,14,30,245,31,54,31,139,31,139,30,97,31,217,31,94,31,94,31,76,31,236,31,115,31,213,31,158,31,96,31,210,31,94,31,70,31,70,30,203,31,169,31,169,30,170,31,170,30,138,31,215,31,82,31,82,30,186,31,51,31,65,31,185,31,107,31,201,31,157,31,157,30,213,31,140,31,65,31,30,31,38,31,38,31,38,30,164,31,185,31,46,31,105,31,105,30,63,31,63,30,63,29,108,31,231,31,90,31,131,31,112,31,125,31,125,30,252,31,36,31,165,31,165,30,6,31,12,31,104,31,70,31,81,31,41,31,255,31,133,31,236,31,105,31,105,30,239,31,255,31,132,31,160,31,160,30,160,29,64,31,64,30,108,31,114,31,190,31,57,31,225,31,80,31,72,31,172,31,44,31,121,31,25,31,18,31,51,31,171,31,171,30,173,31,229,31,12,31,137,31,137,30,4,31,170,31,4,31,134,31,195,31,118,31,231,31,231,30,39,31,167,31,204,31,107,31,103,31,55,31,170,31,23,31,23,30,23,29,23,28,14,31,11,31,33,31,7,31,92,31,42,31,28,31,132,31,132,30,132,29,132,31,142,31,251,31,251,30,61,31,5,31,80,31,212,31,237,31,86,31,11,31,134,31,46,31,70,31,222,31,184,31,83,31,67,31,214,31,6,31,19,31,19,30,122,31,108,31,114,31,47,31,181,31,181,30,202,31,139,31,173,31,152,31,56,31,215,31,123,31,197,31,179,31,179,30,191,31,117,31,117,30,159,31,106,31,57,31,143,31,174,31,92,31,129,31,249,31,70,31,70,30,70,29,68,31,68,30,33,31,116,31,224,31,22,31,148,31,116,31,97,31,65,31,228,31,228,30,127,31,16,31,205,31,49,31,220,31,5,31,187,31,187,30,21,31,32,31,98,31,209,31,66,31,103,31,103,30,148,31,30,31,91,31,19,31,226,31,168,31,252,31,52,31,48,31,156,31,248,31,152,31,55,31,147,31,200,31,200,30,54,31,145,31,26,31,79,31,176,31,235,31,235,30,235,29,235,28,225,31,99,31,99,30,99,29,188,31,188,30,188,29,196,31,196,30,106,31,126,31,133,31,133,30,195,31,66,31,66,30,178,31,87,31,89,31,89,30,241,31,4,31,219,31,211,31,142,31,98,31,192,31,192,30,192,29,53,31,79,31,79,30,79,29,255,31,136,31,136,30,177,31,51,31,152,31,21,31,21,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
