-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 223;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (163,0,245,0,22,0,128,0,215,0,2,0,144,0,251,0,199,0,20,0,94,0,0,0,68,0,210,0,32,0,37,0,155,0,217,0,190,0,240,0,174,0,0,0,0,0,63,0,161,0,0,0,210,0,0,0,157,0,157,0,211,0,25,0,144,0,0,0,148,0,85,0,0,0,127,0,58,0,199,0,46,0,172,0,64,0,7,0,104,0,0,0,217,0,20,0,174,0,85,0,0,0,99,0,73,0,218,0,230,0,73,0,245,0,0,0,40,0,132,0,121,0,250,0,93,0,0,0,20,0,0,0,242,0,174,0,185,0,64,0,60,0,104,0,155,0,167,0,0,0,0,0,205,0,0,0,249,0,23,0,134,0,136,0,49,0,31,0,24,0,110,0,0,0,234,0,227,0,58,0,74,0,75,0,200,0,75,0,222,0,254,0,240,0,0,0,225,0,0,0,68,0,0,0,12,0,202,0,242,0,232,0,189,0,199,0,0,0,166,0,158,0,0,0,26,0,23,0,199,0,225,0,44,0,205,0,0,0,0,0,75,0,242,0,161,0,20,0,195,0,167,0,231,0,207,0,39,0,98,0,188,0,51,0,170,0,40,0,101,0,93,0,239,0,85,0,0,0,17,0,3,0,0,0,0,0,193,0,255,0,113,0,218,0,186,0,65,0,164,0,48,0,135,0,0,0,200,0,167,0,220,0,122,0,0,0,75,0,68,0,241,0,130,0,0,0,0,0,178,0,44,0,225,0,0,0,0,0,219,0,181,0,143,0,145,0,144,0,11,0,165,0,254,0,0,0,133,0,0,0,83,0,166,0,58,0,137,0,252,0,136,0,74,0,27,0,175,0,236,0,186,0,0,0,0,0,151,0,90,0,0,0,184,0,241,0,0,0,8,0,213,0,0,0,40,0,39,0,137,0,236,0,120,0,76,0,65,0,19,0,33,0,202,0,0,0,157,0,16,0,70,0,139,0,136,0,0,0,191,0,0,0,189,0,234,0);
signal scenario_full  : scenario_type := (163,31,245,31,22,31,128,31,215,31,2,31,144,31,251,31,199,31,20,31,94,31,94,30,68,31,210,31,32,31,37,31,155,31,217,31,190,31,240,31,174,31,174,30,174,29,63,31,161,31,161,30,210,31,210,30,157,31,157,31,211,31,25,31,144,31,144,30,148,31,85,31,85,30,127,31,58,31,199,31,46,31,172,31,64,31,7,31,104,31,104,30,217,31,20,31,174,31,85,31,85,30,99,31,73,31,218,31,230,31,73,31,245,31,245,30,40,31,132,31,121,31,250,31,93,31,93,30,20,31,20,30,242,31,174,31,185,31,64,31,60,31,104,31,155,31,167,31,167,30,167,29,205,31,205,30,249,31,23,31,134,31,136,31,49,31,31,31,24,31,110,31,110,30,234,31,227,31,58,31,74,31,75,31,200,31,75,31,222,31,254,31,240,31,240,30,225,31,225,30,68,31,68,30,12,31,202,31,242,31,232,31,189,31,199,31,199,30,166,31,158,31,158,30,26,31,23,31,199,31,225,31,44,31,205,31,205,30,205,29,75,31,242,31,161,31,20,31,195,31,167,31,231,31,207,31,39,31,98,31,188,31,51,31,170,31,40,31,101,31,93,31,239,31,85,31,85,30,17,31,3,31,3,30,3,29,193,31,255,31,113,31,218,31,186,31,65,31,164,31,48,31,135,31,135,30,200,31,167,31,220,31,122,31,122,30,75,31,68,31,241,31,130,31,130,30,130,29,178,31,44,31,225,31,225,30,225,29,219,31,181,31,143,31,145,31,144,31,11,31,165,31,254,31,254,30,133,31,133,30,83,31,166,31,58,31,137,31,252,31,136,31,74,31,27,31,175,31,236,31,186,31,186,30,186,29,151,31,90,31,90,30,184,31,241,31,241,30,8,31,213,31,213,30,40,31,39,31,137,31,236,31,120,31,76,31,65,31,19,31,33,31,202,31,202,30,157,31,16,31,70,31,139,31,136,31,136,30,191,31,191,30,189,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
