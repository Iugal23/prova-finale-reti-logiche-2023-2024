-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 962;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,184,0,142,0,118,0,154,0,70,0,50,0,117,0,101,0,40,0,0,0,0,0,231,0,226,0,181,0,250,0,207,0,36,0,49,0,143,0,103,0,3,0,25,0,7,0,0,0,172,0,233,0,152,0,55,0,245,0,0,0,152,0,218,0,223,0,90,0,37,0,149,0,72,0,219,0,116,0,175,0,44,0,81,0,11,0,206,0,151,0,0,0,114,0,116,0,129,0,171,0,146,0,213,0,184,0,42,0,66,0,180,0,0,0,0,0,207,0,140,0,135,0,81,0,166,0,142,0,13,0,54,0,0,0,71,0,255,0,151,0,152,0,252,0,27,0,158,0,254,0,10,0,123,0,153,0,73,0,22,0,178,0,190,0,175,0,140,0,146,0,250,0,89,0,99,0,0,0,55,0,9,0,0,0,189,0,0,0,74,0,0,0,152,0,34,0,40,0,236,0,220,0,33,0,15,0,232,0,0,0,126,0,171,0,162,0,244,0,188,0,147,0,0,0,43,0,140,0,37,0,146,0,76,0,102,0,129,0,230,0,102,0,246,0,0,0,22,0,0,0,237,0,57,0,0,0,0,0,8,0,100,0,48,0,46,0,0,0,230,0,53,0,0,0,32,0,123,0,114,0,0,0,72,0,66,0,86,0,237,0,153,0,111,0,126,0,127,0,0,0,134,0,0,0,0,0,9,0,253,0,36,0,153,0,214,0,77,0,77,0,0,0,0,0,0,0,74,0,0,0,245,0,199,0,199,0,203,0,117,0,75,0,0,0,179,0,39,0,0,0,88,0,53,0,83,0,13,0,254,0,0,0,0,0,0,0,29,0,142,0,52,0,0,0,0,0,33,0,0,0,0,0,84,0,0,0,101,0,174,0,85,0,0,0,78,0,238,0,203,0,176,0,0,0,0,0,201,0,183,0,154,0,120,0,203,0,98,0,182,0,56,0,209,0,0,0,78,0,157,0,141,0,2,0,109,0,227,0,217,0,190,0,98,0,117,0,28,0,196,0,0,0,91,0,151,0,0,0,237,0,0,0,12,0,162,0,84,0,64,0,113,0,0,0,0,0,183,0,160,0,237,0,155,0,180,0,200,0,103,0,26,0,32,0,131,0,184,0,236,0,198,0,163,0,147,0,0,0,54,0,38,0,168,0,0,0,123,0,157,0,0,0,0,0,55,0,0,0,159,0,71,0,78,0,237,0,8,0,137,0,0,0,1,0,50,0,193,0,119,0,119,0,179,0,0,0,11,0,49,0,200,0,173,0,98,0,156,0,0,0,35,0,251,0,225,0,0,0,0,0,208,0,145,0,202,0,41,0,0,0,49,0,122,0,145,0,179,0,39,0,43,0,33,0,207,0,12,0,38,0,146,0,0,0,62,0,109,0,112,0,159,0,7,0,25,0,45,0,179,0,0,0,136,0,115,0,0,0,75,0,0,0,0,0,176,0,42,0,212,0,158,0,44,0,202,0,0,0,0,0,200,0,230,0,0,0,20,0,131,0,248,0,0,0,18,0,0,0,0,0,0,0,186,0,70,0,57,0,184,0,19,0,0,0,244,0,94,0,255,0,49,0,220,0,41,0,13,0,155,0,79,0,205,0,22,0,0,0,248,0,0,0,151,0,197,0,180,0,87,0,38,0,0,0,105,0,0,0,72,0,215,0,68,0,50,0,188,0,200,0,0,0,227,0,169,0,19,0,254,0,0,0,0,0,205,0,100,0,116,0,96,0,218,0,209,0,3,0,18,0,185,0,132,0,105,0,30,0,184,0,133,0,16,0,0,0,163,0,118,0,233,0,194,0,121,0,0,0,0,0,18,0,0,0,127,0,133,0,0,0,0,0,252,0,181,0,142,0,189,0,239,0,96,0,28,0,111,0,194,0,49,0,55,0,140,0,166,0,63,0,99,0,204,0,157,0,208,0,43,0,102,0,0,0,48,0,88,0,49,0,16,0,0,0,255,0,190,0,0,0,2,0,0,0,117,0,96,0,4,0,0,0,219,0,141,0,122,0,192,0,0,0,0,0,0,0,6,0,0,0,129,0,170,0,54,0,46,0,227,0,125,0,10,0,5,0,25,0,112,0,100,0,255,0,27,0,167,0,91,0,203,0,72,0,80,0,87,0,220,0,254,0,153,0,88,0,129,0,239,0,132,0,212,0,216,0,0,0,189,0,153,0,47,0,0,0,38,0,100,0,60,0,68,0,219,0,216,0,107,0,67,0,0,0,0,0,199,0,150,0,178,0,70,0,6,0,200,0,28,0,74,0,0,0,158,0,121,0,45,0,0,0,97,0,23,0,0,0,148,0,190,0,132,0,109,0,92,0,97,0,243,0,132,0,250,0,59,0,75,0,80,0,133,0,15,0,0,0,224,0,137,0,0,0,217,0,84,0,23,0,39,0,0,0,131,0,216,0,136,0,27,0,116,0,0,0,69,0,166,0,253,0,27,0,0,0,67,0,0,0,82,0,38,0,22,0,0,0,175,0,3,0,0,0,201,0,218,0,136,0,165,0,8,0,255,0,199,0,0,0,32,0,12,0,113,0,0,0,0,0,234,0,0,0,121,0,158,0,122,0,190,0,0,0,0,0,183,0,67,0,76,0,84,0,238,0,189,0,144,0,71,0,249,0,148,0,16,0,89,0,230,0,0,0,218,0,126,0,135,0,125,0,198,0,0,0,16,0,1,0,50,0,51,0,226,0,130,0,39,0,0,0,69,0,0,0,235,0,14,0,186,0,66,0,185,0,216,0,242,0,48,0,161,0,182,0,11,0,30,0,0,0,237,0,106,0,153,0,0,0,0,0,207,0,25,0,8,0,129,0,239,0,70,0,88,0,233,0,117,0,115,0,28,0,240,0,91,0,185,0,97,0,223,0,72,0,19,0,250,0,55,0,0,0,154,0,166,0,218,0,208,0,248,0,225,0,67,0,222,0,225,0,219,0,0,0,227,0,43,0,2,0,7,0,88,0,97,0,49,0,0,0,96,0,238,0,68,0,39,0,0,0,85,0,168,0,0,0,195,0,30,0,233,0,180,0,0,0,164,0,0,0,0,0,0,0,0,0,0,0,0,0,99,0,205,0,206,0,37,0,96,0,9,0,122,0,20,0,69,0,72,0,116,0,140,0,135,0,202,0,196,0,7,0,59,0,0,0,125,0,0,0,125,0,28,0,43,0,27,0,112,0,15,0,0,0,69,0,201,0,33,0,0,0,32,0,3,0,131,0,210,0,123,0,58,0,0,0,145,0,0,0,42,0,121,0,29,0,114,0,32,0,83,0,0,0,31,0,11,0,0,0,184,0,253,0,174,0,160,0,54,0,0,0,140,0,39,0,11,0,215,0,53,0,0,0,0,0,177,0,185,0,180,0,206,0,221,0,117,0,145,0,74,0,47,0,185,0,70,0,54,0,28,0,205,0,208,0,19,0,58,0,114,0,43,0,0,0,0,0,26,0,220,0,69,0,170,0,28,0,87,0,137,0,173,0,93,0,152,0,206,0,172,0,249,0,144,0,166,0,42,0,211,0,206,0,223,0,119,0,108,0,172,0,79,0,55,0,0,0,0,0,14,0,215,0,122,0,0,0,208,0,62,0,144,0,11,0,0,0,0,0,143,0,125,0,0,0,27,0,124,0,198,0,91,0,0,0,66,0,80,0,0,0,36,0,206,0,216,0,74,0,214,0,44,0,0,0,68,0,231,0,198,0,203,0,97,0,139,0,164,0,75,0,0,0,140,0,239,0,206,0,19,0,148,0,6,0,237,0,112,0,0,0,168,0,110,0,74,0,205,0,173,0,0,0,0,0,4,0,0,0,108,0,134,0,0,0,127,0,0,0,48,0,20,0,183,0,107,0,155,0,83,0,3,0,153,0,71,0,119,0,0,0,0,0,154,0,246,0,223,0,143,0,0,0,178,0,134,0,30,0,137,0,252,0,148,0,0,0,218,0,60,0,155,0,198,0,6,0,6,0,29,0,0,0,0,0,0,0,0,0,133,0,146,0,18,0,208,0,155,0,73,0,211,0,20,0,115,0,140,0,43,0,164,0,194,0,225,0,63,0,178,0,230,0,36,0,223,0,156,0,54,0,237,0,140,0,16,0,73,0,206,0,198,0,69,0,79,0,103,0,109,0,177,0,230,0,2,0,5,0,6,0,0,0,17,0,161,0,0,0,0,0,0,0,228,0,121,0,131,0,138,0,204,0,0,0,225,0,1,0,146,0,0,0,183,0,0,0,113,0,241,0,0,0,176,0,165,0,0,0,0,0,195,0,152,0,153,0,0,0,15,0,51,0,0,0,119,0);
signal scenario_full  : scenario_type := (0,0,0,0,184,31,142,31,118,31,154,31,70,31,50,31,117,31,101,31,40,31,40,30,40,29,231,31,226,31,181,31,250,31,207,31,36,31,49,31,143,31,103,31,3,31,25,31,7,31,7,30,172,31,233,31,152,31,55,31,245,31,245,30,152,31,218,31,223,31,90,31,37,31,149,31,72,31,219,31,116,31,175,31,44,31,81,31,11,31,206,31,151,31,151,30,114,31,116,31,129,31,171,31,146,31,213,31,184,31,42,31,66,31,180,31,180,30,180,29,207,31,140,31,135,31,81,31,166,31,142,31,13,31,54,31,54,30,71,31,255,31,151,31,152,31,252,31,27,31,158,31,254,31,10,31,123,31,153,31,73,31,22,31,178,31,190,31,175,31,140,31,146,31,250,31,89,31,99,31,99,30,55,31,9,31,9,30,189,31,189,30,74,31,74,30,152,31,34,31,40,31,236,31,220,31,33,31,15,31,232,31,232,30,126,31,171,31,162,31,244,31,188,31,147,31,147,30,43,31,140,31,37,31,146,31,76,31,102,31,129,31,230,31,102,31,246,31,246,30,22,31,22,30,237,31,57,31,57,30,57,29,8,31,100,31,48,31,46,31,46,30,230,31,53,31,53,30,32,31,123,31,114,31,114,30,72,31,66,31,86,31,237,31,153,31,111,31,126,31,127,31,127,30,134,31,134,30,134,29,9,31,253,31,36,31,153,31,214,31,77,31,77,31,77,30,77,29,77,28,74,31,74,30,245,31,199,31,199,31,203,31,117,31,75,31,75,30,179,31,39,31,39,30,88,31,53,31,83,31,13,31,254,31,254,30,254,29,254,28,29,31,142,31,52,31,52,30,52,29,33,31,33,30,33,29,84,31,84,30,101,31,174,31,85,31,85,30,78,31,238,31,203,31,176,31,176,30,176,29,201,31,183,31,154,31,120,31,203,31,98,31,182,31,56,31,209,31,209,30,78,31,157,31,141,31,2,31,109,31,227,31,217,31,190,31,98,31,117,31,28,31,196,31,196,30,91,31,151,31,151,30,237,31,237,30,12,31,162,31,84,31,64,31,113,31,113,30,113,29,183,31,160,31,237,31,155,31,180,31,200,31,103,31,26,31,32,31,131,31,184,31,236,31,198,31,163,31,147,31,147,30,54,31,38,31,168,31,168,30,123,31,157,31,157,30,157,29,55,31,55,30,159,31,71,31,78,31,237,31,8,31,137,31,137,30,1,31,50,31,193,31,119,31,119,31,179,31,179,30,11,31,49,31,200,31,173,31,98,31,156,31,156,30,35,31,251,31,225,31,225,30,225,29,208,31,145,31,202,31,41,31,41,30,49,31,122,31,145,31,179,31,39,31,43,31,33,31,207,31,12,31,38,31,146,31,146,30,62,31,109,31,112,31,159,31,7,31,25,31,45,31,179,31,179,30,136,31,115,31,115,30,75,31,75,30,75,29,176,31,42,31,212,31,158,31,44,31,202,31,202,30,202,29,200,31,230,31,230,30,20,31,131,31,248,31,248,30,18,31,18,30,18,29,18,28,186,31,70,31,57,31,184,31,19,31,19,30,244,31,94,31,255,31,49,31,220,31,41,31,13,31,155,31,79,31,205,31,22,31,22,30,248,31,248,30,151,31,197,31,180,31,87,31,38,31,38,30,105,31,105,30,72,31,215,31,68,31,50,31,188,31,200,31,200,30,227,31,169,31,19,31,254,31,254,30,254,29,205,31,100,31,116,31,96,31,218,31,209,31,3,31,18,31,185,31,132,31,105,31,30,31,184,31,133,31,16,31,16,30,163,31,118,31,233,31,194,31,121,31,121,30,121,29,18,31,18,30,127,31,133,31,133,30,133,29,252,31,181,31,142,31,189,31,239,31,96,31,28,31,111,31,194,31,49,31,55,31,140,31,166,31,63,31,99,31,204,31,157,31,208,31,43,31,102,31,102,30,48,31,88,31,49,31,16,31,16,30,255,31,190,31,190,30,2,31,2,30,117,31,96,31,4,31,4,30,219,31,141,31,122,31,192,31,192,30,192,29,192,28,6,31,6,30,129,31,170,31,54,31,46,31,227,31,125,31,10,31,5,31,25,31,112,31,100,31,255,31,27,31,167,31,91,31,203,31,72,31,80,31,87,31,220,31,254,31,153,31,88,31,129,31,239,31,132,31,212,31,216,31,216,30,189,31,153,31,47,31,47,30,38,31,100,31,60,31,68,31,219,31,216,31,107,31,67,31,67,30,67,29,199,31,150,31,178,31,70,31,6,31,200,31,28,31,74,31,74,30,158,31,121,31,45,31,45,30,97,31,23,31,23,30,148,31,190,31,132,31,109,31,92,31,97,31,243,31,132,31,250,31,59,31,75,31,80,31,133,31,15,31,15,30,224,31,137,31,137,30,217,31,84,31,23,31,39,31,39,30,131,31,216,31,136,31,27,31,116,31,116,30,69,31,166,31,253,31,27,31,27,30,67,31,67,30,82,31,38,31,22,31,22,30,175,31,3,31,3,30,201,31,218,31,136,31,165,31,8,31,255,31,199,31,199,30,32,31,12,31,113,31,113,30,113,29,234,31,234,30,121,31,158,31,122,31,190,31,190,30,190,29,183,31,67,31,76,31,84,31,238,31,189,31,144,31,71,31,249,31,148,31,16,31,89,31,230,31,230,30,218,31,126,31,135,31,125,31,198,31,198,30,16,31,1,31,50,31,51,31,226,31,130,31,39,31,39,30,69,31,69,30,235,31,14,31,186,31,66,31,185,31,216,31,242,31,48,31,161,31,182,31,11,31,30,31,30,30,237,31,106,31,153,31,153,30,153,29,207,31,25,31,8,31,129,31,239,31,70,31,88,31,233,31,117,31,115,31,28,31,240,31,91,31,185,31,97,31,223,31,72,31,19,31,250,31,55,31,55,30,154,31,166,31,218,31,208,31,248,31,225,31,67,31,222,31,225,31,219,31,219,30,227,31,43,31,2,31,7,31,88,31,97,31,49,31,49,30,96,31,238,31,68,31,39,31,39,30,85,31,168,31,168,30,195,31,30,31,233,31,180,31,180,30,164,31,164,30,164,29,164,28,164,27,164,26,164,25,99,31,205,31,206,31,37,31,96,31,9,31,122,31,20,31,69,31,72,31,116,31,140,31,135,31,202,31,196,31,7,31,59,31,59,30,125,31,125,30,125,31,28,31,43,31,27,31,112,31,15,31,15,30,69,31,201,31,33,31,33,30,32,31,3,31,131,31,210,31,123,31,58,31,58,30,145,31,145,30,42,31,121,31,29,31,114,31,32,31,83,31,83,30,31,31,11,31,11,30,184,31,253,31,174,31,160,31,54,31,54,30,140,31,39,31,11,31,215,31,53,31,53,30,53,29,177,31,185,31,180,31,206,31,221,31,117,31,145,31,74,31,47,31,185,31,70,31,54,31,28,31,205,31,208,31,19,31,58,31,114,31,43,31,43,30,43,29,26,31,220,31,69,31,170,31,28,31,87,31,137,31,173,31,93,31,152,31,206,31,172,31,249,31,144,31,166,31,42,31,211,31,206,31,223,31,119,31,108,31,172,31,79,31,55,31,55,30,55,29,14,31,215,31,122,31,122,30,208,31,62,31,144,31,11,31,11,30,11,29,143,31,125,31,125,30,27,31,124,31,198,31,91,31,91,30,66,31,80,31,80,30,36,31,206,31,216,31,74,31,214,31,44,31,44,30,68,31,231,31,198,31,203,31,97,31,139,31,164,31,75,31,75,30,140,31,239,31,206,31,19,31,148,31,6,31,237,31,112,31,112,30,168,31,110,31,74,31,205,31,173,31,173,30,173,29,4,31,4,30,108,31,134,31,134,30,127,31,127,30,48,31,20,31,183,31,107,31,155,31,83,31,3,31,153,31,71,31,119,31,119,30,119,29,154,31,246,31,223,31,143,31,143,30,178,31,134,31,30,31,137,31,252,31,148,31,148,30,218,31,60,31,155,31,198,31,6,31,6,31,29,31,29,30,29,29,29,28,29,27,133,31,146,31,18,31,208,31,155,31,73,31,211,31,20,31,115,31,140,31,43,31,164,31,194,31,225,31,63,31,178,31,230,31,36,31,223,31,156,31,54,31,237,31,140,31,16,31,73,31,206,31,198,31,69,31,79,31,103,31,109,31,177,31,230,31,2,31,5,31,6,31,6,30,17,31,161,31,161,30,161,29,161,28,228,31,121,31,131,31,138,31,204,31,204,30,225,31,1,31,146,31,146,30,183,31,183,30,113,31,241,31,241,30,176,31,165,31,165,30,165,29,195,31,152,31,153,31,153,30,15,31,51,31,51,30,119,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
