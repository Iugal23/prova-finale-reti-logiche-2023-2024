-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 327;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (129,0,58,0,0,0,70,0,0,0,92,0,202,0,175,0,154,0,0,0,71,0,198,0,204,0,0,0,162,0,0,0,70,0,79,0,228,0,0,0,95,0,0,0,125,0,81,0,203,0,117,0,145,0,194,0,88,0,155,0,254,0,84,0,0,0,97,0,0,0,0,0,245,0,67,0,162,0,212,0,195,0,6,0,47,0,222,0,56,0,229,0,0,0,40,0,59,0,172,0,188,0,0,0,162,0,0,0,42,0,124,0,38,0,222,0,150,0,251,0,154,0,0,0,0,0,250,0,94,0,132,0,92,0,73,0,58,0,0,0,213,0,113,0,142,0,2,0,0,0,0,0,2,0,224,0,196,0,160,0,43,0,136,0,108,0,0,0,186,0,201,0,127,0,190,0,187,0,53,0,228,0,65,0,0,0,0,0,2,0,76,0,71,0,5,0,205,0,233,0,255,0,51,0,242,0,93,0,91,0,215,0,39,0,147,0,0,0,194,0,213,0,238,0,184,0,234,0,0,0,0,0,0,0,212,0,253,0,178,0,132,0,129,0,0,0,0,0,0,0,0,0,248,0,156,0,250,0,124,0,163,0,138,0,94,0,10,0,162,0,158,0,56,0,0,0,0,0,194,0,246,0,221,0,185,0,84,0,246,0,199,0,89,0,161,0,193,0,6,0,44,0,124,0,2,0,115,0,124,0,0,0,42,0,233,0,91,0,23,0,226,0,0,0,146,0,123,0,126,0,0,0,73,0,198,0,176,0,215,0,27,0,82,0,0,0,79,0,171,0,0,0,71,0,68,0,232,0,0,0,213,0,0,0,178,0,235,0,184,0,210,0,0,0,227,0,186,0,63,0,0,0,207,0,11,0,143,0,41,0,235,0,58,0,0,0,224,0,131,0,232,0,188,0,20,0,116,0,73,0,206,0,166,0,170,0,69,0,168,0,218,0,0,0,155,0,231,0,54,0,190,0,151,0,156,0,128,0,0,0,113,0,0,0,183,0,52,0,113,0,34,0,72,0,0,0,86,0,151,0,60,0,42,0,125,0,172,0,162,0,1,0,83,0,43,0,0,0,114,0,209,0,179,0,0,0,33,0,203,0,229,0,73,0,22,0,0,0,46,0,0,0,0,0,217,0,5,0,49,0,50,0,245,0,132,0,56,0,0,0,78,0,208,0,75,0,59,0,170,0,0,0,0,0,203,0,0,0,62,0,207,0,236,0,252,0,111,0,81,0,0,0,178,0,0,0,0,0,125,0,126,0,44,0,161,0,144,0,224,0,118,0,67,0,209,0,155,0,75,0,147,0,192,0,133,0,13,0,0,0,0,0,104,0,141,0,55,0,0,0,159,0,253,0,200,0,27,0,204,0,146,0,203,0,114,0,219,0,191,0,168,0,177,0,0,0,120,0,26,0,99,0,206,0,40,0,10,0,71,0,245,0,7,0,29,0,245,0,26,0,95,0,116,0);
signal scenario_full  : scenario_type := (129,31,58,31,58,30,70,31,70,30,92,31,202,31,175,31,154,31,154,30,71,31,198,31,204,31,204,30,162,31,162,30,70,31,79,31,228,31,228,30,95,31,95,30,125,31,81,31,203,31,117,31,145,31,194,31,88,31,155,31,254,31,84,31,84,30,97,31,97,30,97,29,245,31,67,31,162,31,212,31,195,31,6,31,47,31,222,31,56,31,229,31,229,30,40,31,59,31,172,31,188,31,188,30,162,31,162,30,42,31,124,31,38,31,222,31,150,31,251,31,154,31,154,30,154,29,250,31,94,31,132,31,92,31,73,31,58,31,58,30,213,31,113,31,142,31,2,31,2,30,2,29,2,31,224,31,196,31,160,31,43,31,136,31,108,31,108,30,186,31,201,31,127,31,190,31,187,31,53,31,228,31,65,31,65,30,65,29,2,31,76,31,71,31,5,31,205,31,233,31,255,31,51,31,242,31,93,31,91,31,215,31,39,31,147,31,147,30,194,31,213,31,238,31,184,31,234,31,234,30,234,29,234,28,212,31,253,31,178,31,132,31,129,31,129,30,129,29,129,28,129,27,248,31,156,31,250,31,124,31,163,31,138,31,94,31,10,31,162,31,158,31,56,31,56,30,56,29,194,31,246,31,221,31,185,31,84,31,246,31,199,31,89,31,161,31,193,31,6,31,44,31,124,31,2,31,115,31,124,31,124,30,42,31,233,31,91,31,23,31,226,31,226,30,146,31,123,31,126,31,126,30,73,31,198,31,176,31,215,31,27,31,82,31,82,30,79,31,171,31,171,30,71,31,68,31,232,31,232,30,213,31,213,30,178,31,235,31,184,31,210,31,210,30,227,31,186,31,63,31,63,30,207,31,11,31,143,31,41,31,235,31,58,31,58,30,224,31,131,31,232,31,188,31,20,31,116,31,73,31,206,31,166,31,170,31,69,31,168,31,218,31,218,30,155,31,231,31,54,31,190,31,151,31,156,31,128,31,128,30,113,31,113,30,183,31,52,31,113,31,34,31,72,31,72,30,86,31,151,31,60,31,42,31,125,31,172,31,162,31,1,31,83,31,43,31,43,30,114,31,209,31,179,31,179,30,33,31,203,31,229,31,73,31,22,31,22,30,46,31,46,30,46,29,217,31,5,31,49,31,50,31,245,31,132,31,56,31,56,30,78,31,208,31,75,31,59,31,170,31,170,30,170,29,203,31,203,30,62,31,207,31,236,31,252,31,111,31,81,31,81,30,178,31,178,30,178,29,125,31,126,31,44,31,161,31,144,31,224,31,118,31,67,31,209,31,155,31,75,31,147,31,192,31,133,31,13,31,13,30,13,29,104,31,141,31,55,31,55,30,159,31,253,31,200,31,27,31,204,31,146,31,203,31,114,31,219,31,191,31,168,31,177,31,177,30,120,31,26,31,99,31,206,31,40,31,10,31,71,31,245,31,7,31,29,31,245,31,26,31,95,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
