-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_534 is
end project_tb_534;

architecture project_tb_arch_534 of project_tb_534 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 698;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,0,0,130,0,127,0,0,0,249,0,211,0,17,0,92,0,227,0,252,0,45,0,32,0,94,0,251,0,151,0,202,0,0,0,39,0,186,0,121,0,218,0,80,0,148,0,0,0,101,0,86,0,217,0,114,0,68,0,186,0,215,0,240,0,181,0,133,0,140,0,0,0,163,0,222,0,0,0,248,0,81,0,82,0,3,0,201,0,0,0,221,0,4,0,0,0,228,0,137,0,129,0,7,0,0,0,178,0,185,0,105,0,229,0,162,0,0,0,8,0,0,0,15,0,44,0,192,0,49,0,114,0,20,0,51,0,211,0,243,0,0,0,92,0,23,0,51,0,61,0,48,0,232,0,120,0,28,0,5,0,0,0,116,0,89,0,117,0,237,0,78,0,0,0,114,0,70,0,191,0,100,0,0,0,0,0,44,0,0,0,76,0,79,0,55,0,0,0,0,0,135,0,118,0,92,0,0,0,0,0,165,0,247,0,0,0,21,0,90,0,85,0,121,0,0,0,9,0,15,0,223,0,215,0,69,0,105,0,213,0,0,0,17,0,0,0,35,0,22,0,0,0,21,0,149,0,119,0,33,0,182,0,43,0,132,0,198,0,4,0,17,0,16,0,88,0,9,0,0,0,0,0,25,0,97,0,204,0,111,0,98,0,142,0,0,0,0,0,111,0,31,0,161,0,241,0,169,0,250,0,148,0,0,0,0,0,229,0,24,0,197,0,7,0,20,0,130,0,82,0,99,0,0,0,4,0,126,0,228,0,229,0,90,0,0,0,179,0,13,0,0,0,25,0,35,0,116,0,132,0,141,0,42,0,10,0,0,0,42,0,72,0,207,0,33,0,106,0,0,0,168,0,101,0,71,0,78,0,140,0,191,0,0,0,86,0,229,0,57,0,0,0,15,0,0,0,131,0,96,0,124,0,32,0,154,0,0,0,0,0,67,0,132,0,231,0,69,0,64,0,2,0,227,0,170,0,21,0,253,0,159,0,54,0,89,0,140,0,149,0,66,0,64,0,113,0,80,0,86,0,250,0,0,0,189,0,0,0,207,0,236,0,191,0,254,0,35,0,189,0,77,0,156,0,251,0,22,0,0,0,0,0,11,0,168,0,0,0,94,0,0,0,78,0,203,0,194,0,93,0,83,0,216,0,109,0,0,0,228,0,0,0,236,0,216,0,0,0,34,0,120,0,196,0,81,0,0,0,40,0,0,0,171,0,11,0,94,0,89,0,174,0,237,0,187,0,169,0,0,0,0,0,0,0,55,0,159,0,188,0,72,0,74,0,70,0,0,0,74,0,0,0,0,0,45,0,0,0,223,0,206,0,118,0,122,0,133,0,176,0,143,0,75,0,0,0,215,0,35,0,128,0,142,0,88,0,35,0,23,0,91,0,43,0,60,0,225,0,196,0,0,0,0,0,0,0,0,0,0,0,72,0,241,0,118,0,171,0,0,0,99,0,37,0,0,0,213,0,207,0,221,0,47,0,0,0,0,0,248,0,110,0,234,0,141,0,211,0,0,0,192,0,0,0,113,0,96,0,75,0,0,0,0,0,64,0,0,0,0,0,242,0,183,0,190,0,13,0,113,0,166,0,237,0,53,0,155,0,114,0,0,0,59,0,19,0,140,0,0,0,228,0,0,0,243,0,35,0,202,0,19,0,0,0,128,0,0,0,0,0,171,0,118,0,116,0,0,0,0,0,212,0,136,0,151,0,137,0,172,0,0,0,160,0,185,0,237,0,192,0,117,0,163,0,136,0,0,0,72,0,0,0,181,0,0,0,65,0,0,0,104,0,26,0,228,0,47,0,88,0,37,0,73,0,241,0,0,0,0,0,0,0,0,0,197,0,114,0,238,0,0,0,151,0,152,0,213,0,190,0,160,0,148,0,243,0,36,0,90,0,0,0,220,0,226,0,0,0,215,0,203,0,132,0,65,0,0,0,0,0,136,0,208,0,211,0,12,0,119,0,25,0,47,0,60,0,99,0,128,0,143,0,83,0,157,0,0,0,5,0,52,0,107,0,245,0,173,0,107,0,0,0,212,0,19,0,4,0,0,0,156,0,7,0,149,0,180,0,147,0,59,0,0,0,0,0,10,0,198,0,56,0,60,0,0,0,0,0,67,0,186,0,88,0,116,0,114,0,0,0,41,0,111,0,66,0,0,0,227,0,8,0,120,0,209,0,109,0,0,0,0,0,147,0,0,0,0,0,200,0,79,0,237,0,0,0,80,0,0,0,159,0,0,0,179,0,0,0,94,0,64,0,117,0,66,0,0,0,238,0,211,0,225,0,239,0,31,0,0,0,71,0,233,0,18,0,201,0,232,0,204,0,172,0,223,0,0,0,96,0,89,0,106,0,152,0,161,0,0,0,157,0,0,0,157,0,219,0,216,0,222,0,66,0,2,0,216,0,0,0,82,0,162,0,0,0,172,0,75,0,153,0,0,0,113,0,0,0,184,0,231,0,107,0,237,0,13,0,0,0,253,0,122,0,31,0,243,0,140,0,146,0,12,0,208,0,0,0,64,0,144,0,0,0,200,0,198,0,83,0,0,0,60,0,202,0,212,0,0,0,241,0,193,0,0,0,144,0,48,0,24,0,253,0,201,0,15,0,129,0,69,0,0,0,148,0,28,0,216,0,247,0,213,0,195,0,156,0,67,0,99,0,68,0,0,0,222,0,0,0,88,0,0,0,182,0,141,0,35,0,164,0,245,0,183,0,0,0,3,0,209,0,159,0,228,0,221,0,215,0,251,0,162,0,60,0,253,0,0,0,152,0,14,0,0,0,245,0,0,0,30,0,42,0,55,0,149,0,170,0,0,0,0,0,0,0,82,0,28,0,142,0,0,0,0,0,45,0,0,0,0,0,0,0,174,0,87,0,121,0,134,0,159,0,98,0,230,0,0,0,27,0,4,0,60,0,68,0,237,0,130,0,85,0,198,0,50,0,35,0,0,0,106,0,0,0,0,0,206,0,240,0,175,0,110,0,114,0,207,0,123,0,179,0,97,0,34,0,168,0,104,0,134,0,235,0,0,0,1,0,240,0,0,0,155,0,25,0,0,0,220,0,50,0,0,0,143,0,147,0,203,0,133,0,160,0,214,0,30,0,102,0,0,0);
signal scenario_full  : scenario_type := (197,31,197,30,130,31,127,31,127,30,249,31,211,31,17,31,92,31,227,31,252,31,45,31,32,31,94,31,251,31,151,31,202,31,202,30,39,31,186,31,121,31,218,31,80,31,148,31,148,30,101,31,86,31,217,31,114,31,68,31,186,31,215,31,240,31,181,31,133,31,140,31,140,30,163,31,222,31,222,30,248,31,81,31,82,31,3,31,201,31,201,30,221,31,4,31,4,30,228,31,137,31,129,31,7,31,7,30,178,31,185,31,105,31,229,31,162,31,162,30,8,31,8,30,15,31,44,31,192,31,49,31,114,31,20,31,51,31,211,31,243,31,243,30,92,31,23,31,51,31,61,31,48,31,232,31,120,31,28,31,5,31,5,30,116,31,89,31,117,31,237,31,78,31,78,30,114,31,70,31,191,31,100,31,100,30,100,29,44,31,44,30,76,31,79,31,55,31,55,30,55,29,135,31,118,31,92,31,92,30,92,29,165,31,247,31,247,30,21,31,90,31,85,31,121,31,121,30,9,31,15,31,223,31,215,31,69,31,105,31,213,31,213,30,17,31,17,30,35,31,22,31,22,30,21,31,149,31,119,31,33,31,182,31,43,31,132,31,198,31,4,31,17,31,16,31,88,31,9,31,9,30,9,29,25,31,97,31,204,31,111,31,98,31,142,31,142,30,142,29,111,31,31,31,161,31,241,31,169,31,250,31,148,31,148,30,148,29,229,31,24,31,197,31,7,31,20,31,130,31,82,31,99,31,99,30,4,31,126,31,228,31,229,31,90,31,90,30,179,31,13,31,13,30,25,31,35,31,116,31,132,31,141,31,42,31,10,31,10,30,42,31,72,31,207,31,33,31,106,31,106,30,168,31,101,31,71,31,78,31,140,31,191,31,191,30,86,31,229,31,57,31,57,30,15,31,15,30,131,31,96,31,124,31,32,31,154,31,154,30,154,29,67,31,132,31,231,31,69,31,64,31,2,31,227,31,170,31,21,31,253,31,159,31,54,31,89,31,140,31,149,31,66,31,64,31,113,31,80,31,86,31,250,31,250,30,189,31,189,30,207,31,236,31,191,31,254,31,35,31,189,31,77,31,156,31,251,31,22,31,22,30,22,29,11,31,168,31,168,30,94,31,94,30,78,31,203,31,194,31,93,31,83,31,216,31,109,31,109,30,228,31,228,30,236,31,216,31,216,30,34,31,120,31,196,31,81,31,81,30,40,31,40,30,171,31,11,31,94,31,89,31,174,31,237,31,187,31,169,31,169,30,169,29,169,28,55,31,159,31,188,31,72,31,74,31,70,31,70,30,74,31,74,30,74,29,45,31,45,30,223,31,206,31,118,31,122,31,133,31,176,31,143,31,75,31,75,30,215,31,35,31,128,31,142,31,88,31,35,31,23,31,91,31,43,31,60,31,225,31,196,31,196,30,196,29,196,28,196,27,196,26,72,31,241,31,118,31,171,31,171,30,99,31,37,31,37,30,213,31,207,31,221,31,47,31,47,30,47,29,248,31,110,31,234,31,141,31,211,31,211,30,192,31,192,30,113,31,96,31,75,31,75,30,75,29,64,31,64,30,64,29,242,31,183,31,190,31,13,31,113,31,166,31,237,31,53,31,155,31,114,31,114,30,59,31,19,31,140,31,140,30,228,31,228,30,243,31,35,31,202,31,19,31,19,30,128,31,128,30,128,29,171,31,118,31,116,31,116,30,116,29,212,31,136,31,151,31,137,31,172,31,172,30,160,31,185,31,237,31,192,31,117,31,163,31,136,31,136,30,72,31,72,30,181,31,181,30,65,31,65,30,104,31,26,31,228,31,47,31,88,31,37,31,73,31,241,31,241,30,241,29,241,28,241,27,197,31,114,31,238,31,238,30,151,31,152,31,213,31,190,31,160,31,148,31,243,31,36,31,90,31,90,30,220,31,226,31,226,30,215,31,203,31,132,31,65,31,65,30,65,29,136,31,208,31,211,31,12,31,119,31,25,31,47,31,60,31,99,31,128,31,143,31,83,31,157,31,157,30,5,31,52,31,107,31,245,31,173,31,107,31,107,30,212,31,19,31,4,31,4,30,156,31,7,31,149,31,180,31,147,31,59,31,59,30,59,29,10,31,198,31,56,31,60,31,60,30,60,29,67,31,186,31,88,31,116,31,114,31,114,30,41,31,111,31,66,31,66,30,227,31,8,31,120,31,209,31,109,31,109,30,109,29,147,31,147,30,147,29,200,31,79,31,237,31,237,30,80,31,80,30,159,31,159,30,179,31,179,30,94,31,64,31,117,31,66,31,66,30,238,31,211,31,225,31,239,31,31,31,31,30,71,31,233,31,18,31,201,31,232,31,204,31,172,31,223,31,223,30,96,31,89,31,106,31,152,31,161,31,161,30,157,31,157,30,157,31,219,31,216,31,222,31,66,31,2,31,216,31,216,30,82,31,162,31,162,30,172,31,75,31,153,31,153,30,113,31,113,30,184,31,231,31,107,31,237,31,13,31,13,30,253,31,122,31,31,31,243,31,140,31,146,31,12,31,208,31,208,30,64,31,144,31,144,30,200,31,198,31,83,31,83,30,60,31,202,31,212,31,212,30,241,31,193,31,193,30,144,31,48,31,24,31,253,31,201,31,15,31,129,31,69,31,69,30,148,31,28,31,216,31,247,31,213,31,195,31,156,31,67,31,99,31,68,31,68,30,222,31,222,30,88,31,88,30,182,31,141,31,35,31,164,31,245,31,183,31,183,30,3,31,209,31,159,31,228,31,221,31,215,31,251,31,162,31,60,31,253,31,253,30,152,31,14,31,14,30,245,31,245,30,30,31,42,31,55,31,149,31,170,31,170,30,170,29,170,28,82,31,28,31,142,31,142,30,142,29,45,31,45,30,45,29,45,28,174,31,87,31,121,31,134,31,159,31,98,31,230,31,230,30,27,31,4,31,60,31,68,31,237,31,130,31,85,31,198,31,50,31,35,31,35,30,106,31,106,30,106,29,206,31,240,31,175,31,110,31,114,31,207,31,123,31,179,31,97,31,34,31,168,31,104,31,134,31,235,31,235,30,1,31,240,31,240,30,155,31,25,31,25,30,220,31,50,31,50,30,143,31,147,31,203,31,133,31,160,31,214,31,30,31,102,31,102,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
