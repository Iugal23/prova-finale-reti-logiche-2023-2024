-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 581;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (74,0,191,0,154,0,222,0,249,0,86,0,231,0,0,0,73,0,109,0,38,0,154,0,66,0,245,0,216,0,154,0,0,0,0,0,230,0,61,0,180,0,159,0,0,0,241,0,93,0,193,0,1,0,0,0,0,0,160,0,179,0,137,0,0,0,80,0,220,0,185,0,45,0,205,0,33,0,17,0,179,0,111,0,205,0,253,0,8,0,56,0,0,0,237,0,156,0,0,0,223,0,69,0,63,0,169,0,171,0,80,0,238,0,30,0,178,0,234,0,202,0,148,0,53,0,0,0,116,0,96,0,0,0,212,0,158,0,85,0,105,0,0,0,172,0,0,0,123,0,109,0,131,0,25,0,88,0,14,0,0,0,0,0,136,0,223,0,203,0,12,0,125,0,63,0,209,0,172,0,240,0,64,0,0,0,16,0,210,0,85,0,47,0,228,0,177,0,172,0,145,0,0,0,103,0,41,0,33,0,0,0,62,0,24,0,78,0,0,0,147,0,182,0,86,0,198,0,245,0,131,0,104,0,148,0,64,0,21,0,146,0,114,0,14,0,95,0,168,0,47,0,175,0,215,0,82,0,0,0,0,0,0,0,99,0,35,0,0,0,0,0,64,0,129,0,77,0,203,0,78,0,41,0,99,0,5,0,101,0,218,0,143,0,0,0,0,0,22,0,190,0,0,0,228,0,0,0,244,0,8,0,0,0,200,0,72,0,0,0,176,0,106,0,154,0,118,0,7,0,0,0,247,0,215,0,87,0,140,0,40,0,200,0,46,0,4,0,0,0,163,0,0,0,202,0,159,0,19,0,30,0,5,0,98,0,0,0,1,0,165,0,0,0,145,0,188,0,54,0,0,0,47,0,0,0,18,0,0,0,47,0,0,0,87,0,45,0,101,0,170,0,241,0,20,0,232,0,33,0,235,0,153,0,79,0,145,0,0,0,80,0,165,0,142,0,227,0,0,0,0,0,0,0,108,0,95,0,152,0,0,0,0,0,54,0,35,0,0,0,16,0,192,0,215,0,41,0,69,0,178,0,0,0,53,0,0,0,0,0,74,0,88,0,21,0,86,0,224,0,207,0,199,0,10,0,0,0,44,0,2,0,67,0,0,0,0,0,140,0,26,0,88,0,12,0,113,0,135,0,0,0,244,0,217,0,0,0,2,0,92,0,9,0,80,0,229,0,232,0,77,0,143,0,241,0,216,0,0,0,31,0,47,0,0,0,0,0,217,0,125,0,222,0,5,0,220,0,53,0,0,0,6,0,185,0,0,0,83,0,168,0,62,0,162,0,137,0,219,0,136,0,83,0,247,0,252,0,0,0,149,0,0,0,239,0,242,0,168,0,40,0,150,0,250,0,0,0,131,0,29,0,189,0,0,0,0,0,35,0,200,0,132,0,6,0,30,0,156,0,246,0,160,0,0,0,50,0,237,0,233,0,0,0,177,0,156,0,0,0,199,0,253,0,112,0,165,0,0,0,119,0,75,0,192,0,0,0,18,0,30,0,136,0,209,0,244,0,247,0,151,0,0,0,15,0,0,0,0,0,0,0,118,0,208,0,120,0,220,0,54,0,126,0,127,0,37,0,86,0,0,0,199,0,127,0,8,0,90,0,0,0,0,0,0,0,35,0,201,0,7,0,108,0,236,0,180,0,74,0,238,0,99,0,174,0,41,0,51,0,249,0,86,0,0,0,0,0,68,0,172,0,0,0,197,0,98,0,0,0,73,0,0,0,59,0,0,0,43,0,154,0,189,0,147,0,235,0,87,0,0,0,0,0,230,0,3,0,135,0,28,0,0,0,0,0,213,0,0,0,145,0,52,0,5,0,249,0,113,0,39,0,94,0,232,0,3,0,136,0,15,0,145,0,49,0,27,0,39,0,0,0,138,0,0,0,0,0,123,0,191,0,0,0,82,0,0,0,198,0,157,0,107,0,177,0,0,0,107,0,124,0,0,0,92,0,241,0,151,0,218,0,0,0,0,0,55,0,0,0,181,0,57,0,0,0,115,0,242,0,184,0,31,0,162,0,81,0,0,0,225,0,17,0,26,0,68,0,90,0,16,0,235,0,43,0,0,0,0,0,84,0,0,0,85,0,164,0,0,0,94,0,39,0,25,0,87,0,0,0,232,0,241,0,109,0,254,0,0,0,191,0,23,0,254,0,52,0,25,0,190,0,107,0,63,0,209,0,0,0,21,0,0,0,52,0,0,0,10,0,182,0,42,0,182,0,0,0,99,0,7,0,0,0,105,0,10,0,139,0,0,0,107,0,223,0,27,0,148,0,186,0,68,0,38,0,187,0,210,0,62,0,0,0,0,0,73,0,239,0,81,0,220,0,117,0,163,0,0,0,238,0,0,0,30,0,37,0,111,0,0,0,8,0,56,0,0,0,99,0,222,0,0,0,0,0,107,0,0,0,0,0,17,0,0,0,0,0,120,0,205,0,0,0,32,0,0,0,164,0,17,0,86,0,181,0,218,0,61,0,204,0,208,0,231,0,215,0,29,0,0,0,221,0,73,0,0,0,23,0,1,0,118,0,131,0,121,0,0,0,53,0,0,0,64,0,112,0,96,0,132,0,189,0,84,0,157,0,112,0,100,0);
signal scenario_full  : scenario_type := (74,31,191,31,154,31,222,31,249,31,86,31,231,31,231,30,73,31,109,31,38,31,154,31,66,31,245,31,216,31,154,31,154,30,154,29,230,31,61,31,180,31,159,31,159,30,241,31,93,31,193,31,1,31,1,30,1,29,160,31,179,31,137,31,137,30,80,31,220,31,185,31,45,31,205,31,33,31,17,31,179,31,111,31,205,31,253,31,8,31,56,31,56,30,237,31,156,31,156,30,223,31,69,31,63,31,169,31,171,31,80,31,238,31,30,31,178,31,234,31,202,31,148,31,53,31,53,30,116,31,96,31,96,30,212,31,158,31,85,31,105,31,105,30,172,31,172,30,123,31,109,31,131,31,25,31,88,31,14,31,14,30,14,29,136,31,223,31,203,31,12,31,125,31,63,31,209,31,172,31,240,31,64,31,64,30,16,31,210,31,85,31,47,31,228,31,177,31,172,31,145,31,145,30,103,31,41,31,33,31,33,30,62,31,24,31,78,31,78,30,147,31,182,31,86,31,198,31,245,31,131,31,104,31,148,31,64,31,21,31,146,31,114,31,14,31,95,31,168,31,47,31,175,31,215,31,82,31,82,30,82,29,82,28,99,31,35,31,35,30,35,29,64,31,129,31,77,31,203,31,78,31,41,31,99,31,5,31,101,31,218,31,143,31,143,30,143,29,22,31,190,31,190,30,228,31,228,30,244,31,8,31,8,30,200,31,72,31,72,30,176,31,106,31,154,31,118,31,7,31,7,30,247,31,215,31,87,31,140,31,40,31,200,31,46,31,4,31,4,30,163,31,163,30,202,31,159,31,19,31,30,31,5,31,98,31,98,30,1,31,165,31,165,30,145,31,188,31,54,31,54,30,47,31,47,30,18,31,18,30,47,31,47,30,87,31,45,31,101,31,170,31,241,31,20,31,232,31,33,31,235,31,153,31,79,31,145,31,145,30,80,31,165,31,142,31,227,31,227,30,227,29,227,28,108,31,95,31,152,31,152,30,152,29,54,31,35,31,35,30,16,31,192,31,215,31,41,31,69,31,178,31,178,30,53,31,53,30,53,29,74,31,88,31,21,31,86,31,224,31,207,31,199,31,10,31,10,30,44,31,2,31,67,31,67,30,67,29,140,31,26,31,88,31,12,31,113,31,135,31,135,30,244,31,217,31,217,30,2,31,92,31,9,31,80,31,229,31,232,31,77,31,143,31,241,31,216,31,216,30,31,31,47,31,47,30,47,29,217,31,125,31,222,31,5,31,220,31,53,31,53,30,6,31,185,31,185,30,83,31,168,31,62,31,162,31,137,31,219,31,136,31,83,31,247,31,252,31,252,30,149,31,149,30,239,31,242,31,168,31,40,31,150,31,250,31,250,30,131,31,29,31,189,31,189,30,189,29,35,31,200,31,132,31,6,31,30,31,156,31,246,31,160,31,160,30,50,31,237,31,233,31,233,30,177,31,156,31,156,30,199,31,253,31,112,31,165,31,165,30,119,31,75,31,192,31,192,30,18,31,30,31,136,31,209,31,244,31,247,31,151,31,151,30,15,31,15,30,15,29,15,28,118,31,208,31,120,31,220,31,54,31,126,31,127,31,37,31,86,31,86,30,199,31,127,31,8,31,90,31,90,30,90,29,90,28,35,31,201,31,7,31,108,31,236,31,180,31,74,31,238,31,99,31,174,31,41,31,51,31,249,31,86,31,86,30,86,29,68,31,172,31,172,30,197,31,98,31,98,30,73,31,73,30,59,31,59,30,43,31,154,31,189,31,147,31,235,31,87,31,87,30,87,29,230,31,3,31,135,31,28,31,28,30,28,29,213,31,213,30,145,31,52,31,5,31,249,31,113,31,39,31,94,31,232,31,3,31,136,31,15,31,145,31,49,31,27,31,39,31,39,30,138,31,138,30,138,29,123,31,191,31,191,30,82,31,82,30,198,31,157,31,107,31,177,31,177,30,107,31,124,31,124,30,92,31,241,31,151,31,218,31,218,30,218,29,55,31,55,30,181,31,57,31,57,30,115,31,242,31,184,31,31,31,162,31,81,31,81,30,225,31,17,31,26,31,68,31,90,31,16,31,235,31,43,31,43,30,43,29,84,31,84,30,85,31,164,31,164,30,94,31,39,31,25,31,87,31,87,30,232,31,241,31,109,31,254,31,254,30,191,31,23,31,254,31,52,31,25,31,190,31,107,31,63,31,209,31,209,30,21,31,21,30,52,31,52,30,10,31,182,31,42,31,182,31,182,30,99,31,7,31,7,30,105,31,10,31,139,31,139,30,107,31,223,31,27,31,148,31,186,31,68,31,38,31,187,31,210,31,62,31,62,30,62,29,73,31,239,31,81,31,220,31,117,31,163,31,163,30,238,31,238,30,30,31,37,31,111,31,111,30,8,31,56,31,56,30,99,31,222,31,222,30,222,29,107,31,107,30,107,29,17,31,17,30,17,29,120,31,205,31,205,30,32,31,32,30,164,31,17,31,86,31,181,31,218,31,61,31,204,31,208,31,231,31,215,31,29,31,29,30,221,31,73,31,73,30,23,31,1,31,118,31,131,31,121,31,121,30,53,31,53,30,64,31,112,31,96,31,132,31,189,31,84,31,157,31,112,31,100,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
