-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 803;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (80,0,0,0,228,0,212,0,128,0,0,0,101,0,131,0,0,0,111,0,174,0,0,0,0,0,83,0,215,0,239,0,3,0,181,0,218,0,214,0,51,0,255,0,113,0,0,0,221,0,22,0,207,0,167,0,62,0,0,0,209,0,198,0,88,0,57,0,186,0,0,0,56,0,151,0,20,0,212,0,0,0,242,0,134,0,0,0,99,0,8,0,0,0,0,0,184,0,203,0,175,0,232,0,195,0,0,0,49,0,0,0,158,0,0,0,175,0,32,0,62,0,171,0,52,0,0,0,0,0,176,0,156,0,54,0,227,0,21,0,0,0,8,0,89,0,236,0,147,0,41,0,143,0,129,0,0,0,0,0,75,0,70,0,165,0,82,0,147,0,231,0,227,0,62,0,0,0,0,0,0,0,157,0,20,0,43,0,113,0,0,0,126,0,218,0,10,0,0,0,190,0,3,0,0,0,0,0,0,0,183,0,7,0,0,0,240,0,95,0,0,0,45,0,0,0,123,0,0,0,0,0,192,0,116,0,113,0,0,0,0,0,100,0,0,0,173,0,173,0,0,0,0,0,26,0,89,0,111,0,59,0,0,0,226,0,0,0,0,0,176,0,239,0,209,0,26,0,91,0,15,0,175,0,0,0,73,0,148,0,124,0,209,0,9,0,0,0,0,0,0,0,0,0,0,0,41,0,38,0,184,0,24,0,0,0,0,0,0,0,195,0,175,0,26,0,58,0,86,0,227,0,101,0,98,0,34,0,0,0,197,0,230,0,131,0,149,0,222,0,55,0,189,0,172,0,117,0,0,0,117,0,238,0,199,0,71,0,154,0,164,0,0,0,166,0,23,0,99,0,0,0,0,0,163,0,74,0,139,0,238,0,29,0,223,0,82,0,106,0,193,0,0,0,0,0,0,0,11,0,42,0,77,0,119,0,240,0,99,0,18,0,161,0,221,0,29,0,125,0,165,0,26,0,0,0,0,0,170,0,217,0,103,0,237,0,91,0,85,0,65,0,50,0,126,0,137,0,164,0,244,0,0,0,10,0,152,0,78,0,131,0,10,0,222,0,37,0,86,0,109,0,59,0,156,0,99,0,46,0,0,0,58,0,130,0,56,0,0,0,33,0,193,0,181,0,76,0,0,0,112,0,66,0,0,0,15,0,7,0,25,0,0,0,108,0,219,0,0,0,0,0,159,0,255,0,32,0,221,0,113,0,147,0,43,0,149,0,6,0,5,0,240,0,61,0,0,0,232,0,36,0,75,0,33,0,91,0,84,0,46,0,0,0,140,0,166,0,128,0,24,0,172,0,6,0,0,0,69,0,0,0,205,0,0,0,160,0,127,0,143,0,0,0,0,0,0,0,0,0,240,0,0,0,110,0,250,0,103,0,12,0,89,0,184,0,112,0,138,0,0,0,0,0,108,0,96,0,75,0,170,0,1,0,24,0,24,0,46,0,130,0,157,0,0,0,170,0,99,0,239,0,0,0,100,0,241,0,136,0,0,0,208,0,0,0,60,0,0,0,230,0,64,0,66,0,0,0,5,0,178,0,50,0,0,0,47,0,0,0,35,0,2,0,0,0,0,0,32,0,168,0,0,0,126,0,127,0,20,0,114,0,0,0,138,0,212,0,232,0,192,0,21,0,227,0,41,0,16,0,158,0,170,0,12,0,107,0,0,0,225,0,137,0,95,0,29,0,233,0,62,0,182,0,222,0,118,0,145,0,175,0,184,0,67,0,106,0,207,0,14,0,145,0,106,0,26,0,90,0,11,0,215,0,196,0,90,0,148,0,51,0,15,0,97,0,0,0,0,0,0,0,26,0,220,0,62,0,57,0,53,0,14,0,198,0,13,0,174,0,80,0,218,0,0,0,101,0,208,0,64,0,208,0,138,0,0,0,11,0,217,0,48,0,25,0,0,0,61,0,125,0,166,0,0,0,127,0,64,0,57,0,156,0,0,0,244,0,10,0,156,0,236,0,3,0,18,0,0,0,0,0,175,0,10,0,235,0,0,0,0,0,196,0,15,0,131,0,228,0,89,0,29,0,102,0,42,0,95,0,254,0,21,0,0,0,0,0,176,0,214,0,169,0,12,0,74,0,89,0,8,0,228,0,0,0,111,0,64,0,151,0,199,0,0,0,0,0,193,0,80,0,205,0,139,0,42,0,0,0,75,0,155,0,47,0,106,0,179,0,75,0,6,0,107,0,47,0,124,0,168,0,180,0,39,0,66,0,59,0,135,0,133,0,250,0,168,0,15,0,60,0,227,0,223,0,110,0,22,0,218,0,143,0,108,0,193,0,0,0,78,0,0,0,0,0,161,0,223,0,139,0,0,0,254,0,226,0,0,0,78,0,218,0,56,0,161,0,221,0,131,0,137,0,68,0,28,0,237,0,26,0,35,0,52,0,99,0,29,0,0,0,153,0,185,0,63,0,237,0,222,0,0,0,113,0,144,0,0,0,113,0,228,0,100,0,192,0,97,0,207,0,160,0,0,0,85,0,122,0,0,0,43,0,71,0,109,0,103,0,77,0,69,0,105,0,58,0,202,0,191,0,120,0,102,0,109,0,118,0,162,0,192,0,233,0,168,0,0,0,63,0,227,0,240,0,168,0,21,0,157,0,153,0,85,0,0,0,88,0,70,0,94,0,0,0,90,0,136,0,178,0,18,0,85,0,15,0,217,0,117,0,0,0,152,0,136,0,227,0,0,0,3,0,0,0,188,0,0,0,51,0,42,0,150,0,37,0,4,0,85,0,0,0,108,0,0,0,0,0,46,0,29,0,38,0,32,0,219,0,135,0,179,0,114,0,201,0,237,0,0,0,56,0,210,0,0,0,84,0,95,0,233,0,140,0,228,0,216,0,198,0,0,0,0,0,7,0,27,0,0,0,176,0,43,0,196,0,0,0,176,0,93,0,218,0,224,0,31,0,14,0,46,0,185,0,182,0,254,0,0,0,209,0,135,0,222,0,223,0,0,0,212,0,177,0,171,0,91,0,180,0,55,0,0,0,250,0,152,0,178,0,144,0,154,0,248,0,0,0,248,0,168,0,20,0,0,0,41,0,169,0,0,0,231,0,150,0,96,0,74,0,19,0,45,0,0,0,242,0,99,0,132,0,25,0,67,0,208,0,0,0,51,0,226,0,104,0,0,0,110,0,205,0,54,0,139,0,71,0,0,0,79,0,43,0,28,0,136,0,0,0,217,0,36,0,15,0,254,0,20,0,13,0,177,0,27,0,164,0,13,0,174,0,0,0,213,0,13,0,0,0,25,0,163,0,138,0,174,0,44,0,108,0,148,0,104,0,21,0,10,0,83,0,62,0,98,0,188,0,111,0,206,0,61,0,12,0,127,0,155,0,0,0,68,0,128,0,71,0,6,0,98,0,206,0,20,0,30,0,98,0,88,0,242,0,140,0,59,0,64,0,218,0,254,0,253,0,42,0,199,0,214,0,158,0,244,0,216,0,113,0,0,0,0,0,181,0,193,0,107,0,124,0,202,0,214,0,240,0,44,0,0,0,91,0,0,0,139,0,134,0,0,0,231,0,0,0,115,0,0,0,2,0,65,0,115,0,0,0,43,0,45,0,153,0);
signal scenario_full  : scenario_type := (80,31,80,30,228,31,212,31,128,31,128,30,101,31,131,31,131,30,111,31,174,31,174,30,174,29,83,31,215,31,239,31,3,31,181,31,218,31,214,31,51,31,255,31,113,31,113,30,221,31,22,31,207,31,167,31,62,31,62,30,209,31,198,31,88,31,57,31,186,31,186,30,56,31,151,31,20,31,212,31,212,30,242,31,134,31,134,30,99,31,8,31,8,30,8,29,184,31,203,31,175,31,232,31,195,31,195,30,49,31,49,30,158,31,158,30,175,31,32,31,62,31,171,31,52,31,52,30,52,29,176,31,156,31,54,31,227,31,21,31,21,30,8,31,89,31,236,31,147,31,41,31,143,31,129,31,129,30,129,29,75,31,70,31,165,31,82,31,147,31,231,31,227,31,62,31,62,30,62,29,62,28,157,31,20,31,43,31,113,31,113,30,126,31,218,31,10,31,10,30,190,31,3,31,3,30,3,29,3,28,183,31,7,31,7,30,240,31,95,31,95,30,45,31,45,30,123,31,123,30,123,29,192,31,116,31,113,31,113,30,113,29,100,31,100,30,173,31,173,31,173,30,173,29,26,31,89,31,111,31,59,31,59,30,226,31,226,30,226,29,176,31,239,31,209,31,26,31,91,31,15,31,175,31,175,30,73,31,148,31,124,31,209,31,9,31,9,30,9,29,9,28,9,27,9,26,41,31,38,31,184,31,24,31,24,30,24,29,24,28,195,31,175,31,26,31,58,31,86,31,227,31,101,31,98,31,34,31,34,30,197,31,230,31,131,31,149,31,222,31,55,31,189,31,172,31,117,31,117,30,117,31,238,31,199,31,71,31,154,31,164,31,164,30,166,31,23,31,99,31,99,30,99,29,163,31,74,31,139,31,238,31,29,31,223,31,82,31,106,31,193,31,193,30,193,29,193,28,11,31,42,31,77,31,119,31,240,31,99,31,18,31,161,31,221,31,29,31,125,31,165,31,26,31,26,30,26,29,170,31,217,31,103,31,237,31,91,31,85,31,65,31,50,31,126,31,137,31,164,31,244,31,244,30,10,31,152,31,78,31,131,31,10,31,222,31,37,31,86,31,109,31,59,31,156,31,99,31,46,31,46,30,58,31,130,31,56,31,56,30,33,31,193,31,181,31,76,31,76,30,112,31,66,31,66,30,15,31,7,31,25,31,25,30,108,31,219,31,219,30,219,29,159,31,255,31,32,31,221,31,113,31,147,31,43,31,149,31,6,31,5,31,240,31,61,31,61,30,232,31,36,31,75,31,33,31,91,31,84,31,46,31,46,30,140,31,166,31,128,31,24,31,172,31,6,31,6,30,69,31,69,30,205,31,205,30,160,31,127,31,143,31,143,30,143,29,143,28,143,27,240,31,240,30,110,31,250,31,103,31,12,31,89,31,184,31,112,31,138,31,138,30,138,29,108,31,96,31,75,31,170,31,1,31,24,31,24,31,46,31,130,31,157,31,157,30,170,31,99,31,239,31,239,30,100,31,241,31,136,31,136,30,208,31,208,30,60,31,60,30,230,31,64,31,66,31,66,30,5,31,178,31,50,31,50,30,47,31,47,30,35,31,2,31,2,30,2,29,32,31,168,31,168,30,126,31,127,31,20,31,114,31,114,30,138,31,212,31,232,31,192,31,21,31,227,31,41,31,16,31,158,31,170,31,12,31,107,31,107,30,225,31,137,31,95,31,29,31,233,31,62,31,182,31,222,31,118,31,145,31,175,31,184,31,67,31,106,31,207,31,14,31,145,31,106,31,26,31,90,31,11,31,215,31,196,31,90,31,148,31,51,31,15,31,97,31,97,30,97,29,97,28,26,31,220,31,62,31,57,31,53,31,14,31,198,31,13,31,174,31,80,31,218,31,218,30,101,31,208,31,64,31,208,31,138,31,138,30,11,31,217,31,48,31,25,31,25,30,61,31,125,31,166,31,166,30,127,31,64,31,57,31,156,31,156,30,244,31,10,31,156,31,236,31,3,31,18,31,18,30,18,29,175,31,10,31,235,31,235,30,235,29,196,31,15,31,131,31,228,31,89,31,29,31,102,31,42,31,95,31,254,31,21,31,21,30,21,29,176,31,214,31,169,31,12,31,74,31,89,31,8,31,228,31,228,30,111,31,64,31,151,31,199,31,199,30,199,29,193,31,80,31,205,31,139,31,42,31,42,30,75,31,155,31,47,31,106,31,179,31,75,31,6,31,107,31,47,31,124,31,168,31,180,31,39,31,66,31,59,31,135,31,133,31,250,31,168,31,15,31,60,31,227,31,223,31,110,31,22,31,218,31,143,31,108,31,193,31,193,30,78,31,78,30,78,29,161,31,223,31,139,31,139,30,254,31,226,31,226,30,78,31,218,31,56,31,161,31,221,31,131,31,137,31,68,31,28,31,237,31,26,31,35,31,52,31,99,31,29,31,29,30,153,31,185,31,63,31,237,31,222,31,222,30,113,31,144,31,144,30,113,31,228,31,100,31,192,31,97,31,207,31,160,31,160,30,85,31,122,31,122,30,43,31,71,31,109,31,103,31,77,31,69,31,105,31,58,31,202,31,191,31,120,31,102,31,109,31,118,31,162,31,192,31,233,31,168,31,168,30,63,31,227,31,240,31,168,31,21,31,157,31,153,31,85,31,85,30,88,31,70,31,94,31,94,30,90,31,136,31,178,31,18,31,85,31,15,31,217,31,117,31,117,30,152,31,136,31,227,31,227,30,3,31,3,30,188,31,188,30,51,31,42,31,150,31,37,31,4,31,85,31,85,30,108,31,108,30,108,29,46,31,29,31,38,31,32,31,219,31,135,31,179,31,114,31,201,31,237,31,237,30,56,31,210,31,210,30,84,31,95,31,233,31,140,31,228,31,216,31,198,31,198,30,198,29,7,31,27,31,27,30,176,31,43,31,196,31,196,30,176,31,93,31,218,31,224,31,31,31,14,31,46,31,185,31,182,31,254,31,254,30,209,31,135,31,222,31,223,31,223,30,212,31,177,31,171,31,91,31,180,31,55,31,55,30,250,31,152,31,178,31,144,31,154,31,248,31,248,30,248,31,168,31,20,31,20,30,41,31,169,31,169,30,231,31,150,31,96,31,74,31,19,31,45,31,45,30,242,31,99,31,132,31,25,31,67,31,208,31,208,30,51,31,226,31,104,31,104,30,110,31,205,31,54,31,139,31,71,31,71,30,79,31,43,31,28,31,136,31,136,30,217,31,36,31,15,31,254,31,20,31,13,31,177,31,27,31,164,31,13,31,174,31,174,30,213,31,13,31,13,30,25,31,163,31,138,31,174,31,44,31,108,31,148,31,104,31,21,31,10,31,83,31,62,31,98,31,188,31,111,31,206,31,61,31,12,31,127,31,155,31,155,30,68,31,128,31,71,31,6,31,98,31,206,31,20,31,30,31,98,31,88,31,242,31,140,31,59,31,64,31,218,31,254,31,253,31,42,31,199,31,214,31,158,31,244,31,216,31,113,31,113,30,113,29,181,31,193,31,107,31,124,31,202,31,214,31,240,31,44,31,44,30,91,31,91,30,139,31,134,31,134,30,231,31,231,30,115,31,115,30,2,31,65,31,115,31,115,30,43,31,45,31,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
