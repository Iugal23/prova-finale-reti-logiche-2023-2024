-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 654;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,114,0,175,0,254,0,229,0,249,0,236,0,175,0,73,0,28,0,72,0,123,0,131,0,0,0,254,0,65,0,0,0,171,0,152,0,214,0,250,0,113,0,0,0,125,0,33,0,22,0,176,0,76,0,0,0,248,0,140,0,202,0,234,0,245,0,82,0,0,0,0,0,91,0,67,0,188,0,4,0,205,0,32,0,201,0,234,0,19,0,126,0,188,0,96,0,0,0,0,0,0,0,216,0,0,0,12,0,209,0,205,0,126,0,130,0,216,0,187,0,0,0,0,0,0,0,56,0,158,0,221,0,0,0,36,0,145,0,88,0,160,0,122,0,0,0,0,0,80,0,218,0,211,0,0,0,189,0,148,0,197,0,19,0,23,0,215,0,0,0,75,0,0,0,191,0,0,0,121,0,135,0,90,0,0,0,88,0,0,0,171,0,32,0,143,0,0,0,0,0,145,0,0,0,0,0,192,0,27,0,0,0,173,0,182,0,0,0,56,0,0,0,0,0,0,0,251,0,0,0,0,0,0,0,0,0,67,0,0,0,69,0,63,0,119,0,44,0,57,0,0,0,0,0,93,0,161,0,188,0,106,0,98,0,0,0,126,0,216,0,144,0,83,0,134,0,69,0,192,0,171,0,140,0,121,0,163,0,141,0,70,0,216,0,70,0,99,0,171,0,0,0,138,0,238,0,219,0,21,0,139,0,0,0,74,0,38,0,16,0,0,0,226,0,37,0,97,0,0,0,0,0,248,0,192,0,0,0,0,0,38,0,211,0,165,0,42,0,174,0,225,0,233,0,122,0,64,0,13,0,100,0,0,0,218,0,42,0,80,0,0,0,72,0,30,0,172,0,198,0,5,0,0,0,135,0,7,0,250,0,47,0,125,0,183,0,211,0,140,0,0,0,132,0,0,0,95,0,237,0,0,0,40,0,213,0,0,0,53,0,0,0,33,0,127,0,66,0,142,0,0,0,198,0,156,0,245,0,248,0,43,0,253,0,47,0,146,0,102,0,0,0,184,0,0,0,214,0,46,0,0,0,114,0,124,0,119,0,0,0,251,0,53,0,3,0,114,0,180,0,51,0,0,0,190,0,201,0,95,0,17,0,74,0,63,0,215,0,0,0,28,0,127,0,134,0,43,0,107,0,199,0,0,0,189,0,34,0,88,0,35,0,10,0,43,0,42,0,71,0,168,0,124,0,0,0,0,0,105,0,0,0,80,0,92,0,0,0,67,0,133,0,19,0,66,0,215,0,89,0,253,0,24,0,197,0,90,0,0,0,0,0,166,0,40,0,0,0,158,0,200,0,0,0,29,0,113,0,174,0,218,0,74,0,182,0,116,0,0,0,21,0,115,0,0,0,79,0,2,0,0,0,110,0,0,0,24,0,230,0,122,0,0,0,198,0,119,0,253,0,8,0,199,0,60,0,136,0,0,0,216,0,223,0,0,0,206,0,228,0,190,0,151,0,171,0,64,0,227,0,191,0,250,0,0,0,0,0,0,0,168,0,66,0,0,0,0,0,89,0,130,0,206,0,0,0,54,0,70,0,197,0,0,0,176,0,51,0,81,0,115,0,0,0,185,0,179,0,100,0,115,0,141,0,145,0,77,0,125,0,0,0,214,0,199,0,165,0,226,0,6,0,0,0,75,0,21,0,78,0,0,0,204,0,29,0,38,0,215,0,105,0,182,0,203,0,87,0,0,0,0,0,204,0,1,0,203,0,205,0,57,0,107,0,0,0,0,0,39,0,221,0,65,0,77,0,90,0,0,0,0,0,113,0,43,0,160,0,203,0,90,0,251,0,244,0,60,0,11,0,171,0,212,0,112,0,226,0,11,0,112,0,46,0,207,0,195,0,65,0,79,0,241,0,0,0,85,0,49,0,193,0,25,0,88,0,0,0,17,0,245,0,77,0,176,0,182,0,182,0,35,0,123,0,148,0,252,0,96,0,41,0,63,0,188,0,180,0,36,0,0,0,9,0,152,0,240,0,139,0,239,0,210,0,97,0,209,0,212,0,0,0,0,0,137,0,0,0,200,0,98,0,0,0,0,0,116,0,9,0,41,0,233,0,60,0,47,0,247,0,0,0,30,0,115,0,0,0,128,0,0,0,156,0,8,0,253,0,164,0,56,0,78,0,80,0,161,0,0,0,110,0,181,0,197,0,145,0,128,0,114,0,13,0,133,0,211,0,42,0,0,0,0,0,56,0,58,0,0,0,31,0,111,0,58,0,251,0,230,0,206,0,0,0,0,0,227,0,0,0,201,0,0,0,5,0,238,0,133,0,145,0,55,0,233,0,40,0,187,0,23,0,61,0,162,0,131,0,182,0,231,0,23,0,1,0,204,0,60,0,0,0,0,0,40,0,41,0,0,0,213,0,135,0,0,0,70,0,158,0,99,0,248,0,0,0,188,0,182,0,241,0,85,0,0,0,202,0,244,0,0,0,131,0,28,0,145,0,0,0,52,0,165,0,24,0,17,0,97,0,140,0,93,0,172,0,109,0,80,0,162,0,53,0,183,0,224,0,219,0,124,0,2,0,0,0,62,0,0,0,154,0,0,0,0,0,249,0,238,0,174,0,159,0,117,0,43,0,81,0,68,0,171,0,13,0,0,0,0,0,0,0,10,0,112,0,168,0,182,0,102,0,0,0,220,0,0,0,103,0,0,0,236,0,213,0,0,0,105,0,0,0,2,0,110,0,156,0,153,0,14,0,0,0,214,0,46,0,134,0,0,0,67,0,14,0,112,0,68,0,0,0,61,0,181,0,143,0,110,0,41,0,126,0,0,0,0,0,56,0,69,0,162,0,0,0,118,0,253,0,0,0,229,0,160,0,2,0,0,0,21,0,0,0,177,0,81,0,0,0,153,0,0,0,58,0,241,0,3,0,0,0,0,0,0,0,226,0,0,0,230,0,169,0,0,0);
signal scenario_full  : scenario_type := (0,0,114,31,175,31,254,31,229,31,249,31,236,31,175,31,73,31,28,31,72,31,123,31,131,31,131,30,254,31,65,31,65,30,171,31,152,31,214,31,250,31,113,31,113,30,125,31,33,31,22,31,176,31,76,31,76,30,248,31,140,31,202,31,234,31,245,31,82,31,82,30,82,29,91,31,67,31,188,31,4,31,205,31,32,31,201,31,234,31,19,31,126,31,188,31,96,31,96,30,96,29,96,28,216,31,216,30,12,31,209,31,205,31,126,31,130,31,216,31,187,31,187,30,187,29,187,28,56,31,158,31,221,31,221,30,36,31,145,31,88,31,160,31,122,31,122,30,122,29,80,31,218,31,211,31,211,30,189,31,148,31,197,31,19,31,23,31,215,31,215,30,75,31,75,30,191,31,191,30,121,31,135,31,90,31,90,30,88,31,88,30,171,31,32,31,143,31,143,30,143,29,145,31,145,30,145,29,192,31,27,31,27,30,173,31,182,31,182,30,56,31,56,30,56,29,56,28,251,31,251,30,251,29,251,28,251,27,67,31,67,30,69,31,63,31,119,31,44,31,57,31,57,30,57,29,93,31,161,31,188,31,106,31,98,31,98,30,126,31,216,31,144,31,83,31,134,31,69,31,192,31,171,31,140,31,121,31,163,31,141,31,70,31,216,31,70,31,99,31,171,31,171,30,138,31,238,31,219,31,21,31,139,31,139,30,74,31,38,31,16,31,16,30,226,31,37,31,97,31,97,30,97,29,248,31,192,31,192,30,192,29,38,31,211,31,165,31,42,31,174,31,225,31,233,31,122,31,64,31,13,31,100,31,100,30,218,31,42,31,80,31,80,30,72,31,30,31,172,31,198,31,5,31,5,30,135,31,7,31,250,31,47,31,125,31,183,31,211,31,140,31,140,30,132,31,132,30,95,31,237,31,237,30,40,31,213,31,213,30,53,31,53,30,33,31,127,31,66,31,142,31,142,30,198,31,156,31,245,31,248,31,43,31,253,31,47,31,146,31,102,31,102,30,184,31,184,30,214,31,46,31,46,30,114,31,124,31,119,31,119,30,251,31,53,31,3,31,114,31,180,31,51,31,51,30,190,31,201,31,95,31,17,31,74,31,63,31,215,31,215,30,28,31,127,31,134,31,43,31,107,31,199,31,199,30,189,31,34,31,88,31,35,31,10,31,43,31,42,31,71,31,168,31,124,31,124,30,124,29,105,31,105,30,80,31,92,31,92,30,67,31,133,31,19,31,66,31,215,31,89,31,253,31,24,31,197,31,90,31,90,30,90,29,166,31,40,31,40,30,158,31,200,31,200,30,29,31,113,31,174,31,218,31,74,31,182,31,116,31,116,30,21,31,115,31,115,30,79,31,2,31,2,30,110,31,110,30,24,31,230,31,122,31,122,30,198,31,119,31,253,31,8,31,199,31,60,31,136,31,136,30,216,31,223,31,223,30,206,31,228,31,190,31,151,31,171,31,64,31,227,31,191,31,250,31,250,30,250,29,250,28,168,31,66,31,66,30,66,29,89,31,130,31,206,31,206,30,54,31,70,31,197,31,197,30,176,31,51,31,81,31,115,31,115,30,185,31,179,31,100,31,115,31,141,31,145,31,77,31,125,31,125,30,214,31,199,31,165,31,226,31,6,31,6,30,75,31,21,31,78,31,78,30,204,31,29,31,38,31,215,31,105,31,182,31,203,31,87,31,87,30,87,29,204,31,1,31,203,31,205,31,57,31,107,31,107,30,107,29,39,31,221,31,65,31,77,31,90,31,90,30,90,29,113,31,43,31,160,31,203,31,90,31,251,31,244,31,60,31,11,31,171,31,212,31,112,31,226,31,11,31,112,31,46,31,207,31,195,31,65,31,79,31,241,31,241,30,85,31,49,31,193,31,25,31,88,31,88,30,17,31,245,31,77,31,176,31,182,31,182,31,35,31,123,31,148,31,252,31,96,31,41,31,63,31,188,31,180,31,36,31,36,30,9,31,152,31,240,31,139,31,239,31,210,31,97,31,209,31,212,31,212,30,212,29,137,31,137,30,200,31,98,31,98,30,98,29,116,31,9,31,41,31,233,31,60,31,47,31,247,31,247,30,30,31,115,31,115,30,128,31,128,30,156,31,8,31,253,31,164,31,56,31,78,31,80,31,161,31,161,30,110,31,181,31,197,31,145,31,128,31,114,31,13,31,133,31,211,31,42,31,42,30,42,29,56,31,58,31,58,30,31,31,111,31,58,31,251,31,230,31,206,31,206,30,206,29,227,31,227,30,201,31,201,30,5,31,238,31,133,31,145,31,55,31,233,31,40,31,187,31,23,31,61,31,162,31,131,31,182,31,231,31,23,31,1,31,204,31,60,31,60,30,60,29,40,31,41,31,41,30,213,31,135,31,135,30,70,31,158,31,99,31,248,31,248,30,188,31,182,31,241,31,85,31,85,30,202,31,244,31,244,30,131,31,28,31,145,31,145,30,52,31,165,31,24,31,17,31,97,31,140,31,93,31,172,31,109,31,80,31,162,31,53,31,183,31,224,31,219,31,124,31,2,31,2,30,62,31,62,30,154,31,154,30,154,29,249,31,238,31,174,31,159,31,117,31,43,31,81,31,68,31,171,31,13,31,13,30,13,29,13,28,10,31,112,31,168,31,182,31,102,31,102,30,220,31,220,30,103,31,103,30,236,31,213,31,213,30,105,31,105,30,2,31,110,31,156,31,153,31,14,31,14,30,214,31,46,31,134,31,134,30,67,31,14,31,112,31,68,31,68,30,61,31,181,31,143,31,110,31,41,31,126,31,126,30,126,29,56,31,69,31,162,31,162,30,118,31,253,31,253,30,229,31,160,31,2,31,2,30,21,31,21,30,177,31,81,31,81,30,153,31,153,30,58,31,241,31,3,31,3,30,3,29,3,28,226,31,226,30,230,31,169,31,169,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
