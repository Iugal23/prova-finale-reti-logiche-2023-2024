-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_665 is
end project_tb_665;

architecture project_tb_arch_665 of project_tb_665 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 462;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,0,0,0,0,0,0,117,0,125,0,201,0,132,0,96,0,140,0,158,0,0,0,148,0,26,0,138,0,0,0,209,0,226,0,0,0,0,0,48,0,240,0,17,0,175,0,164,0,54,0,12,0,7,0,232,0,245,0,0,0,173,0,159,0,94,0,80,0,228,0,165,0,82,0,238,0,183,0,148,0,111,0,183,0,0,0,0,0,92,0,0,0,8,0,233,0,0,0,37,0,220,0,23,0,6,0,0,0,214,0,0,0,80,0,0,0,0,0,189,0,207,0,121,0,0,0,0,0,87,0,179,0,243,0,204,0,18,0,0,0,147,0,13,0,242,0,135,0,168,0,145,0,48,0,33,0,0,0,93,0,101,0,219,0,193,0,236,0,166,0,0,0,190,0,153,0,57,0,62,0,140,0,12,0,126,0,47,0,17,0,0,0,0,0,76,0,16,0,63,0,0,0,123,0,32,0,45,0,52,0,73,0,0,0,239,0,0,0,28,0,96,0,0,0,0,0,187,0,196,0,4,0,217,0,177,0,251,0,0,0,204,0,196,0,19,0,18,0,63,0,178,0,46,0,73,0,147,0,18,0,138,0,171,0,0,0,162,0,16,0,0,0,57,0,0,0,194,0,226,0,72,0,22,0,125,0,83,0,0,0,113,0,2,0,227,0,202,0,166,0,92,0,0,0,57,0,0,0,214,0,248,0,70,0,73,0,253,0,10,0,228,0,101,0,74,0,17,0,171,0,105,0,0,0,178,0,233,0,146,0,65,0,237,0,208,0,68,0,187,0,171,0,0,0,0,0,135,0,9,0,191,0,23,0,17,0,155,0,242,0,0,0,28,0,0,0,232,0,40,0,212,0,106,0,0,0,129,0,214,0,0,0,253,0,209,0,162,0,65,0,9,0,73,0,0,0,238,0,0,0,75,0,69,0,68,0,147,0,14,0,233,0,0,0,224,0,190,0,0,0,0,0,156,0,19,0,115,0,11,0,143,0,163,0,0,0,146,0,210,0,153,0,0,0,37,0,0,0,0,0,27,0,16,0,117,0,178,0,179,0,44,0,213,0,0,0,60,0,173,0,205,0,0,0,60,0,171,0,184,0,50,0,232,0,217,0,164,0,111,0,100,0,113,0,149,0,109,0,236,0,56,0,30,0,0,0,108,0,0,0,0,0,0,0,58,0,206,0,99,0,22,0,0,0,139,0,0,0,108,0,22,0,89,0,57,0,248,0,173,0,0,0,142,0,0,0,0,0,237,0,203,0,119,0,46,0,48,0,143,0,143,0,109,0,6,0,66,0,105,0,51,0,209,0,183,0,48,0,200,0,111,0,204,0,0,0,93,0,0,0,0,0,189,0,117,0,196,0,51,0,52,0,156,0,116,0,58,0,36,0,185,0,0,0,183,0,51,0,239,0,1,0,74,0,210,0,251,0,141,0,147,0,0,0,16,0,27,0,0,0,44,0,1,0,72,0,70,0,0,0,247,0,135,0,51,0,0,0,1,0,69,0,134,0,218,0,3,0,102,0,88,0,67,0,65,0,109,0,112,0,0,0,77,0,103,0,62,0,252,0,8,0,0,0,163,0,235,0,0,0,0,0,168,0,173,0,152,0,0,0,0,0,0,0,44,0,56,0,71,0,0,0,190,0,106,0,0,0,184,0,128,0,24,0,203,0,0,0,120,0,234,0,86,0,16,0,142,0,251,0,0,0,64,0,0,0,24,0,100,0,19,0,158,0,179,0,200,0,9,0,213,0,0,0,117,0,0,0,77,0,117,0,134,0,0,0,102,0,144,0,168,0,247,0,94,0,179,0,148,0,50,0,207,0,92,0,22,0,21,0,122,0,203,0,114,0,254,0,156,0,0,0,24,0,83,0,86,0,146,0,252,0,192,0,55,0,20,0,0,0,255,0,195,0,141,0,145,0,157,0,83,0,128,0,162,0,220,0,162,0,0,0,121,0,125,0,137,0,105,0,160,0,0,0,105,0,105,0,253,0,143,0,66,0,232,0,149,0,0,0,126,0,242,0,0,0,167,0,125,0,237,0,112,0,170,0,89,0,123,0,72,0);
signal scenario_full  : scenario_type := (9,31,9,30,9,29,9,28,117,31,125,31,201,31,132,31,96,31,140,31,158,31,158,30,148,31,26,31,138,31,138,30,209,31,226,31,226,30,226,29,48,31,240,31,17,31,175,31,164,31,54,31,12,31,7,31,232,31,245,31,245,30,173,31,159,31,94,31,80,31,228,31,165,31,82,31,238,31,183,31,148,31,111,31,183,31,183,30,183,29,92,31,92,30,8,31,233,31,233,30,37,31,220,31,23,31,6,31,6,30,214,31,214,30,80,31,80,30,80,29,189,31,207,31,121,31,121,30,121,29,87,31,179,31,243,31,204,31,18,31,18,30,147,31,13,31,242,31,135,31,168,31,145,31,48,31,33,31,33,30,93,31,101,31,219,31,193,31,236,31,166,31,166,30,190,31,153,31,57,31,62,31,140,31,12,31,126,31,47,31,17,31,17,30,17,29,76,31,16,31,63,31,63,30,123,31,32,31,45,31,52,31,73,31,73,30,239,31,239,30,28,31,96,31,96,30,96,29,187,31,196,31,4,31,217,31,177,31,251,31,251,30,204,31,196,31,19,31,18,31,63,31,178,31,46,31,73,31,147,31,18,31,138,31,171,31,171,30,162,31,16,31,16,30,57,31,57,30,194,31,226,31,72,31,22,31,125,31,83,31,83,30,113,31,2,31,227,31,202,31,166,31,92,31,92,30,57,31,57,30,214,31,248,31,70,31,73,31,253,31,10,31,228,31,101,31,74,31,17,31,171,31,105,31,105,30,178,31,233,31,146,31,65,31,237,31,208,31,68,31,187,31,171,31,171,30,171,29,135,31,9,31,191,31,23,31,17,31,155,31,242,31,242,30,28,31,28,30,232,31,40,31,212,31,106,31,106,30,129,31,214,31,214,30,253,31,209,31,162,31,65,31,9,31,73,31,73,30,238,31,238,30,75,31,69,31,68,31,147,31,14,31,233,31,233,30,224,31,190,31,190,30,190,29,156,31,19,31,115,31,11,31,143,31,163,31,163,30,146,31,210,31,153,31,153,30,37,31,37,30,37,29,27,31,16,31,117,31,178,31,179,31,44,31,213,31,213,30,60,31,173,31,205,31,205,30,60,31,171,31,184,31,50,31,232,31,217,31,164,31,111,31,100,31,113,31,149,31,109,31,236,31,56,31,30,31,30,30,108,31,108,30,108,29,108,28,58,31,206,31,99,31,22,31,22,30,139,31,139,30,108,31,22,31,89,31,57,31,248,31,173,31,173,30,142,31,142,30,142,29,237,31,203,31,119,31,46,31,48,31,143,31,143,31,109,31,6,31,66,31,105,31,51,31,209,31,183,31,48,31,200,31,111,31,204,31,204,30,93,31,93,30,93,29,189,31,117,31,196,31,51,31,52,31,156,31,116,31,58,31,36,31,185,31,185,30,183,31,51,31,239,31,1,31,74,31,210,31,251,31,141,31,147,31,147,30,16,31,27,31,27,30,44,31,1,31,72,31,70,31,70,30,247,31,135,31,51,31,51,30,1,31,69,31,134,31,218,31,3,31,102,31,88,31,67,31,65,31,109,31,112,31,112,30,77,31,103,31,62,31,252,31,8,31,8,30,163,31,235,31,235,30,235,29,168,31,173,31,152,31,152,30,152,29,152,28,44,31,56,31,71,31,71,30,190,31,106,31,106,30,184,31,128,31,24,31,203,31,203,30,120,31,234,31,86,31,16,31,142,31,251,31,251,30,64,31,64,30,24,31,100,31,19,31,158,31,179,31,200,31,9,31,213,31,213,30,117,31,117,30,77,31,117,31,134,31,134,30,102,31,144,31,168,31,247,31,94,31,179,31,148,31,50,31,207,31,92,31,22,31,21,31,122,31,203,31,114,31,254,31,156,31,156,30,24,31,83,31,86,31,146,31,252,31,192,31,55,31,20,31,20,30,255,31,195,31,141,31,145,31,157,31,83,31,128,31,162,31,220,31,162,31,162,30,121,31,125,31,137,31,105,31,160,31,160,30,105,31,105,31,253,31,143,31,66,31,232,31,149,31,149,30,126,31,242,31,242,30,167,31,125,31,237,31,112,31,170,31,89,31,123,31,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
