-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 873;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,28,0,0,0,71,0,0,0,0,0,241,0,82,0,0,0,147,0,0,0,130,0,228,0,33,0,188,0,37,0,211,0,0,0,0,0,111,0,147,0,107,0,195,0,110,0,0,0,0,0,227,0,0,0,58,0,0,0,147,0,0,0,0,0,68,0,105,0,168,0,27,0,227,0,252,0,63,0,14,0,0,0,217,0,22,0,6,0,168,0,32,0,0,0,32,0,184,0,69,0,230,0,0,0,95,0,0,0,71,0,38,0,220,0,0,0,219,0,0,0,191,0,131,0,0,0,41,0,30,0,145,0,241,0,182,0,200,0,30,0,0,0,209,0,174,0,204,0,3,0,41,0,37,0,2,0,119,0,158,0,14,0,31,0,211,0,194,0,37,0,244,0,0,0,201,0,0,0,176,0,107,0,169,0,40,0,136,0,198,0,0,0,20,0,2,0,134,0,154,0,247,0,114,0,0,0,124,0,97,0,76,0,113,0,0,0,60,0,31,0,223,0,63,0,75,0,172,0,40,0,126,0,76,0,26,0,0,0,229,0,0,0,144,0,25,0,56,0,10,0,37,0,105,0,28,0,57,0,0,0,154,0,151,0,106,0,89,0,51,0,219,0,17,0,0,0,65,0,0,0,217,0,78,0,106,0,59,0,130,0,104,0,201,0,0,0,207,0,177,0,227,0,124,0,180,0,189,0,101,0,120,0,38,0,195,0,0,0,47,0,51,0,174,0,101,0,10,0,0,0,11,0,103,0,0,0,228,0,89,0,128,0,60,0,180,0,0,0,219,0,200,0,152,0,199,0,186,0,0,0,177,0,185,0,100,0,167,0,151,0,138,0,99,0,174,0,0,0,0,0,237,0,10,0,0,0,17,0,170,0,152,0,199,0,83,0,129,0,182,0,0,0,238,0,96,0,158,0,0,0,107,0,90,0,166,0,252,0,64,0,250,0,216,0,208,0,127,0,0,0,0,0,124,0,226,0,30,0,185,0,62,0,0,0,27,0,97,0,162,0,76,0,35,0,143,0,0,0,0,0,37,0,8,0,199,0,135,0,228,0,230,0,214,0,235,0,117,0,110,0,79,0,54,0,186,0,141,0,191,0,0,0,151,0,251,0,1,0,224,0,0,0,157,0,65,0,151,0,0,0,239,0,120,0,228,0,0,0,215,0,143,0,83,0,90,0,34,0,96,0,149,0,79,0,160,0,28,0,247,0,6,0,0,0,7,0,145,0,122,0,160,0,0,0,254,0,61,0,0,0,28,0,0,0,83,0,7,0,109,0,53,0,0,0,97,0,44,0,168,0,0,0,65,0,129,0,162,0,7,0,197,0,0,0,199,0,80,0,83,0,0,0,247,0,64,0,0,0,0,0,19,0,207,0,0,0,97,0,91,0,10,0,16,0,98,0,130,0,0,0,227,0,121,0,0,0,228,0,202,0,236,0,75,0,43,0,0,0,33,0,213,0,0,0,70,0,79,0,172,0,42,0,0,0,84,0,98,0,8,0,18,0,54,0,144,0,0,0,0,0,60,0,116,0,132,0,2,0,211,0,80,0,192,0,139,0,158,0,64,0,112,0,187,0,133,0,251,0,158,0,0,0,160,0,91,0,134,0,152,0,5,0,228,0,205,0,134,0,51,0,75,0,6,0,0,0,153,0,188,0,89,0,17,0,81,0,135,0,73,0,197,0,121,0,86,0,128,0,0,0,116,0,0,0,191,0,129,0,2,0,134,0,60,0,0,0,23,0,0,0,0,0,0,0,238,0,17,0,132,0,0,0,115,0,134,0,18,0,192,0,111,0,156,0,119,0,0,0,254,0,184,0,83,0,158,0,87,0,111,0,33,0,173,0,136,0,97,0,0,0,218,0,140,0,131,0,93,0,0,0,78,0,44,0,46,0,0,0,168,0,154,0,0,0,192,0,0,0,92,0,225,0,134,0,246,0,98,0,97,0,0,0,54,0,193,0,198,0,0,0,17,0,130,0,0,0,181,0,0,0,82,0,134,0,57,0,0,0,0,0,62,0,53,0,247,0,0,0,187,0,76,0,6,0,0,0,211,0,252,0,235,0,108,0,155,0,19,0,151,0,95,0,42,0,96,0,241,0,224,0,28,0,77,0,123,0,0,0,29,0,112,0,0,0,0,0,81,0,74,0,0,0,0,0,175,0,0,0,185,0,18,0,123,0,85,0,81,0,117,0,157,0,0,0,60,0,198,0,21,0,155,0,78,0,49,0,26,0,254,0,90,0,106,0,197,0,7,0,0,0,0,0,101,0,68,0,67,0,0,0,79,0,235,0,103,0,204,0,137,0,227,0,23,0,26,0,55,0,0,0,92,0,239,0,0,0,213,0,33,0,89,0,233,0,11,0,234,0,172,0,0,0,0,0,47,0,121,0,137,0,0,0,114,0,191,0,58,0,49,0,14,0,0,0,8,0,97,0,0,0,0,0,148,0,175,0,74,0,0,0,0,0,0,0,163,0,214,0,173,0,115,0,247,0,54,0,115,0,196,0,22,0,8,0,136,0,213,0,67,0,0,0,0,0,33,0,105,0,213,0,252,0,49,0,91,0,162,0,149,0,237,0,164,0,0,0,145,0,26,0,0,0,157,0,199,0,18,0,130,0,176,0,225,0,126,0,181,0,73,0,254,0,59,0,0,0,46,0,221,0,65,0,201,0,0,0,39,0,237,0,22,0,0,0,124,0,27,0,233,0,99,0,53,0,37,0,201,0,138,0,0,0,0,0,45,0,47,0,17,0,189,0,129,0,230,0,22,0,133,0,0,0,0,0,57,0,34,0,0,0,0,0,115,0,116,0,13,0,159,0,64,0,0,0,154,0,219,0,185,0,108,0,0,0,59,0,227,0,196,0,23,0,159,0,13,0,32,0,139,0,0,0,130,0,142,0,197,0,148,0,80,0,0,0,188,0,0,0,110,0,181,0,0,0,194,0,241,0,64,0,0,0,14,0,0,0,0,0,41,0,0,0,222,0,183,0,0,0,0,0,62,0,100,0,122,0,242,0,63,0,20,0,166,0,225,0,250,0,93,0,239,0,236,0,168,0,53,0,188,0,60,0,85,0,198,0,158,0,71,0,65,0,0,0,87,0,10,0,67,0,0,0,146,0,2,0,49,0,72,0,254,0,0,0,104,0,0,0,3,0,239,0,0,0,48,0,196,0,10,0,15,0,48,0,88,0,59,0,0,0,0,0,68,0,124,0,145,0,158,0,67,0,0,0,169,0,6,0,99,0,0,0,74,0,149,0,129,0,220,0,0,0,153,0,112,0,111,0,126,0,100,0,240,0,6,0,0,0,34,0,45,0,91,0,0,0,114,0,0,0,0,0,212,0,61,0,62,0,90,0,102,0,153,0,38,0,189,0,87,0,68,0,99,0,44,0,0,0,115,0,252,0,77,0,0,0,197,0,141,0,0,0,63,0,184,0,140,0,93,0,4,0,76,0,139,0,78,0,216,0,17,0,86,0,173,0,114,0,75,0,241,0,9,0,21,0,241,0,0,0,16,0,79,0,11,0,214,0,233,0,99,0,112,0,179,0,0,0,33,0,168,0,193,0,109,0,0,0,90,0,132,0,0,0,0,0,242,0,134,0,31,0,0,0,58,0,180,0,243,0,5,0,117,0,153,0,1,0,0,0,184,0,223,0,237,0,226,0,0,0,0,0,51,0,0,0,1,0,195,0,146,0,0,0,208,0,71,0,120,0,6,0,121,0,0,0,132,0,208,0,26,0,158,0,0,0,15,0,239,0,216,0,0,0,61,0,0,0,77,0,85,0,176,0,163,0,245,0,158,0,54,0,0,0,47,0,0,0,0,0,166,0,0,0,239,0,64,0,189,0,47,0,59,0,199,0,0,0,161,0,110,0,30,0,176,0,233,0,114,0,234,0,65,0);
signal scenario_full  : scenario_type := (0,0,28,31,28,30,71,31,71,30,71,29,241,31,82,31,82,30,147,31,147,30,130,31,228,31,33,31,188,31,37,31,211,31,211,30,211,29,111,31,147,31,107,31,195,31,110,31,110,30,110,29,227,31,227,30,58,31,58,30,147,31,147,30,147,29,68,31,105,31,168,31,27,31,227,31,252,31,63,31,14,31,14,30,217,31,22,31,6,31,168,31,32,31,32,30,32,31,184,31,69,31,230,31,230,30,95,31,95,30,71,31,38,31,220,31,220,30,219,31,219,30,191,31,131,31,131,30,41,31,30,31,145,31,241,31,182,31,200,31,30,31,30,30,209,31,174,31,204,31,3,31,41,31,37,31,2,31,119,31,158,31,14,31,31,31,211,31,194,31,37,31,244,31,244,30,201,31,201,30,176,31,107,31,169,31,40,31,136,31,198,31,198,30,20,31,2,31,134,31,154,31,247,31,114,31,114,30,124,31,97,31,76,31,113,31,113,30,60,31,31,31,223,31,63,31,75,31,172,31,40,31,126,31,76,31,26,31,26,30,229,31,229,30,144,31,25,31,56,31,10,31,37,31,105,31,28,31,57,31,57,30,154,31,151,31,106,31,89,31,51,31,219,31,17,31,17,30,65,31,65,30,217,31,78,31,106,31,59,31,130,31,104,31,201,31,201,30,207,31,177,31,227,31,124,31,180,31,189,31,101,31,120,31,38,31,195,31,195,30,47,31,51,31,174,31,101,31,10,31,10,30,11,31,103,31,103,30,228,31,89,31,128,31,60,31,180,31,180,30,219,31,200,31,152,31,199,31,186,31,186,30,177,31,185,31,100,31,167,31,151,31,138,31,99,31,174,31,174,30,174,29,237,31,10,31,10,30,17,31,170,31,152,31,199,31,83,31,129,31,182,31,182,30,238,31,96,31,158,31,158,30,107,31,90,31,166,31,252,31,64,31,250,31,216,31,208,31,127,31,127,30,127,29,124,31,226,31,30,31,185,31,62,31,62,30,27,31,97,31,162,31,76,31,35,31,143,31,143,30,143,29,37,31,8,31,199,31,135,31,228,31,230,31,214,31,235,31,117,31,110,31,79,31,54,31,186,31,141,31,191,31,191,30,151,31,251,31,1,31,224,31,224,30,157,31,65,31,151,31,151,30,239,31,120,31,228,31,228,30,215,31,143,31,83,31,90,31,34,31,96,31,149,31,79,31,160,31,28,31,247,31,6,31,6,30,7,31,145,31,122,31,160,31,160,30,254,31,61,31,61,30,28,31,28,30,83,31,7,31,109,31,53,31,53,30,97,31,44,31,168,31,168,30,65,31,129,31,162,31,7,31,197,31,197,30,199,31,80,31,83,31,83,30,247,31,64,31,64,30,64,29,19,31,207,31,207,30,97,31,91,31,10,31,16,31,98,31,130,31,130,30,227,31,121,31,121,30,228,31,202,31,236,31,75,31,43,31,43,30,33,31,213,31,213,30,70,31,79,31,172,31,42,31,42,30,84,31,98,31,8,31,18,31,54,31,144,31,144,30,144,29,60,31,116,31,132,31,2,31,211,31,80,31,192,31,139,31,158,31,64,31,112,31,187,31,133,31,251,31,158,31,158,30,160,31,91,31,134,31,152,31,5,31,228,31,205,31,134,31,51,31,75,31,6,31,6,30,153,31,188,31,89,31,17,31,81,31,135,31,73,31,197,31,121,31,86,31,128,31,128,30,116,31,116,30,191,31,129,31,2,31,134,31,60,31,60,30,23,31,23,30,23,29,23,28,238,31,17,31,132,31,132,30,115,31,134,31,18,31,192,31,111,31,156,31,119,31,119,30,254,31,184,31,83,31,158,31,87,31,111,31,33,31,173,31,136,31,97,31,97,30,218,31,140,31,131,31,93,31,93,30,78,31,44,31,46,31,46,30,168,31,154,31,154,30,192,31,192,30,92,31,225,31,134,31,246,31,98,31,97,31,97,30,54,31,193,31,198,31,198,30,17,31,130,31,130,30,181,31,181,30,82,31,134,31,57,31,57,30,57,29,62,31,53,31,247,31,247,30,187,31,76,31,6,31,6,30,211,31,252,31,235,31,108,31,155,31,19,31,151,31,95,31,42,31,96,31,241,31,224,31,28,31,77,31,123,31,123,30,29,31,112,31,112,30,112,29,81,31,74,31,74,30,74,29,175,31,175,30,185,31,18,31,123,31,85,31,81,31,117,31,157,31,157,30,60,31,198,31,21,31,155,31,78,31,49,31,26,31,254,31,90,31,106,31,197,31,7,31,7,30,7,29,101,31,68,31,67,31,67,30,79,31,235,31,103,31,204,31,137,31,227,31,23,31,26,31,55,31,55,30,92,31,239,31,239,30,213,31,33,31,89,31,233,31,11,31,234,31,172,31,172,30,172,29,47,31,121,31,137,31,137,30,114,31,191,31,58,31,49,31,14,31,14,30,8,31,97,31,97,30,97,29,148,31,175,31,74,31,74,30,74,29,74,28,163,31,214,31,173,31,115,31,247,31,54,31,115,31,196,31,22,31,8,31,136,31,213,31,67,31,67,30,67,29,33,31,105,31,213,31,252,31,49,31,91,31,162,31,149,31,237,31,164,31,164,30,145,31,26,31,26,30,157,31,199,31,18,31,130,31,176,31,225,31,126,31,181,31,73,31,254,31,59,31,59,30,46,31,221,31,65,31,201,31,201,30,39,31,237,31,22,31,22,30,124,31,27,31,233,31,99,31,53,31,37,31,201,31,138,31,138,30,138,29,45,31,47,31,17,31,189,31,129,31,230,31,22,31,133,31,133,30,133,29,57,31,34,31,34,30,34,29,115,31,116,31,13,31,159,31,64,31,64,30,154,31,219,31,185,31,108,31,108,30,59,31,227,31,196,31,23,31,159,31,13,31,32,31,139,31,139,30,130,31,142,31,197,31,148,31,80,31,80,30,188,31,188,30,110,31,181,31,181,30,194,31,241,31,64,31,64,30,14,31,14,30,14,29,41,31,41,30,222,31,183,31,183,30,183,29,62,31,100,31,122,31,242,31,63,31,20,31,166,31,225,31,250,31,93,31,239,31,236,31,168,31,53,31,188,31,60,31,85,31,198,31,158,31,71,31,65,31,65,30,87,31,10,31,67,31,67,30,146,31,2,31,49,31,72,31,254,31,254,30,104,31,104,30,3,31,239,31,239,30,48,31,196,31,10,31,15,31,48,31,88,31,59,31,59,30,59,29,68,31,124,31,145,31,158,31,67,31,67,30,169,31,6,31,99,31,99,30,74,31,149,31,129,31,220,31,220,30,153,31,112,31,111,31,126,31,100,31,240,31,6,31,6,30,34,31,45,31,91,31,91,30,114,31,114,30,114,29,212,31,61,31,62,31,90,31,102,31,153,31,38,31,189,31,87,31,68,31,99,31,44,31,44,30,115,31,252,31,77,31,77,30,197,31,141,31,141,30,63,31,184,31,140,31,93,31,4,31,76,31,139,31,78,31,216,31,17,31,86,31,173,31,114,31,75,31,241,31,9,31,21,31,241,31,241,30,16,31,79,31,11,31,214,31,233,31,99,31,112,31,179,31,179,30,33,31,168,31,193,31,109,31,109,30,90,31,132,31,132,30,132,29,242,31,134,31,31,31,31,30,58,31,180,31,243,31,5,31,117,31,153,31,1,31,1,30,184,31,223,31,237,31,226,31,226,30,226,29,51,31,51,30,1,31,195,31,146,31,146,30,208,31,71,31,120,31,6,31,121,31,121,30,132,31,208,31,26,31,158,31,158,30,15,31,239,31,216,31,216,30,61,31,61,30,77,31,85,31,176,31,163,31,245,31,158,31,54,31,54,30,47,31,47,30,47,29,166,31,166,30,239,31,64,31,189,31,47,31,59,31,199,31,199,30,161,31,110,31,30,31,176,31,233,31,114,31,234,31,65,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
