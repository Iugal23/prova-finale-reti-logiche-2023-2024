-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_159 is
end project_tb_159;

architecture project_tb_arch_159 of project_tb_159 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 928;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (65,0,205,0,9,0,4,0,2,0,0,0,187,0,238,0,0,0,56,0,184,0,6,0,193,0,28,0,0,0,228,0,121,0,137,0,0,0,253,0,0,0,162,0,211,0,0,0,5,0,248,0,25,0,76,0,194,0,226,0,162,0,12,0,0,0,7,0,166,0,202,0,233,0,0,0,109,0,128,0,143,0,245,0,11,0,14,0,0,0,189,0,134,0,168,0,69,0,4,0,159,0,107,0,133,0,235,0,0,0,60,0,0,0,165,0,189,0,0,0,255,0,194,0,0,0,236,0,0,0,165,0,59,0,186,0,101,0,0,0,0,0,136,0,0,0,0,0,7,0,55,0,0,0,115,0,0,0,19,0,216,0,111,0,156,0,131,0,143,0,111,0,38,0,66,0,0,0,0,0,207,0,18,0,0,0,126,0,10,0,39,0,200,0,0,0,169,0,208,0,190,0,0,0,0,0,176,0,155,0,124,0,109,0,0,0,143,0,14,0,1,0,156,0,232,0,244,0,217,0,32,0,248,0,141,0,0,0,0,0,69,0,117,0,153,0,253,0,213,0,182,0,118,0,45,0,189,0,81,0,94,0,22,0,197,0,28,0,90,0,213,0,203,0,99,0,249,0,21,0,90,0,79,0,0,0,80,0,0,0,124,0,158,0,0,0,145,0,141,0,132,0,225,0,96,0,0,0,75,0,210,0,187,0,74,0,128,0,72,0,223,0,0,0,0,0,84,0,111,0,156,0,97,0,46,0,0,0,220,0,24,0,0,0,181,0,6,0,197,0,0,0,3,0,154,0,0,0,138,0,187,0,105,0,107,0,236,0,137,0,159,0,0,0,0,0,250,0,247,0,215,0,0,0,162,0,247,0,223,0,51,0,57,0,0,0,132,0,174,0,47,0,0,0,136,0,0,0,96,0,216,0,198,0,192,0,0,0,0,0,19,0,234,0,53,0,46,0,221,0,235,0,237,0,83,0,200,0,55,0,109,0,98,0,93,0,73,0,134,0,174,0,111,0,122,0,92,0,245,0,41,0,0,0,2,0,0,0,218,0,0,0,166,0,213,0,9,0,23,0,0,0,243,0,0,0,172,0,187,0,178,0,48,0,30,0,182,0,248,0,24,0,50,0,216,0,212,0,6,0,253,0,203,0,84,0,2,0,145,0,245,0,103,0,166,0,0,0,240,0,94,0,231,0,100,0,156,0,160,0,176,0,144,0,103,0,190,0,1,0,33,0,0,0,218,0,88,0,232,0,21,0,2,0,160,0,114,0,12,0,132,0,252,0,96,0,46,0,139,0,96,0,54,0,141,0,250,0,220,0,45,0,207,0,206,0,244,0,0,0,8,0,44,0,4,0,50,0,20,0,105,0,87,0,0,0,58,0,204,0,0,0,24,0,83,0,200,0,153,0,4,0,232,0,0,0,182,0,254,0,230,0,145,0,170,0,64,0,198,0,187,0,178,0,88,0,16,0,129,0,32,0,15,0,0,0,0,0,221,0,72,0,0,0,96,0,254,0,0,0,15,0,192,0,165,0,56,0,0,0,180,0,0,0,0,0,188,0,111,0,102,0,131,0,0,0,93,0,249,0,0,0,77,0,249,0,35,0,149,0,88,0,70,0,154,0,185,0,73,0,54,0,57,0,184,0,233,0,248,0,147,0,89,0,175,0,201,0,181,0,0,0,0,0,4,0,67,0,3,0,248,0,216,0,155,0,167,0,189,0,165,0,98,0,147,0,149,0,161,0,0,0,227,0,0,0,213,0,0,0,107,0,121,0,170,0,61,0,19,0,136,0,16,0,232,0,247,0,0,0,182,0,30,0,82,0,0,0,200,0,240,0,22,0,48,0,114,0,111,0,121,0,21,0,186,0,0,0,7,0,55,0,43,0,243,0,200,0,161,0,139,0,50,0,0,0,140,0,168,0,178,0,151,0,148,0,223,0,137,0,47,0,14,0,144,0,51,0,134,0,143,0,169,0,54,0,28,0,0,0,254,0,0,0,86,0,85,0,182,0,162,0,0,0,25,0,0,0,0,0,0,0,128,0,0,0,0,0,27,0,13,0,237,0,17,0,151,0,97,0,0,0,49,0,227,0,208,0,0,0,108,0,0,0,128,0,91,0,4,0,9,0,111,0,24,0,0,0,123,0,94,0,186,0,0,0,0,0,219,0,140,0,0,0,87,0,150,0,191,0,0,0,94,0,0,0,178,0,35,0,35,0,3,0,32,0,172,0,32,0,192,0,0,0,221,0,97,0,51,0,39,0,14,0,193,0,104,0,0,0,20,0,0,0,205,0,0,0,149,0,58,0,175,0,96,0,219,0,61,0,186,0,126,0,17,0,70,0,121,0,86,0,0,0,247,0,202,0,71,0,59,0,233,0,121,0,54,0,159,0,225,0,0,0,0,0,82,0,198,0,70,0,153,0,144,0,249,0,165,0,123,0,133,0,143,0,213,0,214,0,233,0,42,0,28,0,181,0,164,0,0,0,81,0,95,0,154,0,186,0,0,0,93,0,77,0,75,0,120,0,18,0,214,0,190,0,0,0,0,0,155,0,120,0,169,0,19,0,0,0,33,0,191,0,133,0,125,0,191,0,0,0,96,0,0,0,93,0,227,0,74,0,0,0,38,0,254,0,0,0,0,0,185,0,0,0,159,0,41,0,0,0,8,0,151,0,24,0,122,0,58,0,0,0,171,0,74,0,145,0,9,0,75,0,156,0,226,0,189,0,224,0,184,0,198,0,91,0,25,0,50,0,124,0,188,0,0,0,15,0,43,0,80,0,222,0,160,0,37,0,197,0,0,0,146,0,0,0,164,0,93,0,0,0,254,0,0,0,179,0,0,0,131,0,95,0,236,0,19,0,26,0,235,0,240,0,92,0,50,0,172,0,43,0,197,0,22,0,85,0,244,0,200,0,0,0,205,0,0,0,201,0,205,0,87,0,130,0,217,0,94,0,0,0,60,0,62,0,163,0,163,0,0,0,0,0,81,0,159,0,131,0,0,0,0,0,122,0,0,0,215,0,31,0,134,0,168,0,0,0,181,0,242,0,0,0,168,0,26,0,214,0,0,0,0,0,88,0,103,0,254,0,0,0,151,0,176,0,102,0,236,0,168,0,179,0,178,0,167,0,245,0,0,0,96,0,69,0,226,0,0,0,35,0,142,0,132,0,75,0,22,0,114,0,0,0,242,0,177,0,0,0,0,0,131,0,219,0,0,0,154,0,140,0,68,0,223,0,88,0,189,0,0,0,243,0,33,0,223,0,213,0,0,0,66,0,186,0,158,0,188,0,92,0,158,0,159,0,226,0,21,0,137,0,42,0,223,0,232,0,247,0,175,0,171,0,76,0,164,0,190,0,105,0,107,0,78,0,3,0,63,0,113,0,133,0,108,0,222,0,0,0,140,0,160,0,191,0,0,0,0,0,50,0,205,0,30,0,51,0,0,0,183,0,153,0,183,0,0,0,95,0,185,0,41,0,5,0,218,0,38,0,0,0,189,0,240,0,74,0,128,0,24,0,76,0,0,0,70,0,147,0,106,0,0,0,229,0,2,0,0,0,97,0,0,0,95,0,0,0,61,0,254,0,79,0,207,0,186,0,232,0,98,0,249,0,35,0,101,0,62,0,0,0,120,0,0,0,188,0,30,0,0,0,90,0,181,0,0,0,129,0,161,0,0,0,0,0,0,0,71,0,119,0,217,0,230,0,0,0,10,0,0,0,17,0,0,0,83,0,173,0,183,0,239,0,168,0,167,0,0,0,83,0,48,0,45,0,176,0,0,0,117,0,150,0,86,0,231,0,4,0,20,0,70,0,0,0,93,0,0,0,148,0,247,0,131,0,0,0,0,0,234,0,0,0,0,0,78,0,234,0,59,0,17,0,0,0,231,0,169,0,135,0,93,0,46,0,68,0,155,0,127,0,146,0,252,0,0,0,0,0,85,0,0,0,223,0,1,0,82,0,0,0,30,0,225,0,177,0,110,0,113,0,51,0,0,0,126,0,121,0,133,0,254,0,120,0,60,0,175,0,119,0,7,0,59,0,201,0,232,0,74,0,0,0,0,0,117,0,12,0,152,0,0,0,54,0,226,0,1,0,0,0,113,0,102,0,0,0,87,0,209,0,125,0,235,0,101,0,207,0,225,0,122,0);
signal scenario_full  : scenario_type := (65,31,205,31,9,31,4,31,2,31,2,30,187,31,238,31,238,30,56,31,184,31,6,31,193,31,28,31,28,30,228,31,121,31,137,31,137,30,253,31,253,30,162,31,211,31,211,30,5,31,248,31,25,31,76,31,194,31,226,31,162,31,12,31,12,30,7,31,166,31,202,31,233,31,233,30,109,31,128,31,143,31,245,31,11,31,14,31,14,30,189,31,134,31,168,31,69,31,4,31,159,31,107,31,133,31,235,31,235,30,60,31,60,30,165,31,189,31,189,30,255,31,194,31,194,30,236,31,236,30,165,31,59,31,186,31,101,31,101,30,101,29,136,31,136,30,136,29,7,31,55,31,55,30,115,31,115,30,19,31,216,31,111,31,156,31,131,31,143,31,111,31,38,31,66,31,66,30,66,29,207,31,18,31,18,30,126,31,10,31,39,31,200,31,200,30,169,31,208,31,190,31,190,30,190,29,176,31,155,31,124,31,109,31,109,30,143,31,14,31,1,31,156,31,232,31,244,31,217,31,32,31,248,31,141,31,141,30,141,29,69,31,117,31,153,31,253,31,213,31,182,31,118,31,45,31,189,31,81,31,94,31,22,31,197,31,28,31,90,31,213,31,203,31,99,31,249,31,21,31,90,31,79,31,79,30,80,31,80,30,124,31,158,31,158,30,145,31,141,31,132,31,225,31,96,31,96,30,75,31,210,31,187,31,74,31,128,31,72,31,223,31,223,30,223,29,84,31,111,31,156,31,97,31,46,31,46,30,220,31,24,31,24,30,181,31,6,31,197,31,197,30,3,31,154,31,154,30,138,31,187,31,105,31,107,31,236,31,137,31,159,31,159,30,159,29,250,31,247,31,215,31,215,30,162,31,247,31,223,31,51,31,57,31,57,30,132,31,174,31,47,31,47,30,136,31,136,30,96,31,216,31,198,31,192,31,192,30,192,29,19,31,234,31,53,31,46,31,221,31,235,31,237,31,83,31,200,31,55,31,109,31,98,31,93,31,73,31,134,31,174,31,111,31,122,31,92,31,245,31,41,31,41,30,2,31,2,30,218,31,218,30,166,31,213,31,9,31,23,31,23,30,243,31,243,30,172,31,187,31,178,31,48,31,30,31,182,31,248,31,24,31,50,31,216,31,212,31,6,31,253,31,203,31,84,31,2,31,145,31,245,31,103,31,166,31,166,30,240,31,94,31,231,31,100,31,156,31,160,31,176,31,144,31,103,31,190,31,1,31,33,31,33,30,218,31,88,31,232,31,21,31,2,31,160,31,114,31,12,31,132,31,252,31,96,31,46,31,139,31,96,31,54,31,141,31,250,31,220,31,45,31,207,31,206,31,244,31,244,30,8,31,44,31,4,31,50,31,20,31,105,31,87,31,87,30,58,31,204,31,204,30,24,31,83,31,200,31,153,31,4,31,232,31,232,30,182,31,254,31,230,31,145,31,170,31,64,31,198,31,187,31,178,31,88,31,16,31,129,31,32,31,15,31,15,30,15,29,221,31,72,31,72,30,96,31,254,31,254,30,15,31,192,31,165,31,56,31,56,30,180,31,180,30,180,29,188,31,111,31,102,31,131,31,131,30,93,31,249,31,249,30,77,31,249,31,35,31,149,31,88,31,70,31,154,31,185,31,73,31,54,31,57,31,184,31,233,31,248,31,147,31,89,31,175,31,201,31,181,31,181,30,181,29,4,31,67,31,3,31,248,31,216,31,155,31,167,31,189,31,165,31,98,31,147,31,149,31,161,31,161,30,227,31,227,30,213,31,213,30,107,31,121,31,170,31,61,31,19,31,136,31,16,31,232,31,247,31,247,30,182,31,30,31,82,31,82,30,200,31,240,31,22,31,48,31,114,31,111,31,121,31,21,31,186,31,186,30,7,31,55,31,43,31,243,31,200,31,161,31,139,31,50,31,50,30,140,31,168,31,178,31,151,31,148,31,223,31,137,31,47,31,14,31,144,31,51,31,134,31,143,31,169,31,54,31,28,31,28,30,254,31,254,30,86,31,85,31,182,31,162,31,162,30,25,31,25,30,25,29,25,28,128,31,128,30,128,29,27,31,13,31,237,31,17,31,151,31,97,31,97,30,49,31,227,31,208,31,208,30,108,31,108,30,128,31,91,31,4,31,9,31,111,31,24,31,24,30,123,31,94,31,186,31,186,30,186,29,219,31,140,31,140,30,87,31,150,31,191,31,191,30,94,31,94,30,178,31,35,31,35,31,3,31,32,31,172,31,32,31,192,31,192,30,221,31,97,31,51,31,39,31,14,31,193,31,104,31,104,30,20,31,20,30,205,31,205,30,149,31,58,31,175,31,96,31,219,31,61,31,186,31,126,31,17,31,70,31,121,31,86,31,86,30,247,31,202,31,71,31,59,31,233,31,121,31,54,31,159,31,225,31,225,30,225,29,82,31,198,31,70,31,153,31,144,31,249,31,165,31,123,31,133,31,143,31,213,31,214,31,233,31,42,31,28,31,181,31,164,31,164,30,81,31,95,31,154,31,186,31,186,30,93,31,77,31,75,31,120,31,18,31,214,31,190,31,190,30,190,29,155,31,120,31,169,31,19,31,19,30,33,31,191,31,133,31,125,31,191,31,191,30,96,31,96,30,93,31,227,31,74,31,74,30,38,31,254,31,254,30,254,29,185,31,185,30,159,31,41,31,41,30,8,31,151,31,24,31,122,31,58,31,58,30,171,31,74,31,145,31,9,31,75,31,156,31,226,31,189,31,224,31,184,31,198,31,91,31,25,31,50,31,124,31,188,31,188,30,15,31,43,31,80,31,222,31,160,31,37,31,197,31,197,30,146,31,146,30,164,31,93,31,93,30,254,31,254,30,179,31,179,30,131,31,95,31,236,31,19,31,26,31,235,31,240,31,92,31,50,31,172,31,43,31,197,31,22,31,85,31,244,31,200,31,200,30,205,31,205,30,201,31,205,31,87,31,130,31,217,31,94,31,94,30,60,31,62,31,163,31,163,31,163,30,163,29,81,31,159,31,131,31,131,30,131,29,122,31,122,30,215,31,31,31,134,31,168,31,168,30,181,31,242,31,242,30,168,31,26,31,214,31,214,30,214,29,88,31,103,31,254,31,254,30,151,31,176,31,102,31,236,31,168,31,179,31,178,31,167,31,245,31,245,30,96,31,69,31,226,31,226,30,35,31,142,31,132,31,75,31,22,31,114,31,114,30,242,31,177,31,177,30,177,29,131,31,219,31,219,30,154,31,140,31,68,31,223,31,88,31,189,31,189,30,243,31,33,31,223,31,213,31,213,30,66,31,186,31,158,31,188,31,92,31,158,31,159,31,226,31,21,31,137,31,42,31,223,31,232,31,247,31,175,31,171,31,76,31,164,31,190,31,105,31,107,31,78,31,3,31,63,31,113,31,133,31,108,31,222,31,222,30,140,31,160,31,191,31,191,30,191,29,50,31,205,31,30,31,51,31,51,30,183,31,153,31,183,31,183,30,95,31,185,31,41,31,5,31,218,31,38,31,38,30,189,31,240,31,74,31,128,31,24,31,76,31,76,30,70,31,147,31,106,31,106,30,229,31,2,31,2,30,97,31,97,30,95,31,95,30,61,31,254,31,79,31,207,31,186,31,232,31,98,31,249,31,35,31,101,31,62,31,62,30,120,31,120,30,188,31,30,31,30,30,90,31,181,31,181,30,129,31,161,31,161,30,161,29,161,28,71,31,119,31,217,31,230,31,230,30,10,31,10,30,17,31,17,30,83,31,173,31,183,31,239,31,168,31,167,31,167,30,83,31,48,31,45,31,176,31,176,30,117,31,150,31,86,31,231,31,4,31,20,31,70,31,70,30,93,31,93,30,148,31,247,31,131,31,131,30,131,29,234,31,234,30,234,29,78,31,234,31,59,31,17,31,17,30,231,31,169,31,135,31,93,31,46,31,68,31,155,31,127,31,146,31,252,31,252,30,252,29,85,31,85,30,223,31,1,31,82,31,82,30,30,31,225,31,177,31,110,31,113,31,51,31,51,30,126,31,121,31,133,31,254,31,120,31,60,31,175,31,119,31,7,31,59,31,201,31,232,31,74,31,74,30,74,29,117,31,12,31,152,31,152,30,54,31,226,31,1,31,1,30,113,31,102,31,102,30,87,31,209,31,125,31,235,31,101,31,207,31,225,31,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
