-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_341 is
end project_tb_341;

architecture project_tb_arch_341 of project_tb_341 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 746;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (164,0,16,0,0,0,213,0,185,0,167,0,0,0,205,0,250,0,133,0,0,0,210,0,0,0,18,0,84,0,154,0,96,0,103,0,186,0,148,0,221,0,0,0,37,0,205,0,118,0,152,0,178,0,178,0,0,0,236,0,153,0,0,0,204,0,99,0,0,0,205,0,205,0,64,0,238,0,205,0,0,0,0,0,80,0,35,0,0,0,10,0,0,0,232,0,0,0,78,0,38,0,139,0,66,0,59,0,247,0,194,0,62,0,217,0,210,0,36,0,235,0,111,0,0,0,91,0,0,0,177,0,161,0,192,0,138,0,60,0,7,0,124,0,19,0,106,0,205,0,85,0,39,0,16,0,0,0,92,0,193,0,217,0,29,0,139,0,254,0,198,0,9,0,0,0,26,0,24,0,192,0,194,0,199,0,41,0,232,0,6,0,0,0,224,0,0,0,0,0,129,0,119,0,0,0,38,0,0,0,173,0,178,0,0,0,136,0,191,0,223,0,13,0,68,0,6,0,0,0,168,0,0,0,246,0,238,0,185,0,50,0,72,0,5,0,72,0,96,0,238,0,118,0,226,0,37,0,195,0,78,0,0,0,179,0,121,0,195,0,0,0,227,0,222,0,235,0,88,0,87,0,212,0,233,0,56,0,0,0,229,0,209,0,0,0,0,0,176,0,161,0,0,0,212,0,22,0,17,0,33,0,121,0,96,0,171,0,242,0,134,0,0,0,153,0,0,0,81,0,0,0,92,0,24,0,75,0,15,0,44,0,99,0,206,0,12,0,81,0,76,0,97,0,0,0,0,0,158,0,241,0,225,0,187,0,148,0,0,0,63,0,247,0,253,0,209,0,150,0,0,0,97,0,67,0,81,0,0,0,220,0,40,0,169,0,28,0,245,0,98,0,203,0,0,0,242,0,0,0,62,0,189,0,0,0,0,0,53,0,99,0,247,0,57,0,0,0,85,0,250,0,0,0,235,0,160,0,249,0,103,0,0,0,0,0,219,0,0,0,58,0,0,0,171,0,210,0,83,0,32,0,185,0,215,0,219,0,201,0,44,0,169,0,223,0,0,0,63,0,104,0,150,0,0,0,0,0,249,0,40,0,0,0,3,0,57,0,253,0,0,0,240,0,246,0,157,0,162,0,177,0,228,0,92,0,5,0,159,0,0,0,0,0,107,0,49,0,0,0,21,0,0,0,0,0,61,0,0,0,212,0,56,0,8,0,206,0,89,0,0,0,155,0,74,0,93,0,5,0,0,0,28,0,89,0,190,0,193,0,52,0,205,0,143,0,132,0,19,0,194,0,0,0,81,0,0,0,221,0,0,0,44,0,0,0,54,0,83,0,120,0,0,0,182,0,0,0,238,0,147,0,130,0,158,0,155,0,237,0,62,0,255,0,74,0,67,0,0,0,0,0,183,0,143,0,0,0,252,0,180,0,78,0,169,0,233,0,64,0,171,0,228,0,88,0,35,0,0,0,103,0,117,0,202,0,25,0,10,0,40,0,13,0,186,0,0,0,32,0,103,0,79,0,0,0,134,0,0,0,0,0,204,0,182,0,169,0,42,0,7,0,199,0,173,0,196,0,152,0,0,0,0,0,0,0,212,0,61,0,233,0,136,0,85,0,174,0,0,0,4,0,100,0,78,0,133,0,240,0,76,0,109,0,0,0,248,0,0,0,13,0,137,0,149,0,14,0,166,0,182,0,147,0,27,0,100,0,138,0,211,0,208,0,40,0,0,0,0,0,223,0,191,0,173,0,0,0,83,0,113,0,214,0,162,0,144,0,73,0,150,0,187,0,105,0,90,0,195,0,91,0,0,0,241,0,14,0,140,0,148,0,247,0,39,0,97,0,162,0,217,0,162,0,203,0,15,0,255,0,189,0,19,0,0,0,81,0,177,0,60,0,0,0,195,0,253,0,179,0,0,0,189,0,0,0,0,0,85,0,0,0,75,0,195,0,87,0,208,0,30,0,217,0,243,0,181,0,213,0,100,0,0,0,186,0,16,0,177,0,200,0,110,0,246,0,37,0,88,0,95,0,0,0,229,0,131,0,34,0,0,0,204,0,0,0,145,0,0,0,243,0,0,0,103,0,0,0,90,0,0,0,0,0,195,0,0,0,127,0,0,0,221,0,116,0,129,0,157,0,31,0,234,0,92,0,0,0,56,0,23,0,30,0,170,0,6,0,102,0,129,0,98,0,24,0,205,0,16,0,48,0,57,0,89,0,5,0,110,0,37,0,0,0,111,0,187,0,185,0,41,0,21,0,0,0,171,0,151,0,247,0,199,0,4,0,25,0,100,0,219,0,173,0,245,0,0,0,225,0,245,0,195,0,7,0,237,0,0,0,242,0,79,0,142,0,2,0,168,0,246,0,0,0,220,0,98,0,243,0,114,0,4,0,240,0,70,0,11,0,161,0,227,0,245,0,26,0,56,0,113,0,175,0,178,0,187,0,4,0,29,0,0,0,245,0,43,0,12,0,248,0,74,0,100,0,145,0,239,0,178,0,101,0,0,0,60,0,138,0,0,0,124,0,186,0,19,0,0,0,131,0,7,0,208,0,180,0,20,0,55,0,122,0,14,0,73,0,31,0,0,0,64,0,166,0,0,0,44,0,202,0,36,0,0,0,110,0,226,0,176,0,0,0,0,0,208,0,170,0,255,0,178,0,214,0,32,0,43,0,160,0,162,0,81,0,0,0,224,0,123,0,78,0,12,0,106,0,11,0,0,0,175,0,210,0,183,0,0,0,133,0,199,0,71,0,0,0,104,0,205,0,159,0,138,0,218,0,167,0,0,0,110,0,66,0,136,0,220,0,186,0,204,0,0,0,120,0,96,0,37,0,10,0,0,0,141,0,142,0,0,0,16,0,77,0,0,0,226,0,0,0,155,0,117,0,42,0,134,0,159,0,0,0,162,0,36,0,83,0,0,0,219,0,111,0,212,0,19,0,252,0,0,0,44,0,127,0,191,0,161,0,200,0,0,0,19,0,199,0,245,0,0,0,208,0,96,0,187,0,0,0,19,0,129,0,204,0,87,0,235,0,0,0,100,0,0,0,0,0,174,0,178,0,0,0,29,0,150,0,23,0,220,0,219,0,0,0,0,0,64,0,241,0,60,0,57,0,156,0,130,0,44,0,0,0,177,0,235,0,190,0,0,0,0,0,0,0,119,0,137,0,219,0,179,0,172,0,72,0,221,0,4,0,205,0,24,0,64,0,62,0,74,0,0,0,0,0,170,0,0,0,129,0,151,0,222,0,224,0,216,0,56,0,111,0,56,0,171,0,148,0,222,0,0,0,25,0,110,0,105,0,175,0,2,0,206,0,220,0,3,0);
signal scenario_full  : scenario_type := (164,31,16,31,16,30,213,31,185,31,167,31,167,30,205,31,250,31,133,31,133,30,210,31,210,30,18,31,84,31,154,31,96,31,103,31,186,31,148,31,221,31,221,30,37,31,205,31,118,31,152,31,178,31,178,31,178,30,236,31,153,31,153,30,204,31,99,31,99,30,205,31,205,31,64,31,238,31,205,31,205,30,205,29,80,31,35,31,35,30,10,31,10,30,232,31,232,30,78,31,38,31,139,31,66,31,59,31,247,31,194,31,62,31,217,31,210,31,36,31,235,31,111,31,111,30,91,31,91,30,177,31,161,31,192,31,138,31,60,31,7,31,124,31,19,31,106,31,205,31,85,31,39,31,16,31,16,30,92,31,193,31,217,31,29,31,139,31,254,31,198,31,9,31,9,30,26,31,24,31,192,31,194,31,199,31,41,31,232,31,6,31,6,30,224,31,224,30,224,29,129,31,119,31,119,30,38,31,38,30,173,31,178,31,178,30,136,31,191,31,223,31,13,31,68,31,6,31,6,30,168,31,168,30,246,31,238,31,185,31,50,31,72,31,5,31,72,31,96,31,238,31,118,31,226,31,37,31,195,31,78,31,78,30,179,31,121,31,195,31,195,30,227,31,222,31,235,31,88,31,87,31,212,31,233,31,56,31,56,30,229,31,209,31,209,30,209,29,176,31,161,31,161,30,212,31,22,31,17,31,33,31,121,31,96,31,171,31,242,31,134,31,134,30,153,31,153,30,81,31,81,30,92,31,24,31,75,31,15,31,44,31,99,31,206,31,12,31,81,31,76,31,97,31,97,30,97,29,158,31,241,31,225,31,187,31,148,31,148,30,63,31,247,31,253,31,209,31,150,31,150,30,97,31,67,31,81,31,81,30,220,31,40,31,169,31,28,31,245,31,98,31,203,31,203,30,242,31,242,30,62,31,189,31,189,30,189,29,53,31,99,31,247,31,57,31,57,30,85,31,250,31,250,30,235,31,160,31,249,31,103,31,103,30,103,29,219,31,219,30,58,31,58,30,171,31,210,31,83,31,32,31,185,31,215,31,219,31,201,31,44,31,169,31,223,31,223,30,63,31,104,31,150,31,150,30,150,29,249,31,40,31,40,30,3,31,57,31,253,31,253,30,240,31,246,31,157,31,162,31,177,31,228,31,92,31,5,31,159,31,159,30,159,29,107,31,49,31,49,30,21,31,21,30,21,29,61,31,61,30,212,31,56,31,8,31,206,31,89,31,89,30,155,31,74,31,93,31,5,31,5,30,28,31,89,31,190,31,193,31,52,31,205,31,143,31,132,31,19,31,194,31,194,30,81,31,81,30,221,31,221,30,44,31,44,30,54,31,83,31,120,31,120,30,182,31,182,30,238,31,147,31,130,31,158,31,155,31,237,31,62,31,255,31,74,31,67,31,67,30,67,29,183,31,143,31,143,30,252,31,180,31,78,31,169,31,233,31,64,31,171,31,228,31,88,31,35,31,35,30,103,31,117,31,202,31,25,31,10,31,40,31,13,31,186,31,186,30,32,31,103,31,79,31,79,30,134,31,134,30,134,29,204,31,182,31,169,31,42,31,7,31,199,31,173,31,196,31,152,31,152,30,152,29,152,28,212,31,61,31,233,31,136,31,85,31,174,31,174,30,4,31,100,31,78,31,133,31,240,31,76,31,109,31,109,30,248,31,248,30,13,31,137,31,149,31,14,31,166,31,182,31,147,31,27,31,100,31,138,31,211,31,208,31,40,31,40,30,40,29,223,31,191,31,173,31,173,30,83,31,113,31,214,31,162,31,144,31,73,31,150,31,187,31,105,31,90,31,195,31,91,31,91,30,241,31,14,31,140,31,148,31,247,31,39,31,97,31,162,31,217,31,162,31,203,31,15,31,255,31,189,31,19,31,19,30,81,31,177,31,60,31,60,30,195,31,253,31,179,31,179,30,189,31,189,30,189,29,85,31,85,30,75,31,195,31,87,31,208,31,30,31,217,31,243,31,181,31,213,31,100,31,100,30,186,31,16,31,177,31,200,31,110,31,246,31,37,31,88,31,95,31,95,30,229,31,131,31,34,31,34,30,204,31,204,30,145,31,145,30,243,31,243,30,103,31,103,30,90,31,90,30,90,29,195,31,195,30,127,31,127,30,221,31,116,31,129,31,157,31,31,31,234,31,92,31,92,30,56,31,23,31,30,31,170,31,6,31,102,31,129,31,98,31,24,31,205,31,16,31,48,31,57,31,89,31,5,31,110,31,37,31,37,30,111,31,187,31,185,31,41,31,21,31,21,30,171,31,151,31,247,31,199,31,4,31,25,31,100,31,219,31,173,31,245,31,245,30,225,31,245,31,195,31,7,31,237,31,237,30,242,31,79,31,142,31,2,31,168,31,246,31,246,30,220,31,98,31,243,31,114,31,4,31,240,31,70,31,11,31,161,31,227,31,245,31,26,31,56,31,113,31,175,31,178,31,187,31,4,31,29,31,29,30,245,31,43,31,12,31,248,31,74,31,100,31,145,31,239,31,178,31,101,31,101,30,60,31,138,31,138,30,124,31,186,31,19,31,19,30,131,31,7,31,208,31,180,31,20,31,55,31,122,31,14,31,73,31,31,31,31,30,64,31,166,31,166,30,44,31,202,31,36,31,36,30,110,31,226,31,176,31,176,30,176,29,208,31,170,31,255,31,178,31,214,31,32,31,43,31,160,31,162,31,81,31,81,30,224,31,123,31,78,31,12,31,106,31,11,31,11,30,175,31,210,31,183,31,183,30,133,31,199,31,71,31,71,30,104,31,205,31,159,31,138,31,218,31,167,31,167,30,110,31,66,31,136,31,220,31,186,31,204,31,204,30,120,31,96,31,37,31,10,31,10,30,141,31,142,31,142,30,16,31,77,31,77,30,226,31,226,30,155,31,117,31,42,31,134,31,159,31,159,30,162,31,36,31,83,31,83,30,219,31,111,31,212,31,19,31,252,31,252,30,44,31,127,31,191,31,161,31,200,31,200,30,19,31,199,31,245,31,245,30,208,31,96,31,187,31,187,30,19,31,129,31,204,31,87,31,235,31,235,30,100,31,100,30,100,29,174,31,178,31,178,30,29,31,150,31,23,31,220,31,219,31,219,30,219,29,64,31,241,31,60,31,57,31,156,31,130,31,44,31,44,30,177,31,235,31,190,31,190,30,190,29,190,28,119,31,137,31,219,31,179,31,172,31,72,31,221,31,4,31,205,31,24,31,64,31,62,31,74,31,74,30,74,29,170,31,170,30,129,31,151,31,222,31,224,31,216,31,56,31,111,31,56,31,171,31,148,31,222,31,222,30,25,31,110,31,105,31,175,31,2,31,206,31,220,31,3,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
