-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 636;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (38,0,255,0,97,0,112,0,64,0,178,0,0,0,108,0,11,0,0,0,16,0,230,0,88,0,70,0,112,0,243,0,246,0,250,0,39,0,0,0,114,0,0,0,39,0,181,0,0,0,205,0,198,0,95,0,175,0,7,0,119,0,0,0,220,0,225,0,0,0,200,0,0,0,95,0,0,0,0,0,6,0,239,0,207,0,0,0,244,0,91,0,96,0,144,0,82,0,18,0,110,0,127,0,81,0,157,0,30,0,166,0,223,0,121,0,188,0,220,0,121,0,0,0,0,0,235,0,7,0,220,0,63,0,0,0,165,0,201,0,28,0,239,0,76,0,17,0,14,0,238,0,0,0,0,0,32,0,0,0,2,0,0,0,116,0,206,0,24,0,204,0,45,0,33,0,79,0,0,0,70,0,247,0,0,0,82,0,81,0,246,0,21,0,156,0,151,0,241,0,77,0,0,0,218,0,35,0,0,0,121,0,0,0,171,0,153,0,0,0,0,0,0,0,0,0,112,0,140,0,211,0,1,0,51,0,166,0,114,0,240,0,52,0,53,0,60,0,193,0,201,0,148,0,160,0,241,0,175,0,237,0,0,0,0,0,101,0,195,0,0,0,76,0,237,0,189,0,128,0,14,0,48,0,125,0,0,0,0,0,0,0,137,0,0,0,142,0,174,0,3,0,151,0,214,0,0,0,0,0,121,0,252,0,250,0,48,0,194,0,211,0,189,0,197,0,241,0,77,0,99,0,221,0,0,0,53,0,15,0,30,0,50,0,177,0,241,0,243,0,27,0,0,0,107,0,0,0,23,0,31,0,76,0,168,0,25,0,0,0,55,0,196,0,47,0,15,0,187,0,202,0,237,0,16,0,172,0,67,0,0,0,0,0,241,0,0,0,0,0,0,0,120,0,247,0,116,0,151,0,233,0,102,0,84,0,139,0,152,0,158,0,4,0,171,0,2,0,25,0,3,0,144,0,0,0,30,0,125,0,134,0,0,0,77,0,147,0,244,0,145,0,92,0,24,0,80,0,93,0,153,0,178,0,157,0,81,0,181,0,215,0,230,0,188,0,0,0,169,0,222,0,9,0,38,0,0,0,161,0,160,0,171,0,34,0,0,0,37,0,0,0,193,0,176,0,43,0,145,0,47,0,104,0,166,0,216,0,0,0,50,0,108,0,0,0,0,0,181,0,44,0,0,0,132,0,126,0,77,0,254,0,7,0,221,0,158,0,46,0,174,0,80,0,0,0,14,0,98,0,244,0,237,0,165,0,0,0,1,0,126,0,137,0,242,0,28,0,118,0,67,0,159,0,0,0,0,0,252,0,138,0,0,0,80,0,251,0,119,0,0,0,141,0,204,0,125,0,190,0,148,0,153,0,188,0,75,0,188,0,196,0,214,0,0,0,118,0,149,0,58,0,215,0,153,0,0,0,0,0,6,0,76,0,0,0,46,0,121,0,14,0,0,0,34,0,160,0,0,0,0,0,251,0,45,0,109,0,0,0,0,0,36,0,0,0,79,0,93,0,143,0,178,0,0,0,223,0,6,0,247,0,184,0,9,0,147,0,198,0,57,0,164,0,152,0,170,0,0,0,176,0,83,0,85,0,110,0,134,0,249,0,83,0,134,0,61,0,14,0,110,0,7,0,191,0,88,0,0,0,132,0,167,0,37,0,80,0,17,0,237,0,0,0,216,0,82,0,0,0,153,0,100,0,188,0,252,0,0,0,96,0,225,0,180,0,232,0,237,0,165,0,218,0,165,0,128,0,11,0,129,0,0,0,85,0,0,0,154,0,0,0,95,0,0,0,0,0,204,0,211,0,0,0,189,0,22,0,76,0,208,0,110,0,172,0,0,0,158,0,95,0,0,0,163,0,54,0,151,0,14,0,55,0,190,0,26,0,0,0,210,0,227,0,0,0,111,0,104,0,35,0,0,0,35,0,97,0,57,0,93,0,224,0,0,0,213,0,250,0,241,0,197,0,88,0,79,0,0,0,0,0,84,0,0,0,85,0,211,0,93,0,109,0,16,0,6,0,135,0,108,0,241,0,0,0,0,0,39,0,12,0,115,0,55,0,0,0,0,0,187,0,253,0,187,0,179,0,219,0,0,0,175,0,21,0,0,0,0,0,151,0,57,0,227,0,0,0,236,0,125,0,213,0,0,0,97,0,1,0,39,0,89,0,100,0,184,0,129,0,0,0,170,0,193,0,92,0,5,0,33,0,0,0,167,0,35,0,46,0,151,0,153,0,0,0,0,0,133,0,220,0,81,0,210,0,65,0,39,0,0,0,173,0,53,0,0,0,125,0,89,0,0,0,220,0,120,0,180,0,109,0,26,0,193,0,64,0,0,0,173,0,15,0,63,0,26,0,84,0,0,0,69,0,39,0,219,0,0,0,252,0,57,0,219,0,0,0,203,0,171,0,0,0,198,0,0,0,0,0,99,0,44,0,99,0,0,0,246,0,226,0,96,0,0,0,107,0,175,0,130,0,187,0,118,0,146,0,0,0,132,0,108,0,193,0,53,0,182,0,44,0,210,0,26,0,210,0,115,0,136,0,189,0,181,0,0,0,0,0,243,0,0,0,68,0,0,0,239,0,250,0,14,0,0,0,34,0,239,0,37,0,62,0,231,0,5,0,198,0,244,0,203,0,68,0,189,0,170,0,0,0,114,0,107,0,136,0,104,0,190,0,0,0,181,0,0,0,98,0,197,0,187,0,0,0,159,0,6,0,43,0,0,0,188,0,159,0,0,0,62,0,103,0,194,0,206,0,172,0,250,0,162,0,228,0,27,0,0,0,74,0,205,0,27,0,19,0,78,0,119,0,0,0,53,0,241,0,22,0,118,0);
signal scenario_full  : scenario_type := (38,31,255,31,97,31,112,31,64,31,178,31,178,30,108,31,11,31,11,30,16,31,230,31,88,31,70,31,112,31,243,31,246,31,250,31,39,31,39,30,114,31,114,30,39,31,181,31,181,30,205,31,198,31,95,31,175,31,7,31,119,31,119,30,220,31,225,31,225,30,200,31,200,30,95,31,95,30,95,29,6,31,239,31,207,31,207,30,244,31,91,31,96,31,144,31,82,31,18,31,110,31,127,31,81,31,157,31,30,31,166,31,223,31,121,31,188,31,220,31,121,31,121,30,121,29,235,31,7,31,220,31,63,31,63,30,165,31,201,31,28,31,239,31,76,31,17,31,14,31,238,31,238,30,238,29,32,31,32,30,2,31,2,30,116,31,206,31,24,31,204,31,45,31,33,31,79,31,79,30,70,31,247,31,247,30,82,31,81,31,246,31,21,31,156,31,151,31,241,31,77,31,77,30,218,31,35,31,35,30,121,31,121,30,171,31,153,31,153,30,153,29,153,28,153,27,112,31,140,31,211,31,1,31,51,31,166,31,114,31,240,31,52,31,53,31,60,31,193,31,201,31,148,31,160,31,241,31,175,31,237,31,237,30,237,29,101,31,195,31,195,30,76,31,237,31,189,31,128,31,14,31,48,31,125,31,125,30,125,29,125,28,137,31,137,30,142,31,174,31,3,31,151,31,214,31,214,30,214,29,121,31,252,31,250,31,48,31,194,31,211,31,189,31,197,31,241,31,77,31,99,31,221,31,221,30,53,31,15,31,30,31,50,31,177,31,241,31,243,31,27,31,27,30,107,31,107,30,23,31,31,31,76,31,168,31,25,31,25,30,55,31,196,31,47,31,15,31,187,31,202,31,237,31,16,31,172,31,67,31,67,30,67,29,241,31,241,30,241,29,241,28,120,31,247,31,116,31,151,31,233,31,102,31,84,31,139,31,152,31,158,31,4,31,171,31,2,31,25,31,3,31,144,31,144,30,30,31,125,31,134,31,134,30,77,31,147,31,244,31,145,31,92,31,24,31,80,31,93,31,153,31,178,31,157,31,81,31,181,31,215,31,230,31,188,31,188,30,169,31,222,31,9,31,38,31,38,30,161,31,160,31,171,31,34,31,34,30,37,31,37,30,193,31,176,31,43,31,145,31,47,31,104,31,166,31,216,31,216,30,50,31,108,31,108,30,108,29,181,31,44,31,44,30,132,31,126,31,77,31,254,31,7,31,221,31,158,31,46,31,174,31,80,31,80,30,14,31,98,31,244,31,237,31,165,31,165,30,1,31,126,31,137,31,242,31,28,31,118,31,67,31,159,31,159,30,159,29,252,31,138,31,138,30,80,31,251,31,119,31,119,30,141,31,204,31,125,31,190,31,148,31,153,31,188,31,75,31,188,31,196,31,214,31,214,30,118,31,149,31,58,31,215,31,153,31,153,30,153,29,6,31,76,31,76,30,46,31,121,31,14,31,14,30,34,31,160,31,160,30,160,29,251,31,45,31,109,31,109,30,109,29,36,31,36,30,79,31,93,31,143,31,178,31,178,30,223,31,6,31,247,31,184,31,9,31,147,31,198,31,57,31,164,31,152,31,170,31,170,30,176,31,83,31,85,31,110,31,134,31,249,31,83,31,134,31,61,31,14,31,110,31,7,31,191,31,88,31,88,30,132,31,167,31,37,31,80,31,17,31,237,31,237,30,216,31,82,31,82,30,153,31,100,31,188,31,252,31,252,30,96,31,225,31,180,31,232,31,237,31,165,31,218,31,165,31,128,31,11,31,129,31,129,30,85,31,85,30,154,31,154,30,95,31,95,30,95,29,204,31,211,31,211,30,189,31,22,31,76,31,208,31,110,31,172,31,172,30,158,31,95,31,95,30,163,31,54,31,151,31,14,31,55,31,190,31,26,31,26,30,210,31,227,31,227,30,111,31,104,31,35,31,35,30,35,31,97,31,57,31,93,31,224,31,224,30,213,31,250,31,241,31,197,31,88,31,79,31,79,30,79,29,84,31,84,30,85,31,211,31,93,31,109,31,16,31,6,31,135,31,108,31,241,31,241,30,241,29,39,31,12,31,115,31,55,31,55,30,55,29,187,31,253,31,187,31,179,31,219,31,219,30,175,31,21,31,21,30,21,29,151,31,57,31,227,31,227,30,236,31,125,31,213,31,213,30,97,31,1,31,39,31,89,31,100,31,184,31,129,31,129,30,170,31,193,31,92,31,5,31,33,31,33,30,167,31,35,31,46,31,151,31,153,31,153,30,153,29,133,31,220,31,81,31,210,31,65,31,39,31,39,30,173,31,53,31,53,30,125,31,89,31,89,30,220,31,120,31,180,31,109,31,26,31,193,31,64,31,64,30,173,31,15,31,63,31,26,31,84,31,84,30,69,31,39,31,219,31,219,30,252,31,57,31,219,31,219,30,203,31,171,31,171,30,198,31,198,30,198,29,99,31,44,31,99,31,99,30,246,31,226,31,96,31,96,30,107,31,175,31,130,31,187,31,118,31,146,31,146,30,132,31,108,31,193,31,53,31,182,31,44,31,210,31,26,31,210,31,115,31,136,31,189,31,181,31,181,30,181,29,243,31,243,30,68,31,68,30,239,31,250,31,14,31,14,30,34,31,239,31,37,31,62,31,231,31,5,31,198,31,244,31,203,31,68,31,189,31,170,31,170,30,114,31,107,31,136,31,104,31,190,31,190,30,181,31,181,30,98,31,197,31,187,31,187,30,159,31,6,31,43,31,43,30,188,31,159,31,159,30,62,31,103,31,194,31,206,31,172,31,250,31,162,31,228,31,27,31,27,30,74,31,205,31,27,31,19,31,78,31,119,31,119,30,53,31,241,31,22,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
