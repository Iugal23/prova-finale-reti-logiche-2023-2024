-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 719;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,240,0,241,0,161,0,116,0,84,0,0,0,81,0,214,0,232,0,198,0,0,0,125,0,0,0,247,0,86,0,94,0,0,0,254,0,133,0,251,0,148,0,128,0,172,0,0,0,72,0,214,0,0,0,96,0,231,0,178,0,0,0,106,0,189,0,135,0,101,0,0,0,188,0,220,0,215,0,221,0,63,0,0,0,193,0,125,0,192,0,249,0,0,0,253,0,165,0,220,0,199,0,156,0,97,0,0,0,161,0,0,0,0,0,201,0,0,0,0,0,30,0,54,0,0,0,168,0,242,0,135,0,222,0,97,0,95,0,203,0,0,0,0,0,19,0,105,0,241,0,4,0,0,0,4,0,159,0,159,0,106,0,146,0,50,0,135,0,196,0,188,0,0,0,23,0,68,0,252,0,148,0,0,0,117,0,84,0,2,0,59,0,0,0,0,0,175,0,65,0,0,0,171,0,164,0,96,0,217,0,69,0,223,0,64,0,95,0,121,0,124,0,69,0,200,0,0,0,236,0,181,0,39,0,215,0,73,0,0,0,0,0,192,0,0,0,18,0,180,0,87,0,127,0,89,0,144,0,165,0,117,0,91,0,15,0,98,0,0,0,104,0,0,0,0,0,0,0,175,0,199,0,80,0,161,0,0,0,116,0,218,0,177,0,0,0,200,0,102,0,170,0,113,0,3,0,0,0,0,0,0,0,0,0,227,0,50,0,115,0,50,0,208,0,67,0,142,0,0,0,100,0,180,0,0,0,0,0,157,0,159,0,245,0,32,0,110,0,115,0,79,0,211,0,65,0,212,0,29,0,68,0,195,0,224,0,170,0,131,0,59,0,209,0,166,0,139,0,63,0,28,0,0,0,30,0,61,0,69,0,0,0,151,0,161,0,229,0,157,0,84,0,0,0,0,0,134,0,232,0,0,0,12,0,10,0,25,0,45,0,170,0,198,0,40,0,98,0,179,0,197,0,0,0,84,0,206,0,169,0,142,0,250,0,78,0,91,0,54,0,10,0,0,0,0,0,95,0,121,0,0,0,167,0,255,0,31,0,187,0,22,0,227,0,190,0,155,0,189,0,179,0,87,0,72,0,228,0,214,0,237,0,149,0,212,0,159,0,32,0,77,0,177,0,159,0,0,0,112,0,98,0,0,0,7,0,215,0,158,0,87,0,0,0,211,0,82,0,229,0,197,0,254,0,130,0,0,0,0,0,0,0,135,0,106,0,163,0,91,0,93,0,0,0,7,0,178,0,115,0,0,0,61,0,168,0,115,0,81,0,128,0,224,0,100,0,202,0,54,0,105,0,85,0,148,0,119,0,54,0,41,0,247,0,0,0,96,0,76,0,143,0,0,0,194,0,58,0,84,0,0,0,130,0,0,0,29,0,10,0,72,0,103,0,200,0,136,0,24,0,168,0,129,0,45,0,172,0,203,0,141,0,238,0,216,0,196,0,33,0,47,0,75,0,201,0,95,0,206,0,0,0,0,0,104,0,0,0,219,0,119,0,0,0,0,0,201,0,146,0,0,0,0,0,152,0,133,0,0,0,168,0,121,0,0,0,170,0,75,0,233,0,0,0,121,0,186,0,85,0,15,0,67,0,33,0,8,0,0,0,73,0,69,0,253,0,0,0,29,0,211,0,0,0,0,0,147,0,139,0,23,0,58,0,0,0,62,0,193,0,10,0,0,0,0,0,65,0,64,0,98,0,1,0,89,0,141,0,160,0,0,0,156,0,115,0,106,0,200,0,182,0,0,0,43,0,174,0,0,0,84,0,147,0,195,0,145,0,0,0,0,0,0,0,192,0,104,0,77,0,238,0,157,0,18,0,173,0,0,0,106,0,76,0,0,0,0,0,209,0,81,0,63,0,0,0,36,0,139,0,198,0,159,0,0,0,0,0,138,0,153,0,57,0,0,0,10,0,185,0,53,0,168,0,103,0,0,0,0,0,117,0,46,0,94,0,106,0,136,0,0,0,0,0,0,0,190,0,238,0,4,0,169,0,0,0,61,0,186,0,71,0,0,0,125,0,0,0,20,0,182,0,62,0,24,0,0,0,0,0,84,0,247,0,102,0,0,0,216,0,30,0,169,0,25,0,0,0,225,0,0,0,180,0,0,0,165,0,134,0,227,0,73,0,13,0,66,0,0,0,9,0,219,0,108,0,0,0,79,0,0,0,0,0,249,0,0,0,56,0,57,0,32,0,0,0,107,0,58,0,220,0,0,0,130,0,0,0,34,0,213,0,45,0,169,0,244,0,16,0,0,0,68,0,83,0,61,0,30,0,21,0,1,0,26,0,25,0,146,0,189,0,97,0,0,0,242,0,0,0,3,0,225,0,39,0,0,0,55,0,0,0,202,0,0,0,247,0,0,0,71,0,195,0,238,0,173,0,158,0,239,0,103,0,112,0,189,0,0,0,30,0,18,0,205,0,207,0,18,0,215,0,245,0,14,0,240,0,195,0,119,0,216,0,60,0,0,0,81,0,251,0,247,0,20,0,0,0,138,0,0,0,228,0,0,0,63,0,187,0,45,0,81,0,0,0,0,0,105,0,236,0,124,0,0,0,120,0,182,0,249,0,48,0,111,0,46,0,4,0,2,0,208,0,45,0,33,0,33,0,242,0,95,0,203,0,51,0,113,0,142,0,45,0,85,0,7,0,34,0,10,0,63,0,50,0,163,0,144,0,110,0,53,0,30,0,52,0,0,0,201,0,70,0,255,0,153,0,146,0,140,0,146,0,60,0,8,0,186,0,6,0,36,0,187,0,79,0,0,0,74,0,37,0,0,0,111,0,239,0,66,0,222,0,0,0,0,0,100,0,218,0,80,0,0,0,113,0,0,0,0,0,229,0,0,0,242,0,49,0,44,0,102,0,0,0,242,0,0,0,0,0,0,0,52,0,176,0,232,0,243,0,2,0,117,0,0,0,170,0,0,0,169,0,142,0,101,0,0,0,95,0,0,0,107,0,0,0,0,0,242,0,235,0,10,0,127,0,15,0,247,0,193,0,142,0,23,0,200,0,125,0,42,0,210,0,106,0,139,0,179,0,106,0,174,0,70,0,0,0,204,0,195,0,0,0,60,0,202,0,236,0,197,0,41,0,140,0,24,0,250,0,242,0,211,0,40,0,101,0,63,0,57,0,0,0,178,0,142,0,140,0,189,0,75,0,81,0,23,0,108,0,121,0,39,0,0,0,250,0,1,0,109,0,234,0);
signal scenario_full  : scenario_type := (135,31,240,31,241,31,161,31,116,31,84,31,84,30,81,31,214,31,232,31,198,31,198,30,125,31,125,30,247,31,86,31,94,31,94,30,254,31,133,31,251,31,148,31,128,31,172,31,172,30,72,31,214,31,214,30,96,31,231,31,178,31,178,30,106,31,189,31,135,31,101,31,101,30,188,31,220,31,215,31,221,31,63,31,63,30,193,31,125,31,192,31,249,31,249,30,253,31,165,31,220,31,199,31,156,31,97,31,97,30,161,31,161,30,161,29,201,31,201,30,201,29,30,31,54,31,54,30,168,31,242,31,135,31,222,31,97,31,95,31,203,31,203,30,203,29,19,31,105,31,241,31,4,31,4,30,4,31,159,31,159,31,106,31,146,31,50,31,135,31,196,31,188,31,188,30,23,31,68,31,252,31,148,31,148,30,117,31,84,31,2,31,59,31,59,30,59,29,175,31,65,31,65,30,171,31,164,31,96,31,217,31,69,31,223,31,64,31,95,31,121,31,124,31,69,31,200,31,200,30,236,31,181,31,39,31,215,31,73,31,73,30,73,29,192,31,192,30,18,31,180,31,87,31,127,31,89,31,144,31,165,31,117,31,91,31,15,31,98,31,98,30,104,31,104,30,104,29,104,28,175,31,199,31,80,31,161,31,161,30,116,31,218,31,177,31,177,30,200,31,102,31,170,31,113,31,3,31,3,30,3,29,3,28,3,27,227,31,50,31,115,31,50,31,208,31,67,31,142,31,142,30,100,31,180,31,180,30,180,29,157,31,159,31,245,31,32,31,110,31,115,31,79,31,211,31,65,31,212,31,29,31,68,31,195,31,224,31,170,31,131,31,59,31,209,31,166,31,139,31,63,31,28,31,28,30,30,31,61,31,69,31,69,30,151,31,161,31,229,31,157,31,84,31,84,30,84,29,134,31,232,31,232,30,12,31,10,31,25,31,45,31,170,31,198,31,40,31,98,31,179,31,197,31,197,30,84,31,206,31,169,31,142,31,250,31,78,31,91,31,54,31,10,31,10,30,10,29,95,31,121,31,121,30,167,31,255,31,31,31,187,31,22,31,227,31,190,31,155,31,189,31,179,31,87,31,72,31,228,31,214,31,237,31,149,31,212,31,159,31,32,31,77,31,177,31,159,31,159,30,112,31,98,31,98,30,7,31,215,31,158,31,87,31,87,30,211,31,82,31,229,31,197,31,254,31,130,31,130,30,130,29,130,28,135,31,106,31,163,31,91,31,93,31,93,30,7,31,178,31,115,31,115,30,61,31,168,31,115,31,81,31,128,31,224,31,100,31,202,31,54,31,105,31,85,31,148,31,119,31,54,31,41,31,247,31,247,30,96,31,76,31,143,31,143,30,194,31,58,31,84,31,84,30,130,31,130,30,29,31,10,31,72,31,103,31,200,31,136,31,24,31,168,31,129,31,45,31,172,31,203,31,141,31,238,31,216,31,196,31,33,31,47,31,75,31,201,31,95,31,206,31,206,30,206,29,104,31,104,30,219,31,119,31,119,30,119,29,201,31,146,31,146,30,146,29,152,31,133,31,133,30,168,31,121,31,121,30,170,31,75,31,233,31,233,30,121,31,186,31,85,31,15,31,67,31,33,31,8,31,8,30,73,31,69,31,253,31,253,30,29,31,211,31,211,30,211,29,147,31,139,31,23,31,58,31,58,30,62,31,193,31,10,31,10,30,10,29,65,31,64,31,98,31,1,31,89,31,141,31,160,31,160,30,156,31,115,31,106,31,200,31,182,31,182,30,43,31,174,31,174,30,84,31,147,31,195,31,145,31,145,30,145,29,145,28,192,31,104,31,77,31,238,31,157,31,18,31,173,31,173,30,106,31,76,31,76,30,76,29,209,31,81,31,63,31,63,30,36,31,139,31,198,31,159,31,159,30,159,29,138,31,153,31,57,31,57,30,10,31,185,31,53,31,168,31,103,31,103,30,103,29,117,31,46,31,94,31,106,31,136,31,136,30,136,29,136,28,190,31,238,31,4,31,169,31,169,30,61,31,186,31,71,31,71,30,125,31,125,30,20,31,182,31,62,31,24,31,24,30,24,29,84,31,247,31,102,31,102,30,216,31,30,31,169,31,25,31,25,30,225,31,225,30,180,31,180,30,165,31,134,31,227,31,73,31,13,31,66,31,66,30,9,31,219,31,108,31,108,30,79,31,79,30,79,29,249,31,249,30,56,31,57,31,32,31,32,30,107,31,58,31,220,31,220,30,130,31,130,30,34,31,213,31,45,31,169,31,244,31,16,31,16,30,68,31,83,31,61,31,30,31,21,31,1,31,26,31,25,31,146,31,189,31,97,31,97,30,242,31,242,30,3,31,225,31,39,31,39,30,55,31,55,30,202,31,202,30,247,31,247,30,71,31,195,31,238,31,173,31,158,31,239,31,103,31,112,31,189,31,189,30,30,31,18,31,205,31,207,31,18,31,215,31,245,31,14,31,240,31,195,31,119,31,216,31,60,31,60,30,81,31,251,31,247,31,20,31,20,30,138,31,138,30,228,31,228,30,63,31,187,31,45,31,81,31,81,30,81,29,105,31,236,31,124,31,124,30,120,31,182,31,249,31,48,31,111,31,46,31,4,31,2,31,208,31,45,31,33,31,33,31,242,31,95,31,203,31,51,31,113,31,142,31,45,31,85,31,7,31,34,31,10,31,63,31,50,31,163,31,144,31,110,31,53,31,30,31,52,31,52,30,201,31,70,31,255,31,153,31,146,31,140,31,146,31,60,31,8,31,186,31,6,31,36,31,187,31,79,31,79,30,74,31,37,31,37,30,111,31,239,31,66,31,222,31,222,30,222,29,100,31,218,31,80,31,80,30,113,31,113,30,113,29,229,31,229,30,242,31,49,31,44,31,102,31,102,30,242,31,242,30,242,29,242,28,52,31,176,31,232,31,243,31,2,31,117,31,117,30,170,31,170,30,169,31,142,31,101,31,101,30,95,31,95,30,107,31,107,30,107,29,242,31,235,31,10,31,127,31,15,31,247,31,193,31,142,31,23,31,200,31,125,31,42,31,210,31,106,31,139,31,179,31,106,31,174,31,70,31,70,30,204,31,195,31,195,30,60,31,202,31,236,31,197,31,41,31,140,31,24,31,250,31,242,31,211,31,40,31,101,31,63,31,57,31,57,30,178,31,142,31,140,31,189,31,75,31,81,31,23,31,108,31,121,31,39,31,39,30,250,31,1,31,109,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
