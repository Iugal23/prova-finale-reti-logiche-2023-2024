-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 769;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (156,0,176,0,76,0,0,0,0,0,0,0,67,0,44,0,38,0,32,0,106,0,94,0,107,0,0,0,185,0,123,0,82,0,1,0,100,0,0,0,205,0,86,0,51,0,101,0,130,0,228,0,0,0,0,0,218,0,0,0,204,0,28,0,251,0,131,0,243,0,80,0,0,0,130,0,128,0,144,0,38,0,210,0,160,0,161,0,252,0,103,0,0,0,141,0,92,0,175,0,143,0,178,0,63,0,13,0,0,0,160,0,78,0,6,0,116,0,2,0,1,0,23,0,139,0,0,0,218,0,193,0,153,0,238,0,67,0,209,0,59,0,84,0,232,0,0,0,87,0,163,0,244,0,205,0,125,0,0,0,73,0,131,0,125,0,201,0,0,0,54,0,0,0,231,0,8,0,134,0,0,0,188,0,181,0,209,0,0,0,158,0,0,0,140,0,216,0,41,0,0,0,75,0,151,0,73,0,227,0,213,0,75,0,2,0,220,0,105,0,63,0,0,0,65,0,251,0,77,0,141,0,10,0,211,0,63,0,0,0,68,0,233,0,121,0,127,0,131,0,226,0,201,0,230,0,122,0,0,0,107,0,106,0,153,0,210,0,122,0,103,0,101,0,0,0,6,0,121,0,237,0,0,0,24,0,212,0,109,0,5,0,44,0,53,0,154,0,148,0,154,0,246,0,16,0,28,0,0,0,43,0,64,0,248,0,115,0,104,0,252,0,101,0,0,0,193,0,22,0,0,0,0,0,180,0,0,0,79,0,148,0,66,0,101,0,45,0,0,0,145,0,0,0,133,0,207,0,158,0,0,0,0,0,162,0,0,0,0,0,60,0,80,0,221,0,112,0,0,0,172,0,217,0,250,0,137,0,105,0,0,0,168,0,169,0,1,0,5,0,168,0,16,0,52,0,92,0,15,0,133,0,166,0,237,0,213,0,199,0,223,0,0,0,189,0,164,0,130,0,0,0,227,0,0,0,91,0,34,0,0,0,183,0,196,0,59,0,141,0,29,0,0,0,0,0,65,0,0,0,217,0,52,0,86,0,65,0,219,0,33,0,177,0,55,0,160,0,0,0,75,0,0,0,35,0,0,0,74,0,68,0,185,0,90,0,87,0,118,0,169,0,222,0,210,0,232,0,239,0,155,0,171,0,136,0,194,0,0,0,173,0,34,0,4,0,200,0,0,0,68,0,53,0,212,0,0,0,252,0,114,0,0,0,0,0,252,0,100,0,0,0,119,0,178,0,194,0,29,0,178,0,185,0,0,0,0,0,129,0,34,0,54,0,155,0,9,0,152,0,0,0,176,0,227,0,179,0,183,0,0,0,0,0,205,0,187,0,29,0,16,0,0,0,117,0,0,0,11,0,82,0,186,0,95,0,0,0,167,0,121,0,0,0,16,0,212,0,116,0,15,0,82,0,167,0,67,0,0,0,16,0,0,0,231,0,6,0,14,0,253,0,243,0,10,0,35,0,234,0,124,0,176,0,159,0,44,0,176,0,237,0,240,0,211,0,117,0,193,0,214,0,182,0,75,0,168,0,83,0,5,0,211,0,243,0,205,0,128,0,0,0,0,0,79,0,0,0,89,0,205,0,154,0,166,0,25,0,138,0,8,0,250,0,61,0,94,0,192,0,135,0,213,0,82,0,140,0,153,0,105,0,215,0,192,0,164,0,22,0,33,0,113,0,176,0,73,0,174,0,0,0,147,0,102,0,130,0,42,0,94,0,86,0,214,0,0,0,0,0,148,0,124,0,22,0,152,0,241,0,23,0,86,0,247,0,209,0,0,0,40,0,68,0,210,0,176,0,76,0,88,0,0,0,110,0,6,0,181,0,213,0,105,0,0,0,0,0,122,0,114,0,0,0,102,0,207,0,0,0,3,0,0,0,58,0,0,0,128,0,235,0,130,0,0,0,101,0,79,0,171,0,193,0,211,0,230,0,132,0,186,0,0,0,0,0,233,0,81,0,55,0,113,0,102,0,0,0,134,0,124,0,0,0,0,0,184,0,173,0,81,0,55,0,0,0,144,0,156,0,191,0,103,0,18,0,236,0,143,0,33,0,90,0,179,0,113,0,114,0,143,0,213,0,27,0,177,0,194,0,144,0,253,0,86,0,0,0,75,0,107,0,67,0,237,0,0,0,58,0,137,0,7,0,105,0,24,0,35,0,0,0,228,0,14,0,123,0,207,0,60,0,42,0,224,0,234,0,84,0,66,0,223,0,0,0,216,0,0,0,0,0,199,0,0,0,24,0,184,0,0,0,227,0,27,0,0,0,251,0,26,0,0,0,0,0,79,0,89,0,56,0,0,0,231,0,79,0,0,0,0,0,219,0,0,0,12,0,0,0,200,0,0,0,0,0,42,0,146,0,235,0,22,0,22,0,45,0,64,0,0,0,0,0,106,0,243,0,1,0,0,0,74,0,231,0,120,0,189,0,115,0,0,0,194,0,15,0,57,0,60,0,147,0,253,0,28,0,165,0,172,0,43,0,0,0,77,0,0,0,242,0,166,0,72,0,181,0,183,0,0,0,11,0,0,0,0,0,235,0,107,0,0,0,196,0,8,0,0,0,0,0,0,0,220,0,0,0,0,0,74,0,210,0,15,0,133,0,120,0,190,0,9,0,173,0,188,0,185,0,66,0,150,0,33,0,230,0,96,0,68,0,15,0,159,0,26,0,146,0,42,0,41,0,144,0,151,0,219,0,210,0,149,0,201,0,100,0,0,0,99,0,109,0,233,0,130,0,248,0,76,0,2,0,229,0,84,0,92,0,231,0,0,0,146,0,0,0,120,0,178,0,242,0,111,0,149,0,234,0,115,0,0,0,187,0,153,0,0,0,95,0,152,0,39,0,211,0,172,0,42,0,230,0,29,0,85,0,171,0,53,0,102,0,241,0,54,0,0,0,0,0,239,0,0,0,111,0,88,0,108,0,0,0,97,0,0,0,243,0,50,0,31,0,201,0,98,0,213,0,109,0,221,0,23,0,178,0,73,0,204,0,121,0,139,0,156,0,0,0,32,0,55,0,0,0,227,0,19,0,90,0,102,0,196,0,82,0,25,0,111,0,24,0,0,0,53,0,239,0,76,0,0,0,0,0,73,0,0,0,240,0,54,0,165,0,0,0,207,0,197,0,55,0,117,0,0,0,0,0,144,0,141,0,0,0,12,0,50,0,0,0,137,0,0,0,102,0,40,0,79,0,253,0,165,0,216,0,19,0,0,0,135,0,203,0,239,0,0,0,0,0,0,0,88,0,141,0,31,0,126,0,0,0,123,0,128,0,87,0,54,0,69,0,49,0,85,0,0,0,205,0,146,0,82,0,0,0,91,0,163,0,3,0,248,0,162,0,0,0,226,0,0,0,217,0,0,0,0,0,214,0,90,0,191,0,68,0,21,0,103,0,161,0,146,0,150,0,134,0,31,0,70,0,0,0,5,0);
signal scenario_full  : scenario_type := (156,31,176,31,76,31,76,30,76,29,76,28,67,31,44,31,38,31,32,31,106,31,94,31,107,31,107,30,185,31,123,31,82,31,1,31,100,31,100,30,205,31,86,31,51,31,101,31,130,31,228,31,228,30,228,29,218,31,218,30,204,31,28,31,251,31,131,31,243,31,80,31,80,30,130,31,128,31,144,31,38,31,210,31,160,31,161,31,252,31,103,31,103,30,141,31,92,31,175,31,143,31,178,31,63,31,13,31,13,30,160,31,78,31,6,31,116,31,2,31,1,31,23,31,139,31,139,30,218,31,193,31,153,31,238,31,67,31,209,31,59,31,84,31,232,31,232,30,87,31,163,31,244,31,205,31,125,31,125,30,73,31,131,31,125,31,201,31,201,30,54,31,54,30,231,31,8,31,134,31,134,30,188,31,181,31,209,31,209,30,158,31,158,30,140,31,216,31,41,31,41,30,75,31,151,31,73,31,227,31,213,31,75,31,2,31,220,31,105,31,63,31,63,30,65,31,251,31,77,31,141,31,10,31,211,31,63,31,63,30,68,31,233,31,121,31,127,31,131,31,226,31,201,31,230,31,122,31,122,30,107,31,106,31,153,31,210,31,122,31,103,31,101,31,101,30,6,31,121,31,237,31,237,30,24,31,212,31,109,31,5,31,44,31,53,31,154,31,148,31,154,31,246,31,16,31,28,31,28,30,43,31,64,31,248,31,115,31,104,31,252,31,101,31,101,30,193,31,22,31,22,30,22,29,180,31,180,30,79,31,148,31,66,31,101,31,45,31,45,30,145,31,145,30,133,31,207,31,158,31,158,30,158,29,162,31,162,30,162,29,60,31,80,31,221,31,112,31,112,30,172,31,217,31,250,31,137,31,105,31,105,30,168,31,169,31,1,31,5,31,168,31,16,31,52,31,92,31,15,31,133,31,166,31,237,31,213,31,199,31,223,31,223,30,189,31,164,31,130,31,130,30,227,31,227,30,91,31,34,31,34,30,183,31,196,31,59,31,141,31,29,31,29,30,29,29,65,31,65,30,217,31,52,31,86,31,65,31,219,31,33,31,177,31,55,31,160,31,160,30,75,31,75,30,35,31,35,30,74,31,68,31,185,31,90,31,87,31,118,31,169,31,222,31,210,31,232,31,239,31,155,31,171,31,136,31,194,31,194,30,173,31,34,31,4,31,200,31,200,30,68,31,53,31,212,31,212,30,252,31,114,31,114,30,114,29,252,31,100,31,100,30,119,31,178,31,194,31,29,31,178,31,185,31,185,30,185,29,129,31,34,31,54,31,155,31,9,31,152,31,152,30,176,31,227,31,179,31,183,31,183,30,183,29,205,31,187,31,29,31,16,31,16,30,117,31,117,30,11,31,82,31,186,31,95,31,95,30,167,31,121,31,121,30,16,31,212,31,116,31,15,31,82,31,167,31,67,31,67,30,16,31,16,30,231,31,6,31,14,31,253,31,243,31,10,31,35,31,234,31,124,31,176,31,159,31,44,31,176,31,237,31,240,31,211,31,117,31,193,31,214,31,182,31,75,31,168,31,83,31,5,31,211,31,243,31,205,31,128,31,128,30,128,29,79,31,79,30,89,31,205,31,154,31,166,31,25,31,138,31,8,31,250,31,61,31,94,31,192,31,135,31,213,31,82,31,140,31,153,31,105,31,215,31,192,31,164,31,22,31,33,31,113,31,176,31,73,31,174,31,174,30,147,31,102,31,130,31,42,31,94,31,86,31,214,31,214,30,214,29,148,31,124,31,22,31,152,31,241,31,23,31,86,31,247,31,209,31,209,30,40,31,68,31,210,31,176,31,76,31,88,31,88,30,110,31,6,31,181,31,213,31,105,31,105,30,105,29,122,31,114,31,114,30,102,31,207,31,207,30,3,31,3,30,58,31,58,30,128,31,235,31,130,31,130,30,101,31,79,31,171,31,193,31,211,31,230,31,132,31,186,31,186,30,186,29,233,31,81,31,55,31,113,31,102,31,102,30,134,31,124,31,124,30,124,29,184,31,173,31,81,31,55,31,55,30,144,31,156,31,191,31,103,31,18,31,236,31,143,31,33,31,90,31,179,31,113,31,114,31,143,31,213,31,27,31,177,31,194,31,144,31,253,31,86,31,86,30,75,31,107,31,67,31,237,31,237,30,58,31,137,31,7,31,105,31,24,31,35,31,35,30,228,31,14,31,123,31,207,31,60,31,42,31,224,31,234,31,84,31,66,31,223,31,223,30,216,31,216,30,216,29,199,31,199,30,24,31,184,31,184,30,227,31,27,31,27,30,251,31,26,31,26,30,26,29,79,31,89,31,56,31,56,30,231,31,79,31,79,30,79,29,219,31,219,30,12,31,12,30,200,31,200,30,200,29,42,31,146,31,235,31,22,31,22,31,45,31,64,31,64,30,64,29,106,31,243,31,1,31,1,30,74,31,231,31,120,31,189,31,115,31,115,30,194,31,15,31,57,31,60,31,147,31,253,31,28,31,165,31,172,31,43,31,43,30,77,31,77,30,242,31,166,31,72,31,181,31,183,31,183,30,11,31,11,30,11,29,235,31,107,31,107,30,196,31,8,31,8,30,8,29,8,28,220,31,220,30,220,29,74,31,210,31,15,31,133,31,120,31,190,31,9,31,173,31,188,31,185,31,66,31,150,31,33,31,230,31,96,31,68,31,15,31,159,31,26,31,146,31,42,31,41,31,144,31,151,31,219,31,210,31,149,31,201,31,100,31,100,30,99,31,109,31,233,31,130,31,248,31,76,31,2,31,229,31,84,31,92,31,231,31,231,30,146,31,146,30,120,31,178,31,242,31,111,31,149,31,234,31,115,31,115,30,187,31,153,31,153,30,95,31,152,31,39,31,211,31,172,31,42,31,230,31,29,31,85,31,171,31,53,31,102,31,241,31,54,31,54,30,54,29,239,31,239,30,111,31,88,31,108,31,108,30,97,31,97,30,243,31,50,31,31,31,201,31,98,31,213,31,109,31,221,31,23,31,178,31,73,31,204,31,121,31,139,31,156,31,156,30,32,31,55,31,55,30,227,31,19,31,90,31,102,31,196,31,82,31,25,31,111,31,24,31,24,30,53,31,239,31,76,31,76,30,76,29,73,31,73,30,240,31,54,31,165,31,165,30,207,31,197,31,55,31,117,31,117,30,117,29,144,31,141,31,141,30,12,31,50,31,50,30,137,31,137,30,102,31,40,31,79,31,253,31,165,31,216,31,19,31,19,30,135,31,203,31,239,31,239,30,239,29,239,28,88,31,141,31,31,31,126,31,126,30,123,31,128,31,87,31,54,31,69,31,49,31,85,31,85,30,205,31,146,31,82,31,82,30,91,31,163,31,3,31,248,31,162,31,162,30,226,31,226,30,217,31,217,30,217,29,214,31,90,31,191,31,68,31,21,31,103,31,161,31,146,31,150,31,134,31,31,31,70,31,70,30,5,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
