-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_185 is
end project_tb_185;

architecture project_tb_arch_185 of project_tb_185 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 545;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (46,0,0,0,68,0,93,0,86,0,0,0,59,0,60,0,54,0,241,0,0,0,57,0,0,0,148,0,0,0,0,0,8,0,52,0,119,0,161,0,194,0,18,0,185,0,17,0,178,0,214,0,249,0,0,0,109,0,244,0,169,0,248,0,238,0,167,0,27,0,121,0,148,0,49,0,0,0,240,0,0,0,20,0,249,0,23,0,103,0,0,0,0,0,0,0,238,0,104,0,58,0,49,0,24,0,177,0,21,0,8,0,0,0,216,0,171,0,199,0,195,0,0,0,161,0,101,0,78,0,235,0,102,0,148,0,121,0,0,0,208,0,81,0,36,0,0,0,219,0,40,0,255,0,210,0,0,0,148,0,238,0,28,0,36,0,0,0,196,0,22,0,68,0,0,0,0,0,41,0,19,0,14,0,30,0,32,0,79,0,118,0,0,0,208,0,0,0,185,0,14,0,240,0,184,0,66,0,0,0,0,0,252,0,209,0,0,0,0,0,209,0,89,0,158,0,90,0,197,0,48,0,249,0,33,0,55,0,244,0,172,0,59,0,0,0,0,0,72,0,197,0,24,0,244,0,24,0,0,0,115,0,226,0,121,0,25,0,0,0,44,0,59,0,0,0,0,0,72,0,106,0,0,0,85,0,146,0,136,0,0,0,49,0,18,0,43,0,245,0,0,0,0,0,30,0,0,0,118,0,5,0,249,0,0,0,85,0,227,0,0,0,0,0,75,0,121,0,4,0,0,0,52,0,150,0,0,0,20,0,225,0,0,0,118,0,87,0,96,0,189,0,252,0,0,0,0,0,120,0,28,0,54,0,150,0,190,0,137,0,112,0,84,0,18,0,0,0,68,0,37,0,245,0,47,0,127,0,0,0,67,0,125,0,53,0,0,0,36,0,0,0,249,0,100,0,24,0,250,0,0,0,0,0,27,0,198,0,72,0,0,0,200,0,0,0,101,0,123,0,33,0,0,0,175,0,2,0,5,0,99,0,0,0,250,0,69,0,166,0,57,0,68,0,118,0,184,0,96,0,36,0,0,0,93,0,135,0,61,0,137,0,67,0,163,0,0,0,201,0,66,0,158,0,14,0,90,0,60,0,6,0,5,0,75,0,171,0,159,0,0,0,14,0,249,0,35,0,217,0,0,0,0,0,98,0,0,0,108,0,0,0,162,0,218,0,47,0,200,0,71,0,220,0,215,0,242,0,144,0,167,0,135,0,129,0,151,0,0,0,0,0,209,0,1,0,0,0,187,0,0,0,25,0,0,0,19,0,160,0,100,0,0,0,253,0,214,0,128,0,3,0,41,0,0,0,239,0,0,0,184,0,140,0,230,0,134,0,32,0,114,0,28,0,89,0,162,0,175,0,123,0,168,0,204,0,86,0,0,0,43,0,0,0,135,0,115,0,89,0,194,0,0,0,77,0,106,0,163,0,235,0,99,0,227,0,103,0,77,0,0,0,108,0,211,0,177,0,89,0,112,0,20,0,10,0,43,0,167,0,0,0,10,0,226,0,212,0,0,0,0,0,82,0,213,0,188,0,85,0,239,0,0,0,205,0,0,0,223,0,0,0,124,0,0,0,231,0,113,0,163,0,0,0,55,0,0,0,65,0,178,0,0,0,60,0,221,0,24,0,28,0,118,0,218,0,63,0,0,0,0,0,222,0,227,0,0,0,0,0,217,0,211,0,133,0,0,0,69,0,164,0,77,0,51,0,124,0,0,0,191,0,133,0,0,0,0,0,189,0,142,0,220,0,253,0,147,0,0,0,176,0,0,0,9,0,25,0,0,0,0,0,104,0,111,0,7,0,105,0,16,0,183,0,52,0,96,0,127,0,209,0,88,0,0,0,0,0,101,0,126,0,199,0,223,0,232,0,203,0,176,0,239,0,0,0,206,0,166,0,57,0,47,0,73,0,113,0,96,0,0,0,165,0,254,0,4,0,0,0,202,0,0,0,16,0,11,0,0,0,66,0,23,0,0,0,248,0,126,0,204,0,26,0,0,0,109,0,82,0,134,0,187,0,128,0,181,0,99,0,179,0,0,0,1,0,0,0,29,0,0,0,120,0,0,0,6,0,0,0,136,0,0,0,0,0,0,0,0,0,0,0,213,0,117,0,25,0,101,0,0,0,222,0,131,0,28,0,71,0,29,0,203,0,164,0,188,0,250,0,210,0,138,0,197,0,175,0,231,0,63,0,153,0,80,0,140,0,130,0,168,0,20,0,247,0,185,0,92,0,231,0,0,0,69,0,148,0,23,0,56,0,244,0,55,0,108,0,171,0,0,0,0,0,209,0,253,0,10,0,226,0,57,0,0,0,92,0,110,0,67,0,91,0,131,0,0,0,232,0,215,0,0,0,156,0,92,0,19,0,0,0,83,0,193,0,180,0,144,0,174,0,234,0,159,0,174,0,56,0,194,0,12,0,164,0,0,0,66,0);
signal scenario_full  : scenario_type := (46,31,46,30,68,31,93,31,86,31,86,30,59,31,60,31,54,31,241,31,241,30,57,31,57,30,148,31,148,30,148,29,8,31,52,31,119,31,161,31,194,31,18,31,185,31,17,31,178,31,214,31,249,31,249,30,109,31,244,31,169,31,248,31,238,31,167,31,27,31,121,31,148,31,49,31,49,30,240,31,240,30,20,31,249,31,23,31,103,31,103,30,103,29,103,28,238,31,104,31,58,31,49,31,24,31,177,31,21,31,8,31,8,30,216,31,171,31,199,31,195,31,195,30,161,31,101,31,78,31,235,31,102,31,148,31,121,31,121,30,208,31,81,31,36,31,36,30,219,31,40,31,255,31,210,31,210,30,148,31,238,31,28,31,36,31,36,30,196,31,22,31,68,31,68,30,68,29,41,31,19,31,14,31,30,31,32,31,79,31,118,31,118,30,208,31,208,30,185,31,14,31,240,31,184,31,66,31,66,30,66,29,252,31,209,31,209,30,209,29,209,31,89,31,158,31,90,31,197,31,48,31,249,31,33,31,55,31,244,31,172,31,59,31,59,30,59,29,72,31,197,31,24,31,244,31,24,31,24,30,115,31,226,31,121,31,25,31,25,30,44,31,59,31,59,30,59,29,72,31,106,31,106,30,85,31,146,31,136,31,136,30,49,31,18,31,43,31,245,31,245,30,245,29,30,31,30,30,118,31,5,31,249,31,249,30,85,31,227,31,227,30,227,29,75,31,121,31,4,31,4,30,52,31,150,31,150,30,20,31,225,31,225,30,118,31,87,31,96,31,189,31,252,31,252,30,252,29,120,31,28,31,54,31,150,31,190,31,137,31,112,31,84,31,18,31,18,30,68,31,37,31,245,31,47,31,127,31,127,30,67,31,125,31,53,31,53,30,36,31,36,30,249,31,100,31,24,31,250,31,250,30,250,29,27,31,198,31,72,31,72,30,200,31,200,30,101,31,123,31,33,31,33,30,175,31,2,31,5,31,99,31,99,30,250,31,69,31,166,31,57,31,68,31,118,31,184,31,96,31,36,31,36,30,93,31,135,31,61,31,137,31,67,31,163,31,163,30,201,31,66,31,158,31,14,31,90,31,60,31,6,31,5,31,75,31,171,31,159,31,159,30,14,31,249,31,35,31,217,31,217,30,217,29,98,31,98,30,108,31,108,30,162,31,218,31,47,31,200,31,71,31,220,31,215,31,242,31,144,31,167,31,135,31,129,31,151,31,151,30,151,29,209,31,1,31,1,30,187,31,187,30,25,31,25,30,19,31,160,31,100,31,100,30,253,31,214,31,128,31,3,31,41,31,41,30,239,31,239,30,184,31,140,31,230,31,134,31,32,31,114,31,28,31,89,31,162,31,175,31,123,31,168,31,204,31,86,31,86,30,43,31,43,30,135,31,115,31,89,31,194,31,194,30,77,31,106,31,163,31,235,31,99,31,227,31,103,31,77,31,77,30,108,31,211,31,177,31,89,31,112,31,20,31,10,31,43,31,167,31,167,30,10,31,226,31,212,31,212,30,212,29,82,31,213,31,188,31,85,31,239,31,239,30,205,31,205,30,223,31,223,30,124,31,124,30,231,31,113,31,163,31,163,30,55,31,55,30,65,31,178,31,178,30,60,31,221,31,24,31,28,31,118,31,218,31,63,31,63,30,63,29,222,31,227,31,227,30,227,29,217,31,211,31,133,31,133,30,69,31,164,31,77,31,51,31,124,31,124,30,191,31,133,31,133,30,133,29,189,31,142,31,220,31,253,31,147,31,147,30,176,31,176,30,9,31,25,31,25,30,25,29,104,31,111,31,7,31,105,31,16,31,183,31,52,31,96,31,127,31,209,31,88,31,88,30,88,29,101,31,126,31,199,31,223,31,232,31,203,31,176,31,239,31,239,30,206,31,166,31,57,31,47,31,73,31,113,31,96,31,96,30,165,31,254,31,4,31,4,30,202,31,202,30,16,31,11,31,11,30,66,31,23,31,23,30,248,31,126,31,204,31,26,31,26,30,109,31,82,31,134,31,187,31,128,31,181,31,99,31,179,31,179,30,1,31,1,30,29,31,29,30,120,31,120,30,6,31,6,30,136,31,136,30,136,29,136,28,136,27,136,26,213,31,117,31,25,31,101,31,101,30,222,31,131,31,28,31,71,31,29,31,203,31,164,31,188,31,250,31,210,31,138,31,197,31,175,31,231,31,63,31,153,31,80,31,140,31,130,31,168,31,20,31,247,31,185,31,92,31,231,31,231,30,69,31,148,31,23,31,56,31,244,31,55,31,108,31,171,31,171,30,171,29,209,31,253,31,10,31,226,31,57,31,57,30,92,31,110,31,67,31,91,31,131,31,131,30,232,31,215,31,215,30,156,31,92,31,19,31,19,30,83,31,193,31,180,31,144,31,174,31,234,31,159,31,174,31,56,31,194,31,12,31,164,31,164,30,66,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
