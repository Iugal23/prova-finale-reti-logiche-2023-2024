-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_151 is
end project_tb_151;

architecture project_tb_arch_151 of project_tb_151 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 293;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (44,0,0,0,0,0,110,0,0,0,20,0,155,0,81,0,0,0,87,0,75,0,165,0,138,0,101,0,248,0,105,0,0,0,52,0,61,0,9,0,115,0,80,0,245,0,220,0,65,0,55,0,0,0,71,0,49,0,80,0,64,0,87,0,8,0,245,0,0,0,212,0,195,0,90,0,71,0,141,0,53,0,23,0,128,0,142,0,165,0,43,0,84,0,13,0,137,0,147,0,0,0,143,0,197,0,191,0,143,0,0,0,70,0,0,0,0,0,197,0,206,0,175,0,177,0,81,0,210,0,183,0,0,0,81,0,42,0,106,0,0,0,125,0,249,0,171,0,97,0,223,0,177,0,79,0,209,0,0,0,136,0,7,0,8,0,207,0,253,0,6,0,214,0,168,0,77,0,231,0,138,0,242,0,0,0,88,0,0,0,186,0,252,0,217,0,130,0,136,0,48,0,199,0,73,0,201,0,238,0,136,0,0,0,32,0,209,0,218,0,11,0,113,0,108,0,0,0,244,0,250,0,209,0,218,0,0,0,156,0,212,0,144,0,224,0,91,0,141,0,175,0,7,0,42,0,144,0,0,0,120,0,29,0,116,0,0,0,106,0,121,0,157,0,0,0,195,0,0,0,178,0,230,0,208,0,252,0,87,0,197,0,61,0,113,0,141,0,4,0,152,0,228,0,0,0,50,0,92,0,150,0,0,0,49,0,225,0,202,0,127,0,83,0,0,0,114,0,115,0,118,0,148,0,69,0,70,0,91,0,190,0,52,0,0,0,217,0,250,0,41,0,0,0,134,0,34,0,177,0,130,0,0,0,34,0,127,0,78,0,159,0,0,0,0,0,230,0,0,0,55,0,71,0,99,0,193,0,4,0,205,0,187,0,208,0,6,0,94,0,13,0,166,0,111,0,105,0,218,0,1,0,212,0,0,0,9,0,153,0,0,0,67,0,42,0,35,0,136,0,181,0,101,0,226,0,98,0,230,0,196,0,0,0,188,0,72,0,0,0,158,0,136,0,115,0,0,0,0,0,175,0,79,0,158,0,94,0,89,0,143,0,107,0,204,0,38,0,101,0,97,0,121,0,59,0,216,0,19,0,216,0,85,0,66,0,45,0,0,0,226,0,0,0,11,0,164,0,216,0,0,0,165,0,241,0,102,0,0,0,194,0,0,0,53,0,135,0,164,0,149,0,70,0,121,0,0,0,0,0,42,0,16,0,207,0,102,0,0,0,22,0,235,0,70,0,122,0,0,0,114,0,181,0,186,0,242,0,0,0,11,0,0,0,114,0,144,0,213,0,175,0,202,0,167,0);
signal scenario_full  : scenario_type := (44,31,44,30,44,29,110,31,110,30,20,31,155,31,81,31,81,30,87,31,75,31,165,31,138,31,101,31,248,31,105,31,105,30,52,31,61,31,9,31,115,31,80,31,245,31,220,31,65,31,55,31,55,30,71,31,49,31,80,31,64,31,87,31,8,31,245,31,245,30,212,31,195,31,90,31,71,31,141,31,53,31,23,31,128,31,142,31,165,31,43,31,84,31,13,31,137,31,147,31,147,30,143,31,197,31,191,31,143,31,143,30,70,31,70,30,70,29,197,31,206,31,175,31,177,31,81,31,210,31,183,31,183,30,81,31,42,31,106,31,106,30,125,31,249,31,171,31,97,31,223,31,177,31,79,31,209,31,209,30,136,31,7,31,8,31,207,31,253,31,6,31,214,31,168,31,77,31,231,31,138,31,242,31,242,30,88,31,88,30,186,31,252,31,217,31,130,31,136,31,48,31,199,31,73,31,201,31,238,31,136,31,136,30,32,31,209,31,218,31,11,31,113,31,108,31,108,30,244,31,250,31,209,31,218,31,218,30,156,31,212,31,144,31,224,31,91,31,141,31,175,31,7,31,42,31,144,31,144,30,120,31,29,31,116,31,116,30,106,31,121,31,157,31,157,30,195,31,195,30,178,31,230,31,208,31,252,31,87,31,197,31,61,31,113,31,141,31,4,31,152,31,228,31,228,30,50,31,92,31,150,31,150,30,49,31,225,31,202,31,127,31,83,31,83,30,114,31,115,31,118,31,148,31,69,31,70,31,91,31,190,31,52,31,52,30,217,31,250,31,41,31,41,30,134,31,34,31,177,31,130,31,130,30,34,31,127,31,78,31,159,31,159,30,159,29,230,31,230,30,55,31,71,31,99,31,193,31,4,31,205,31,187,31,208,31,6,31,94,31,13,31,166,31,111,31,105,31,218,31,1,31,212,31,212,30,9,31,153,31,153,30,67,31,42,31,35,31,136,31,181,31,101,31,226,31,98,31,230,31,196,31,196,30,188,31,72,31,72,30,158,31,136,31,115,31,115,30,115,29,175,31,79,31,158,31,94,31,89,31,143,31,107,31,204,31,38,31,101,31,97,31,121,31,59,31,216,31,19,31,216,31,85,31,66,31,45,31,45,30,226,31,226,30,11,31,164,31,216,31,216,30,165,31,241,31,102,31,102,30,194,31,194,30,53,31,135,31,164,31,149,31,70,31,121,31,121,30,121,29,42,31,16,31,207,31,102,31,102,30,22,31,235,31,70,31,122,31,122,30,114,31,181,31,186,31,242,31,242,30,11,31,11,30,114,31,144,31,213,31,175,31,202,31,167,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
