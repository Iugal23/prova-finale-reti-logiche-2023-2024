-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 606;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (228,0,108,0,47,0,185,0,0,0,226,0,139,0,73,0,48,0,248,0,174,0,24,0,5,0,160,0,184,0,41,0,15,0,125,0,24,0,0,0,219,0,21,0,0,0,252,0,183,0,232,0,18,0,0,0,79,0,0,0,109,0,0,0,0,0,17,0,167,0,92,0,12,0,7,0,92,0,40,0,188,0,0,0,32,0,156,0,6,0,189,0,0,0,131,0,161,0,157,0,5,0,163,0,159,0,0,0,145,0,36,0,150,0,207,0,247,0,3,0,218,0,214,0,0,0,204,0,24,0,19,0,247,0,241,0,229,0,247,0,60,0,101,0,44,0,234,0,155,0,106,0,154,0,124,0,69,0,152,0,222,0,108,0,0,0,0,0,245,0,48,0,0,0,0,0,0,0,88,0,0,0,213,0,184,0,206,0,51,0,20,0,179,0,0,0,62,0,35,0,0,0,0,0,0,0,6,0,226,0,2,0,37,0,136,0,0,0,71,0,66,0,74,0,0,0,109,0,148,0,141,0,7,0,48,0,64,0,247,0,117,0,133,0,27,0,5,0,92,0,70,0,34,0,0,0,226,0,47,0,144,0,159,0,0,0,194,0,249,0,143,0,78,0,0,0,0,0,53,0,218,0,0,0,0,0,0,0,217,0,0,0,0,0,0,0,96,0,68,0,84,0,130,0,157,0,0,0,240,0,53,0,214,0,29,0,45,0,41,0,243,0,61,0,225,0,198,0,155,0,158,0,97,0,127,0,58,0,119,0,102,0,103,0,193,0,198,0,0,0,119,0,154,0,206,0,0,0,33,0,103,0,236,0,106,0,88,0,152,0,88,0,18,0,0,0,9,0,89,0,147,0,214,0,222,0,142,0,223,0,93,0,121,0,147,0,207,0,0,0,0,0,20,0,102,0,194,0,103,0,0,0,0,0,0,0,44,0,207,0,11,0,70,0,34,0,252,0,193,0,234,0,249,0,46,0,0,0,214,0,192,0,235,0,228,0,56,0,0,0,101,0,0,0,71,0,62,0,19,0,244,0,203,0,128,0,163,0,0,0,60,0,207,0,220,0,212,0,214,0,0,0,199,0,225,0,9,0,133,0,155,0,114,0,0,0,201,0,180,0,48,0,190,0,236,0,138,0,151,0,252,0,181,0,114,0,142,0,29,0,0,0,4,0,238,0,0,0,0,0,51,0,0,0,0,0,0,0,200,0,36,0,0,0,1,0,25,0,199,0,160,0,69,0,0,0,101,0,232,0,81,0,59,0,90,0,202,0,5,0,0,0,0,0,154,0,102,0,75,0,248,0,32,0,100,0,106,0,112,0,150,0,41,0,110,0,151,0,0,0,168,0,21,0,0,0,225,0,3,0,167,0,0,0,0,0,0,0,128,0,58,0,0,0,117,0,199,0,0,0,48,0,0,0,70,0,23,0,0,0,201,0,230,0,51,0,0,0,0,0,0,0,87,0,0,0,195,0,220,0,57,0,171,0,178,0,119,0,252,0,113,0,4,0,57,0,212,0,213,0,135,0,166,0,79,0,246,0,226,0,18,0,155,0,71,0,179,0,0,0,39,0,74,0,163,0,236,0,202,0,187,0,0,0,0,0,27,0,0,0,246,0,68,0,0,0,147,0,0,0,77,0,125,0,162,0,0,0,125,0,149,0,96,0,33,0,0,0,22,0,91,0,0,0,237,0,76,0,17,0,10,0,246,0,50,0,160,0,172,0,31,0,0,0,216,0,83,0,239,0,179,0,75,0,38,0,200,0,211,0,229,0,18,0,0,0,0,0,204,0,238,0,53,0,184,0,96,0,248,0,0,0,255,0,18,0,165,0,0,0,118,0,122,0,177,0,229,0,172,0,254,0,0,0,0,0,63,0,235,0,0,0,247,0,31,0,62,0,0,0,94,0,0,0,0,0,14,0,0,0,152,0,22,0,231,0,0,0,95,0,211,0,122,0,196,0,52,0,30,0,32,0,204,0,0,0,160,0,176,0,167,0,61,0,49,0,0,0,104,0,65,0,124,0,166,0,195,0,166,0,62,0,0,0,230,0,234,0,94,0,251,0,102,0,239,0,94,0,57,0,28,0,0,0,0,0,0,0,0,0,177,0,159,0,0,0,27,0,21,0,216,0,170,0,8,0,113,0,28,0,0,0,137,0,244,0,194,0,0,0,245,0,0,0,163,0,0,0,42,0,89,0,102,0,183,0,65,0,135,0,225,0,218,0,97,0,25,0,80,0,255,0,226,0,123,0,111,0,0,0,7,0,0,0,6,0,40,0,23,0,0,0,11,0,15,0,253,0,0,0,51,0,237,0,214,0,166,0,110,0,253,0,0,0,232,0,76,0,138,0,0,0,229,0,147,0,0,0,196,0,71,0,0,0,84,0,209,0,76,0,144,0,0,0,28,0,0,0,40,0,188,0,112,0,126,0,123,0,91,0,161,0,0,0,176,0,254,0,182,0,175,0,196,0,0,0,116,0,136,0,241,0,2,0,142,0,9,0,79,0,131,0,164,0,90,0,203,0,192,0,0,0,55,0,32,0,55,0,20,0,96,0,60,0,0,0,113,0,221,0,0,0,27,0,218,0,57,0,141,0,57,0,0,0,134,0,0,0,58,0,231,0,51,0,114,0,17,0,255,0,55,0,134,0,171,0,0,0,3,0,0,0,0,0,150,0,5,0,190,0,0,0,0,0,201,0,59,0,233,0,0,0);
signal scenario_full  : scenario_type := (228,31,108,31,47,31,185,31,185,30,226,31,139,31,73,31,48,31,248,31,174,31,24,31,5,31,160,31,184,31,41,31,15,31,125,31,24,31,24,30,219,31,21,31,21,30,252,31,183,31,232,31,18,31,18,30,79,31,79,30,109,31,109,30,109,29,17,31,167,31,92,31,12,31,7,31,92,31,40,31,188,31,188,30,32,31,156,31,6,31,189,31,189,30,131,31,161,31,157,31,5,31,163,31,159,31,159,30,145,31,36,31,150,31,207,31,247,31,3,31,218,31,214,31,214,30,204,31,24,31,19,31,247,31,241,31,229,31,247,31,60,31,101,31,44,31,234,31,155,31,106,31,154,31,124,31,69,31,152,31,222,31,108,31,108,30,108,29,245,31,48,31,48,30,48,29,48,28,88,31,88,30,213,31,184,31,206,31,51,31,20,31,179,31,179,30,62,31,35,31,35,30,35,29,35,28,6,31,226,31,2,31,37,31,136,31,136,30,71,31,66,31,74,31,74,30,109,31,148,31,141,31,7,31,48,31,64,31,247,31,117,31,133,31,27,31,5,31,92,31,70,31,34,31,34,30,226,31,47,31,144,31,159,31,159,30,194,31,249,31,143,31,78,31,78,30,78,29,53,31,218,31,218,30,218,29,218,28,217,31,217,30,217,29,217,28,96,31,68,31,84,31,130,31,157,31,157,30,240,31,53,31,214,31,29,31,45,31,41,31,243,31,61,31,225,31,198,31,155,31,158,31,97,31,127,31,58,31,119,31,102,31,103,31,193,31,198,31,198,30,119,31,154,31,206,31,206,30,33,31,103,31,236,31,106,31,88,31,152,31,88,31,18,31,18,30,9,31,89,31,147,31,214,31,222,31,142,31,223,31,93,31,121,31,147,31,207,31,207,30,207,29,20,31,102,31,194,31,103,31,103,30,103,29,103,28,44,31,207,31,11,31,70,31,34,31,252,31,193,31,234,31,249,31,46,31,46,30,214,31,192,31,235,31,228,31,56,31,56,30,101,31,101,30,71,31,62,31,19,31,244,31,203,31,128,31,163,31,163,30,60,31,207,31,220,31,212,31,214,31,214,30,199,31,225,31,9,31,133,31,155,31,114,31,114,30,201,31,180,31,48,31,190,31,236,31,138,31,151,31,252,31,181,31,114,31,142,31,29,31,29,30,4,31,238,31,238,30,238,29,51,31,51,30,51,29,51,28,200,31,36,31,36,30,1,31,25,31,199,31,160,31,69,31,69,30,101,31,232,31,81,31,59,31,90,31,202,31,5,31,5,30,5,29,154,31,102,31,75,31,248,31,32,31,100,31,106,31,112,31,150,31,41,31,110,31,151,31,151,30,168,31,21,31,21,30,225,31,3,31,167,31,167,30,167,29,167,28,128,31,58,31,58,30,117,31,199,31,199,30,48,31,48,30,70,31,23,31,23,30,201,31,230,31,51,31,51,30,51,29,51,28,87,31,87,30,195,31,220,31,57,31,171,31,178,31,119,31,252,31,113,31,4,31,57,31,212,31,213,31,135,31,166,31,79,31,246,31,226,31,18,31,155,31,71,31,179,31,179,30,39,31,74,31,163,31,236,31,202,31,187,31,187,30,187,29,27,31,27,30,246,31,68,31,68,30,147,31,147,30,77,31,125,31,162,31,162,30,125,31,149,31,96,31,33,31,33,30,22,31,91,31,91,30,237,31,76,31,17,31,10,31,246,31,50,31,160,31,172,31,31,31,31,30,216,31,83,31,239,31,179,31,75,31,38,31,200,31,211,31,229,31,18,31,18,30,18,29,204,31,238,31,53,31,184,31,96,31,248,31,248,30,255,31,18,31,165,31,165,30,118,31,122,31,177,31,229,31,172,31,254,31,254,30,254,29,63,31,235,31,235,30,247,31,31,31,62,31,62,30,94,31,94,30,94,29,14,31,14,30,152,31,22,31,231,31,231,30,95,31,211,31,122,31,196,31,52,31,30,31,32,31,204,31,204,30,160,31,176,31,167,31,61,31,49,31,49,30,104,31,65,31,124,31,166,31,195,31,166,31,62,31,62,30,230,31,234,31,94,31,251,31,102,31,239,31,94,31,57,31,28,31,28,30,28,29,28,28,28,27,177,31,159,31,159,30,27,31,21,31,216,31,170,31,8,31,113,31,28,31,28,30,137,31,244,31,194,31,194,30,245,31,245,30,163,31,163,30,42,31,89,31,102,31,183,31,65,31,135,31,225,31,218,31,97,31,25,31,80,31,255,31,226,31,123,31,111,31,111,30,7,31,7,30,6,31,40,31,23,31,23,30,11,31,15,31,253,31,253,30,51,31,237,31,214,31,166,31,110,31,253,31,253,30,232,31,76,31,138,31,138,30,229,31,147,31,147,30,196,31,71,31,71,30,84,31,209,31,76,31,144,31,144,30,28,31,28,30,40,31,188,31,112,31,126,31,123,31,91,31,161,31,161,30,176,31,254,31,182,31,175,31,196,31,196,30,116,31,136,31,241,31,2,31,142,31,9,31,79,31,131,31,164,31,90,31,203,31,192,31,192,30,55,31,32,31,55,31,20,31,96,31,60,31,60,30,113,31,221,31,221,30,27,31,218,31,57,31,141,31,57,31,57,30,134,31,134,30,58,31,231,31,51,31,114,31,17,31,255,31,55,31,134,31,171,31,171,30,3,31,3,30,3,29,150,31,5,31,190,31,190,30,190,29,201,31,59,31,233,31,233,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
