-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_466 is
end project_tb_466;

architecture project_tb_arch_466 of project_tb_466 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 701;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (33,0,227,0,134,0,209,0,117,0,198,0,39,0,70,0,68,0,0,0,0,0,112,0,240,0,61,0,254,0,4,0,143,0,205,0,123,0,166,0,0,0,151,0,96,0,244,0,178,0,166,0,64,0,60,0,168,0,0,0,0,0,0,0,118,0,0,0,224,0,216,0,16,0,56,0,85,0,159,0,1,0,122,0,0,0,63,0,23,0,159,0,255,0,137,0,0,0,0,0,196,0,61,0,154,0,101,0,0,0,77,0,20,0,0,0,0,0,143,0,100,0,5,0,20,0,0,0,228,0,181,0,101,0,111,0,29,0,125,0,30,0,216,0,81,0,54,0,192,0,54,0,7,0,7,0,222,0,241,0,91,0,157,0,0,0,151,0,0,0,104,0,0,0,14,0,0,0,171,0,134,0,12,0,171,0,69,0,0,0,102,0,225,0,242,0,20,0,138,0,82,0,61,0,99,0,168,0,89,0,203,0,0,0,0,0,211,0,42,0,195,0,132,0,193,0,215,0,165,0,142,0,0,0,57,0,110,0,251,0,47,0,0,0,227,0,0,0,0,0,173,0,84,0,69,0,134,0,0,0,108,0,107,0,105,0,0,0,122,0,0,0,33,0,150,0,0,0,22,0,111,0,171,0,58,0,0,0,177,0,79,0,0,0,0,0,0,0,66,0,242,0,159,0,205,0,0,0,0,0,134,0,158,0,0,0,83,0,191,0,16,0,185,0,116,0,144,0,0,0,0,0,40,0,192,0,193,0,150,0,0,0,0,0,0,0,255,0,31,0,251,0,206,0,0,0,163,0,0,0,55,0,138,0,57,0,14,0,12,0,49,0,157,0,0,0,48,0,44,0,0,0,110,0,43,0,131,0,75,0,214,0,135,0,236,0,217,0,104,0,59,0,181,0,209,0,246,0,56,0,145,0,0,0,0,0,89,0,221,0,236,0,0,0,59,0,0,0,41,0,0,0,0,0,142,0,46,0,121,0,0,0,109,0,0,0,128,0,129,0,111,0,48,0,108,0,197,0,160,0,81,0,8,0,25,0,128,0,246,0,122,0,128,0,0,0,173,0,127,0,139,0,222,0,4,0,0,0,131,0,21,0,0,0,36,0,201,0,176,0,131,0,245,0,0,0,176,0,176,0,147,0,159,0,70,0,187,0,210,0,155,0,85,0,25,0,3,0,148,0,0,0,96,0,112,0,115,0,170,0,23,0,48,0,221,0,2,0,58,0,0,0,247,0,172,0,130,0,69,0,0,0,58,0,69,0,254,0,0,0,60,0,108,0,177,0,23,0,62,0,10,0,205,0,160,0,31,0,174,0,0,0,28,0,23,0,200,0,0,0,117,0,91,0,191,0,0,0,117,0,63,0,142,0,216,0,0,0,183,0,0,0,103,0,30,0,183,0,214,0,119,0,11,0,0,0,208,0,0,0,97,0,0,0,0,0,60,0,28,0,206,0,0,0,101,0,107,0,0,0,98,0,75,0,178,0,99,0,251,0,0,0,118,0,98,0,0,0,0,0,0,0,31,0,189,0,163,0,0,0,195,0,200,0,172,0,255,0,228,0,206,0,199,0,80,0,88,0,34,0,131,0,65,0,167,0,68,0,193,0,229,0,152,0,57,0,0,0,204,0,0,0,135,0,41,0,0,0,0,0,212,0,8,0,32,0,0,0,0,0,150,0,0,0,0,0,19,0,164,0,16,0,207,0,125,0,129,0,16,0,79,0,174,0,0,0,79,0,235,0,132,0,70,0,131,0,16,0,137,0,0,0,104,0,120,0,127,0,157,0,113,0,13,0,68,0,204,0,227,0,145,0,49,0,0,0,0,0,191,0,240,0,0,0,206,0,117,0,37,0,112,0,119,0,145,0,123,0,132,0,130,0,81,0,35,0,3,0,0,0,154,0,138,0,14,0,106,0,11,0,0,0,34,0,70,0,252,0,43,0,5,0,32,0,247,0,97,0,67,0,0,0,251,0,199,0,66,0,0,0,225,0,170,0,119,0,75,0,252,0,0,0,209,0,242,0,0,0,70,0,0,0,20,0,139,0,0,0,0,0,231,0,5,0,93,0,101,0,150,0,188,0,0,0,239,0,228,0,75,0,130,0,16,0,25,0,70,0,214,0,218,0,168,0,155,0,0,0,169,0,164,0,129,0,0,0,246,0,205,0,157,0,225,0,90,0,144,0,157,0,148,0,20,0,200,0,247,0,181,0,17,0,140,0,105,0,222,0,0,0,36,0,135,0,65,0,116,0,130,0,247,0,144,0,32,0,240,0,0,0,185,0,0,0,200,0,10,0,239,0,98,0,145,0,155,0,181,0,0,0,85,0,71,0,139,0,208,0,198,0,17,0,59,0,0,0,0,0,110,0,63,0,43,0,0,0,0,0,102,0,197,0,55,0,14,0,51,0,223,0,3,0,126,0,48,0,215,0,102,0,182,0,239,0,85,0,111,0,16,0,240,0,148,0,0,0,221,0,255,0,0,0,39,0,44,0,15,0,54,0,107,0,14,0,0,0,0,0,220,0,154,0,13,0,105,0,158,0,150,0,166,0,163,0,19,0,184,0,74,0,17,0,0,0,85,0,0,0,0,0,172,0,0,0,36,0,232,0,194,0,149,0,253,0,168,0,222,0,143,0,29,0,35,0,97,0,0,0,32,0,82,0,0,0,0,0,0,0,206,0,19,0,71,0,255,0,0,0,0,0,0,0,206,0,237,0,115,0,0,0,0,0,0,0,187,0,0,0,32,0,0,0,0,0,10,0,214,0,5,0,39,0,200,0,237,0,91,0,174,0,155,0,139,0,0,0,4,0,50,0,5,0,0,0,120,0,108,0,185,0,184,0,239,0,247,0,59,0,251,0,0,0,200,0,0,0,49,0,247,0,97,0,251,0,82,0,186,0,23,0,246,0,147,0,110,0,201,0,0,0,135,0,91,0,192,0,19,0,247,0,74,0,164,0,0,0,39,0,0,0,36,0,161,0,8,0,103,0,233,0,1,0,0,0,0,0,0,0,16,0,207,0,125,0,219,0,210,0,36,0,0,0,0,0,15,0,64,0,201,0,150,0,14,0,247,0,177,0,0,0,90,0,37,0,119,0,77,0,78,0,113,0,183,0,114,0,0,0,0,0,19,0);
signal scenario_full  : scenario_type := (33,31,227,31,134,31,209,31,117,31,198,31,39,31,70,31,68,31,68,30,68,29,112,31,240,31,61,31,254,31,4,31,143,31,205,31,123,31,166,31,166,30,151,31,96,31,244,31,178,31,166,31,64,31,60,31,168,31,168,30,168,29,168,28,118,31,118,30,224,31,216,31,16,31,56,31,85,31,159,31,1,31,122,31,122,30,63,31,23,31,159,31,255,31,137,31,137,30,137,29,196,31,61,31,154,31,101,31,101,30,77,31,20,31,20,30,20,29,143,31,100,31,5,31,20,31,20,30,228,31,181,31,101,31,111,31,29,31,125,31,30,31,216,31,81,31,54,31,192,31,54,31,7,31,7,31,222,31,241,31,91,31,157,31,157,30,151,31,151,30,104,31,104,30,14,31,14,30,171,31,134,31,12,31,171,31,69,31,69,30,102,31,225,31,242,31,20,31,138,31,82,31,61,31,99,31,168,31,89,31,203,31,203,30,203,29,211,31,42,31,195,31,132,31,193,31,215,31,165,31,142,31,142,30,57,31,110,31,251,31,47,31,47,30,227,31,227,30,227,29,173,31,84,31,69,31,134,31,134,30,108,31,107,31,105,31,105,30,122,31,122,30,33,31,150,31,150,30,22,31,111,31,171,31,58,31,58,30,177,31,79,31,79,30,79,29,79,28,66,31,242,31,159,31,205,31,205,30,205,29,134,31,158,31,158,30,83,31,191,31,16,31,185,31,116,31,144,31,144,30,144,29,40,31,192,31,193,31,150,31,150,30,150,29,150,28,255,31,31,31,251,31,206,31,206,30,163,31,163,30,55,31,138,31,57,31,14,31,12,31,49,31,157,31,157,30,48,31,44,31,44,30,110,31,43,31,131,31,75,31,214,31,135,31,236,31,217,31,104,31,59,31,181,31,209,31,246,31,56,31,145,31,145,30,145,29,89,31,221,31,236,31,236,30,59,31,59,30,41,31,41,30,41,29,142,31,46,31,121,31,121,30,109,31,109,30,128,31,129,31,111,31,48,31,108,31,197,31,160,31,81,31,8,31,25,31,128,31,246,31,122,31,128,31,128,30,173,31,127,31,139,31,222,31,4,31,4,30,131,31,21,31,21,30,36,31,201,31,176,31,131,31,245,31,245,30,176,31,176,31,147,31,159,31,70,31,187,31,210,31,155,31,85,31,25,31,3,31,148,31,148,30,96,31,112,31,115,31,170,31,23,31,48,31,221,31,2,31,58,31,58,30,247,31,172,31,130,31,69,31,69,30,58,31,69,31,254,31,254,30,60,31,108,31,177,31,23,31,62,31,10,31,205,31,160,31,31,31,174,31,174,30,28,31,23,31,200,31,200,30,117,31,91,31,191,31,191,30,117,31,63,31,142,31,216,31,216,30,183,31,183,30,103,31,30,31,183,31,214,31,119,31,11,31,11,30,208,31,208,30,97,31,97,30,97,29,60,31,28,31,206,31,206,30,101,31,107,31,107,30,98,31,75,31,178,31,99,31,251,31,251,30,118,31,98,31,98,30,98,29,98,28,31,31,189,31,163,31,163,30,195,31,200,31,172,31,255,31,228,31,206,31,199,31,80,31,88,31,34,31,131,31,65,31,167,31,68,31,193,31,229,31,152,31,57,31,57,30,204,31,204,30,135,31,41,31,41,30,41,29,212,31,8,31,32,31,32,30,32,29,150,31,150,30,150,29,19,31,164,31,16,31,207,31,125,31,129,31,16,31,79,31,174,31,174,30,79,31,235,31,132,31,70,31,131,31,16,31,137,31,137,30,104,31,120,31,127,31,157,31,113,31,13,31,68,31,204,31,227,31,145,31,49,31,49,30,49,29,191,31,240,31,240,30,206,31,117,31,37,31,112,31,119,31,145,31,123,31,132,31,130,31,81,31,35,31,3,31,3,30,154,31,138,31,14,31,106,31,11,31,11,30,34,31,70,31,252,31,43,31,5,31,32,31,247,31,97,31,67,31,67,30,251,31,199,31,66,31,66,30,225,31,170,31,119,31,75,31,252,31,252,30,209,31,242,31,242,30,70,31,70,30,20,31,139,31,139,30,139,29,231,31,5,31,93,31,101,31,150,31,188,31,188,30,239,31,228,31,75,31,130,31,16,31,25,31,70,31,214,31,218,31,168,31,155,31,155,30,169,31,164,31,129,31,129,30,246,31,205,31,157,31,225,31,90,31,144,31,157,31,148,31,20,31,200,31,247,31,181,31,17,31,140,31,105,31,222,31,222,30,36,31,135,31,65,31,116,31,130,31,247,31,144,31,32,31,240,31,240,30,185,31,185,30,200,31,10,31,239,31,98,31,145,31,155,31,181,31,181,30,85,31,71,31,139,31,208,31,198,31,17,31,59,31,59,30,59,29,110,31,63,31,43,31,43,30,43,29,102,31,197,31,55,31,14,31,51,31,223,31,3,31,126,31,48,31,215,31,102,31,182,31,239,31,85,31,111,31,16,31,240,31,148,31,148,30,221,31,255,31,255,30,39,31,44,31,15,31,54,31,107,31,14,31,14,30,14,29,220,31,154,31,13,31,105,31,158,31,150,31,166,31,163,31,19,31,184,31,74,31,17,31,17,30,85,31,85,30,85,29,172,31,172,30,36,31,232,31,194,31,149,31,253,31,168,31,222,31,143,31,29,31,35,31,97,31,97,30,32,31,82,31,82,30,82,29,82,28,206,31,19,31,71,31,255,31,255,30,255,29,255,28,206,31,237,31,115,31,115,30,115,29,115,28,187,31,187,30,32,31,32,30,32,29,10,31,214,31,5,31,39,31,200,31,237,31,91,31,174,31,155,31,139,31,139,30,4,31,50,31,5,31,5,30,120,31,108,31,185,31,184,31,239,31,247,31,59,31,251,31,251,30,200,31,200,30,49,31,247,31,97,31,251,31,82,31,186,31,23,31,246,31,147,31,110,31,201,31,201,30,135,31,91,31,192,31,19,31,247,31,74,31,164,31,164,30,39,31,39,30,36,31,161,31,8,31,103,31,233,31,1,31,1,30,1,29,1,28,16,31,207,31,125,31,219,31,210,31,36,31,36,30,36,29,15,31,64,31,201,31,150,31,14,31,247,31,177,31,177,30,90,31,37,31,119,31,77,31,78,31,113,31,183,31,114,31,114,30,114,29,19,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
