-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 960;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (193,0,133,0,0,0,9,0,0,0,198,0,121,0,252,0,170,0,14,0,171,0,15,0,6,0,104,0,188,0,0,0,170,0,87,0,167,0,214,0,47,0,0,0,213,0,69,0,0,0,34,0,120,0,120,0,0,0,89,0,0,0,146,0,25,0,175,0,232,0,81,0,113,0,68,0,212,0,175,0,20,0,188,0,0,0,0,0,188,0,20,0,21,0,36,0,4,0,8,0,0,0,80,0,53,0,0,0,168,0,0,0,15,0,243,0,91,0,191,0,164,0,89,0,197,0,247,0,218,0,73,0,141,0,0,0,0,0,55,0,192,0,120,0,58,0,198,0,75,0,98,0,0,0,95,0,219,0,209,0,10,0,178,0,0,0,150,0,32,0,65,0,21,0,244,0,82,0,66,0,134,0,91,0,0,0,0,0,94,0,0,0,0,0,254,0,114,0,9,0,16,0,186,0,155,0,62,0,162,0,214,0,183,0,56,0,0,0,0,0,191,0,158,0,210,0,24,0,28,0,254,0,193,0,177,0,113,0,55,0,6,0,135,0,232,0,62,0,207,0,0,0,64,0,113,0,0,0,51,0,100,0,0,0,197,0,0,0,209,0,74,0,16,0,153,0,96,0,74,0,144,0,122,0,79,0,195,0,75,0,18,0,159,0,0,0,159,0,21,0,0,0,0,0,95,0,170,0,239,0,52,0,4,0,119,0,39,0,32,0,69,0,0,0,9,0,243,0,114,0,111,0,88,0,249,0,75,0,0,0,202,0,34,0,0,0,60,0,221,0,0,0,166,0,0,0,60,0,7,0,146,0,168,0,166,0,82,0,207,0,249,0,52,0,30,0,0,0,167,0,217,0,1,0,97,0,37,0,49,0,245,0,140,0,168,0,179,0,68,0,97,0,145,0,149,0,141,0,122,0,106,0,81,0,40,0,182,0,0,0,0,0,40,0,36,0,247,0,0,0,5,0,22,0,184,0,24,0,61,0,165,0,138,0,30,0,49,0,181,0,106,0,210,0,0,0,89,0,0,0,107,0,87,0,0,0,157,0,211,0,139,0,33,0,55,0,122,0,250,0,56,0,114,0,190,0,142,0,6,0,25,0,73,0,69,0,21,0,255,0,0,0,43,0,38,0,0,0,0,0,0,0,194,0,14,0,0,0,193,0,85,0,224,0,94,0,0,0,103,0,103,0,116,0,79,0,228,0,27,0,0,0,155,0,121,0,0,0,0,0,0,0,0,0,0,0,62,0,131,0,105,0,0,0,0,0,129,0,144,0,29,0,0,0,19,0,89,0,0,0,20,0,0,0,187,0,131,0,82,0,20,0,170,0,0,0,0,0,0,0,230,0,234,0,113,0,90,0,0,0,0,0,157,0,218,0,224,0,22,0,93,0,19,0,154,0,37,0,45,0,9,0,33,0,100,0,31,0,149,0,183,0,115,0,15,0,188,0,143,0,172,0,10,0,120,0,198,0,172,0,20,0,25,0,79,0,125,0,117,0,32,0,56,0,0,0,47,0,128,0,248,0,10,0,115,0,149,0,198,0,29,0,0,0,5,0,123,0,157,0,198,0,230,0,0,0,231,0,0,0,0,0,90,0,0,0,187,0,222,0,0,0,138,0,0,0,215,0,96,0,252,0,86,0,0,0,71,0,4,0,241,0,170,0,65,0,0,0,45,0,237,0,0,0,108,0,0,0,0,0,0,0,41,0,136,0,0,0,209,0,14,0,238,0,52,0,148,0,103,0,208,0,56,0,184,0,31,0,107,0,149,0,151,0,15,0,174,0,48,0,156,0,195,0,0,0,218,0,0,0,84,0,188,0,0,0,236,0,217,0,152,0,66,0,85,0,147,0,0,0,242,0,0,0,208,0,0,0,70,0,53,0,0,0,58,0,62,0,75,0,10,0,179,0,170,0,0,0,150,0,0,0,110,0,251,0,0,0,199,0,188,0,0,0,74,0,133,0,97,0,75,0,188,0,40,0,4,0,143,0,180,0,0,0,67,0,2,0,21,0,152,0,209,0,218,0,0,0,57,0,147,0,253,0,0,0,0,0,61,0,102,0,152,0,244,0,109,0,92,0,112,0,19,0,73,0,236,0,157,0,161,0,167,0,202,0,176,0,0,0,0,0,164,0,220,0,94,0,78,0,148,0,128,0,116,0,132,0,105,0,161,0,218,0,0,0,145,0,135,0,59,0,0,0,185,0,220,0,0,0,214,0,0,0,0,0,121,0,0,0,195,0,171,0,236,0,117,0,148,0,0,0,132,0,55,0,174,0,18,0,69,0,241,0,218,0,174,0,66,0,5,0,170,0,173,0,0,0,0,0,170,0,187,0,22,0,33,0,135,0,149,0,177,0,0,0,125,0,0,0,70,0,210,0,9,0,237,0,252,0,0,0,34,0,0,0,183,0,70,0,108,0,96,0,0,0,213,0,195,0,0,0,41,0,0,0,234,0,11,0,0,0,236,0,217,0,0,0,0,0,190,0,250,0,0,0,33,0,0,0,97,0,191,0,232,0,0,0,0,0,238,0,0,0,145,0,237,0,0,0,56,0,0,0,114,0,247,0,164,0,0,0,149,0,151,0,0,0,177,0,0,0,37,0,174,0,76,0,190,0,0,0,174,0,111,0,0,0,205,0,0,0,247,0,0,0,0,0,191,0,33,0,0,0,0,0,0,0,225,0,106,0,119,0,0,0,0,0,152,0,65,0,8,0,95,0,0,0,0,0,18,0,0,0,0,0,29,0,0,0,121,0,244,0,0,0,120,0,183,0,0,0,129,0,62,0,216,0,151,0,42,0,128,0,70,0,112,0,0,0,148,0,80,0,0,0,129,0,0,0,39,0,0,0,241,0,57,0,0,0,37,0,29,0,180,0,0,0,62,0,47,0,102,0,108,0,11,0,0,0,154,0,67,0,204,0,161,0,245,0,249,0,169,0,116,0,159,0,0,0,6,0,118,0,90,0,195,0,162,0,180,0,178,0,19,0,212,0,0,0,141,0,0,0,248,0,55,0,0,0,175,0,150,0,0,0,0,0,185,0,184,0,48,0,102,0,147,0,0,0,41,0,0,0,8,0,4,0,251,0,64,0,162,0,120,0,144,0,184,0,0,0,48,0,175,0,151,0,220,0,45,0,0,0,151,0,164,0,87,0,50,0,209,0,127,0,211,0,105,0,11,0,244,0,216,0,161,0,0,0,6,0,0,0,224,0,105,0,0,0,226,0,0,0,70,0,94,0,131,0,176,0,0,0,3,0,87,0,235,0,178,0,247,0,28,0,4,0,0,0,0,0,152,0,78,0,205,0,59,0,51,0,225,0,176,0,181,0,154,0,119,0,227,0,0,0,0,0,246,0,102,0,0,0,26,0,53,0,25,0,38,0,73,0,9,0,0,0,68,0,0,0,138,0,130,0,204,0,101,0,20,0,0,0,128,0,241,0,0,0,29,0,0,0,193,0,16,0,104,0,246,0,0,0,198,0,166,0,169,0,0,0,34,0,112,0,154,0,46,0,188,0,225,0,117,0,51,0,245,0,216,0,188,0,28,0,0,0,158,0,249,0,76,0,0,0,255,0,111,0,184,0,0,0,186,0,197,0,168,0,113,0,231,0,65,0,28,0,0,0,0,0,3,0,247,0,0,0,174,0,107,0,95,0,122,0,224,0,157,0,0,0,0,0,47,0,241,0,88,0,219,0,56,0,59,0,0,0,155,0,192,0,207,0,50,0,168,0,112,0,40,0,238,0,48,0,0,0,0,0,88,0,57,0,12,0,200,0,40,0,0,0,66,0,0,0,207,0,0,0,44,0,126,0,104,0,160,0,100,0,87,0,151,0,229,0,197,0,250,0,233,0,161,0,2,0,241,0,111,0,205,0,59,0,80,0,0,0,0,0,61,0,67,0,201,0,167,0,252,0,81,0,53,0,181,0,0,0,130,0,239,0,0,0,46,0,70,0,183,0,0,0,123,0,60,0,111,0,140,0,0,0,75,0,6,0,0,0,201,0,0,0,128,0,217,0,95,0,0,0,133,0,100,0,222,0,23,0,190,0,0,0,0,0,99,0,31,0,4,0,0,0,86,0,213,0,191,0,176,0,169,0,178,0,0,0,67,0,217,0,30,0,187,0,177,0,208,0,54,0,247,0,16,0,75,0,209,0,109,0,55,0,129,0,58,0,42,0,0,0,63,0,24,0,62,0,0,0,208,0,0,0,27,0,204,0,52,0,143,0,67,0,0,0,0,0,116,0,187,0,0,0,238,0,7,0,0,0,0,0,247,0,13,0,0,0,43,0,43,0);
signal scenario_full  : scenario_type := (193,31,133,31,133,30,9,31,9,30,198,31,121,31,252,31,170,31,14,31,171,31,15,31,6,31,104,31,188,31,188,30,170,31,87,31,167,31,214,31,47,31,47,30,213,31,69,31,69,30,34,31,120,31,120,31,120,30,89,31,89,30,146,31,25,31,175,31,232,31,81,31,113,31,68,31,212,31,175,31,20,31,188,31,188,30,188,29,188,31,20,31,21,31,36,31,4,31,8,31,8,30,80,31,53,31,53,30,168,31,168,30,15,31,243,31,91,31,191,31,164,31,89,31,197,31,247,31,218,31,73,31,141,31,141,30,141,29,55,31,192,31,120,31,58,31,198,31,75,31,98,31,98,30,95,31,219,31,209,31,10,31,178,31,178,30,150,31,32,31,65,31,21,31,244,31,82,31,66,31,134,31,91,31,91,30,91,29,94,31,94,30,94,29,254,31,114,31,9,31,16,31,186,31,155,31,62,31,162,31,214,31,183,31,56,31,56,30,56,29,191,31,158,31,210,31,24,31,28,31,254,31,193,31,177,31,113,31,55,31,6,31,135,31,232,31,62,31,207,31,207,30,64,31,113,31,113,30,51,31,100,31,100,30,197,31,197,30,209,31,74,31,16,31,153,31,96,31,74,31,144,31,122,31,79,31,195,31,75,31,18,31,159,31,159,30,159,31,21,31,21,30,21,29,95,31,170,31,239,31,52,31,4,31,119,31,39,31,32,31,69,31,69,30,9,31,243,31,114,31,111,31,88,31,249,31,75,31,75,30,202,31,34,31,34,30,60,31,221,31,221,30,166,31,166,30,60,31,7,31,146,31,168,31,166,31,82,31,207,31,249,31,52,31,30,31,30,30,167,31,217,31,1,31,97,31,37,31,49,31,245,31,140,31,168,31,179,31,68,31,97,31,145,31,149,31,141,31,122,31,106,31,81,31,40,31,182,31,182,30,182,29,40,31,36,31,247,31,247,30,5,31,22,31,184,31,24,31,61,31,165,31,138,31,30,31,49,31,181,31,106,31,210,31,210,30,89,31,89,30,107,31,87,31,87,30,157,31,211,31,139,31,33,31,55,31,122,31,250,31,56,31,114,31,190,31,142,31,6,31,25,31,73,31,69,31,21,31,255,31,255,30,43,31,38,31,38,30,38,29,38,28,194,31,14,31,14,30,193,31,85,31,224,31,94,31,94,30,103,31,103,31,116,31,79,31,228,31,27,31,27,30,155,31,121,31,121,30,121,29,121,28,121,27,121,26,62,31,131,31,105,31,105,30,105,29,129,31,144,31,29,31,29,30,19,31,89,31,89,30,20,31,20,30,187,31,131,31,82,31,20,31,170,31,170,30,170,29,170,28,230,31,234,31,113,31,90,31,90,30,90,29,157,31,218,31,224,31,22,31,93,31,19,31,154,31,37,31,45,31,9,31,33,31,100,31,31,31,149,31,183,31,115,31,15,31,188,31,143,31,172,31,10,31,120,31,198,31,172,31,20,31,25,31,79,31,125,31,117,31,32,31,56,31,56,30,47,31,128,31,248,31,10,31,115,31,149,31,198,31,29,31,29,30,5,31,123,31,157,31,198,31,230,31,230,30,231,31,231,30,231,29,90,31,90,30,187,31,222,31,222,30,138,31,138,30,215,31,96,31,252,31,86,31,86,30,71,31,4,31,241,31,170,31,65,31,65,30,45,31,237,31,237,30,108,31,108,30,108,29,108,28,41,31,136,31,136,30,209,31,14,31,238,31,52,31,148,31,103,31,208,31,56,31,184,31,31,31,107,31,149,31,151,31,15,31,174,31,48,31,156,31,195,31,195,30,218,31,218,30,84,31,188,31,188,30,236,31,217,31,152,31,66,31,85,31,147,31,147,30,242,31,242,30,208,31,208,30,70,31,53,31,53,30,58,31,62,31,75,31,10,31,179,31,170,31,170,30,150,31,150,30,110,31,251,31,251,30,199,31,188,31,188,30,74,31,133,31,97,31,75,31,188,31,40,31,4,31,143,31,180,31,180,30,67,31,2,31,21,31,152,31,209,31,218,31,218,30,57,31,147,31,253,31,253,30,253,29,61,31,102,31,152,31,244,31,109,31,92,31,112,31,19,31,73,31,236,31,157,31,161,31,167,31,202,31,176,31,176,30,176,29,164,31,220,31,94,31,78,31,148,31,128,31,116,31,132,31,105,31,161,31,218,31,218,30,145,31,135,31,59,31,59,30,185,31,220,31,220,30,214,31,214,30,214,29,121,31,121,30,195,31,171,31,236,31,117,31,148,31,148,30,132,31,55,31,174,31,18,31,69,31,241,31,218,31,174,31,66,31,5,31,170,31,173,31,173,30,173,29,170,31,187,31,22,31,33,31,135,31,149,31,177,31,177,30,125,31,125,30,70,31,210,31,9,31,237,31,252,31,252,30,34,31,34,30,183,31,70,31,108,31,96,31,96,30,213,31,195,31,195,30,41,31,41,30,234,31,11,31,11,30,236,31,217,31,217,30,217,29,190,31,250,31,250,30,33,31,33,30,97,31,191,31,232,31,232,30,232,29,238,31,238,30,145,31,237,31,237,30,56,31,56,30,114,31,247,31,164,31,164,30,149,31,151,31,151,30,177,31,177,30,37,31,174,31,76,31,190,31,190,30,174,31,111,31,111,30,205,31,205,30,247,31,247,30,247,29,191,31,33,31,33,30,33,29,33,28,225,31,106,31,119,31,119,30,119,29,152,31,65,31,8,31,95,31,95,30,95,29,18,31,18,30,18,29,29,31,29,30,121,31,244,31,244,30,120,31,183,31,183,30,129,31,62,31,216,31,151,31,42,31,128,31,70,31,112,31,112,30,148,31,80,31,80,30,129,31,129,30,39,31,39,30,241,31,57,31,57,30,37,31,29,31,180,31,180,30,62,31,47,31,102,31,108,31,11,31,11,30,154,31,67,31,204,31,161,31,245,31,249,31,169,31,116,31,159,31,159,30,6,31,118,31,90,31,195,31,162,31,180,31,178,31,19,31,212,31,212,30,141,31,141,30,248,31,55,31,55,30,175,31,150,31,150,30,150,29,185,31,184,31,48,31,102,31,147,31,147,30,41,31,41,30,8,31,4,31,251,31,64,31,162,31,120,31,144,31,184,31,184,30,48,31,175,31,151,31,220,31,45,31,45,30,151,31,164,31,87,31,50,31,209,31,127,31,211,31,105,31,11,31,244,31,216,31,161,31,161,30,6,31,6,30,224,31,105,31,105,30,226,31,226,30,70,31,94,31,131,31,176,31,176,30,3,31,87,31,235,31,178,31,247,31,28,31,4,31,4,30,4,29,152,31,78,31,205,31,59,31,51,31,225,31,176,31,181,31,154,31,119,31,227,31,227,30,227,29,246,31,102,31,102,30,26,31,53,31,25,31,38,31,73,31,9,31,9,30,68,31,68,30,138,31,130,31,204,31,101,31,20,31,20,30,128,31,241,31,241,30,29,31,29,30,193,31,16,31,104,31,246,31,246,30,198,31,166,31,169,31,169,30,34,31,112,31,154,31,46,31,188,31,225,31,117,31,51,31,245,31,216,31,188,31,28,31,28,30,158,31,249,31,76,31,76,30,255,31,111,31,184,31,184,30,186,31,197,31,168,31,113,31,231,31,65,31,28,31,28,30,28,29,3,31,247,31,247,30,174,31,107,31,95,31,122,31,224,31,157,31,157,30,157,29,47,31,241,31,88,31,219,31,56,31,59,31,59,30,155,31,192,31,207,31,50,31,168,31,112,31,40,31,238,31,48,31,48,30,48,29,88,31,57,31,12,31,200,31,40,31,40,30,66,31,66,30,207,31,207,30,44,31,126,31,104,31,160,31,100,31,87,31,151,31,229,31,197,31,250,31,233,31,161,31,2,31,241,31,111,31,205,31,59,31,80,31,80,30,80,29,61,31,67,31,201,31,167,31,252,31,81,31,53,31,181,31,181,30,130,31,239,31,239,30,46,31,70,31,183,31,183,30,123,31,60,31,111,31,140,31,140,30,75,31,6,31,6,30,201,31,201,30,128,31,217,31,95,31,95,30,133,31,100,31,222,31,23,31,190,31,190,30,190,29,99,31,31,31,4,31,4,30,86,31,213,31,191,31,176,31,169,31,178,31,178,30,67,31,217,31,30,31,187,31,177,31,208,31,54,31,247,31,16,31,75,31,209,31,109,31,55,31,129,31,58,31,42,31,42,30,63,31,24,31,62,31,62,30,208,31,208,30,27,31,204,31,52,31,143,31,67,31,67,30,67,29,116,31,187,31,187,30,238,31,7,31,7,30,7,29,247,31,13,31,13,30,43,31,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
