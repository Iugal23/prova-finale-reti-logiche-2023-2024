-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 786;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,215,0,93,0,0,0,59,0,0,0,16,0,57,0,172,0,79,0,34,0,177,0,0,0,188,0,8,0,147,0,178,0,30,0,12,0,83,0,0,0,0,0,195,0,40,0,0,0,0,0,113,0,0,0,205,0,199,0,125,0,216,0,0,0,162,0,55,0,210,0,203,0,225,0,73,0,245,0,211,0,230,0,73,0,0,0,0,0,16,0,30,0,41,0,138,0,58,0,155,0,47,0,35,0,187,0,209,0,0,0,75,0,47,0,121,0,50,0,48,0,148,0,218,0,93,0,220,0,114,0,0,0,49,0,0,0,13,0,26,0,10,0,0,0,78,0,0,0,175,0,7,0,22,0,64,0,221,0,0,0,200,0,18,0,8,0,141,0,83,0,38,0,0,0,0,0,73,0,120,0,227,0,200,0,0,0,16,0,156,0,110,0,177,0,99,0,48,0,190,0,0,0,89,0,0,0,65,0,193,0,48,0,0,0,197,0,10,0,223,0,200,0,0,0,249,0,226,0,208,0,215,0,0,0,41,0,160,0,0,0,37,0,214,0,186,0,58,0,0,0,125,0,226,0,0,0,145,0,0,0,0,0,130,0,99,0,0,0,147,0,0,0,157,0,38,0,111,0,0,0,82,0,0,0,47,0,155,0,245,0,55,0,0,0,103,0,218,0,97,0,122,0,175,0,0,0,151,0,169,0,77,0,150,0,72,0,190,0,106,0,239,0,218,0,74,0,200,0,106,0,188,0,0,0,166,0,0,0,80,0,157,0,0,0,50,0,149,0,235,0,66,0,149,0,241,0,209,0,107,0,47,0,0,0,83,0,188,0,26,0,243,0,239,0,78,0,60,0,112,0,0,0,219,0,96,0,102,0,82,0,246,0,114,0,0,0,141,0,198,0,0,0,0,0,74,0,166,0,24,0,1,0,0,0,162,0,117,0,124,0,35,0,204,0,55,0,119,0,0,0,5,0,130,0,0,0,0,0,0,0,95,0,68,0,38,0,245,0,157,0,0,0,87,0,97,0,103,0,92,0,212,0,203,0,119,0,0,0,0,0,82,0,217,0,176,0,251,0,194,0,245,0,106,0,132,0,56,0,58,0,109,0,139,0,0,0,135,0,0,0,186,0,182,0,117,0,45,0,34,0,0,0,153,0,194,0,0,0,89,0,0,0,189,0,146,0,134,0,75,0,227,0,138,0,0,0,191,0,0,0,216,0,19,0,38,0,200,0,235,0,59,0,216,0,106,0,218,0,0,0,159,0,71,0,12,0,252,0,105,0,40,0,2,0,3,0,38,0,199,0,234,0,35,0,0,0,167,0,250,0,12,0,133,0,0,0,33,0,0,0,4,0,119,0,177,0,73,0,30,0,225,0,91,0,230,0,149,0,110,0,50,0,39,0,243,0,75,0,111,0,200,0,0,0,217,0,146,0,72,0,20,0,0,0,154,0,187,0,191,0,193,0,151,0,0,0,19,0,0,0,25,0,138,0,62,0,0,0,191,0,146,0,76,0,25,0,117,0,74,0,242,0,2,0,87,0,246,0,54,0,0,0,85,0,20,0,38,0,229,0,13,0,117,0,173,0,198,0,87,0,101,0,229,0,243,0,0,0,0,0,0,0,19,0,137,0,0,0,1,0,185,0,142,0,228,0,148,0,52,0,101,0,0,0,126,0,213,0,0,0,234,0,0,0,156,0,0,0,45,0,215,0,97,0,158,0,38,0,87,0,221,0,205,0,70,0,59,0,36,0,104,0,0,0,0,0,102,0,0,0,11,0,127,0,134,0,26,0,0,0,59,0,39,0,3,0,98,0,0,0,157,0,38,0,0,0,216,0,48,0,112,0,154,0,0,0,122,0,245,0,0,0,195,0,0,0,199,0,123,0,196,0,154,0,44,0,37,0,96,0,161,0,224,0,0,0,209,0,0,0,98,0,12,0,130,0,0,0,0,0,167,0,205,0,36,0,57,0,114,0,0,0,17,0,100,0,0,0,118,0,42,0,225,0,36,0,17,0,144,0,220,0,135,0,158,0,90,0,0,0,113,0,11,0,166,0,19,0,34,0,11,0,0,0,174,0,70,0,0,0,255,0,198,0,138,0,0,0,75,0,155,0,198,0,90,0,102,0,2,0,222,0,74,0,0,0,191,0,0,0,56,0,82,0,30,0,0,0,64,0,12,0,101,0,0,0,79,0,74,0,0,0,87,0,241,0,135,0,0,0,0,0,9,0,216,0,0,0,224,0,19,0,36,0,243,0,41,0,93,0,7,0,187,0,0,0,130,0,136,0,39,0,126,0,89,0,158,0,45,0,82,0,148,0,110,0,21,0,175,0,184,0,0,0,161,0,52,0,0,0,167,0,169,0,245,0,76,0,84,0,106,0,0,0,205,0,9,0,40,0,200,0,24,0,101,0,0,0,0,0,145,0,149,0,21,0,0,0,0,0,0,0,0,0,30,0,0,0,0,0,186,0,0,0,229,0,243,0,0,0,47,0,245,0,173,0,202,0,90,0,43,0,157,0,194,0,16,0,0,0,0,0,0,0,152,0,233,0,135,0,117,0,145,0,193,0,55,0,45,0,244,0,0,0,0,0,204,0,17,0,87,0,19,0,181,0,22,0,92,0,221,0,100,0,196,0,0,0,0,0,226,0,30,0,254,0,181,0,107,0,13,0,232,0,0,0,0,0,166,0,67,0,41,0,0,0,211,0,171,0,214,0,39,0,0,0,86,0,0,0,195,0,244,0,109,0,0,0,240,0,243,0,115,0,119,0,209,0,96,0,248,0,144,0,144,0,246,0,191,0,136,0,61,0,242,0,16,0,152,0,63,0,218,0,0,0,186,0,0,0,7,0,0,0,66,0,114,0,161,0,253,0,155,0,214,0,179,0,252,0,0,0,63,0,22,0,224,0,196,0,0,0,0,0,180,0,0,0,6,0,25,0,79,0,223,0,219,0,232,0,92,0,185,0,225,0,55,0,136,0,192,0,0,0,47,0,0,0,25,0,0,0,246,0,0,0,246,0,214,0,58,0,0,0,237,0,235,0,193,0,183,0,18,0,69,0,29,0,13,0,0,0,159,0,109,0,74,0,153,0,209,0,186,0,0,0,133,0,0,0,216,0,18,0,245,0,48,0,0,0,0,0,56,0,0,0,22,0,82,0,210,0,224,0,17,0,212,0,161,0,0,0,144,0,233,0,104,0,122,0,75,0,66,0,134,0,0,0,18,0,3,0,0,0,224,0,13,0,95,0,252,0,29,0,196,0,136,0,36,0,35,0,243,0,142,0,18,0,139,0,0,0,242,0,175,0,130,0,46,0,99,0,80,0,172,0,150,0,196,0,0,0,0,0,130,0,229,0,180,0,104,0,0,0,169,0,68,0,0,0,0,0,204,0,161,0,104,0,76,0,48,0,0,0,0,0,212,0,113,0,0,0,177,0,0,0,0,0,185,0,154,0,160,0,0,0,0,0,207,0,163,0,98,0,135,0,130,0,3,0,152,0,25,0,243,0,0,0,0,0);
signal scenario_full  : scenario_type := (219,31,215,31,93,31,93,30,59,31,59,30,16,31,57,31,172,31,79,31,34,31,177,31,177,30,188,31,8,31,147,31,178,31,30,31,12,31,83,31,83,30,83,29,195,31,40,31,40,30,40,29,113,31,113,30,205,31,199,31,125,31,216,31,216,30,162,31,55,31,210,31,203,31,225,31,73,31,245,31,211,31,230,31,73,31,73,30,73,29,16,31,30,31,41,31,138,31,58,31,155,31,47,31,35,31,187,31,209,31,209,30,75,31,47,31,121,31,50,31,48,31,148,31,218,31,93,31,220,31,114,31,114,30,49,31,49,30,13,31,26,31,10,31,10,30,78,31,78,30,175,31,7,31,22,31,64,31,221,31,221,30,200,31,18,31,8,31,141,31,83,31,38,31,38,30,38,29,73,31,120,31,227,31,200,31,200,30,16,31,156,31,110,31,177,31,99,31,48,31,190,31,190,30,89,31,89,30,65,31,193,31,48,31,48,30,197,31,10,31,223,31,200,31,200,30,249,31,226,31,208,31,215,31,215,30,41,31,160,31,160,30,37,31,214,31,186,31,58,31,58,30,125,31,226,31,226,30,145,31,145,30,145,29,130,31,99,31,99,30,147,31,147,30,157,31,38,31,111,31,111,30,82,31,82,30,47,31,155,31,245,31,55,31,55,30,103,31,218,31,97,31,122,31,175,31,175,30,151,31,169,31,77,31,150,31,72,31,190,31,106,31,239,31,218,31,74,31,200,31,106,31,188,31,188,30,166,31,166,30,80,31,157,31,157,30,50,31,149,31,235,31,66,31,149,31,241,31,209,31,107,31,47,31,47,30,83,31,188,31,26,31,243,31,239,31,78,31,60,31,112,31,112,30,219,31,96,31,102,31,82,31,246,31,114,31,114,30,141,31,198,31,198,30,198,29,74,31,166,31,24,31,1,31,1,30,162,31,117,31,124,31,35,31,204,31,55,31,119,31,119,30,5,31,130,31,130,30,130,29,130,28,95,31,68,31,38,31,245,31,157,31,157,30,87,31,97,31,103,31,92,31,212,31,203,31,119,31,119,30,119,29,82,31,217,31,176,31,251,31,194,31,245,31,106,31,132,31,56,31,58,31,109,31,139,31,139,30,135,31,135,30,186,31,182,31,117,31,45,31,34,31,34,30,153,31,194,31,194,30,89,31,89,30,189,31,146,31,134,31,75,31,227,31,138,31,138,30,191,31,191,30,216,31,19,31,38,31,200,31,235,31,59,31,216,31,106,31,218,31,218,30,159,31,71,31,12,31,252,31,105,31,40,31,2,31,3,31,38,31,199,31,234,31,35,31,35,30,167,31,250,31,12,31,133,31,133,30,33,31,33,30,4,31,119,31,177,31,73,31,30,31,225,31,91,31,230,31,149,31,110,31,50,31,39,31,243,31,75,31,111,31,200,31,200,30,217,31,146,31,72,31,20,31,20,30,154,31,187,31,191,31,193,31,151,31,151,30,19,31,19,30,25,31,138,31,62,31,62,30,191,31,146,31,76,31,25,31,117,31,74,31,242,31,2,31,87,31,246,31,54,31,54,30,85,31,20,31,38,31,229,31,13,31,117,31,173,31,198,31,87,31,101,31,229,31,243,31,243,30,243,29,243,28,19,31,137,31,137,30,1,31,185,31,142,31,228,31,148,31,52,31,101,31,101,30,126,31,213,31,213,30,234,31,234,30,156,31,156,30,45,31,215,31,97,31,158,31,38,31,87,31,221,31,205,31,70,31,59,31,36,31,104,31,104,30,104,29,102,31,102,30,11,31,127,31,134,31,26,31,26,30,59,31,39,31,3,31,98,31,98,30,157,31,38,31,38,30,216,31,48,31,112,31,154,31,154,30,122,31,245,31,245,30,195,31,195,30,199,31,123,31,196,31,154,31,44,31,37,31,96,31,161,31,224,31,224,30,209,31,209,30,98,31,12,31,130,31,130,30,130,29,167,31,205,31,36,31,57,31,114,31,114,30,17,31,100,31,100,30,118,31,42,31,225,31,36,31,17,31,144,31,220,31,135,31,158,31,90,31,90,30,113,31,11,31,166,31,19,31,34,31,11,31,11,30,174,31,70,31,70,30,255,31,198,31,138,31,138,30,75,31,155,31,198,31,90,31,102,31,2,31,222,31,74,31,74,30,191,31,191,30,56,31,82,31,30,31,30,30,64,31,12,31,101,31,101,30,79,31,74,31,74,30,87,31,241,31,135,31,135,30,135,29,9,31,216,31,216,30,224,31,19,31,36,31,243,31,41,31,93,31,7,31,187,31,187,30,130,31,136,31,39,31,126,31,89,31,158,31,45,31,82,31,148,31,110,31,21,31,175,31,184,31,184,30,161,31,52,31,52,30,167,31,169,31,245,31,76,31,84,31,106,31,106,30,205,31,9,31,40,31,200,31,24,31,101,31,101,30,101,29,145,31,149,31,21,31,21,30,21,29,21,28,21,27,30,31,30,30,30,29,186,31,186,30,229,31,243,31,243,30,47,31,245,31,173,31,202,31,90,31,43,31,157,31,194,31,16,31,16,30,16,29,16,28,152,31,233,31,135,31,117,31,145,31,193,31,55,31,45,31,244,31,244,30,244,29,204,31,17,31,87,31,19,31,181,31,22,31,92,31,221,31,100,31,196,31,196,30,196,29,226,31,30,31,254,31,181,31,107,31,13,31,232,31,232,30,232,29,166,31,67,31,41,31,41,30,211,31,171,31,214,31,39,31,39,30,86,31,86,30,195,31,244,31,109,31,109,30,240,31,243,31,115,31,119,31,209,31,96,31,248,31,144,31,144,31,246,31,191,31,136,31,61,31,242,31,16,31,152,31,63,31,218,31,218,30,186,31,186,30,7,31,7,30,66,31,114,31,161,31,253,31,155,31,214,31,179,31,252,31,252,30,63,31,22,31,224,31,196,31,196,30,196,29,180,31,180,30,6,31,25,31,79,31,223,31,219,31,232,31,92,31,185,31,225,31,55,31,136,31,192,31,192,30,47,31,47,30,25,31,25,30,246,31,246,30,246,31,214,31,58,31,58,30,237,31,235,31,193,31,183,31,18,31,69,31,29,31,13,31,13,30,159,31,109,31,74,31,153,31,209,31,186,31,186,30,133,31,133,30,216,31,18,31,245,31,48,31,48,30,48,29,56,31,56,30,22,31,82,31,210,31,224,31,17,31,212,31,161,31,161,30,144,31,233,31,104,31,122,31,75,31,66,31,134,31,134,30,18,31,3,31,3,30,224,31,13,31,95,31,252,31,29,31,196,31,136,31,36,31,35,31,243,31,142,31,18,31,139,31,139,30,242,31,175,31,130,31,46,31,99,31,80,31,172,31,150,31,196,31,196,30,196,29,130,31,229,31,180,31,104,31,104,30,169,31,68,31,68,30,68,29,204,31,161,31,104,31,76,31,48,31,48,30,48,29,212,31,113,31,113,30,177,31,177,30,177,29,185,31,154,31,160,31,160,30,160,29,207,31,163,31,98,31,135,31,130,31,3,31,152,31,25,31,243,31,243,30,243,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
