-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 836;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,154,0,57,0,0,0,131,0,3,0,53,0,0,0,136,0,50,0,62,0,10,0,34,0,37,0,59,0,226,0,55,0,0,0,157,0,230,0,39,0,0,0,0,0,87,0,0,0,6,0,56,0,123,0,0,0,0,0,53,0,171,0,232,0,0,0,0,0,60,0,191,0,4,0,217,0,0,0,168,0,191,0,50,0,194,0,140,0,179,0,204,0,161,0,179,0,199,0,5,0,96,0,190,0,144,0,0,0,149,0,228,0,212,0,103,0,69,0,12,0,249,0,229,0,0,0,54,0,137,0,0,0,232,0,191,0,219,0,108,0,0,0,0,0,148,0,233,0,15,0,225,0,242,0,33,0,67,0,0,0,165,0,0,0,0,0,200,0,156,0,221,0,244,0,52,0,75,0,93,0,187,0,35,0,128,0,126,0,156,0,64,0,0,0,54,0,73,0,0,0,55,0,14,0,0,0,226,0,183,0,69,0,116,0,0,0,224,0,221,0,61,0,165,0,248,0,176,0,209,0,195,0,2,0,141,0,231,0,0,0,75,0,102,0,107,0,131,0,131,0,0,0,198,0,212,0,165,0,180,0,0,0,243,0,96,0,71,0,94,0,99,0,41,0,34,0,159,0,249,0,109,0,54,0,97,0,0,0,0,0,238,0,19,0,197,0,141,0,91,0,134,0,172,0,150,0,99,0,21,0,0,0,185,0,15,0,171,0,69,0,44,0,103,0,0,0,187,0,106,0,101,0,207,0,177,0,173,0,120,0,148,0,0,0,0,0,194,0,77,0,123,0,20,0,0,0,0,0,143,0,40,0,120,0,135,0,132,0,220,0,240,0,0,0,112,0,108,0,203,0,0,0,221,0,200,0,47,0,201,0,0,0,39,0,32,0,0,0,208,0,243,0,164,0,222,0,145,0,102,0,0,0,239,0,42,0,123,0,99,0,0,0,40,0,159,0,250,0,0,0,185,0,53,0,0,0,0,0,46,0,186,0,255,0,156,0,6,0,193,0,0,0,209,0,0,0,49,0,0,0,233,0,82,0,166,0,49,0,152,0,125,0,0,0,53,0,192,0,254,0,253,0,0,0,42,0,46,0,25,0,49,0,68,0,191,0,144,0,198,0,84,0,72,0,159,0,196,0,234,0,0,0,85,0,0,0,133,0,247,0,95,0,97,0,253,0,239,0,0,0,0,0,0,0,41,0,40,0,12,0,188,0,0,0,68,0,0,0,181,0,72,0,47,0,149,0,72,0,255,0,119,0,0,0,0,0,0,0,163,0,196,0,84,0,201,0,0,0,230,0,71,0,45,0,236,0,212,0,112,0,31,0,0,0,132,0,115,0,129,0,60,0,0,0,241,0,202,0,11,0,244,0,89,0,249,0,182,0,0,0,124,0,22,0,0,0,156,0,5,0,200,0,148,0,33,0,198,0,163,0,0,0,253,0,0,0,0,0,0,0,205,0,0,0,2,0,80,0,191,0,31,0,0,0,205,0,0,0,0,0,143,0,160,0,59,0,99,0,0,0,90,0,21,0,118,0,218,0,10,0,136,0,0,0,31,0,133,0,0,0,73,0,211,0,102,0,0,0,77,0,0,0,127,0,194,0,15,0,254,0,0,0,0,0,142,0,234,0,63,0,0,0,162,0,213,0,251,0,237,0,151,0,121,0,158,0,27,0,218,0,7,0,16,0,124,0,70,0,5,0,222,0,12,0,0,0,119,0,137,0,116,0,4,0,17,0,254,0,106,0,204,0,0,0,0,0,188,0,183,0,75,0,187,0,59,0,242,0,0,0,0,0,136,0,222,0,21,0,208,0,120,0,203,0,128,0,143,0,7,0,235,0,69,0,23,0,245,0,1,0,97,0,166,0,38,0,130,0,55,0,155,0,103,0,39,0,166,0,0,0,0,0,0,0,23,0,160,0,96,0,55,0,232,0,222,0,0,0,246,0,0,0,132,0,0,0,68,0,192,0,0,0,63,0,0,0,8,0,94,0,114,0,221,0,122,0,14,0,74,0,143,0,116,0,76,0,200,0,202,0,0,0,0,0,98,0,209,0,99,0,114,0,8,0,94,0,246,0,180,0,192,0,128,0,24,0,0,0,2,0,114,0,28,0,160,0,190,0,171,0,198,0,186,0,105,0,48,0,45,0,0,0,136,0,0,0,161,0,40,0,122,0,46,0,124,0,15,0,0,0,105,0,139,0,238,0,0,0,212,0,1,0,0,0,126,0,155,0,2,0,0,0,55,0,90,0,182,0,12,0,0,0,215,0,34,0,0,0,194,0,58,0,33,0,0,0,0,0,26,0,52,0,96,0,112,0,0,0,253,0,98,0,111,0,58,0,246,0,236,0,231,0,119,0,16,0,6,0,74,0,254,0,108,0,8,0,181,0,217,0,137,0,55,0,30,0,55,0,34,0,113,0,0,0,0,0,239,0,215,0,230,0,167,0,208,0,10,0,44,0,209,0,78,0,197,0,239,0,79,0,172,0,0,0,40,0,203,0,174,0,110,0,200,0,0,0,0,0,197,0,210,0,161,0,0,0,25,0,40,0,124,0,158,0,0,0,193,0,55,0,56,0,0,0,74,0,164,0,0,0,0,0,240,0,0,0,23,0,212,0,0,0,24,0,0,0,36,0,213,0,0,0,65,0,92,0,92,0,0,0,0,0,202,0,239,0,86,0,163,0,10,0,54,0,0,0,105,0,0,0,120,0,0,0,245,0,169,0,212,0,230,0,0,0,133,0,188,0,0,0,0,0,224,0,114,0,172,0,153,0,94,0,163,0,128,0,179,0,76,0,188,0,62,0,41,0,164,0,61,0,235,0,106,0,186,0,245,0,0,0,163,0,185,0,94,0,0,0,128,0,95,0,0,0,54,0,0,0,0,0,89,0,203,0,150,0,0,0,59,0,72,0,227,0,147,0,115,0,53,0,172,0,0,0,42,0,177,0,0,0,0,0,48,0,210,0,238,0,60,0,61,0,70,0,233,0,205,0,191,0,59,0,33,0,142,0,66,0,0,0,0,0,79,0,220,0,0,0,0,0,206,0,80,0,0,0,31,0,160,0,163,0,234,0,244,0,208,0,106,0,100,0,251,0,6,0,0,0,65,0,187,0,103,0,51,0,214,0,167,0,0,0,242,0,183,0,250,0,128,0,229,0,0,0,181,0,0,0,0,0,0,0,24,0,219,0,23,0,67,0,73,0,0,0,92,0,66,0,0,0,0,0,85,0,248,0,42,0,240,0,0,0,94,0,227,0,0,0,66,0,227,0,23,0,240,0,0,0,247,0,210,0,210,0,4,0,220,0,0,0,0,0,223,0,57,0,0,0,218,0,0,0,40,0,81,0,188,0,230,0,99,0,0,0,38,0,49,0,252,0,239,0,49,0,0,0,154,0,224,0,156,0,219,0,147,0,41,0,91,0,112,0,214,0,53,0,73,0,102,0,238,0,206,0,104,0,111,0,74,0,142,0,206,0,116,0,140,0,0,0,0,0,253,0,0,0,255,0,0,0,144,0,23,0,77,0,0,0,103,0,54,0,23,0,0,0,246,0,95,0,153,0,168,0,148,0,46,0,0,0,202,0,190,0,148,0,26,0,0,0,12,0,228,0,14,0,123,0,0,0,14,0,254,0,243,0,0,0,4,0,124,0,175,0,84,0,0,0,178,0,103,0,124,0,0,0,53,0,0,0,223,0,154,0,72,0,45,0,184,0,140,0,196,0,101,0,0,0,195,0);
signal scenario_full  : scenario_type := (0,0,154,31,57,31,57,30,131,31,3,31,53,31,53,30,136,31,50,31,62,31,10,31,34,31,37,31,59,31,226,31,55,31,55,30,157,31,230,31,39,31,39,30,39,29,87,31,87,30,6,31,56,31,123,31,123,30,123,29,53,31,171,31,232,31,232,30,232,29,60,31,191,31,4,31,217,31,217,30,168,31,191,31,50,31,194,31,140,31,179,31,204,31,161,31,179,31,199,31,5,31,96,31,190,31,144,31,144,30,149,31,228,31,212,31,103,31,69,31,12,31,249,31,229,31,229,30,54,31,137,31,137,30,232,31,191,31,219,31,108,31,108,30,108,29,148,31,233,31,15,31,225,31,242,31,33,31,67,31,67,30,165,31,165,30,165,29,200,31,156,31,221,31,244,31,52,31,75,31,93,31,187,31,35,31,128,31,126,31,156,31,64,31,64,30,54,31,73,31,73,30,55,31,14,31,14,30,226,31,183,31,69,31,116,31,116,30,224,31,221,31,61,31,165,31,248,31,176,31,209,31,195,31,2,31,141,31,231,31,231,30,75,31,102,31,107,31,131,31,131,31,131,30,198,31,212,31,165,31,180,31,180,30,243,31,96,31,71,31,94,31,99,31,41,31,34,31,159,31,249,31,109,31,54,31,97,31,97,30,97,29,238,31,19,31,197,31,141,31,91,31,134,31,172,31,150,31,99,31,21,31,21,30,185,31,15,31,171,31,69,31,44,31,103,31,103,30,187,31,106,31,101,31,207,31,177,31,173,31,120,31,148,31,148,30,148,29,194,31,77,31,123,31,20,31,20,30,20,29,143,31,40,31,120,31,135,31,132,31,220,31,240,31,240,30,112,31,108,31,203,31,203,30,221,31,200,31,47,31,201,31,201,30,39,31,32,31,32,30,208,31,243,31,164,31,222,31,145,31,102,31,102,30,239,31,42,31,123,31,99,31,99,30,40,31,159,31,250,31,250,30,185,31,53,31,53,30,53,29,46,31,186,31,255,31,156,31,6,31,193,31,193,30,209,31,209,30,49,31,49,30,233,31,82,31,166,31,49,31,152,31,125,31,125,30,53,31,192,31,254,31,253,31,253,30,42,31,46,31,25,31,49,31,68,31,191,31,144,31,198,31,84,31,72,31,159,31,196,31,234,31,234,30,85,31,85,30,133,31,247,31,95,31,97,31,253,31,239,31,239,30,239,29,239,28,41,31,40,31,12,31,188,31,188,30,68,31,68,30,181,31,72,31,47,31,149,31,72,31,255,31,119,31,119,30,119,29,119,28,163,31,196,31,84,31,201,31,201,30,230,31,71,31,45,31,236,31,212,31,112,31,31,31,31,30,132,31,115,31,129,31,60,31,60,30,241,31,202,31,11,31,244,31,89,31,249,31,182,31,182,30,124,31,22,31,22,30,156,31,5,31,200,31,148,31,33,31,198,31,163,31,163,30,253,31,253,30,253,29,253,28,205,31,205,30,2,31,80,31,191,31,31,31,31,30,205,31,205,30,205,29,143,31,160,31,59,31,99,31,99,30,90,31,21,31,118,31,218,31,10,31,136,31,136,30,31,31,133,31,133,30,73,31,211,31,102,31,102,30,77,31,77,30,127,31,194,31,15,31,254,31,254,30,254,29,142,31,234,31,63,31,63,30,162,31,213,31,251,31,237,31,151,31,121,31,158,31,27,31,218,31,7,31,16,31,124,31,70,31,5,31,222,31,12,31,12,30,119,31,137,31,116,31,4,31,17,31,254,31,106,31,204,31,204,30,204,29,188,31,183,31,75,31,187,31,59,31,242,31,242,30,242,29,136,31,222,31,21,31,208,31,120,31,203,31,128,31,143,31,7,31,235,31,69,31,23,31,245,31,1,31,97,31,166,31,38,31,130,31,55,31,155,31,103,31,39,31,166,31,166,30,166,29,166,28,23,31,160,31,96,31,55,31,232,31,222,31,222,30,246,31,246,30,132,31,132,30,68,31,192,31,192,30,63,31,63,30,8,31,94,31,114,31,221,31,122,31,14,31,74,31,143,31,116,31,76,31,200,31,202,31,202,30,202,29,98,31,209,31,99,31,114,31,8,31,94,31,246,31,180,31,192,31,128,31,24,31,24,30,2,31,114,31,28,31,160,31,190,31,171,31,198,31,186,31,105,31,48,31,45,31,45,30,136,31,136,30,161,31,40,31,122,31,46,31,124,31,15,31,15,30,105,31,139,31,238,31,238,30,212,31,1,31,1,30,126,31,155,31,2,31,2,30,55,31,90,31,182,31,12,31,12,30,215,31,34,31,34,30,194,31,58,31,33,31,33,30,33,29,26,31,52,31,96,31,112,31,112,30,253,31,98,31,111,31,58,31,246,31,236,31,231,31,119,31,16,31,6,31,74,31,254,31,108,31,8,31,181,31,217,31,137,31,55,31,30,31,55,31,34,31,113,31,113,30,113,29,239,31,215,31,230,31,167,31,208,31,10,31,44,31,209,31,78,31,197,31,239,31,79,31,172,31,172,30,40,31,203,31,174,31,110,31,200,31,200,30,200,29,197,31,210,31,161,31,161,30,25,31,40,31,124,31,158,31,158,30,193,31,55,31,56,31,56,30,74,31,164,31,164,30,164,29,240,31,240,30,23,31,212,31,212,30,24,31,24,30,36,31,213,31,213,30,65,31,92,31,92,31,92,30,92,29,202,31,239,31,86,31,163,31,10,31,54,31,54,30,105,31,105,30,120,31,120,30,245,31,169,31,212,31,230,31,230,30,133,31,188,31,188,30,188,29,224,31,114,31,172,31,153,31,94,31,163,31,128,31,179,31,76,31,188,31,62,31,41,31,164,31,61,31,235,31,106,31,186,31,245,31,245,30,163,31,185,31,94,31,94,30,128,31,95,31,95,30,54,31,54,30,54,29,89,31,203,31,150,31,150,30,59,31,72,31,227,31,147,31,115,31,53,31,172,31,172,30,42,31,177,31,177,30,177,29,48,31,210,31,238,31,60,31,61,31,70,31,233,31,205,31,191,31,59,31,33,31,142,31,66,31,66,30,66,29,79,31,220,31,220,30,220,29,206,31,80,31,80,30,31,31,160,31,163,31,234,31,244,31,208,31,106,31,100,31,251,31,6,31,6,30,65,31,187,31,103,31,51,31,214,31,167,31,167,30,242,31,183,31,250,31,128,31,229,31,229,30,181,31,181,30,181,29,181,28,24,31,219,31,23,31,67,31,73,31,73,30,92,31,66,31,66,30,66,29,85,31,248,31,42,31,240,31,240,30,94,31,227,31,227,30,66,31,227,31,23,31,240,31,240,30,247,31,210,31,210,31,4,31,220,31,220,30,220,29,223,31,57,31,57,30,218,31,218,30,40,31,81,31,188,31,230,31,99,31,99,30,38,31,49,31,252,31,239,31,49,31,49,30,154,31,224,31,156,31,219,31,147,31,41,31,91,31,112,31,214,31,53,31,73,31,102,31,238,31,206,31,104,31,111,31,74,31,142,31,206,31,116,31,140,31,140,30,140,29,253,31,253,30,255,31,255,30,144,31,23,31,77,31,77,30,103,31,54,31,23,31,23,30,246,31,95,31,153,31,168,31,148,31,46,31,46,30,202,31,190,31,148,31,26,31,26,30,12,31,228,31,14,31,123,31,123,30,14,31,254,31,243,31,243,30,4,31,124,31,175,31,84,31,84,30,178,31,103,31,124,31,124,30,53,31,53,30,223,31,154,31,72,31,45,31,184,31,140,31,196,31,101,31,101,30,195,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
