-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 283;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,78,0,151,0,0,0,0,0,61,0,85,0,34,0,90,0,24,0,6,0,227,0,1,0,215,0,154,0,0,0,228,0,22,0,197,0,0,0,76,0,0,0,14,0,147,0,0,0,5,0,0,0,215,0,185,0,212,0,124,0,0,0,249,0,221,0,168,0,88,0,97,0,222,0,248,0,62,0,134,0,3,0,123,0,169,0,52,0,0,0,0,0,161,0,151,0,147,0,31,0,66,0,255,0,9,0,0,0,0,0,0,0,144,0,0,0,234,0,42,0,139,0,45,0,213,0,209,0,119,0,121,0,95,0,110,0,148,0,0,0,0,0,214,0,70,0,0,0,249,0,25,0,170,0,22,0,99,0,127,0,68,0,47,0,230,0,157,0,0,0,104,0,189,0,240,0,73,0,79,0,134,0,0,0,228,0,191,0,27,0,99,0,0,0,134,0,176,0,116,0,18,0,206,0,0,0,151,0,125,0,154,0,194,0,70,0,116,0,43,0,52,0,199,0,208,0,14,0,155,0,72,0,120,0,251,0,181,0,97,0,213,0,86,0,38,0,245,0,73,0,193,0,120,0,130,0,0,0,193,0,0,0,0,0,0,0,175,0,8,0,12,0,175,0,58,0,168,0,169,0,0,0,81,0,117,0,225,0,240,0,225,0,0,0,96,0,204,0,140,0,213,0,58,0,70,0,113,0,94,0,144,0,0,0,236,0,106,0,255,0,237,0,108,0,128,0,112,0,0,0,33,0,169,0,19,0,92,0,80,0,0,0,2,0,151,0,234,0,85,0,0,0,227,0,0,0,0,0,207,0,0,0,19,0,62,0,21,0,192,0,195,0,255,0,198,0,74,0,203,0,117,0,139,0,133,0,95,0,0,0,196,0,203,0,157,0,227,0,232,0,28,0,13,0,45,0,161,0,146,0,116,0,26,0,0,0,214,0,0,0,36,0,62,0,70,0,62,0,52,0,255,0,106,0,0,0,210,0,226,0,206,0,226,0,0,0,164,0,0,0,250,0,0,0,239,0,0,0,54,0,135,0,20,0,223,0,0,0,123,0,206,0,73,0,30,0,112,0,191,0,199,0,157,0,252,0,106,0,0,0,174,0,240,0,12,0,80,0,1,0,245,0,238,0,0,0,165,0,53,0,74,0,205,0,131,0,0,0,240,0,109,0,88,0,0,0,228,0,27,0,82,0,0,0,249,0,0,0,60,0,68,0,170,0,46,0,38,0,0,0,26,0,50,0,83,0,194,0,0,0,248,0,51,0);
signal scenario_full  : scenario_type := (0,0,78,31,151,31,151,30,151,29,61,31,85,31,34,31,90,31,24,31,6,31,227,31,1,31,215,31,154,31,154,30,228,31,22,31,197,31,197,30,76,31,76,30,14,31,147,31,147,30,5,31,5,30,215,31,185,31,212,31,124,31,124,30,249,31,221,31,168,31,88,31,97,31,222,31,248,31,62,31,134,31,3,31,123,31,169,31,52,31,52,30,52,29,161,31,151,31,147,31,31,31,66,31,255,31,9,31,9,30,9,29,9,28,144,31,144,30,234,31,42,31,139,31,45,31,213,31,209,31,119,31,121,31,95,31,110,31,148,31,148,30,148,29,214,31,70,31,70,30,249,31,25,31,170,31,22,31,99,31,127,31,68,31,47,31,230,31,157,31,157,30,104,31,189,31,240,31,73,31,79,31,134,31,134,30,228,31,191,31,27,31,99,31,99,30,134,31,176,31,116,31,18,31,206,31,206,30,151,31,125,31,154,31,194,31,70,31,116,31,43,31,52,31,199,31,208,31,14,31,155,31,72,31,120,31,251,31,181,31,97,31,213,31,86,31,38,31,245,31,73,31,193,31,120,31,130,31,130,30,193,31,193,30,193,29,193,28,175,31,8,31,12,31,175,31,58,31,168,31,169,31,169,30,81,31,117,31,225,31,240,31,225,31,225,30,96,31,204,31,140,31,213,31,58,31,70,31,113,31,94,31,144,31,144,30,236,31,106,31,255,31,237,31,108,31,128,31,112,31,112,30,33,31,169,31,19,31,92,31,80,31,80,30,2,31,151,31,234,31,85,31,85,30,227,31,227,30,227,29,207,31,207,30,19,31,62,31,21,31,192,31,195,31,255,31,198,31,74,31,203,31,117,31,139,31,133,31,95,31,95,30,196,31,203,31,157,31,227,31,232,31,28,31,13,31,45,31,161,31,146,31,116,31,26,31,26,30,214,31,214,30,36,31,62,31,70,31,62,31,52,31,255,31,106,31,106,30,210,31,226,31,206,31,226,31,226,30,164,31,164,30,250,31,250,30,239,31,239,30,54,31,135,31,20,31,223,31,223,30,123,31,206,31,73,31,30,31,112,31,191,31,199,31,157,31,252,31,106,31,106,30,174,31,240,31,12,31,80,31,1,31,245,31,238,31,238,30,165,31,53,31,74,31,205,31,131,31,131,30,240,31,109,31,88,31,88,30,228,31,27,31,82,31,82,30,249,31,249,30,60,31,68,31,170,31,46,31,38,31,38,30,26,31,50,31,83,31,194,31,194,30,248,31,51,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
