-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_117 is
end project_tb_117;

architecture project_tb_arch_117 of project_tb_117 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 708;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (104,0,48,0,124,0,174,0,182,0,138,0,150,0,0,0,0,0,0,0,0,0,0,0,24,0,143,0,122,0,226,0,204,0,168,0,153,0,145,0,82,0,65,0,0,0,172,0,116,0,0,0,75,0,158,0,0,0,19,0,0,0,229,0,245,0,145,0,121,0,61,0,17,0,241,0,111,0,176,0,168,0,20,0,182,0,0,0,25,0,0,0,0,0,0,0,230,0,204,0,99,0,33,0,183,0,182,0,152,0,77,0,31,0,148,0,75,0,244,0,237,0,234,0,7,0,48,0,103,0,53,0,0,0,230,0,95,0,109,0,0,0,187,0,194,0,11,0,203,0,11,0,95,0,122,0,0,0,166,0,204,0,217,0,172,0,98,0,241,0,82,0,19,0,16,0,0,0,0,0,96,0,0,0,169,0,109,0,0,0,134,0,70,0,196,0,206,0,30,0,232,0,104,0,223,0,201,0,233,0,252,0,220,0,155,0,111,0,25,0,24,0,0,0,0,0,85,0,0,0,0,0,191,0,144,0,0,0,135,0,0,0,140,0,200,0,52,0,244,0,103,0,171,0,218,0,55,0,135,0,28,0,183,0,101,0,19,0,131,0,113,0,219,0,23,0,0,0,129,0,66,0,158,0,20,0,205,0,42,0,190,0,0,0,119,0,142,0,48,0,36,0,71,0,0,0,110,0,153,0,0,0,176,0,172,0,153,0,13,0,0,0,190,0,39,0,137,0,0,0,164,0,244,0,0,0,224,0,124,0,96,0,199,0,0,0,231,0,211,0,165,0,0,0,0,0,123,0,0,0,100,0,0,0,198,0,222,0,130,0,233,0,27,0,189,0,68,0,179,0,112,0,0,0,232,0,130,0,252,0,159,0,5,0,9,0,66,0,181,0,95,0,185,0,36,0,243,0,19,0,244,0,221,0,5,0,244,0,112,0,0,0,108,0,125,0,251,0,187,0,128,0,107,0,8,0,0,0,73,0,82,0,18,0,6,0,248,0,83,0,238,0,24,0,178,0,207,0,13,0,50,0,180,0,0,0,0,0,1,0,0,0,143,0,89,0,46,0,155,0,237,0,103,0,19,0,0,0,168,0,0,0,226,0,117,0,113,0,27,0,204,0,230,0,238,0,0,0,0,0,0,0,174,0,141,0,129,0,213,0,0,0,226,0,225,0,0,0,141,0,175,0,0,0,36,0,0,0,0,0,167,0,213,0,116,0,162,0,8,0,68,0,0,0,239,0,11,0,0,0,159,0,116,0,238,0,174,0,37,0,239,0,253,0,14,0,72,0,220,0,185,0,227,0,12,0,102,0,91,0,150,0,0,0,157,0,201,0,95,0,185,0,219,0,0,0,0,0,107,0,73,0,21,0,70,0,183,0,51,0,180,0,0,0,120,0,241,0,143,0,185,0,198,0,50,0,159,0,170,0,94,0,0,0,76,0,0,0,67,0,0,0,187,0,243,0,114,0,51,0,160,0,143,0,94,0,42,0,0,0,9,0,91,0,75,0,0,0,23,0,162,0,248,0,206,0,0,0,0,0,55,0,182,0,64,0,107,0,0,0,113,0,0,0,103,0,140,0,205,0,218,0,0,0,203,0,119,0,9,0,213,0,0,0,204,0,116,0,55,0,117,0,40,0,186,0,17,0,222,0,0,0,214,0,239,0,0,0,237,0,0,0,16,0,0,0,0,0,0,0,24,0,111,0,131,0,40,0,166,0,0,0,158,0,138,0,176,0,0,0,17,0,231,0,232,0,224,0,62,0,8,0,9,0,168,0,222,0,143,0,10,0,237,0,0,0,238,0,0,0,116,0,113,0,0,0,178,0,0,0,136,0,0,0,30,0,103,0,197,0,0,0,27,0,50,0,191,0,209,0,142,0,0,0,26,0,6,0,103,0,122,0,19,0,94,0,6,0,0,0,148,0,0,0,0,0,188,0,10,0,0,0,129,0,255,0,2,0,32,0,223,0,0,0,244,0,63,0,149,0,96,0,251,0,83,0,185,0,156,0,177,0,231,0,12,0,0,0,29,0,37,0,67,0,160,0,0,0,0,0,0,0,249,0,106,0,213,0,0,0,121,0,106,0,105,0,74,0,9,0,133,0,42,0,99,0,4,0,31,0,130,0,150,0,0,0,0,0,184,0,198,0,211,0,33,0,0,0,0,0,16,0,242,0,11,0,202,0,59,0,196,0,76,0,148,0,81,0,0,0,239,0,190,0,186,0,0,0,228,0,211,0,253,0,153,0,195,0,5,0,9,0,111,0,26,0,175,0,160,0,117,0,121,0,198,0,196,0,16,0,151,0,196,0,0,0,32,0,8,0,168,0,77,0,37,0,247,0,52,0,162,0,0,0,0,0,236,0,21,0,63,0,103,0,162,0,75,0,0,0,45,0,77,0,175,0,110,0,68,0,240,0,206,0,254,0,188,0,139,0,219,0,80,0,0,0,79,0,189,0,108,0,111,0,136,0,89,0,146,0,221,0,145,0,0,0,0,0,155,0,237,0,218,0,173,0,68,0,241,0,8,0,112,0,47,0,172,0,16,0,219,0,115,0,69,0,60,0,0,0,13,0,48,0,0,0,106,0,86,0,7,0,161,0,75,0,243,0,235,0,11,0,0,0,18,0,14,0,0,0,45,0,0,0,0,0,245,0,0,0,178,0,173,0,34,0,243,0,127,0,51,0,125,0,115,0,42,0,0,0,109,0,148,0,156,0,124,0,109,0,1,0,93,0,186,0,66,0,132,0,248,0,171,0,4,0,0,0,0,0,72,0,0,0,193,0,162,0,167,0,140,0,166,0,212,0,20,0,78,0,32,0,61,0,211,0,50,0,64,0,249,0,26,0,33,0,65,0,0,0,97,0,72,0,6,0,216,0,209,0,8,0,186,0,0,0,206,0,71,0,94,0,219,0,0,0,0,0,0,0,137,0,22,0,141,0,185,0,241,0,92,0,53,0,117,0,0,0,64,0,0,0,0,0,27,0,9,0,0,0,6,0,2,0,125,0,170,0,90,0,0,0,216,0,244,0,51,0,39,0,38,0,183,0,0,0,230,0,7,0,3,0,101,0,170,0,114,0,66,0,3,0,155,0,104,0,148,0,253,0,111,0,0,0,121,0,0,0,54,0,0,0,149,0,0,0,0,0,83,0,0,0,103,0,0,0);
signal scenario_full  : scenario_type := (104,31,48,31,124,31,174,31,182,31,138,31,150,31,150,30,150,29,150,28,150,27,150,26,24,31,143,31,122,31,226,31,204,31,168,31,153,31,145,31,82,31,65,31,65,30,172,31,116,31,116,30,75,31,158,31,158,30,19,31,19,30,229,31,245,31,145,31,121,31,61,31,17,31,241,31,111,31,176,31,168,31,20,31,182,31,182,30,25,31,25,30,25,29,25,28,230,31,204,31,99,31,33,31,183,31,182,31,152,31,77,31,31,31,148,31,75,31,244,31,237,31,234,31,7,31,48,31,103,31,53,31,53,30,230,31,95,31,109,31,109,30,187,31,194,31,11,31,203,31,11,31,95,31,122,31,122,30,166,31,204,31,217,31,172,31,98,31,241,31,82,31,19,31,16,31,16,30,16,29,96,31,96,30,169,31,109,31,109,30,134,31,70,31,196,31,206,31,30,31,232,31,104,31,223,31,201,31,233,31,252,31,220,31,155,31,111,31,25,31,24,31,24,30,24,29,85,31,85,30,85,29,191,31,144,31,144,30,135,31,135,30,140,31,200,31,52,31,244,31,103,31,171,31,218,31,55,31,135,31,28,31,183,31,101,31,19,31,131,31,113,31,219,31,23,31,23,30,129,31,66,31,158,31,20,31,205,31,42,31,190,31,190,30,119,31,142,31,48,31,36,31,71,31,71,30,110,31,153,31,153,30,176,31,172,31,153,31,13,31,13,30,190,31,39,31,137,31,137,30,164,31,244,31,244,30,224,31,124,31,96,31,199,31,199,30,231,31,211,31,165,31,165,30,165,29,123,31,123,30,100,31,100,30,198,31,222,31,130,31,233,31,27,31,189,31,68,31,179,31,112,31,112,30,232,31,130,31,252,31,159,31,5,31,9,31,66,31,181,31,95,31,185,31,36,31,243,31,19,31,244,31,221,31,5,31,244,31,112,31,112,30,108,31,125,31,251,31,187,31,128,31,107,31,8,31,8,30,73,31,82,31,18,31,6,31,248,31,83,31,238,31,24,31,178,31,207,31,13,31,50,31,180,31,180,30,180,29,1,31,1,30,143,31,89,31,46,31,155,31,237,31,103,31,19,31,19,30,168,31,168,30,226,31,117,31,113,31,27,31,204,31,230,31,238,31,238,30,238,29,238,28,174,31,141,31,129,31,213,31,213,30,226,31,225,31,225,30,141,31,175,31,175,30,36,31,36,30,36,29,167,31,213,31,116,31,162,31,8,31,68,31,68,30,239,31,11,31,11,30,159,31,116,31,238,31,174,31,37,31,239,31,253,31,14,31,72,31,220,31,185,31,227,31,12,31,102,31,91,31,150,31,150,30,157,31,201,31,95,31,185,31,219,31,219,30,219,29,107,31,73,31,21,31,70,31,183,31,51,31,180,31,180,30,120,31,241,31,143,31,185,31,198,31,50,31,159,31,170,31,94,31,94,30,76,31,76,30,67,31,67,30,187,31,243,31,114,31,51,31,160,31,143,31,94,31,42,31,42,30,9,31,91,31,75,31,75,30,23,31,162,31,248,31,206,31,206,30,206,29,55,31,182,31,64,31,107,31,107,30,113,31,113,30,103,31,140,31,205,31,218,31,218,30,203,31,119,31,9,31,213,31,213,30,204,31,116,31,55,31,117,31,40,31,186,31,17,31,222,31,222,30,214,31,239,31,239,30,237,31,237,30,16,31,16,30,16,29,16,28,24,31,111,31,131,31,40,31,166,31,166,30,158,31,138,31,176,31,176,30,17,31,231,31,232,31,224,31,62,31,8,31,9,31,168,31,222,31,143,31,10,31,237,31,237,30,238,31,238,30,116,31,113,31,113,30,178,31,178,30,136,31,136,30,30,31,103,31,197,31,197,30,27,31,50,31,191,31,209,31,142,31,142,30,26,31,6,31,103,31,122,31,19,31,94,31,6,31,6,30,148,31,148,30,148,29,188,31,10,31,10,30,129,31,255,31,2,31,32,31,223,31,223,30,244,31,63,31,149,31,96,31,251,31,83,31,185,31,156,31,177,31,231,31,12,31,12,30,29,31,37,31,67,31,160,31,160,30,160,29,160,28,249,31,106,31,213,31,213,30,121,31,106,31,105,31,74,31,9,31,133,31,42,31,99,31,4,31,31,31,130,31,150,31,150,30,150,29,184,31,198,31,211,31,33,31,33,30,33,29,16,31,242,31,11,31,202,31,59,31,196,31,76,31,148,31,81,31,81,30,239,31,190,31,186,31,186,30,228,31,211,31,253,31,153,31,195,31,5,31,9,31,111,31,26,31,175,31,160,31,117,31,121,31,198,31,196,31,16,31,151,31,196,31,196,30,32,31,8,31,168,31,77,31,37,31,247,31,52,31,162,31,162,30,162,29,236,31,21,31,63,31,103,31,162,31,75,31,75,30,45,31,77,31,175,31,110,31,68,31,240,31,206,31,254,31,188,31,139,31,219,31,80,31,80,30,79,31,189,31,108,31,111,31,136,31,89,31,146,31,221,31,145,31,145,30,145,29,155,31,237,31,218,31,173,31,68,31,241,31,8,31,112,31,47,31,172,31,16,31,219,31,115,31,69,31,60,31,60,30,13,31,48,31,48,30,106,31,86,31,7,31,161,31,75,31,243,31,235,31,11,31,11,30,18,31,14,31,14,30,45,31,45,30,45,29,245,31,245,30,178,31,173,31,34,31,243,31,127,31,51,31,125,31,115,31,42,31,42,30,109,31,148,31,156,31,124,31,109,31,1,31,93,31,186,31,66,31,132,31,248,31,171,31,4,31,4,30,4,29,72,31,72,30,193,31,162,31,167,31,140,31,166,31,212,31,20,31,78,31,32,31,61,31,211,31,50,31,64,31,249,31,26,31,33,31,65,31,65,30,97,31,72,31,6,31,216,31,209,31,8,31,186,31,186,30,206,31,71,31,94,31,219,31,219,30,219,29,219,28,137,31,22,31,141,31,185,31,241,31,92,31,53,31,117,31,117,30,64,31,64,30,64,29,27,31,9,31,9,30,6,31,2,31,125,31,170,31,90,31,90,30,216,31,244,31,51,31,39,31,38,31,183,31,183,30,230,31,7,31,3,31,101,31,170,31,114,31,66,31,3,31,155,31,104,31,148,31,253,31,111,31,111,30,121,31,121,30,54,31,54,30,149,31,149,30,149,29,83,31,83,30,103,31,103,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
