-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 715;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (199,0,206,0,87,0,49,0,240,0,174,0,40,0,11,0,0,0,173,0,38,0,0,0,198,0,240,0,10,0,190,0,14,0,120,0,17,0,64,0,163,0,133,0,218,0,169,0,165,0,103,0,223,0,97,0,4,0,83,0,0,0,196,0,64,0,81,0,65,0,0,0,159,0,0,0,144,0,10,0,103,0,59,0,126,0,247,0,0,0,43,0,127,0,124,0,192,0,0,0,84,0,245,0,32,0,199,0,102,0,0,0,255,0,67,0,71,0,213,0,218,0,0,0,244,0,10,0,176,0,235,0,109,0,106,0,0,0,197,0,38,0,198,0,115,0,33,0,95,0,172,0,210,0,0,0,204,0,144,0,186,0,0,0,24,0,18,0,0,0,163,0,203,0,94,0,238,0,110,0,207,0,161,0,134,0,149,0,184,0,0,0,167,0,181,0,22,0,58,0,183,0,0,0,153,0,0,0,138,0,188,0,0,0,83,0,0,0,226,0,253,0,0,0,84,0,190,0,102,0,0,0,218,0,96,0,48,0,150,0,151,0,44,0,114,0,101,0,181,0,199,0,33,0,132,0,88,0,211,0,160,0,0,0,251,0,246,0,0,0,116,0,0,0,112,0,96,0,0,0,0,0,36,0,0,0,4,0,14,0,187,0,230,0,89,0,214,0,77,0,128,0,198,0,21,0,133,0,120,0,33,0,77,0,60,0,242,0,213,0,23,0,0,0,99,0,0,0,0,0,217,0,35,0,221,0,152,0,14,0,136,0,213,0,65,0,96,0,0,0,43,0,59,0,176,0,167,0,85,0,10,0,136,0,217,0,182,0,0,0,106,0,134,0,243,0,0,0,89,0,113,0,237,0,140,0,14,0,94,0,166,0,218,0,132,0,138,0,0,0,149,0,27,0,151,0,0,0,144,0,56,0,83,0,18,0,15,0,207,0,232,0,23,0,198,0,107,0,55,0,35,0,230,0,171,0,168,0,243,0,59,0,215,0,137,0,211,0,253,0,44,0,193,0,62,0,61,0,141,0,250,0,253,0,89,0,66,0,133,0,226,0,0,0,61,0,0,0,72,0,18,0,117,0,154,0,0,0,0,0,13,0,0,0,0,0,52,0,8,0,215,0,248,0,6,0,16,0,183,0,126,0,197,0,206,0,182,0,2,0,8,0,95,0,104,0,161,0,189,0,119,0,232,0,68,0,0,0,241,0,192,0,69,0,129,0,110,0,0,0,191,0,186,0,85,0,234,0,0,0,156,0,55,0,145,0,183,0,19,0,186,0,140,0,77,0,58,0,199,0,98,0,179,0,234,0,23,0,41,0,23,0,219,0,0,0,166,0,0,0,150,0,0,0,177,0,149,0,19,0,199,0,177,0,194,0,0,0,230,0,49,0,56,0,86,0,49,0,212,0,223,0,213,0,43,0,229,0,0,0,68,0,211,0,0,0,148,0,153,0,166,0,126,0,70,0,153,0,150,0,0,0,0,0,127,0,185,0,209,0,161,0,55,0,200,0,100,0,223,0,0,0,232,0,72,0,161,0,103,0,244,0,163,0,214,0,69,0,0,0,222,0,23,0,168,0,239,0,57,0,108,0,38,0,97,0,0,0,193,0,15,0,0,0,114,0,58,0,59,0,76,0,106,0,214,0,144,0,0,0,59,0,214,0,95,0,43,0,228,0,196,0,58,0,8,0,100,0,220,0,233,0,186,0,202,0,0,0,28,0,218,0,161,0,0,0,88,0,93,0,56,0,0,0,12,0,224,0,0,0,0,0,15,0,250,0,176,0,17,0,0,0,247,0,202,0,224,0,0,0,46,0,176,0,119,0,0,0,137,0,118,0,0,0,52,0,193,0,149,0,0,0,189,0,170,0,0,0,171,0,114,0,0,0,0,0,83,0,0,0,193,0,16,0,0,0,0,0,0,0,189,0,86,0,0,0,29,0,182,0,90,0,0,0,141,0,117,0,58,0,171,0,0,0,66,0,95,0,169,0,226,0,0,0,116,0,13,0,216,0,47,0,230,0,76,0,217,0,37,0,218,0,255,0,252,0,221,0,110,0,64,0,0,0,151,0,0,0,179,0,82,0,111,0,57,0,0,0,25,0,138,0,211,0,138,0,44,0,229,0,110,0,134,0,0,0,0,0,227,0,222,0,235,0,0,0,86,0,206,0,35,0,216,0,11,0,110,0,161,0,104,0,160,0,150,0,0,0,95,0,113,0,0,0,183,0,122,0,97,0,122,0,185,0,39,0,105,0,6,0,0,0,93,0,190,0,75,0,226,0,0,0,154,0,36,0,0,0,170,0,88,0,0,0,229,0,13,0,190,0,202,0,229,0,55,0,0,0,181,0,0,0,222,0,0,0,165,0,222,0,231,0,0,0,164,0,242,0,124,0,222,0,42,0,68,0,229,0,0,0,206,0,0,0,182,0,216,0,100,0,44,0,203,0,50,0,203,0,111,0,207,0,229,0,106,0,12,0,80,0,143,0,0,0,174,0,98,0,135,0,0,0,224,0,125,0,81,0,182,0,162,0,0,0,77,0,211,0,207,0,104,0,67,0,6,0,66,0,150,0,119,0,0,0,48,0,114,0,147,0,0,0,195,0,172,0,12,0,148,0,59,0,69,0,118,0,77,0,0,0,113,0,113,0,150,0,0,0,209,0,235,0,98,0,63,0,0,0,146,0,255,0,0,0,80,0,225,0,134,0,0,0,178,0,152,0,0,0,0,0,134,0,216,0,0,0,25,0,200,0,171,0,0,0,243,0,45,0,119,0,249,0,167,0,212,0,174,0,118,0,227,0,245,0,54,0,82,0,80,0,172,0,0,0,196,0,86,0,100,0,161,0,152,0,222,0,105,0,69,0,248,0,176,0,0,0,111,0,39,0,210,0,55,0,155,0,0,0,210,0,154,0,175,0,249,0,57,0,112,0,94,0,61,0,210,0,2,0,243,0,25,0,60,0,0,0,72,0,183,0,193,0,41,0,97,0,97,0,0,0,242,0,58,0,0,0,67,0,5,0,85,0,47,0,230,0,99,0,0,0,155,0,146,0,137,0,0,0,209,0,213,0,46,0,78,0,178,0,250,0,75,0,220,0,112,0,244,0,125,0,0,0,192,0,19,0,221,0,6,0,157,0,79,0,0,0,0,0,127,0,149,0,7,0,202,0,134,0,116,0,157,0,251,0,160,0,27,0,99,0);
signal scenario_full  : scenario_type := (199,31,206,31,87,31,49,31,240,31,174,31,40,31,11,31,11,30,173,31,38,31,38,30,198,31,240,31,10,31,190,31,14,31,120,31,17,31,64,31,163,31,133,31,218,31,169,31,165,31,103,31,223,31,97,31,4,31,83,31,83,30,196,31,64,31,81,31,65,31,65,30,159,31,159,30,144,31,10,31,103,31,59,31,126,31,247,31,247,30,43,31,127,31,124,31,192,31,192,30,84,31,245,31,32,31,199,31,102,31,102,30,255,31,67,31,71,31,213,31,218,31,218,30,244,31,10,31,176,31,235,31,109,31,106,31,106,30,197,31,38,31,198,31,115,31,33,31,95,31,172,31,210,31,210,30,204,31,144,31,186,31,186,30,24,31,18,31,18,30,163,31,203,31,94,31,238,31,110,31,207,31,161,31,134,31,149,31,184,31,184,30,167,31,181,31,22,31,58,31,183,31,183,30,153,31,153,30,138,31,188,31,188,30,83,31,83,30,226,31,253,31,253,30,84,31,190,31,102,31,102,30,218,31,96,31,48,31,150,31,151,31,44,31,114,31,101,31,181,31,199,31,33,31,132,31,88,31,211,31,160,31,160,30,251,31,246,31,246,30,116,31,116,30,112,31,96,31,96,30,96,29,36,31,36,30,4,31,14,31,187,31,230,31,89,31,214,31,77,31,128,31,198,31,21,31,133,31,120,31,33,31,77,31,60,31,242,31,213,31,23,31,23,30,99,31,99,30,99,29,217,31,35,31,221,31,152,31,14,31,136,31,213,31,65,31,96,31,96,30,43,31,59,31,176,31,167,31,85,31,10,31,136,31,217,31,182,31,182,30,106,31,134,31,243,31,243,30,89,31,113,31,237,31,140,31,14,31,94,31,166,31,218,31,132,31,138,31,138,30,149,31,27,31,151,31,151,30,144,31,56,31,83,31,18,31,15,31,207,31,232,31,23,31,198,31,107,31,55,31,35,31,230,31,171,31,168,31,243,31,59,31,215,31,137,31,211,31,253,31,44,31,193,31,62,31,61,31,141,31,250,31,253,31,89,31,66,31,133,31,226,31,226,30,61,31,61,30,72,31,18,31,117,31,154,31,154,30,154,29,13,31,13,30,13,29,52,31,8,31,215,31,248,31,6,31,16,31,183,31,126,31,197,31,206,31,182,31,2,31,8,31,95,31,104,31,161,31,189,31,119,31,232,31,68,31,68,30,241,31,192,31,69,31,129,31,110,31,110,30,191,31,186,31,85,31,234,31,234,30,156,31,55,31,145,31,183,31,19,31,186,31,140,31,77,31,58,31,199,31,98,31,179,31,234,31,23,31,41,31,23,31,219,31,219,30,166,31,166,30,150,31,150,30,177,31,149,31,19,31,199,31,177,31,194,31,194,30,230,31,49,31,56,31,86,31,49,31,212,31,223,31,213,31,43,31,229,31,229,30,68,31,211,31,211,30,148,31,153,31,166,31,126,31,70,31,153,31,150,31,150,30,150,29,127,31,185,31,209,31,161,31,55,31,200,31,100,31,223,31,223,30,232,31,72,31,161,31,103,31,244,31,163,31,214,31,69,31,69,30,222,31,23,31,168,31,239,31,57,31,108,31,38,31,97,31,97,30,193,31,15,31,15,30,114,31,58,31,59,31,76,31,106,31,214,31,144,31,144,30,59,31,214,31,95,31,43,31,228,31,196,31,58,31,8,31,100,31,220,31,233,31,186,31,202,31,202,30,28,31,218,31,161,31,161,30,88,31,93,31,56,31,56,30,12,31,224,31,224,30,224,29,15,31,250,31,176,31,17,31,17,30,247,31,202,31,224,31,224,30,46,31,176,31,119,31,119,30,137,31,118,31,118,30,52,31,193,31,149,31,149,30,189,31,170,31,170,30,171,31,114,31,114,30,114,29,83,31,83,30,193,31,16,31,16,30,16,29,16,28,189,31,86,31,86,30,29,31,182,31,90,31,90,30,141,31,117,31,58,31,171,31,171,30,66,31,95,31,169,31,226,31,226,30,116,31,13,31,216,31,47,31,230,31,76,31,217,31,37,31,218,31,255,31,252,31,221,31,110,31,64,31,64,30,151,31,151,30,179,31,82,31,111,31,57,31,57,30,25,31,138,31,211,31,138,31,44,31,229,31,110,31,134,31,134,30,134,29,227,31,222,31,235,31,235,30,86,31,206,31,35,31,216,31,11,31,110,31,161,31,104,31,160,31,150,31,150,30,95,31,113,31,113,30,183,31,122,31,97,31,122,31,185,31,39,31,105,31,6,31,6,30,93,31,190,31,75,31,226,31,226,30,154,31,36,31,36,30,170,31,88,31,88,30,229,31,13,31,190,31,202,31,229,31,55,31,55,30,181,31,181,30,222,31,222,30,165,31,222,31,231,31,231,30,164,31,242,31,124,31,222,31,42,31,68,31,229,31,229,30,206,31,206,30,182,31,216,31,100,31,44,31,203,31,50,31,203,31,111,31,207,31,229,31,106,31,12,31,80,31,143,31,143,30,174,31,98,31,135,31,135,30,224,31,125,31,81,31,182,31,162,31,162,30,77,31,211,31,207,31,104,31,67,31,6,31,66,31,150,31,119,31,119,30,48,31,114,31,147,31,147,30,195,31,172,31,12,31,148,31,59,31,69,31,118,31,77,31,77,30,113,31,113,31,150,31,150,30,209,31,235,31,98,31,63,31,63,30,146,31,255,31,255,30,80,31,225,31,134,31,134,30,178,31,152,31,152,30,152,29,134,31,216,31,216,30,25,31,200,31,171,31,171,30,243,31,45,31,119,31,249,31,167,31,212,31,174,31,118,31,227,31,245,31,54,31,82,31,80,31,172,31,172,30,196,31,86,31,100,31,161,31,152,31,222,31,105,31,69,31,248,31,176,31,176,30,111,31,39,31,210,31,55,31,155,31,155,30,210,31,154,31,175,31,249,31,57,31,112,31,94,31,61,31,210,31,2,31,243,31,25,31,60,31,60,30,72,31,183,31,193,31,41,31,97,31,97,31,97,30,242,31,58,31,58,30,67,31,5,31,85,31,47,31,230,31,99,31,99,30,155,31,146,31,137,31,137,30,209,31,213,31,46,31,78,31,178,31,250,31,75,31,220,31,112,31,244,31,125,31,125,30,192,31,19,31,221,31,6,31,157,31,79,31,79,30,79,29,127,31,149,31,7,31,202,31,134,31,116,31,157,31,251,31,160,31,27,31,99,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
