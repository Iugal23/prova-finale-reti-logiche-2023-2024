-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 906;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (112,0,0,0,145,0,154,0,79,0,73,0,0,0,238,0,63,0,51,0,93,0,193,0,4,0,1,0,119,0,223,0,0,0,45,0,196,0,19,0,122,0,83,0,0,0,194,0,22,0,184,0,0,0,245,0,219,0,62,0,204,0,139,0,240,0,0,0,6,0,89,0,101,0,250,0,18,0,144,0,182,0,226,0,0,0,53,0,69,0,200,0,106,0,34,0,121,0,117,0,0,0,254,0,63,0,217,0,0,0,0,0,0,0,243,0,237,0,0,0,15,0,125,0,204,0,66,0,123,0,134,0,132,0,154,0,75,0,0,0,166,0,252,0,171,0,0,0,0,0,204,0,19,0,17,0,215,0,69,0,9,0,115,0,0,0,245,0,0,0,0,0,187,0,156,0,24,0,229,0,126,0,221,0,0,0,84,0,131,0,0,0,28,0,215,0,0,0,56,0,4,0,20,0,83,0,145,0,73,0,168,0,246,0,43,0,48,0,103,0,0,0,0,0,230,0,214,0,215,0,0,0,0,0,0,0,146,0,33,0,108,0,154,0,0,0,242,0,86,0,108,0,206,0,53,0,0,0,69,0,0,0,87,0,0,0,237,0,212,0,97,0,217,0,0,0,195,0,0,0,0,0,0,0,172,0,0,0,114,0,153,0,78,0,18,0,0,0,76,0,0,0,91,0,119,0,52,0,241,0,244,0,0,0,180,0,109,0,190,0,97,0,86,0,9,0,0,0,229,0,209,0,30,0,0,0,0,0,195,0,191,0,82,0,0,0,0,0,202,0,14,0,205,0,107,0,140,0,235,0,50,0,185,0,49,0,68,0,0,0,0,0,31,0,202,0,0,0,81,0,174,0,0,0,123,0,0,0,154,0,99,0,10,0,29,0,219,0,173,0,175,0,192,0,164,0,199,0,0,0,56,0,81,0,0,0,91,0,127,0,0,0,252,0,215,0,244,0,92,0,121,0,240,0,111,0,203,0,109,0,95,0,0,0,112,0,139,0,132,0,10,0,24,0,203,0,187,0,102,0,0,0,165,0,0,0,215,0,82,0,173,0,118,0,0,0,51,0,31,0,159,0,34,0,0,0,178,0,168,0,0,0,22,0,36,0,182,0,103,0,0,0,60,0,0,0,0,0,0,0,107,0,179,0,231,0,240,0,119,0,212,0,130,0,0,0,203,0,0,0,87,0,25,0,158,0,157,0,3,0,0,0,13,0,225,0,0,0,0,0,0,0,84,0,7,0,0,0,0,0,14,0,0,0,8,0,94,0,250,0,11,0,227,0,179,0,21,0,174,0,245,0,60,0,130,0,109,0,20,0,155,0,79,0,82,0,0,0,146,0,55,0,0,0,255,0,185,0,23,0,218,0,131,0,7,0,91,0,24,0,138,0,155,0,0,0,129,0,232,0,0,0,41,0,207,0,233,0,246,0,10,0,0,0,29,0,231,0,222,0,8,0,15,0,3,0,0,0,145,0,107,0,56,0,0,0,49,0,217,0,0,0,214,0,147,0,0,0,119,0,13,0,63,0,59,0,0,0,179,0,0,0,0,0,148,0,0,0,83,0,0,0,110,0,55,0,0,0,122,0,0,0,0,0,161,0,192,0,157,0,0,0,249,0,0,0,195,0,81,0,194,0,169,0,55,0,182,0,123,0,88,0,176,0,182,0,0,0,69,0,101,0,204,0,94,0,103,0,77,0,0,0,42,0,5,0,3,0,67,0,43,0,238,0,0,0,112,0,158,0,240,0,168,0,4,0,110,0,254,0,0,0,173,0,86,0,245,0,2,0,57,0,79,0,181,0,1,0,107,0,137,0,90,0,0,0,228,0,191,0,136,0,0,0,62,0,145,0,0,0,0,0,186,0,188,0,0,0,214,0,58,0,128,0,28,0,108,0,133,0,133,0,3,0,51,0,171,0,103,0,209,0,63,0,0,0,0,0,61,0,48,0,168,0,0,0,0,0,139,0,220,0,78,0,0,0,4,0,99,0,70,0,242,0,25,0,58,0,20,0,0,0,129,0,227,0,25,0,0,0,215,0,51,0,140,0,0,0,203,0,203,0,0,0,0,0,245,0,172,0,0,0,0,0,67,0,122,0,35,0,149,0,0,0,91,0,167,0,41,0,58,0,0,0,0,0,90,0,6,0,22,0,144,0,225,0,47,0,255,0,231,0,0,0,0,0,0,0,250,0,144,0,10,0,86,0,73,0,146,0,96,0,157,0,119,0,238,0,0,0,92,0,0,0,0,0,61,0,74,0,53,0,0,0,7,0,152,0,223,0,162,0,102,0,72,0,73,0,140,0,0,0,0,0,24,0,83,0,4,0,64,0,19,0,16,0,0,0,105,0,206,0,140,0,83,0,0,0,248,0,171,0,149,0,101,0,244,0,66,0,64,0,70,0,175,0,33,0,0,0,225,0,126,0,203,0,148,0,187,0,90,0,242,0,25,0,33,0,0,0,0,0,0,0,0,0,211,0,101,0,45,0,160,0,11,0,16,0,201,0,0,0,0,0,13,0,119,0,202,0,179,0,243,0,0,0,19,0,121,0,116,0,154,0,48,0,228,0,164,0,0,0,9,0,0,0,67,0,111,0,0,0,0,0,77,0,192,0,181,0,226,0,75,0,126,0,17,0,178,0,130,0,0,0,0,0,0,0,44,0,220,0,101,0,0,0,138,0,214,0,242,0,0,0,100,0,7,0,240,0,168,0,15,0,149,0,101,0,40,0,241,0,0,0,108,0,200,0,14,0,118,0,8,0,15,0,246,0,178,0,20,0,150,0,213,0,0,0,95,0,222,0,68,0,190,0,0,0,0,0,233,0,96,0,234,0,133,0,0,0,205,0,207,0,28,0,32,0,238,0,165,0,237,0,56,0,187,0,249,0,0,0,12,0,195,0,125,0,0,0,0,0,254,0,0,0,41,0,0,0,0,0,0,0,0,0,163,0,174,0,183,0,0,0,0,0,0,0,130,0,8,0,62,0,0,0,146,0,89,0,127,0,0,0,41,0,166,0,178,0,144,0,0,0,178,0,254,0,4,0,0,0,0,0,0,0,0,0,159,0,63,0,225,0,124,0,224,0,77,0,120,0,52,0,0,0,152,0,214,0,97,0,242,0,216,0,197,0,41,0,182,0,180,0,137,0,133,0,182,0,56,0,187,0,0,0,0,0,72,0,121,0,126,0,105,0,0,0,0,0,0,0,33,0,185,0,56,0,128,0,172,0,22,0,221,0,0,0,188,0,216,0,10,0,185,0,197,0,180,0,132,0,86,0,0,0,5,0,0,0,121,0,59,0,211,0,210,0,170,0,120,0,44,0,87,0,113,0,98,0,166,0,56,0,249,0,0,0,131,0,54,0,0,0,117,0,67,0,222,0,0,0,103,0,177,0,0,0,130,0,53,0,0,0,68,0,26,0,155,0,168,0,0,0,0,0,0,0,72,0,209,0,135,0,170,0,247,0,0,0,83,0,239,0,42,0,39,0,222,0,153,0,135,0,19,0,8,0,236,0,115,0,22,0,44,0,68,0,51,0,165,0,118,0,59,0,107,0,120,0,0,0,0,0,93,0,168,0,0,0,0,0,145,0,134,0,182,0,223,0,4,0,182,0,94,0,214,0,199,0,197,0,0,0,81,0,0,0,221,0,228,0,255,0,0,0,39,0,171,0,71,0,187,0,19,0,84,0,250,0,0,0,20,0,0,0,240,0,210,0,0,0,0,0,0,0,193,0,116,0,0,0,33,0,0,0,0,0,0,0,226,0,102,0,201,0,162,0,142,0,34,0,125,0,0,0,46,0,0,0,11,0,33,0,121,0,39,0,0,0,254,0,0,0,247,0,185,0,176,0,0,0,188,0,0,0,125,0,68,0,0,0,102,0,142,0,181,0,112,0,202,0,24,0,225,0,43,0,188,0,249,0,158,0,63,0,133,0,18,0,0,0,65,0,0,0,245,0,183,0,156,0,100,0,211,0,153,0,247,0,0,0,217,0,49,0,196,0,0,0,0,0,243,0,226,0,27,0,0,0,2,0,116,0,78,0,0,0,24,0,74,0);
signal scenario_full  : scenario_type := (112,31,112,30,145,31,154,31,79,31,73,31,73,30,238,31,63,31,51,31,93,31,193,31,4,31,1,31,119,31,223,31,223,30,45,31,196,31,19,31,122,31,83,31,83,30,194,31,22,31,184,31,184,30,245,31,219,31,62,31,204,31,139,31,240,31,240,30,6,31,89,31,101,31,250,31,18,31,144,31,182,31,226,31,226,30,53,31,69,31,200,31,106,31,34,31,121,31,117,31,117,30,254,31,63,31,217,31,217,30,217,29,217,28,243,31,237,31,237,30,15,31,125,31,204,31,66,31,123,31,134,31,132,31,154,31,75,31,75,30,166,31,252,31,171,31,171,30,171,29,204,31,19,31,17,31,215,31,69,31,9,31,115,31,115,30,245,31,245,30,245,29,187,31,156,31,24,31,229,31,126,31,221,31,221,30,84,31,131,31,131,30,28,31,215,31,215,30,56,31,4,31,20,31,83,31,145,31,73,31,168,31,246,31,43,31,48,31,103,31,103,30,103,29,230,31,214,31,215,31,215,30,215,29,215,28,146,31,33,31,108,31,154,31,154,30,242,31,86,31,108,31,206,31,53,31,53,30,69,31,69,30,87,31,87,30,237,31,212,31,97,31,217,31,217,30,195,31,195,30,195,29,195,28,172,31,172,30,114,31,153,31,78,31,18,31,18,30,76,31,76,30,91,31,119,31,52,31,241,31,244,31,244,30,180,31,109,31,190,31,97,31,86,31,9,31,9,30,229,31,209,31,30,31,30,30,30,29,195,31,191,31,82,31,82,30,82,29,202,31,14,31,205,31,107,31,140,31,235,31,50,31,185,31,49,31,68,31,68,30,68,29,31,31,202,31,202,30,81,31,174,31,174,30,123,31,123,30,154,31,99,31,10,31,29,31,219,31,173,31,175,31,192,31,164,31,199,31,199,30,56,31,81,31,81,30,91,31,127,31,127,30,252,31,215,31,244,31,92,31,121,31,240,31,111,31,203,31,109,31,95,31,95,30,112,31,139,31,132,31,10,31,24,31,203,31,187,31,102,31,102,30,165,31,165,30,215,31,82,31,173,31,118,31,118,30,51,31,31,31,159,31,34,31,34,30,178,31,168,31,168,30,22,31,36,31,182,31,103,31,103,30,60,31,60,30,60,29,60,28,107,31,179,31,231,31,240,31,119,31,212,31,130,31,130,30,203,31,203,30,87,31,25,31,158,31,157,31,3,31,3,30,13,31,225,31,225,30,225,29,225,28,84,31,7,31,7,30,7,29,14,31,14,30,8,31,94,31,250,31,11,31,227,31,179,31,21,31,174,31,245,31,60,31,130,31,109,31,20,31,155,31,79,31,82,31,82,30,146,31,55,31,55,30,255,31,185,31,23,31,218,31,131,31,7,31,91,31,24,31,138,31,155,31,155,30,129,31,232,31,232,30,41,31,207,31,233,31,246,31,10,31,10,30,29,31,231,31,222,31,8,31,15,31,3,31,3,30,145,31,107,31,56,31,56,30,49,31,217,31,217,30,214,31,147,31,147,30,119,31,13,31,63,31,59,31,59,30,179,31,179,30,179,29,148,31,148,30,83,31,83,30,110,31,55,31,55,30,122,31,122,30,122,29,161,31,192,31,157,31,157,30,249,31,249,30,195,31,81,31,194,31,169,31,55,31,182,31,123,31,88,31,176,31,182,31,182,30,69,31,101,31,204,31,94,31,103,31,77,31,77,30,42,31,5,31,3,31,67,31,43,31,238,31,238,30,112,31,158,31,240,31,168,31,4,31,110,31,254,31,254,30,173,31,86,31,245,31,2,31,57,31,79,31,181,31,1,31,107,31,137,31,90,31,90,30,228,31,191,31,136,31,136,30,62,31,145,31,145,30,145,29,186,31,188,31,188,30,214,31,58,31,128,31,28,31,108,31,133,31,133,31,3,31,51,31,171,31,103,31,209,31,63,31,63,30,63,29,61,31,48,31,168,31,168,30,168,29,139,31,220,31,78,31,78,30,4,31,99,31,70,31,242,31,25,31,58,31,20,31,20,30,129,31,227,31,25,31,25,30,215,31,51,31,140,31,140,30,203,31,203,31,203,30,203,29,245,31,172,31,172,30,172,29,67,31,122,31,35,31,149,31,149,30,91,31,167,31,41,31,58,31,58,30,58,29,90,31,6,31,22,31,144,31,225,31,47,31,255,31,231,31,231,30,231,29,231,28,250,31,144,31,10,31,86,31,73,31,146,31,96,31,157,31,119,31,238,31,238,30,92,31,92,30,92,29,61,31,74,31,53,31,53,30,7,31,152,31,223,31,162,31,102,31,72,31,73,31,140,31,140,30,140,29,24,31,83,31,4,31,64,31,19,31,16,31,16,30,105,31,206,31,140,31,83,31,83,30,248,31,171,31,149,31,101,31,244,31,66,31,64,31,70,31,175,31,33,31,33,30,225,31,126,31,203,31,148,31,187,31,90,31,242,31,25,31,33,31,33,30,33,29,33,28,33,27,211,31,101,31,45,31,160,31,11,31,16,31,201,31,201,30,201,29,13,31,119,31,202,31,179,31,243,31,243,30,19,31,121,31,116,31,154,31,48,31,228,31,164,31,164,30,9,31,9,30,67,31,111,31,111,30,111,29,77,31,192,31,181,31,226,31,75,31,126,31,17,31,178,31,130,31,130,30,130,29,130,28,44,31,220,31,101,31,101,30,138,31,214,31,242,31,242,30,100,31,7,31,240,31,168,31,15,31,149,31,101,31,40,31,241,31,241,30,108,31,200,31,14,31,118,31,8,31,15,31,246,31,178,31,20,31,150,31,213,31,213,30,95,31,222,31,68,31,190,31,190,30,190,29,233,31,96,31,234,31,133,31,133,30,205,31,207,31,28,31,32,31,238,31,165,31,237,31,56,31,187,31,249,31,249,30,12,31,195,31,125,31,125,30,125,29,254,31,254,30,41,31,41,30,41,29,41,28,41,27,163,31,174,31,183,31,183,30,183,29,183,28,130,31,8,31,62,31,62,30,146,31,89,31,127,31,127,30,41,31,166,31,178,31,144,31,144,30,178,31,254,31,4,31,4,30,4,29,4,28,4,27,159,31,63,31,225,31,124,31,224,31,77,31,120,31,52,31,52,30,152,31,214,31,97,31,242,31,216,31,197,31,41,31,182,31,180,31,137,31,133,31,182,31,56,31,187,31,187,30,187,29,72,31,121,31,126,31,105,31,105,30,105,29,105,28,33,31,185,31,56,31,128,31,172,31,22,31,221,31,221,30,188,31,216,31,10,31,185,31,197,31,180,31,132,31,86,31,86,30,5,31,5,30,121,31,59,31,211,31,210,31,170,31,120,31,44,31,87,31,113,31,98,31,166,31,56,31,249,31,249,30,131,31,54,31,54,30,117,31,67,31,222,31,222,30,103,31,177,31,177,30,130,31,53,31,53,30,68,31,26,31,155,31,168,31,168,30,168,29,168,28,72,31,209,31,135,31,170,31,247,31,247,30,83,31,239,31,42,31,39,31,222,31,153,31,135,31,19,31,8,31,236,31,115,31,22,31,44,31,68,31,51,31,165,31,118,31,59,31,107,31,120,31,120,30,120,29,93,31,168,31,168,30,168,29,145,31,134,31,182,31,223,31,4,31,182,31,94,31,214,31,199,31,197,31,197,30,81,31,81,30,221,31,228,31,255,31,255,30,39,31,171,31,71,31,187,31,19,31,84,31,250,31,250,30,20,31,20,30,240,31,210,31,210,30,210,29,210,28,193,31,116,31,116,30,33,31,33,30,33,29,33,28,226,31,102,31,201,31,162,31,142,31,34,31,125,31,125,30,46,31,46,30,11,31,33,31,121,31,39,31,39,30,254,31,254,30,247,31,185,31,176,31,176,30,188,31,188,30,125,31,68,31,68,30,102,31,142,31,181,31,112,31,202,31,24,31,225,31,43,31,188,31,249,31,158,31,63,31,133,31,18,31,18,30,65,31,65,30,245,31,183,31,156,31,100,31,211,31,153,31,247,31,247,30,217,31,49,31,196,31,196,30,196,29,243,31,226,31,27,31,27,30,2,31,116,31,78,31,78,30,24,31,74,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
