-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 877;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (193,0,0,0,137,0,111,0,34,0,0,0,239,0,216,0,0,0,185,0,183,0,228,0,197,0,119,0,45,0,0,0,67,0,0,0,0,0,12,0,0,0,75,0,0,0,235,0,0,0,175,0,0,0,28,0,23,0,0,0,0,0,214,0,184,0,0,0,111,0,0,0,222,0,102,0,39,0,0,0,61,0,100,0,118,0,73,0,204,0,0,0,0,0,75,0,218,0,185,0,109,0,81,0,226,0,0,0,0,0,134,0,30,0,247,0,18,0,0,0,60,0,229,0,114,0,195,0,0,0,23,0,24,0,167,0,67,0,189,0,0,0,182,0,3,0,0,0,119,0,0,0,0,0,190,0,207,0,125,0,202,0,0,0,80,0,99,0,40,0,108,0,59,0,52,0,25,0,164,0,100,0,0,0,251,0,37,0,63,0,204,0,184,0,141,0,0,0,93,0,216,0,165,0,170,0,59,0,94,0,12,0,165,0,157,0,0,0,45,0,69,0,45,0,163,0,165,0,36,0,52,0,48,0,0,0,103,0,178,0,138,0,100,0,1,0,211,0,147,0,107,0,217,0,183,0,0,0,47,0,94,0,121,0,78,0,0,0,92,0,0,0,65,0,182,0,86,0,123,0,214,0,0,0,40,0,138,0,125,0,57,0,0,0,0,0,43,0,29,0,175,0,0,0,86,0,245,0,167,0,0,0,215,0,26,0,15,0,0,0,0,0,52,0,215,0,28,0,61,0,214,0,0,0,78,0,182,0,22,0,138,0,0,0,171,0,67,0,35,0,85,0,67,0,0,0,24,0,90,0,0,0,203,0,116,0,0,0,65,0,0,0,50,0,0,0,25,0,0,0,244,0,195,0,0,0,241,0,17,0,233,0,55,0,82,0,0,0,0,0,0,0,237,0,34,0,12,0,41,0,0,0,129,0,104,0,114,0,121,0,121,0,157,0,35,0,0,0,0,0,174,0,16,0,12,0,121,0,146,0,1,0,0,0,135,0,53,0,115,0,0,0,219,0,202,0,49,0,77,0,27,0,60,0,0,0,149,0,43,0,87,0,0,0,85,0,250,0,250,0,159,0,104,0,130,0,216,0,97,0,0,0,141,0,0,0,101,0,118,0,6,0,0,0,194,0,212,0,206,0,244,0,231,0,0,0,30,0,55,0,204,0,110,0,0,0,41,0,182,0,81,0,149,0,101,0,0,0,9,0,151,0,52,0,0,0,65,0,117,0,93,0,153,0,248,0,145,0,143,0,237,0,90,0,149,0,32,0,0,0,0,0,102,0,0,0,126,0,239,0,150,0,0,0,109,0,4,0,0,0,11,0,188,0,9,0,0,0,4,0,124,0,66,0,0,0,172,0,167,0,1,0,158,0,85,0,0,0,235,0,97,0,14,0,0,0,0,0,169,0,252,0,68,0,69,0,0,0,37,0,95,0,30,0,0,0,0,0,194,0,66,0,0,0,60,0,212,0,43,0,33,0,228,0,248,0,0,0,216,0,0,0,228,0,46,0,141,0,63,0,0,0,244,0,92,0,122,0,169,0,249,0,71,0,214,0,123,0,163,0,0,0,11,0,147,0,0,0,158,0,0,0,123,0,106,0,206,0,159,0,168,0,213,0,22,0,163,0,188,0,0,0,183,0,71,0,105,0,175,0,64,0,0,0,1,0,0,0,190,0,54,0,108,0,0,0,152,0,95,0,45,0,209,0,145,0,63,0,0,0,38,0,0,0,28,0,16,0,237,0,0,0,10,0,177,0,219,0,0,0,21,0,0,0,0,0,0,0,38,0,185,0,173,0,41,0,116,0,36,0,0,0,35,0,245,0,130,0,28,0,0,0,159,0,91,0,153,0,204,0,131,0,45,0,102,0,134,0,106,0,84,0,247,0,0,0,186,0,44,0,4,0,191,0,241,0,0,0,31,0,239,0,22,0,0,0,253,0,0,0,0,0,0,0,244,0,254,0,91,0,131,0,0,0,113,0,126,0,0,0,243,0,0,0,94,0,149,0,110,0,155,0,253,0,142,0,0,0,0,0,21,0,216,0,15,0,247,0,199,0,87,0,81,0,60,0,0,0,28,0,25,0,20,0,86,0,129,0,0,0,226,0,216,0,0,0,0,0,189,0,0,0,105,0,45,0,55,0,0,0,156,0,195,0,131,0,0,0,179,0,118,0,0,0,77,0,125,0,142,0,148,0,26,0,217,0,74,0,109,0,140,0,89,0,145,0,107,0,0,0,0,0,66,0,252,0,202,0,118,0,89,0,0,0,210,0,106,0,0,0,137,0,83,0,41,0,40,0,81,0,250,0,243,0,13,0,51,0,203,0,0,0,68,0,8,0,113,0,254,0,0,0,50,0,177,0,0,0,1,0,63,0,82,0,220,0,20,0,0,0,0,0,162,0,88,0,1,0,30,0,28,0,181,0,133,0,3,0,6,0,44,0,14,0,177,0,179,0,0,0,144,0,253,0,222,0,136,0,0,0,73,0,51,0,209,0,154,0,52,0,220,0,231,0,173,0,19,0,21,0,13,0,238,0,110,0,0,0,69,0,0,0,243,0,162,0,44,0,184,0,0,0,37,0,57,0,18,0,255,0,0,0,178,0,178,0,22,0,199,0,0,0,95,0,132,0,238,0,94,0,119,0,112,0,159,0,203,0,221,0,192,0,0,0,138,0,0,0,229,0,213,0,62,0,28,0,179,0,0,0,115,0,179,0,102,0,84,0,30,0,186,0,0,0,164,0,111,0,0,0,214,0,154,0,0,0,44,0,148,0,0,0,0,0,58,0,0,0,98,0,191,0,127,0,238,0,57,0,60,0,66,0,100,0,226,0,163,0,17,0,204,0,0,0,0,0,177,0,83,0,44,0,0,0,0,0,142,0,33,0,207,0,153,0,0,0,0,0,217,0,50,0,1,0,169,0,128,0,85,0,81,0,50,0,22,0,44,0,49,0,192,0,75,0,0,0,158,0,0,0,77,0,176,0,183,0,184,0,124,0,91,0,151,0,150,0,0,0,0,0,168,0,186,0,55,0,36,0,150,0,0,0,77,0,207,0,187,0,167,0,228,0,0,0,18,0,0,0,0,0,73,0,205,0,1,0,132,0,166,0,0,0,0,0,0,0,0,0,64,0,177,0,227,0,172,0,43,0,84,0,179,0,0,0,34,0,150,0,137,0,56,0,87,0,17,0,54,0,41,0,97,0,21,0,103,0,80,0,153,0,162,0,130,0,111,0,59,0,176,0,0,0,181,0,123,0,116,0,44,0,0,0,219,0,140,0,38,0,0,0,162,0,0,0,247,0,21,0,162,0,17,0,0,0,52,0,250,0,175,0,39,0,220,0,164,0,14,0,0,0,83,0,53,0,176,0,0,0,224,0,4,0,29,0,75,0,89,0,216,0,52,0,87,0,124,0,152,0,0,0,0,0,10,0,162,0,18,0,239,0,234,0,42,0,242,0,196,0,164,0,0,0,138,0,201,0,0,0,74,0,170,0,58,0,219,0,0,0,0,0,150,0,243,0,91,0,0,0,186,0,100,0,56,0,138,0,241,0,162,0,54,0,237,0,129,0,196,0,28,0,117,0,0,0,123,0,164,0,36,0,60,0,1,0,46,0,0,0,27,0,74,0,95,0,175,0,132,0,211,0,15,0,246,0,0,0,206,0,0,0,0,0,0,0,203,0,45,0,171,0,0,0,62,0,188,0,111,0,140,0,0,0,0,0,112,0,0,0,247,0,0,0,175,0,14,0,34,0,0,0,112,0,204,0,0,0,170,0,0,0,123,0,71,0,54,0,190,0,52,0,250,0,0,0,25,0,23,0,230,0,95,0,175,0,255,0,227,0,222,0,62,0,0,0,0,0,70,0,0,0,75,0,105,0,21,0,0,0,2,0,15,0,255,0,0,0,213,0,0,0,77,0,67,0);
signal scenario_full  : scenario_type := (193,31,193,30,137,31,111,31,34,31,34,30,239,31,216,31,216,30,185,31,183,31,228,31,197,31,119,31,45,31,45,30,67,31,67,30,67,29,12,31,12,30,75,31,75,30,235,31,235,30,175,31,175,30,28,31,23,31,23,30,23,29,214,31,184,31,184,30,111,31,111,30,222,31,102,31,39,31,39,30,61,31,100,31,118,31,73,31,204,31,204,30,204,29,75,31,218,31,185,31,109,31,81,31,226,31,226,30,226,29,134,31,30,31,247,31,18,31,18,30,60,31,229,31,114,31,195,31,195,30,23,31,24,31,167,31,67,31,189,31,189,30,182,31,3,31,3,30,119,31,119,30,119,29,190,31,207,31,125,31,202,31,202,30,80,31,99,31,40,31,108,31,59,31,52,31,25,31,164,31,100,31,100,30,251,31,37,31,63,31,204,31,184,31,141,31,141,30,93,31,216,31,165,31,170,31,59,31,94,31,12,31,165,31,157,31,157,30,45,31,69,31,45,31,163,31,165,31,36,31,52,31,48,31,48,30,103,31,178,31,138,31,100,31,1,31,211,31,147,31,107,31,217,31,183,31,183,30,47,31,94,31,121,31,78,31,78,30,92,31,92,30,65,31,182,31,86,31,123,31,214,31,214,30,40,31,138,31,125,31,57,31,57,30,57,29,43,31,29,31,175,31,175,30,86,31,245,31,167,31,167,30,215,31,26,31,15,31,15,30,15,29,52,31,215,31,28,31,61,31,214,31,214,30,78,31,182,31,22,31,138,31,138,30,171,31,67,31,35,31,85,31,67,31,67,30,24,31,90,31,90,30,203,31,116,31,116,30,65,31,65,30,50,31,50,30,25,31,25,30,244,31,195,31,195,30,241,31,17,31,233,31,55,31,82,31,82,30,82,29,82,28,237,31,34,31,12,31,41,31,41,30,129,31,104,31,114,31,121,31,121,31,157,31,35,31,35,30,35,29,174,31,16,31,12,31,121,31,146,31,1,31,1,30,135,31,53,31,115,31,115,30,219,31,202,31,49,31,77,31,27,31,60,31,60,30,149,31,43,31,87,31,87,30,85,31,250,31,250,31,159,31,104,31,130,31,216,31,97,31,97,30,141,31,141,30,101,31,118,31,6,31,6,30,194,31,212,31,206,31,244,31,231,31,231,30,30,31,55,31,204,31,110,31,110,30,41,31,182,31,81,31,149,31,101,31,101,30,9,31,151,31,52,31,52,30,65,31,117,31,93,31,153,31,248,31,145,31,143,31,237,31,90,31,149,31,32,31,32,30,32,29,102,31,102,30,126,31,239,31,150,31,150,30,109,31,4,31,4,30,11,31,188,31,9,31,9,30,4,31,124,31,66,31,66,30,172,31,167,31,1,31,158,31,85,31,85,30,235,31,97,31,14,31,14,30,14,29,169,31,252,31,68,31,69,31,69,30,37,31,95,31,30,31,30,30,30,29,194,31,66,31,66,30,60,31,212,31,43,31,33,31,228,31,248,31,248,30,216,31,216,30,228,31,46,31,141,31,63,31,63,30,244,31,92,31,122,31,169,31,249,31,71,31,214,31,123,31,163,31,163,30,11,31,147,31,147,30,158,31,158,30,123,31,106,31,206,31,159,31,168,31,213,31,22,31,163,31,188,31,188,30,183,31,71,31,105,31,175,31,64,31,64,30,1,31,1,30,190,31,54,31,108,31,108,30,152,31,95,31,45,31,209,31,145,31,63,31,63,30,38,31,38,30,28,31,16,31,237,31,237,30,10,31,177,31,219,31,219,30,21,31,21,30,21,29,21,28,38,31,185,31,173,31,41,31,116,31,36,31,36,30,35,31,245,31,130,31,28,31,28,30,159,31,91,31,153,31,204,31,131,31,45,31,102,31,134,31,106,31,84,31,247,31,247,30,186,31,44,31,4,31,191,31,241,31,241,30,31,31,239,31,22,31,22,30,253,31,253,30,253,29,253,28,244,31,254,31,91,31,131,31,131,30,113,31,126,31,126,30,243,31,243,30,94,31,149,31,110,31,155,31,253,31,142,31,142,30,142,29,21,31,216,31,15,31,247,31,199,31,87,31,81,31,60,31,60,30,28,31,25,31,20,31,86,31,129,31,129,30,226,31,216,31,216,30,216,29,189,31,189,30,105,31,45,31,55,31,55,30,156,31,195,31,131,31,131,30,179,31,118,31,118,30,77,31,125,31,142,31,148,31,26,31,217,31,74,31,109,31,140,31,89,31,145,31,107,31,107,30,107,29,66,31,252,31,202,31,118,31,89,31,89,30,210,31,106,31,106,30,137,31,83,31,41,31,40,31,81,31,250,31,243,31,13,31,51,31,203,31,203,30,68,31,8,31,113,31,254,31,254,30,50,31,177,31,177,30,1,31,63,31,82,31,220,31,20,31,20,30,20,29,162,31,88,31,1,31,30,31,28,31,181,31,133,31,3,31,6,31,44,31,14,31,177,31,179,31,179,30,144,31,253,31,222,31,136,31,136,30,73,31,51,31,209,31,154,31,52,31,220,31,231,31,173,31,19,31,21,31,13,31,238,31,110,31,110,30,69,31,69,30,243,31,162,31,44,31,184,31,184,30,37,31,57,31,18,31,255,31,255,30,178,31,178,31,22,31,199,31,199,30,95,31,132,31,238,31,94,31,119,31,112,31,159,31,203,31,221,31,192,31,192,30,138,31,138,30,229,31,213,31,62,31,28,31,179,31,179,30,115,31,179,31,102,31,84,31,30,31,186,31,186,30,164,31,111,31,111,30,214,31,154,31,154,30,44,31,148,31,148,30,148,29,58,31,58,30,98,31,191,31,127,31,238,31,57,31,60,31,66,31,100,31,226,31,163,31,17,31,204,31,204,30,204,29,177,31,83,31,44,31,44,30,44,29,142,31,33,31,207,31,153,31,153,30,153,29,217,31,50,31,1,31,169,31,128,31,85,31,81,31,50,31,22,31,44,31,49,31,192,31,75,31,75,30,158,31,158,30,77,31,176,31,183,31,184,31,124,31,91,31,151,31,150,31,150,30,150,29,168,31,186,31,55,31,36,31,150,31,150,30,77,31,207,31,187,31,167,31,228,31,228,30,18,31,18,30,18,29,73,31,205,31,1,31,132,31,166,31,166,30,166,29,166,28,166,27,64,31,177,31,227,31,172,31,43,31,84,31,179,31,179,30,34,31,150,31,137,31,56,31,87,31,17,31,54,31,41,31,97,31,21,31,103,31,80,31,153,31,162,31,130,31,111,31,59,31,176,31,176,30,181,31,123,31,116,31,44,31,44,30,219,31,140,31,38,31,38,30,162,31,162,30,247,31,21,31,162,31,17,31,17,30,52,31,250,31,175,31,39,31,220,31,164,31,14,31,14,30,83,31,53,31,176,31,176,30,224,31,4,31,29,31,75,31,89,31,216,31,52,31,87,31,124,31,152,31,152,30,152,29,10,31,162,31,18,31,239,31,234,31,42,31,242,31,196,31,164,31,164,30,138,31,201,31,201,30,74,31,170,31,58,31,219,31,219,30,219,29,150,31,243,31,91,31,91,30,186,31,100,31,56,31,138,31,241,31,162,31,54,31,237,31,129,31,196,31,28,31,117,31,117,30,123,31,164,31,36,31,60,31,1,31,46,31,46,30,27,31,74,31,95,31,175,31,132,31,211,31,15,31,246,31,246,30,206,31,206,30,206,29,206,28,203,31,45,31,171,31,171,30,62,31,188,31,111,31,140,31,140,30,140,29,112,31,112,30,247,31,247,30,175,31,14,31,34,31,34,30,112,31,204,31,204,30,170,31,170,30,123,31,71,31,54,31,190,31,52,31,250,31,250,30,25,31,23,31,230,31,95,31,175,31,255,31,227,31,222,31,62,31,62,30,62,29,70,31,70,30,75,31,105,31,21,31,21,30,2,31,15,31,255,31,255,30,213,31,213,30,77,31,67,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
