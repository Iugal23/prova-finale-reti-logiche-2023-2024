-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 557;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (140,0,114,0,25,0,228,0,252,0,129,0,103,0,174,0,0,0,49,0,28,0,186,0,99,0,96,0,0,0,0,0,182,0,72,0,66,0,94,0,127,0,200,0,29,0,149,0,152,0,18,0,0,0,205,0,237,0,160,0,19,0,62,0,38,0,5,0,57,0,0,0,112,0,95,0,86,0,14,0,159,0,0,0,122,0,154,0,36,0,55,0,143,0,53,0,0,0,8,0,61,0,0,0,121,0,242,0,6,0,0,0,224,0,0,0,77,0,112,0,120,0,88,0,61,0,128,0,123,0,35,0,14,0,0,0,203,0,220,0,178,0,0,0,7,0,249,0,83,0,43,0,102,0,236,0,0,0,79,0,185,0,176,0,180,0,99,0,52,0,183,0,56,0,0,0,182,0,96,0,15,0,206,0,102,0,245,0,0,0,50,0,84,0,0,0,116,0,225,0,167,0,59,0,144,0,62,0,0,0,249,0,118,0,250,0,3,0,13,0,125,0,28,0,0,0,242,0,172,0,171,0,146,0,138,0,25,0,108,0,22,0,55,0,124,0,156,0,122,0,40,0,0,0,143,0,54,0,132,0,0,0,0,0,0,0,92,0,0,0,19,0,138,0,36,0,106,0,0,0,181,0,196,0,37,0,184,0,14,0,0,0,167,0,94,0,0,0,89,0,36,0,0,0,163,0,237,0,178,0,0,0,0,0,102,0,148,0,74,0,0,0,104,0,140,0,0,0,21,0,113,0,83,0,0,0,60,0,193,0,191,0,95,0,162,0,108,0,195,0,149,0,47,0,87,0,51,0,17,0,135,0,46,0,0,0,172,0,60,0,119,0,58,0,19,0,23,0,52,0,225,0,242,0,71,0,157,0,152,0,0,0,121,0,14,0,0,0,0,0,0,0,172,0,88,0,0,0,33,0,37,0,92,0,191,0,37,0,111,0,5,0,76,0,0,0,20,0,161,0,222,0,141,0,0,0,62,0,30,0,208,0,246,0,75,0,90,0,129,0,48,0,50,0,0,0,125,0,67,0,63,0,137,0,0,0,9,0,0,0,159,0,253,0,247,0,81,0,53,0,238,0,5,0,153,0,138,0,0,0,0,0,58,0,106,0,0,0,0,0,168,0,253,0,216,0,0,0,119,0,174,0,30,0,18,0,46,0,0,0,230,0,32,0,146,0,23,0,100,0,61,0,0,0,253,0,232,0,246,0,141,0,8,0,0,0,24,0,27,0,202,0,0,0,0,0,0,0,149,0,137,0,92,0,149,0,0,0,78,0,202,0,225,0,66,0,0,0,30,0,164,0,0,0,120,0,141,0,55,0,207,0,140,0,0,0,70,0,80,0,0,0,216,0,46,0,85,0,158,0,253,0,47,0,0,0,162,0,91,0,0,0,249,0,0,0,213,0,74,0,33,0,0,0,206,0,79,0,184,0,156,0,63,0,156,0,244,0,0,0,103,0,138,0,94,0,8,0,116,0,248,0,35,0,229,0,0,0,91,0,57,0,123,0,218,0,51,0,177,0,210,0,54,0,24,0,0,0,123,0,120,0,209,0,0,0,116,0,0,0,194,0,0,0,52,0,166,0,0,0,0,0,216,0,215,0,154,0,219,0,96,0,135,0,0,0,186,0,113,0,231,0,105,0,165,0,191,0,0,0,0,0,215,0,0,0,0,0,106,0,58,0,0,0,0,0,0,0,60,0,145,0,129,0,15,0,21,0,0,0,16,0,6,0,224,0,0,0,68,0,149,0,216,0,192,0,75,0,0,0,37,0,108,0,228,0,144,0,218,0,169,0,46,0,55,0,25,0,212,0,254,0,102,0,21,0,150,0,43,0,253,0,247,0,36,0,147,0,111,0,10,0,116,0,241,0,162,0,129,0,66,0,116,0,198,0,251,0,0,0,69,0,133,0,188,0,217,0,0,0,58,0,241,0,107,0,195,0,90,0,0,0,137,0,97,0,133,0,247,0,18,0,219,0,0,0,134,0,89,0,142,0,148,0,218,0,193,0,173,0,91,0,162,0,62,0,0,0,0,0,226,0,50,0,76,0,124,0,32,0,239,0,8,0,0,0,196,0,0,0,224,0,0,0,87,0,197,0,4,0,201,0,59,0,22,0,0,0,0,0,161,0,119,0,0,0,132,0,119,0,142,0,0,0,59,0,0,0,0,0,224,0,0,0,192,0,5,0,165,0,44,0,74,0,62,0,68,0,7,0,211,0,0,0,86,0,8,0,59,0,9,0,147,0,59,0,199,0,104,0,56,0,97,0,72,0,106,0,101,0,0,0,0,0,0,0,0,0,176,0,0,0,92,0,176,0,151,0,0,0,120,0,141,0,182,0,116,0,12,0,121,0,51,0,126,0,216,0,61,0,78,0,0,0,20,0,197,0,208,0,97,0,159,0,180,0,71,0,106,0,0,0,0,0,176,0,212,0,0,0,93,0,114,0,205,0,223,0,223,0,21,0,71,0,61,0,0,0,160,0,0,0,0,0);
signal scenario_full  : scenario_type := (140,31,114,31,25,31,228,31,252,31,129,31,103,31,174,31,174,30,49,31,28,31,186,31,99,31,96,31,96,30,96,29,182,31,72,31,66,31,94,31,127,31,200,31,29,31,149,31,152,31,18,31,18,30,205,31,237,31,160,31,19,31,62,31,38,31,5,31,57,31,57,30,112,31,95,31,86,31,14,31,159,31,159,30,122,31,154,31,36,31,55,31,143,31,53,31,53,30,8,31,61,31,61,30,121,31,242,31,6,31,6,30,224,31,224,30,77,31,112,31,120,31,88,31,61,31,128,31,123,31,35,31,14,31,14,30,203,31,220,31,178,31,178,30,7,31,249,31,83,31,43,31,102,31,236,31,236,30,79,31,185,31,176,31,180,31,99,31,52,31,183,31,56,31,56,30,182,31,96,31,15,31,206,31,102,31,245,31,245,30,50,31,84,31,84,30,116,31,225,31,167,31,59,31,144,31,62,31,62,30,249,31,118,31,250,31,3,31,13,31,125,31,28,31,28,30,242,31,172,31,171,31,146,31,138,31,25,31,108,31,22,31,55,31,124,31,156,31,122,31,40,31,40,30,143,31,54,31,132,31,132,30,132,29,132,28,92,31,92,30,19,31,138,31,36,31,106,31,106,30,181,31,196,31,37,31,184,31,14,31,14,30,167,31,94,31,94,30,89,31,36,31,36,30,163,31,237,31,178,31,178,30,178,29,102,31,148,31,74,31,74,30,104,31,140,31,140,30,21,31,113,31,83,31,83,30,60,31,193,31,191,31,95,31,162,31,108,31,195,31,149,31,47,31,87,31,51,31,17,31,135,31,46,31,46,30,172,31,60,31,119,31,58,31,19,31,23,31,52,31,225,31,242,31,71,31,157,31,152,31,152,30,121,31,14,31,14,30,14,29,14,28,172,31,88,31,88,30,33,31,37,31,92,31,191,31,37,31,111,31,5,31,76,31,76,30,20,31,161,31,222,31,141,31,141,30,62,31,30,31,208,31,246,31,75,31,90,31,129,31,48,31,50,31,50,30,125,31,67,31,63,31,137,31,137,30,9,31,9,30,159,31,253,31,247,31,81,31,53,31,238,31,5,31,153,31,138,31,138,30,138,29,58,31,106,31,106,30,106,29,168,31,253,31,216,31,216,30,119,31,174,31,30,31,18,31,46,31,46,30,230,31,32,31,146,31,23,31,100,31,61,31,61,30,253,31,232,31,246,31,141,31,8,31,8,30,24,31,27,31,202,31,202,30,202,29,202,28,149,31,137,31,92,31,149,31,149,30,78,31,202,31,225,31,66,31,66,30,30,31,164,31,164,30,120,31,141,31,55,31,207,31,140,31,140,30,70,31,80,31,80,30,216,31,46,31,85,31,158,31,253,31,47,31,47,30,162,31,91,31,91,30,249,31,249,30,213,31,74,31,33,31,33,30,206,31,79,31,184,31,156,31,63,31,156,31,244,31,244,30,103,31,138,31,94,31,8,31,116,31,248,31,35,31,229,31,229,30,91,31,57,31,123,31,218,31,51,31,177,31,210,31,54,31,24,31,24,30,123,31,120,31,209,31,209,30,116,31,116,30,194,31,194,30,52,31,166,31,166,30,166,29,216,31,215,31,154,31,219,31,96,31,135,31,135,30,186,31,113,31,231,31,105,31,165,31,191,31,191,30,191,29,215,31,215,30,215,29,106,31,58,31,58,30,58,29,58,28,60,31,145,31,129,31,15,31,21,31,21,30,16,31,6,31,224,31,224,30,68,31,149,31,216,31,192,31,75,31,75,30,37,31,108,31,228,31,144,31,218,31,169,31,46,31,55,31,25,31,212,31,254,31,102,31,21,31,150,31,43,31,253,31,247,31,36,31,147,31,111,31,10,31,116,31,241,31,162,31,129,31,66,31,116,31,198,31,251,31,251,30,69,31,133,31,188,31,217,31,217,30,58,31,241,31,107,31,195,31,90,31,90,30,137,31,97,31,133,31,247,31,18,31,219,31,219,30,134,31,89,31,142,31,148,31,218,31,193,31,173,31,91,31,162,31,62,31,62,30,62,29,226,31,50,31,76,31,124,31,32,31,239,31,8,31,8,30,196,31,196,30,224,31,224,30,87,31,197,31,4,31,201,31,59,31,22,31,22,30,22,29,161,31,119,31,119,30,132,31,119,31,142,31,142,30,59,31,59,30,59,29,224,31,224,30,192,31,5,31,165,31,44,31,74,31,62,31,68,31,7,31,211,31,211,30,86,31,8,31,59,31,9,31,147,31,59,31,199,31,104,31,56,31,97,31,72,31,106,31,101,31,101,30,101,29,101,28,101,27,176,31,176,30,92,31,176,31,151,31,151,30,120,31,141,31,182,31,116,31,12,31,121,31,51,31,126,31,216,31,61,31,78,31,78,30,20,31,197,31,208,31,97,31,159,31,180,31,71,31,106,31,106,30,106,29,176,31,212,31,212,30,93,31,114,31,205,31,223,31,223,31,21,31,71,31,61,31,61,30,160,31,160,30,160,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
