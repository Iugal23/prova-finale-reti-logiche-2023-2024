-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_847 is
end project_tb_847;

architecture project_tb_arch_847 of project_tb_847 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 770;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,78,0,134,0,0,0,117,0,66,0,190,0,52,0,0,0,197,0,116,0,241,0,52,0,57,0,157,0,217,0,0,0,16,0,144,0,211,0,136,0,0,0,169,0,0,0,248,0,0,0,140,0,222,0,163,0,51,0,236,0,132,0,0,0,237,0,100,0,2,0,47,0,50,0,0,0,97,0,58,0,5,0,168,0,119,0,175,0,45,0,0,0,56,0,144,0,110,0,127,0,198,0,116,0,152,0,203,0,166,0,43,0,234,0,201,0,180,0,71,0,204,0,19,0,39,0,194,0,0,0,114,0,168,0,186,0,171,0,23,0,128,0,116,0,0,0,0,0,59,0,134,0,28,0,100,0,14,0,121,0,11,0,34,0,123,0,26,0,167,0,21,0,79,0,239,0,249,0,146,0,16,0,88,0,219,0,106,0,8,0,57,0,107,0,0,0,0,0,195,0,102,0,0,0,54,0,172,0,251,0,0,0,38,0,235,0,225,0,217,0,0,0,101,0,0,0,214,0,0,0,116,0,0,0,143,0,188,0,247,0,51,0,220,0,35,0,0,0,0,0,52,0,0,0,0,0,89,0,73,0,11,0,250,0,177,0,0,0,0,0,64,0,246,0,23,0,0,0,0,0,215,0,2,0,165,0,76,0,21,0,232,0,38,0,91,0,225,0,201,0,172,0,94,0,0,0,103,0,137,0,142,0,76,0,131,0,192,0,157,0,0,0,143,0,63,0,13,0,113,0,70,0,150,0,147,0,0,0,55,0,82,0,88,0,162,0,109,0,90,0,103,0,250,0,0,0,180,0,244,0,222,0,205,0,235,0,21,0,202,0,125,0,0,0,80,0,54,0,96,0,112,0,0,0,87,0,1,0,45,0,16,0,54,0,170,0,0,0,10,0,135,0,55,0,107,0,200,0,95,0,191,0,173,0,198,0,212,0,227,0,0,0,108,0,245,0,183,0,22,0,14,0,189,0,41,0,57,0,163,0,181,0,0,0,0,0,4,0,155,0,94,0,0,0,172,0,93,0,236,0,243,0,245,0,43,0,38,0,84,0,0,0,139,0,107,0,254,0,98,0,124,0,0,0,81,0,79,0,0,0,191,0,14,0,50,0,71,0,218,0,198,0,0,0,104,0,161,0,131,0,0,0,0,0,0,0,0,0,29,0,51,0,211,0,22,0,45,0,0,0,18,0,125,0,215,0,128,0,0,0,0,0,74,0,196,0,249,0,0,0,184,0,67,0,46,0,169,0,109,0,80,0,120,0,0,0,206,0,155,0,60,0,84,0,200,0,170,0,173,0,235,0,222,0,85,0,170,0,161,0,159,0,226,0,145,0,44,0,18,0,0,0,26,0,11,0,17,0,123,0,12,0,226,0,151,0,182,0,98,0,244,0,173,0,230,0,171,0,94,0,185,0,110,0,141,0,203,0,27,0,145,0,11,0,161,0,175,0,0,0,151,0,129,0,39,0,63,0,65,0,0,0,113,0,3,0,136,0,8,0,248,0,252,0,17,0,187,0,237,0,0,0,67,0,89,0,246,0,42,0,221,0,62,0,104,0,133,0,76,0,0,0,68,0,69,0,0,0,0,0,167,0,10,0,104,0,0,0,135,0,57,0,238,0,228,0,0,0,164,0,175,0,20,0,117,0,61,0,43,0,138,0,166,0,0,0,0,0,226,0,172,0,0,0,232,0,30,0,91,0,255,0,170,0,149,0,243,0,0,0,13,0,174,0,20,0,160,0,166,0,152,0,0,0,0,0,197,0,224,0,169,0,134,0,235,0,178,0,72,0,0,0,0,0,249,0,185,0,122,0,203,0,123,0,184,0,251,0,57,0,152,0,0,0,98,0,0,0,85,0,246,0,184,0,136,0,156,0,0,0,217,0,250,0,139,0,205,0,242,0,0,0,0,0,0,0,249,0,139,0,175,0,194,0,250,0,93,0,0,0,219,0,0,0,0,0,14,0,103,0,52,0,23,0,0,0,0,0,97,0,244,0,184,0,180,0,8,0,50,0,143,0,26,0,21,0,69,0,84,0,0,0,159,0,186,0,10,0,0,0,37,0,29,0,251,0,237,0,80,0,0,0,20,0,251,0,213,0,6,0,0,0,155,0,0,0,26,0,202,0,129,0,0,0,104,0,189,0,41,0,0,0,109,0,57,0,159,0,253,0,237,0,186,0,0,0,106,0,212,0,91,0,196,0,0,0,118,0,0,0,110,0,217,0,121,0,212,0,98,0,131,0,161,0,180,0,0,0,212,0,139,0,60,0,120,0,0,0,0,0,0,0,0,0,92,0,102,0,55,0,145,0,164,0,108,0,0,0,95,0,1,0,0,0,223,0,154,0,175,0,235,0,45,0,178,0,5,0,0,0,198,0,36,0,53,0,32,0,248,0,84,0,156,0,22,0,113,0,137,0,233,0,0,0,18,0,205,0,45,0,40,0,0,0,110,0,75,0,0,0,0,0,246,0,224,0,182,0,0,0,108,0,47,0,124,0,232,0,31,0,175,0,112,0,209,0,1,0,185,0,90,0,40,0,0,0,137,0,79,0,74,0,0,0,0,0,28,0,213,0,0,0,109,0,26,0,0,0,91,0,125,0,217,0,126,0,121,0,215,0,0,0,141,0,123,0,0,0,68,0,179,0,228,0,52,0,175,0,83,0,140,0,19,0,42,0,0,0,165,0,35,0,30,0,128,0,91,0,117,0,250,0,18,0,0,0,18,0,116,0,119,0,68,0,206,0,56,0,0,0,244,0,65,0,150,0,231,0,205,0,4,0,110,0,254,0,195,0,58,0,250,0,16,0,0,0,170,0,0,0,52,0,63,0,197,0,105,0,137,0,60,0,168,0,94,0,198,0,152,0,0,0,0,0,0,0,79,0,58,0,252,0,16,0,193,0,0,0,235,0,249,0,186,0,99,0,8,0,186,0,0,0,171,0,161,0,254,0,190,0,105,0,157,0,134,0,110,0,238,0,24,0,25,0,229,0,217,0,184,0,233,0,11,0,176,0,166,0,218,0,194,0,224,0,114,0,0,0,78,0,0,0,190,0,171,0,0,0,53,0,169,0,224,0,154,0,48,0,49,0,89,0,0,0,94,0,221,0,128,0,51,0,79,0,231,0,254,0,138,0,49,0,25,0,83,0,0,0,248,0,84,0,33,0,0,0,243,0,98,0,132,0,69,0,82,0,6,0,0,0,63,0,154,0,140,0,61,0,206,0,226,0,193,0,0,0,65,0,0,0,0,0,239,0,0,0,0,0,252,0,0,0,215,0,0,0,157,0,230,0,0,0,147,0,18,0,107,0,152,0,0,0,162,0,61,0,180,0,123,0,99,0,150,0,69,0,176,0,23,0,0,0,0,0,0,0,71,0,232,0,213,0,31,0,114,0,40,0,0,0,0,0,150,0,18,0,56,0,173,0,194,0,14,0,96,0,0,0);
signal scenario_full  : scenario_type := (0,0,78,31,134,31,134,30,117,31,66,31,190,31,52,31,52,30,197,31,116,31,241,31,52,31,57,31,157,31,217,31,217,30,16,31,144,31,211,31,136,31,136,30,169,31,169,30,248,31,248,30,140,31,222,31,163,31,51,31,236,31,132,31,132,30,237,31,100,31,2,31,47,31,50,31,50,30,97,31,58,31,5,31,168,31,119,31,175,31,45,31,45,30,56,31,144,31,110,31,127,31,198,31,116,31,152,31,203,31,166,31,43,31,234,31,201,31,180,31,71,31,204,31,19,31,39,31,194,31,194,30,114,31,168,31,186,31,171,31,23,31,128,31,116,31,116,30,116,29,59,31,134,31,28,31,100,31,14,31,121,31,11,31,34,31,123,31,26,31,167,31,21,31,79,31,239,31,249,31,146,31,16,31,88,31,219,31,106,31,8,31,57,31,107,31,107,30,107,29,195,31,102,31,102,30,54,31,172,31,251,31,251,30,38,31,235,31,225,31,217,31,217,30,101,31,101,30,214,31,214,30,116,31,116,30,143,31,188,31,247,31,51,31,220,31,35,31,35,30,35,29,52,31,52,30,52,29,89,31,73,31,11,31,250,31,177,31,177,30,177,29,64,31,246,31,23,31,23,30,23,29,215,31,2,31,165,31,76,31,21,31,232,31,38,31,91,31,225,31,201,31,172,31,94,31,94,30,103,31,137,31,142,31,76,31,131,31,192,31,157,31,157,30,143,31,63,31,13,31,113,31,70,31,150,31,147,31,147,30,55,31,82,31,88,31,162,31,109,31,90,31,103,31,250,31,250,30,180,31,244,31,222,31,205,31,235,31,21,31,202,31,125,31,125,30,80,31,54,31,96,31,112,31,112,30,87,31,1,31,45,31,16,31,54,31,170,31,170,30,10,31,135,31,55,31,107,31,200,31,95,31,191,31,173,31,198,31,212,31,227,31,227,30,108,31,245,31,183,31,22,31,14,31,189,31,41,31,57,31,163,31,181,31,181,30,181,29,4,31,155,31,94,31,94,30,172,31,93,31,236,31,243,31,245,31,43,31,38,31,84,31,84,30,139,31,107,31,254,31,98,31,124,31,124,30,81,31,79,31,79,30,191,31,14,31,50,31,71,31,218,31,198,31,198,30,104,31,161,31,131,31,131,30,131,29,131,28,131,27,29,31,51,31,211,31,22,31,45,31,45,30,18,31,125,31,215,31,128,31,128,30,128,29,74,31,196,31,249,31,249,30,184,31,67,31,46,31,169,31,109,31,80,31,120,31,120,30,206,31,155,31,60,31,84,31,200,31,170,31,173,31,235,31,222,31,85,31,170,31,161,31,159,31,226,31,145,31,44,31,18,31,18,30,26,31,11,31,17,31,123,31,12,31,226,31,151,31,182,31,98,31,244,31,173,31,230,31,171,31,94,31,185,31,110,31,141,31,203,31,27,31,145,31,11,31,161,31,175,31,175,30,151,31,129,31,39,31,63,31,65,31,65,30,113,31,3,31,136,31,8,31,248,31,252,31,17,31,187,31,237,31,237,30,67,31,89,31,246,31,42,31,221,31,62,31,104,31,133,31,76,31,76,30,68,31,69,31,69,30,69,29,167,31,10,31,104,31,104,30,135,31,57,31,238,31,228,31,228,30,164,31,175,31,20,31,117,31,61,31,43,31,138,31,166,31,166,30,166,29,226,31,172,31,172,30,232,31,30,31,91,31,255,31,170,31,149,31,243,31,243,30,13,31,174,31,20,31,160,31,166,31,152,31,152,30,152,29,197,31,224,31,169,31,134,31,235,31,178,31,72,31,72,30,72,29,249,31,185,31,122,31,203,31,123,31,184,31,251,31,57,31,152,31,152,30,98,31,98,30,85,31,246,31,184,31,136,31,156,31,156,30,217,31,250,31,139,31,205,31,242,31,242,30,242,29,242,28,249,31,139,31,175,31,194,31,250,31,93,31,93,30,219,31,219,30,219,29,14,31,103,31,52,31,23,31,23,30,23,29,97,31,244,31,184,31,180,31,8,31,50,31,143,31,26,31,21,31,69,31,84,31,84,30,159,31,186,31,10,31,10,30,37,31,29,31,251,31,237,31,80,31,80,30,20,31,251,31,213,31,6,31,6,30,155,31,155,30,26,31,202,31,129,31,129,30,104,31,189,31,41,31,41,30,109,31,57,31,159,31,253,31,237,31,186,31,186,30,106,31,212,31,91,31,196,31,196,30,118,31,118,30,110,31,217,31,121,31,212,31,98,31,131,31,161,31,180,31,180,30,212,31,139,31,60,31,120,31,120,30,120,29,120,28,120,27,92,31,102,31,55,31,145,31,164,31,108,31,108,30,95,31,1,31,1,30,223,31,154,31,175,31,235,31,45,31,178,31,5,31,5,30,198,31,36,31,53,31,32,31,248,31,84,31,156,31,22,31,113,31,137,31,233,31,233,30,18,31,205,31,45,31,40,31,40,30,110,31,75,31,75,30,75,29,246,31,224,31,182,31,182,30,108,31,47,31,124,31,232,31,31,31,175,31,112,31,209,31,1,31,185,31,90,31,40,31,40,30,137,31,79,31,74,31,74,30,74,29,28,31,213,31,213,30,109,31,26,31,26,30,91,31,125,31,217,31,126,31,121,31,215,31,215,30,141,31,123,31,123,30,68,31,179,31,228,31,52,31,175,31,83,31,140,31,19,31,42,31,42,30,165,31,35,31,30,31,128,31,91,31,117,31,250,31,18,31,18,30,18,31,116,31,119,31,68,31,206,31,56,31,56,30,244,31,65,31,150,31,231,31,205,31,4,31,110,31,254,31,195,31,58,31,250,31,16,31,16,30,170,31,170,30,52,31,63,31,197,31,105,31,137,31,60,31,168,31,94,31,198,31,152,31,152,30,152,29,152,28,79,31,58,31,252,31,16,31,193,31,193,30,235,31,249,31,186,31,99,31,8,31,186,31,186,30,171,31,161,31,254,31,190,31,105,31,157,31,134,31,110,31,238,31,24,31,25,31,229,31,217,31,184,31,233,31,11,31,176,31,166,31,218,31,194,31,224,31,114,31,114,30,78,31,78,30,190,31,171,31,171,30,53,31,169,31,224,31,154,31,48,31,49,31,89,31,89,30,94,31,221,31,128,31,51,31,79,31,231,31,254,31,138,31,49,31,25,31,83,31,83,30,248,31,84,31,33,31,33,30,243,31,98,31,132,31,69,31,82,31,6,31,6,30,63,31,154,31,140,31,61,31,206,31,226,31,193,31,193,30,65,31,65,30,65,29,239,31,239,30,239,29,252,31,252,30,215,31,215,30,157,31,230,31,230,30,147,31,18,31,107,31,152,31,152,30,162,31,61,31,180,31,123,31,99,31,150,31,69,31,176,31,23,31,23,30,23,29,23,28,71,31,232,31,213,31,31,31,114,31,40,31,40,30,40,29,150,31,18,31,56,31,173,31,194,31,14,31,96,31,96,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
