-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 983;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (17,0,36,0,16,0,112,0,129,0,144,0,8,0,0,0,204,0,187,0,0,0,114,0,0,0,184,0,236,0,94,0,0,0,4,0,153,0,38,0,152,0,39,0,0,0,0,0,73,0,207,0,205,0,45,0,0,0,98,0,0,0,107,0,156,0,179,0,255,0,87,0,0,0,237,0,73,0,7,0,212,0,51,0,160,0,176,0,122,0,52,0,224,0,157,0,145,0,237,0,163,0,0,0,0,0,74,0,75,0,0,0,51,0,0,0,173,0,4,0,30,0,220,0,210,0,116,0,208,0,228,0,150,0,135,0,195,0,0,0,191,0,0,0,205,0,19,0,13,0,122,0,134,0,77,0,38,0,91,0,39,0,0,0,120,0,34,0,36,0,207,0,27,0,0,0,79,0,248,0,116,0,227,0,244,0,0,0,16,0,52,0,82,0,199,0,57,0,169,0,0,0,33,0,106,0,178,0,72,0,236,0,0,0,242,0,235,0,0,0,101,0,5,0,83,0,15,0,161,0,0,0,0,0,95,0,182,0,112,0,0,0,204,0,113,0,21,0,95,0,0,0,0,0,179,0,91,0,129,0,0,0,85,0,62,0,195,0,198,0,197,0,117,0,0,0,103,0,210,0,194,0,105,0,205,0,156,0,109,0,51,0,110,0,33,0,204,0,240,0,0,0,142,0,8,0,2,0,188,0,40,0,105,0,97,0,214,0,236,0,0,0,0,0,0,0,44,0,182,0,168,0,242,0,22,0,130,0,0,0,0,0,0,0,180,0,232,0,172,0,145,0,200,0,133,0,7,0,0,0,0,0,131,0,196,0,0,0,197,0,0,0,171,0,33,0,71,0,0,0,0,0,150,0,16,0,0,0,26,0,0,0,0,0,222,0,255,0,168,0,130,0,42,0,161,0,170,0,74,0,0,0,36,0,245,0,144,0,133,0,251,0,71,0,196,0,0,0,49,0,44,0,194,0,3,0,148,0,250,0,53,0,0,0,53,0,113,0,154,0,0,0,151,0,0,0,128,0,200,0,147,0,24,0,0,0,211,0,0,0,0,0,79,0,105,0,114,0,0,0,0,0,0,0,7,0,113,0,211,0,0,0,233,0,24,0,0,0,227,0,31,0,192,0,166,0,0,0,141,0,121,0,97,0,125,0,32,0,243,0,244,0,131,0,9,0,36,0,78,0,145,0,0,0,216,0,72,0,86,0,11,0,0,0,168,0,0,0,53,0,197,0,34,0,75,0,0,0,120,0,79,0,0,0,221,0,83,0,207,0,115,0,122,0,231,0,172,0,82,0,237,0,244,0,0,0,29,0,132,0,0,0,52,0,24,0,82,0,48,0,40,0,252,0,117,0,20,0,210,0,94,0,137,0,0,0,115,0,37,0,71,0,151,0,234,0,4,0,41,0,230,0,161,0,0,0,7,0,65,0,149,0,43,0,6,0,102,0,186,0,245,0,127,0,98,0,21,0,17,0,37,0,156,0,203,0,0,0,43,0,196,0,84,0,151,0,96,0,71,0,70,0,0,0,5,0,22,0,206,0,6,0,0,0,95,0,0,0,36,0,48,0,15,0,158,0,156,0,247,0,116,0,70,0,82,0,0,0,0,0,8,0,249,0,0,0,0,0,174,0,221,0,139,0,246,0,119,0,137,0,180,0,47,0,193,0,107,0,171,0,50,0,220,0,0,0,190,0,0,0,152,0,140,0,123,0,0,0,66,0,81,0,110,0,108,0,85,0,44,0,227,0,146,0,137,0,0,0,193,0,14,0,0,0,0,0,149,0,167,0,171,0,5,0,0,0,71,0,22,0,170,0,174,0,84,0,98,0,189,0,0,0,165,0,246,0,55,0,152,0,0,0,0,0,162,0,54,0,245,0,0,0,0,0,0,0,48,0,135,0,0,0,0,0,151,0,70,0,81,0,88,0,160,0,13,0,237,0,178,0,170,0,0,0,100,0,103,0,92,0,5,0,0,0,0,0,96,0,227,0,0,0,183,0,192,0,0,0,126,0,0,0,0,0,108,0,0,0,0,0,38,0,173,0,61,0,0,0,242,0,83,0,0,0,0,0,0,0,206,0,97,0,98,0,236,0,163,0,102,0,254,0,0,0,19,0,153,0,137,0,214,0,0,0,96,0,1,0,0,0,196,0,206,0,91,0,133,0,0,0,202,0,117,0,173,0,138,0,146,0,182,0,233,0,243,0,30,0,170,0,74,0,189,0,187,0,0,0,214,0,40,0,21,0,84,0,255,0,145,0,40,0,244,0,119,0,21,0,0,0,209,0,129,0,93,0,207,0,101,0,0,0,127,0,110,0,255,0,254,0,7,0,9,0,181,0,49,0,88,0,230,0,0,0,0,0,0,0,88,0,0,0,0,0,32,0,111,0,47,0,183,0,133,0,101,0,100,0,76,0,203,0,111,0,63,0,159,0,196,0,56,0,219,0,89,0,174,0,0,0,119,0,41,0,74,0,15,0,204,0,220,0,21,0,145,0,201,0,44,0,0,0,0,0,192,0,211,0,0,0,59,0,129,0,0,0,129,0,58,0,140,0,234,0,0,0,0,0,94,0,52,0,195,0,180,0,77,0,95,0,17,0,130,0,164,0,0,0,0,0,66,0,80,0,132,0,12,0,222,0,244,0,114,0,0,0,94,0,177,0,64,0,0,0,211,0,173,0,110,0,145,0,44,0,202,0,218,0,0,0,30,0,140,0,212,0,0,0,0,0,254,0,0,0,28,0,118,0,0,0,0,0,0,0,63,0,194,0,20,0,172,0,216,0,217,0,151,0,0,0,48,0,24,0,21,0,230,0,215,0,205,0,155,0,55,0,222,0,0,0,234,0,0,0,0,0,52,0,108,0,6,0,37,0,176,0,122,0,232,0,189,0,222,0,171,0,221,0,243,0,226,0,160,0,21,0,86,0,13,0,29,0,16,0,28,0,0,0,227,0,0,0,0,0,13,0,0,0,109,0,97,0,126,0,1,0,0,0,81,0,208,0,209,0,0,0,95,0,88,0,0,0,44,0,155,0,13,0,45,0,0,0,162,0,1,0,0,0,155,0,191,0,0,0,93,0,195,0,180,0,34,0,19,0,0,0,31,0,125,0,177,0,210,0,57,0,206,0,6,0,52,0,171,0,0,0,0,0,0,0,32,0,42,0,120,0,167,0,103,0,91,0,76,0,247,0,99,0,38,0,20,0,109,0,0,0,163,0,0,0,154,0,36,0,24,0,0,0,239,0,204,0,172,0,6,0,251,0,0,0,173,0,252,0,41,0,163,0,32,0,196,0,246,0,87,0,52,0,0,0,0,0,69,0,81,0,107,0,168,0,186,0,37,0,76,0,65,0,12,0,231,0,0,0,0,0,139,0,90,0,136,0,82,0,22,0,10,0,135,0,120,0,53,0,117,0,0,0,0,0,116,0,145,0,178,0,33,0,203,0,111,0,0,0,246,0,171,0,191,0,0,0,28,0,191,0,0,0,8,0,0,0,43,0,31,0,0,0,114,0,0,0,153,0,53,0,250,0,0,0,0,0,0,0,196,0,62,0,230,0,148,0,27,0,0,0,0,0,0,0,234,0,212,0,178,0,60,0,35,0,14,0,54,0,37,0,194,0,0,0,150,0,0,0,97,0,83,0,168,0,206,0,222,0,56,0,0,0,98,0,87,0,61,0,181,0,0,0,0,0,91,0,117,0,29,0,128,0,223,0,0,0,0,0,198,0,138,0,124,0,53,0,0,0,0,0,170,0,68,0,10,0,48,0,0,0,189,0,250,0,28,0,120,0,58,0,0,0,203,0,0,0,38,0,38,0,87,0,113,0,255,0,0,0,32,0,0,0,12,0,182,0,72,0,170,0,254,0,32,0,90,0,198,0,94,0,0,0,196,0,248,0,5,0,0,0,255,0,62,0,161,0,5,0,83,0,90,0,126,0,0,0,205,0,1,0,112,0,218,0,62,0,223,0,255,0,120,0,128,0,0,0,239,0,229,0,71,0,41,0,0,0,250,0,208,0,129,0,80,0,179,0,245,0,0,0,155,0,9,0,164,0,120,0,176,0,12,0,70,0,172,0,77,0,144,0,0,0,230,0,215,0,0,0,0,0,197,0,250,0,0,0,25,0,199,0,35,0,29,0,168,0,186,0,202,0,56,0,200,0,218,0,28,0,0,0,59,0,0,0,55,0,0,0,77,0,135,0,167,0,149,0,122,0,220,0,219,0,77,0,0,0,0,0,0,0,0,0,139,0,137,0,0,0,0,0,206,0,0,0,124,0,26,0,52,0,0,0,0,0,0,0,36,0,35,0,136,0,0,0,102,0,240,0,73,0,211,0,97,0,42,0,0,0,0,0,20,0,35,0,0,0,202,0,76,0,240,0,90,0,0,0,136,0,67,0);
signal scenario_full  : scenario_type := (17,31,36,31,16,31,112,31,129,31,144,31,8,31,8,30,204,31,187,31,187,30,114,31,114,30,184,31,236,31,94,31,94,30,4,31,153,31,38,31,152,31,39,31,39,30,39,29,73,31,207,31,205,31,45,31,45,30,98,31,98,30,107,31,156,31,179,31,255,31,87,31,87,30,237,31,73,31,7,31,212,31,51,31,160,31,176,31,122,31,52,31,224,31,157,31,145,31,237,31,163,31,163,30,163,29,74,31,75,31,75,30,51,31,51,30,173,31,4,31,30,31,220,31,210,31,116,31,208,31,228,31,150,31,135,31,195,31,195,30,191,31,191,30,205,31,19,31,13,31,122,31,134,31,77,31,38,31,91,31,39,31,39,30,120,31,34,31,36,31,207,31,27,31,27,30,79,31,248,31,116,31,227,31,244,31,244,30,16,31,52,31,82,31,199,31,57,31,169,31,169,30,33,31,106,31,178,31,72,31,236,31,236,30,242,31,235,31,235,30,101,31,5,31,83,31,15,31,161,31,161,30,161,29,95,31,182,31,112,31,112,30,204,31,113,31,21,31,95,31,95,30,95,29,179,31,91,31,129,31,129,30,85,31,62,31,195,31,198,31,197,31,117,31,117,30,103,31,210,31,194,31,105,31,205,31,156,31,109,31,51,31,110,31,33,31,204,31,240,31,240,30,142,31,8,31,2,31,188,31,40,31,105,31,97,31,214,31,236,31,236,30,236,29,236,28,44,31,182,31,168,31,242,31,22,31,130,31,130,30,130,29,130,28,180,31,232,31,172,31,145,31,200,31,133,31,7,31,7,30,7,29,131,31,196,31,196,30,197,31,197,30,171,31,33,31,71,31,71,30,71,29,150,31,16,31,16,30,26,31,26,30,26,29,222,31,255,31,168,31,130,31,42,31,161,31,170,31,74,31,74,30,36,31,245,31,144,31,133,31,251,31,71,31,196,31,196,30,49,31,44,31,194,31,3,31,148,31,250,31,53,31,53,30,53,31,113,31,154,31,154,30,151,31,151,30,128,31,200,31,147,31,24,31,24,30,211,31,211,30,211,29,79,31,105,31,114,31,114,30,114,29,114,28,7,31,113,31,211,31,211,30,233,31,24,31,24,30,227,31,31,31,192,31,166,31,166,30,141,31,121,31,97,31,125,31,32,31,243,31,244,31,131,31,9,31,36,31,78,31,145,31,145,30,216,31,72,31,86,31,11,31,11,30,168,31,168,30,53,31,197,31,34,31,75,31,75,30,120,31,79,31,79,30,221,31,83,31,207,31,115,31,122,31,231,31,172,31,82,31,237,31,244,31,244,30,29,31,132,31,132,30,52,31,24,31,82,31,48,31,40,31,252,31,117,31,20,31,210,31,94,31,137,31,137,30,115,31,37,31,71,31,151,31,234,31,4,31,41,31,230,31,161,31,161,30,7,31,65,31,149,31,43,31,6,31,102,31,186,31,245,31,127,31,98,31,21,31,17,31,37,31,156,31,203,31,203,30,43,31,196,31,84,31,151,31,96,31,71,31,70,31,70,30,5,31,22,31,206,31,6,31,6,30,95,31,95,30,36,31,48,31,15,31,158,31,156,31,247,31,116,31,70,31,82,31,82,30,82,29,8,31,249,31,249,30,249,29,174,31,221,31,139,31,246,31,119,31,137,31,180,31,47,31,193,31,107,31,171,31,50,31,220,31,220,30,190,31,190,30,152,31,140,31,123,31,123,30,66,31,81,31,110,31,108,31,85,31,44,31,227,31,146,31,137,31,137,30,193,31,14,31,14,30,14,29,149,31,167,31,171,31,5,31,5,30,71,31,22,31,170,31,174,31,84,31,98,31,189,31,189,30,165,31,246,31,55,31,152,31,152,30,152,29,162,31,54,31,245,31,245,30,245,29,245,28,48,31,135,31,135,30,135,29,151,31,70,31,81,31,88,31,160,31,13,31,237,31,178,31,170,31,170,30,100,31,103,31,92,31,5,31,5,30,5,29,96,31,227,31,227,30,183,31,192,31,192,30,126,31,126,30,126,29,108,31,108,30,108,29,38,31,173,31,61,31,61,30,242,31,83,31,83,30,83,29,83,28,206,31,97,31,98,31,236,31,163,31,102,31,254,31,254,30,19,31,153,31,137,31,214,31,214,30,96,31,1,31,1,30,196,31,206,31,91,31,133,31,133,30,202,31,117,31,173,31,138,31,146,31,182,31,233,31,243,31,30,31,170,31,74,31,189,31,187,31,187,30,214,31,40,31,21,31,84,31,255,31,145,31,40,31,244,31,119,31,21,31,21,30,209,31,129,31,93,31,207,31,101,31,101,30,127,31,110,31,255,31,254,31,7,31,9,31,181,31,49,31,88,31,230,31,230,30,230,29,230,28,88,31,88,30,88,29,32,31,111,31,47,31,183,31,133,31,101,31,100,31,76,31,203,31,111,31,63,31,159,31,196,31,56,31,219,31,89,31,174,31,174,30,119,31,41,31,74,31,15,31,204,31,220,31,21,31,145,31,201,31,44,31,44,30,44,29,192,31,211,31,211,30,59,31,129,31,129,30,129,31,58,31,140,31,234,31,234,30,234,29,94,31,52,31,195,31,180,31,77,31,95,31,17,31,130,31,164,31,164,30,164,29,66,31,80,31,132,31,12,31,222,31,244,31,114,31,114,30,94,31,177,31,64,31,64,30,211,31,173,31,110,31,145,31,44,31,202,31,218,31,218,30,30,31,140,31,212,31,212,30,212,29,254,31,254,30,28,31,118,31,118,30,118,29,118,28,63,31,194,31,20,31,172,31,216,31,217,31,151,31,151,30,48,31,24,31,21,31,230,31,215,31,205,31,155,31,55,31,222,31,222,30,234,31,234,30,234,29,52,31,108,31,6,31,37,31,176,31,122,31,232,31,189,31,222,31,171,31,221,31,243,31,226,31,160,31,21,31,86,31,13,31,29,31,16,31,28,31,28,30,227,31,227,30,227,29,13,31,13,30,109,31,97,31,126,31,1,31,1,30,81,31,208,31,209,31,209,30,95,31,88,31,88,30,44,31,155,31,13,31,45,31,45,30,162,31,1,31,1,30,155,31,191,31,191,30,93,31,195,31,180,31,34,31,19,31,19,30,31,31,125,31,177,31,210,31,57,31,206,31,6,31,52,31,171,31,171,30,171,29,171,28,32,31,42,31,120,31,167,31,103,31,91,31,76,31,247,31,99,31,38,31,20,31,109,31,109,30,163,31,163,30,154,31,36,31,24,31,24,30,239,31,204,31,172,31,6,31,251,31,251,30,173,31,252,31,41,31,163,31,32,31,196,31,246,31,87,31,52,31,52,30,52,29,69,31,81,31,107,31,168,31,186,31,37,31,76,31,65,31,12,31,231,31,231,30,231,29,139,31,90,31,136,31,82,31,22,31,10,31,135,31,120,31,53,31,117,31,117,30,117,29,116,31,145,31,178,31,33,31,203,31,111,31,111,30,246,31,171,31,191,31,191,30,28,31,191,31,191,30,8,31,8,30,43,31,31,31,31,30,114,31,114,30,153,31,53,31,250,31,250,30,250,29,250,28,196,31,62,31,230,31,148,31,27,31,27,30,27,29,27,28,234,31,212,31,178,31,60,31,35,31,14,31,54,31,37,31,194,31,194,30,150,31,150,30,97,31,83,31,168,31,206,31,222,31,56,31,56,30,98,31,87,31,61,31,181,31,181,30,181,29,91,31,117,31,29,31,128,31,223,31,223,30,223,29,198,31,138,31,124,31,53,31,53,30,53,29,170,31,68,31,10,31,48,31,48,30,189,31,250,31,28,31,120,31,58,31,58,30,203,31,203,30,38,31,38,31,87,31,113,31,255,31,255,30,32,31,32,30,12,31,182,31,72,31,170,31,254,31,32,31,90,31,198,31,94,31,94,30,196,31,248,31,5,31,5,30,255,31,62,31,161,31,5,31,83,31,90,31,126,31,126,30,205,31,1,31,112,31,218,31,62,31,223,31,255,31,120,31,128,31,128,30,239,31,229,31,71,31,41,31,41,30,250,31,208,31,129,31,80,31,179,31,245,31,245,30,155,31,9,31,164,31,120,31,176,31,12,31,70,31,172,31,77,31,144,31,144,30,230,31,215,31,215,30,215,29,197,31,250,31,250,30,25,31,199,31,35,31,29,31,168,31,186,31,202,31,56,31,200,31,218,31,28,31,28,30,59,31,59,30,55,31,55,30,77,31,135,31,167,31,149,31,122,31,220,31,219,31,77,31,77,30,77,29,77,28,77,27,139,31,137,31,137,30,137,29,206,31,206,30,124,31,26,31,52,31,52,30,52,29,52,28,36,31,35,31,136,31,136,30,102,31,240,31,73,31,211,31,97,31,42,31,42,30,42,29,20,31,35,31,35,30,202,31,76,31,240,31,90,31,90,30,136,31,67,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
