-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 192;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,252,0,105,0,146,0,192,0,14,0,152,0,247,0,140,0,58,0,97,0,130,0,39,0,247,0,17,0,69,0,235,0,144,0,38,0,0,0,223,0,228,0,109,0,61,0,117,0,50,0,0,0,0,0,184,0,165,0,52,0,77,0,199,0,58,0,7,0,126,0,17,0,90,0,199,0,230,0,19,0,144,0,101,0,36,0,54,0,225,0,162,0,165,0,0,0,103,0,0,0,241,0,254,0,121,0,47,0,74,0,172,0,35,0,161,0,93,0,130,0,99,0,101,0,7,0,0,0,26,0,29,0,89,0,84,0,201,0,26,0,156,0,211,0,203,0,56,0,169,0,0,0,241,0,0,0,19,0,13,0,96,0,158,0,0,0,229,0,47,0,93,0,72,0,0,0,0,0,35,0,10,0,192,0,251,0,9,0,251,0,50,0,87,0,127,0,200,0,129,0,0,0,0,0,0,0,0,0,31,0,221,0,30,0,74,0,0,0,0,0,84,0,187,0,117,0,174,0,224,0,206,0,167,0,94,0,162,0,210,0,0,0,17,0,142,0,0,0,191,0,68,0,56,0,41,0,118,0,180,0,0,0,198,0,127,0,93,0,38,0,0,0,0,0,125,0,78,0,248,0,251,0,233,0,0,0,12,0,9,0,84,0,0,0,195,0,142,0,147,0,153,0,0,0,69,0,172,0,4,0,35,0,0,0,197,0,251,0,178,0,46,0,160,0,84,0,74,0,0,0,0,0,52,0,0,0,140,0,56,0,52,0,94,0,130,0,253,0,242,0,228,0,150,0,49,0,0,0,207,0,26,0,33,0,0,0,55,0,236,0,112,0,247,0,170,0,105,0,146,0,212,0);
signal scenario_full  : scenario_type := (109,31,252,31,105,31,146,31,192,31,14,31,152,31,247,31,140,31,58,31,97,31,130,31,39,31,247,31,17,31,69,31,235,31,144,31,38,31,38,30,223,31,228,31,109,31,61,31,117,31,50,31,50,30,50,29,184,31,165,31,52,31,77,31,199,31,58,31,7,31,126,31,17,31,90,31,199,31,230,31,19,31,144,31,101,31,36,31,54,31,225,31,162,31,165,31,165,30,103,31,103,30,241,31,254,31,121,31,47,31,74,31,172,31,35,31,161,31,93,31,130,31,99,31,101,31,7,31,7,30,26,31,29,31,89,31,84,31,201,31,26,31,156,31,211,31,203,31,56,31,169,31,169,30,241,31,241,30,19,31,13,31,96,31,158,31,158,30,229,31,47,31,93,31,72,31,72,30,72,29,35,31,10,31,192,31,251,31,9,31,251,31,50,31,87,31,127,31,200,31,129,31,129,30,129,29,129,28,129,27,31,31,221,31,30,31,74,31,74,30,74,29,84,31,187,31,117,31,174,31,224,31,206,31,167,31,94,31,162,31,210,31,210,30,17,31,142,31,142,30,191,31,68,31,56,31,41,31,118,31,180,31,180,30,198,31,127,31,93,31,38,31,38,30,38,29,125,31,78,31,248,31,251,31,233,31,233,30,12,31,9,31,84,31,84,30,195,31,142,31,147,31,153,31,153,30,69,31,172,31,4,31,35,31,35,30,197,31,251,31,178,31,46,31,160,31,84,31,74,31,74,30,74,29,52,31,52,30,140,31,56,31,52,31,94,31,130,31,253,31,242,31,228,31,150,31,49,31,49,30,207,31,26,31,33,31,33,30,55,31,236,31,112,31,247,31,170,31,105,31,146,31,212,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
