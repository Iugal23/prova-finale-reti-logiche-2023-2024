-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_919 is
end project_tb_919;

architecture project_tb_arch_919 of project_tb_919 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 899;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,43,0,35,0,68,0,120,0,244,0,137,0,194,0,95,0,152,0,205,0,251,0,97,0,152,0,231,0,0,0,155,0,0,0,8,0,0,0,134,0,27,0,114,0,122,0,0,0,106,0,187,0,242,0,0,0,0,0,69,0,175,0,67,0,71,0,136,0,150,0,0,0,132,0,141,0,148,0,152,0,226,0,0,0,138,0,217,0,8,0,33,0,151,0,167,0,111,0,20,0,199,0,123,0,0,0,132,0,0,0,201,0,26,0,45,0,0,0,90,0,45,0,0,0,206,0,1,0,0,0,51,0,177,0,138,0,181,0,79,0,50,0,0,0,165,0,108,0,107,0,28,0,61,0,176,0,79,0,102,0,249,0,230,0,146,0,187,0,88,0,11,0,0,0,78,0,111,0,240,0,227,0,36,0,168,0,163,0,0,0,231,0,150,0,70,0,174,0,0,0,132,0,24,0,134,0,0,0,0,0,250,0,143,0,184,0,0,0,0,0,108,0,0,0,73,0,217,0,243,0,174,0,133,0,211,0,177,0,195,0,0,0,0,0,0,0,129,0,56,0,0,0,240,0,1,0,81,0,154,0,44,0,0,0,227,0,31,0,230,0,0,0,39,0,61,0,0,0,228,0,145,0,127,0,210,0,71,0,208,0,0,0,135,0,144,0,37,0,0,0,46,0,169,0,115,0,41,0,0,0,129,0,36,0,222,0,134,0,247,0,32,0,0,0,59,0,0,0,1,0,66,0,131,0,94,0,201,0,71,0,82,0,151,0,24,0,233,0,102,0,0,0,73,0,0,0,208,0,113,0,143,0,200,0,0,0,84,0,106,0,0,0,39,0,121,0,61,0,0,0,34,0,217,0,99,0,45,0,122,0,9,0,2,0,229,0,216,0,119,0,10,0,0,0,0,0,129,0,91,0,228,0,113,0,0,0,0,0,0,0,0,0,211,0,21,0,0,0,114,0,50,0,152,0,215,0,0,0,0,0,73,0,21,0,31,0,186,0,138,0,165,0,0,0,0,0,249,0,121,0,103,0,0,0,30,0,210,0,128,0,46,0,121,0,238,0,245,0,250,0,43,0,217,0,0,0,146,0,196,0,11,0,159,0,0,0,59,0,201,0,146,0,0,0,107,0,253,0,0,0,103,0,1,0,199,0,172,0,7,0,24,0,120,0,80,0,150,0,0,0,172,0,213,0,0,0,57,0,237,0,62,0,73,0,87,0,1,0,163,0,200,0,242,0,144,0,233,0,0,0,177,0,34,0,0,0,235,0,215,0,209,0,123,0,228,0,133,0,10,0,0,0,139,0,193,0,237,0,194,0,70,0,235,0,32,0,138,0,155,0,0,0,239,0,187,0,53,0,170,0,225,0,102,0,0,0,201,0,103,0,151,0,41,0,36,0,140,0,21,0,223,0,50,0,218,0,215,0,104,0,0,0,162,0,0,0,4,0,224,0,2,0,207,0,0,0,102,0,152,0,176,0,97,0,60,0,194,0,0,0,78,0,247,0,154,0,0,0,138,0,212,0,252,0,0,0,0,0,182,0,0,0,198,0,68,0,35,0,237,0,116,0,63,0,27,0,127,0,0,0,14,0,102,0,91,0,162,0,81,0,139,0,0,0,125,0,0,0,245,0,158,0,46,0,0,0,0,0,0,0,0,0,141,0,220,0,86,0,101,0,95,0,176,0,254,0,214,0,199,0,180,0,109,0,1,0,133,0,224,0,0,0,94,0,36,0,149,0,0,0,96,0,0,0,94,0,204,0,223,0,0,0,142,0,141,0,2,0,0,0,127,0,0,0,0,0,101,0,13,0,222,0,136,0,230,0,202,0,66,0,0,0,137,0,181,0,230,0,203,0,30,0,0,0,190,0,88,0,150,0,191,0,42,0,227,0,0,0,249,0,76,0,0,0,76,0,93,0,0,0,101,0,87,0,127,0,255,0,115,0,0,0,0,0,119,0,0,0,49,0,0,0,72,0,0,0,73,0,0,0,0,0,0,0,183,0,173,0,65,0,164,0,231,0,210,0,201,0,13,0,127,0,199,0,0,0,198,0,54,0,225,0,178,0,12,0,175,0,103,0,142,0,176,0,143,0,13,0,22,0,251,0,0,0,141,0,243,0,238,0,155,0,163,0,64,0,90,0,230,0,205,0,107,0,98,0,3,0,36,0,90,0,0,0,158,0,158,0,174,0,40,0,210,0,60,0,61,0,207,0,0,0,47,0,156,0,177,0,64,0,111,0,0,0,228,0,232,0,138,0,234,0,146,0,17,0,0,0,0,0,0,0,0,0,217,0,240,0,153,0,71,0,74,0,119,0,0,0,120,0,54,0,236,0,45,0,0,0,0,0,56,0,0,0,21,0,148,0,103,0,202,0,11,0,168,0,94,0,102,0,191,0,33,0,216,0,61,0,241,0,188,0,168,0,193,0,17,0,0,0,13,0,0,0,0,0,244,0,24,0,237,0,55,0,50,0,178,0,0,0,202,0,109,0,0,0,215,0,63,0,24,0,0,0,0,0,244,0,54,0,107,0,231,0,39,0,15,0,203,0,134,0,0,0,120,0,58,0,16,0,25,0,0,0,182,0,154,0,78,0,0,0,0,0,115,0,19,0,0,0,219,0,0,0,237,0,14,0,31,0,0,0,49,0,28,0,168,0,0,0,136,0,242,0,153,0,220,0,0,0,108,0,203,0,89,0,201,0,41,0,0,0,221,0,0,0,151,0,0,0,157,0,0,0,18,0,0,0,125,0,207,0,95,0,0,0,180,0,67,0,29,0,96,0,99,0,238,0,225,0,50,0,33,0,0,0,37,0,20,0,106,0,13,0,21,0,121,0,239,0,250,0,254,0,200,0,0,0,191,0,86,0,111,0,18,0,101,0,124,0,197,0,0,0,200,0,37,0,0,0,158,0,19,0,0,0,24,0,51,0,64,0,212,0,116,0,133,0,132,0,160,0,0,0,155,0,9,0,87,0,11,0,198,0,207,0,180,0,202,0,89,0,187,0,173,0,92,0,71,0,33,0,185,0,88,0,188,0,0,0,98,0,244,0,0,0,0,0,28,0,0,0,0,0,6,0,1,0,0,0,111,0,248,0,77,0,30,0,0,0,0,0,193,0,155,0,0,0,2,0,152,0,0,0,124,0,75,0,0,0,0,0,54,0,178,0,110,0,53,0,95,0,0,0,87,0,72,0,186,0,106,0,0,0,0,0,0,0,243,0,119,0,91,0,92,0,0,0,209,0,0,0,0,0,59,0,6,0,148,0,191,0,148,0,34,0,0,0,30,0,202,0,65,0,149,0,67,0,0,0,0,0,85,0,228,0,157,0,246,0,119,0,203,0,181,0,0,0,93,0,17,0,148,0,224,0,87,0,32,0,178,0,239,0,116,0,237,0,71,0,98,0,216,0,28,0,147,0,78,0,137,0,192,0,134,0,220,0,0,0,21,0,0,0,0,0,39,0,182,0,134,0,153,0,69,0,103,0,147,0,0,0,82,0,238,0,203,0,66,0,28,0,0,0,11,0,240,0,231,0,184,0,216,0,151,0,0,0,0,0,41,0,30,0,81,0,208,0,0,0,0,0,172,0,0,0,200,0,14,0,110,0,0,0,0,0,156,0,0,0,65,0,241,0,214,0,88,0,0,0,3,0,62,0,242,0,26,0,91,0,19,0,72,0,0,0,0,0,158,0,194,0,77,0,179,0,217,0,27,0,244,0,192,0,103,0,155,0,234,0,187,0,0,0,245,0,124,0,203,0,158,0,0,0,44,0,0,0,249,0,66,0,106,0,170,0,82,0,76,0,5,0,0,0,205,0,100,0,177,0,122,0,161,0,107,0,40,0,143,0,170,0,125,0,150,0,73,0,75,0,0,0,44,0,10,0,140,0,0,0,224,0,13,0,138,0,147,0,0,0,0,0,1,0,162,0,53,0,40,0,136,0,55,0,0,0,189,0,155,0,254,0,121,0,218,0,28,0,20,0,222,0,0,0,156,0,135,0,175,0,0,0,45,0,146,0);
signal scenario_full  : scenario_type := (201,31,43,31,35,31,68,31,120,31,244,31,137,31,194,31,95,31,152,31,205,31,251,31,97,31,152,31,231,31,231,30,155,31,155,30,8,31,8,30,134,31,27,31,114,31,122,31,122,30,106,31,187,31,242,31,242,30,242,29,69,31,175,31,67,31,71,31,136,31,150,31,150,30,132,31,141,31,148,31,152,31,226,31,226,30,138,31,217,31,8,31,33,31,151,31,167,31,111,31,20,31,199,31,123,31,123,30,132,31,132,30,201,31,26,31,45,31,45,30,90,31,45,31,45,30,206,31,1,31,1,30,51,31,177,31,138,31,181,31,79,31,50,31,50,30,165,31,108,31,107,31,28,31,61,31,176,31,79,31,102,31,249,31,230,31,146,31,187,31,88,31,11,31,11,30,78,31,111,31,240,31,227,31,36,31,168,31,163,31,163,30,231,31,150,31,70,31,174,31,174,30,132,31,24,31,134,31,134,30,134,29,250,31,143,31,184,31,184,30,184,29,108,31,108,30,73,31,217,31,243,31,174,31,133,31,211,31,177,31,195,31,195,30,195,29,195,28,129,31,56,31,56,30,240,31,1,31,81,31,154,31,44,31,44,30,227,31,31,31,230,31,230,30,39,31,61,31,61,30,228,31,145,31,127,31,210,31,71,31,208,31,208,30,135,31,144,31,37,31,37,30,46,31,169,31,115,31,41,31,41,30,129,31,36,31,222,31,134,31,247,31,32,31,32,30,59,31,59,30,1,31,66,31,131,31,94,31,201,31,71,31,82,31,151,31,24,31,233,31,102,31,102,30,73,31,73,30,208,31,113,31,143,31,200,31,200,30,84,31,106,31,106,30,39,31,121,31,61,31,61,30,34,31,217,31,99,31,45,31,122,31,9,31,2,31,229,31,216,31,119,31,10,31,10,30,10,29,129,31,91,31,228,31,113,31,113,30,113,29,113,28,113,27,211,31,21,31,21,30,114,31,50,31,152,31,215,31,215,30,215,29,73,31,21,31,31,31,186,31,138,31,165,31,165,30,165,29,249,31,121,31,103,31,103,30,30,31,210,31,128,31,46,31,121,31,238,31,245,31,250,31,43,31,217,31,217,30,146,31,196,31,11,31,159,31,159,30,59,31,201,31,146,31,146,30,107,31,253,31,253,30,103,31,1,31,199,31,172,31,7,31,24,31,120,31,80,31,150,31,150,30,172,31,213,31,213,30,57,31,237,31,62,31,73,31,87,31,1,31,163,31,200,31,242,31,144,31,233,31,233,30,177,31,34,31,34,30,235,31,215,31,209,31,123,31,228,31,133,31,10,31,10,30,139,31,193,31,237,31,194,31,70,31,235,31,32,31,138,31,155,31,155,30,239,31,187,31,53,31,170,31,225,31,102,31,102,30,201,31,103,31,151,31,41,31,36,31,140,31,21,31,223,31,50,31,218,31,215,31,104,31,104,30,162,31,162,30,4,31,224,31,2,31,207,31,207,30,102,31,152,31,176,31,97,31,60,31,194,31,194,30,78,31,247,31,154,31,154,30,138,31,212,31,252,31,252,30,252,29,182,31,182,30,198,31,68,31,35,31,237,31,116,31,63,31,27,31,127,31,127,30,14,31,102,31,91,31,162,31,81,31,139,31,139,30,125,31,125,30,245,31,158,31,46,31,46,30,46,29,46,28,46,27,141,31,220,31,86,31,101,31,95,31,176,31,254,31,214,31,199,31,180,31,109,31,1,31,133,31,224,31,224,30,94,31,36,31,149,31,149,30,96,31,96,30,94,31,204,31,223,31,223,30,142,31,141,31,2,31,2,30,127,31,127,30,127,29,101,31,13,31,222,31,136,31,230,31,202,31,66,31,66,30,137,31,181,31,230,31,203,31,30,31,30,30,190,31,88,31,150,31,191,31,42,31,227,31,227,30,249,31,76,31,76,30,76,31,93,31,93,30,101,31,87,31,127,31,255,31,115,31,115,30,115,29,119,31,119,30,49,31,49,30,72,31,72,30,73,31,73,30,73,29,73,28,183,31,173,31,65,31,164,31,231,31,210,31,201,31,13,31,127,31,199,31,199,30,198,31,54,31,225,31,178,31,12,31,175,31,103,31,142,31,176,31,143,31,13,31,22,31,251,31,251,30,141,31,243,31,238,31,155,31,163,31,64,31,90,31,230,31,205,31,107,31,98,31,3,31,36,31,90,31,90,30,158,31,158,31,174,31,40,31,210,31,60,31,61,31,207,31,207,30,47,31,156,31,177,31,64,31,111,31,111,30,228,31,232,31,138,31,234,31,146,31,17,31,17,30,17,29,17,28,17,27,217,31,240,31,153,31,71,31,74,31,119,31,119,30,120,31,54,31,236,31,45,31,45,30,45,29,56,31,56,30,21,31,148,31,103,31,202,31,11,31,168,31,94,31,102,31,191,31,33,31,216,31,61,31,241,31,188,31,168,31,193,31,17,31,17,30,13,31,13,30,13,29,244,31,24,31,237,31,55,31,50,31,178,31,178,30,202,31,109,31,109,30,215,31,63,31,24,31,24,30,24,29,244,31,54,31,107,31,231,31,39,31,15,31,203,31,134,31,134,30,120,31,58,31,16,31,25,31,25,30,182,31,154,31,78,31,78,30,78,29,115,31,19,31,19,30,219,31,219,30,237,31,14,31,31,31,31,30,49,31,28,31,168,31,168,30,136,31,242,31,153,31,220,31,220,30,108,31,203,31,89,31,201,31,41,31,41,30,221,31,221,30,151,31,151,30,157,31,157,30,18,31,18,30,125,31,207,31,95,31,95,30,180,31,67,31,29,31,96,31,99,31,238,31,225,31,50,31,33,31,33,30,37,31,20,31,106,31,13,31,21,31,121,31,239,31,250,31,254,31,200,31,200,30,191,31,86,31,111,31,18,31,101,31,124,31,197,31,197,30,200,31,37,31,37,30,158,31,19,31,19,30,24,31,51,31,64,31,212,31,116,31,133,31,132,31,160,31,160,30,155,31,9,31,87,31,11,31,198,31,207,31,180,31,202,31,89,31,187,31,173,31,92,31,71,31,33,31,185,31,88,31,188,31,188,30,98,31,244,31,244,30,244,29,28,31,28,30,28,29,6,31,1,31,1,30,111,31,248,31,77,31,30,31,30,30,30,29,193,31,155,31,155,30,2,31,152,31,152,30,124,31,75,31,75,30,75,29,54,31,178,31,110,31,53,31,95,31,95,30,87,31,72,31,186,31,106,31,106,30,106,29,106,28,243,31,119,31,91,31,92,31,92,30,209,31,209,30,209,29,59,31,6,31,148,31,191,31,148,31,34,31,34,30,30,31,202,31,65,31,149,31,67,31,67,30,67,29,85,31,228,31,157,31,246,31,119,31,203,31,181,31,181,30,93,31,17,31,148,31,224,31,87,31,32,31,178,31,239,31,116,31,237,31,71,31,98,31,216,31,28,31,147,31,78,31,137,31,192,31,134,31,220,31,220,30,21,31,21,30,21,29,39,31,182,31,134,31,153,31,69,31,103,31,147,31,147,30,82,31,238,31,203,31,66,31,28,31,28,30,11,31,240,31,231,31,184,31,216,31,151,31,151,30,151,29,41,31,30,31,81,31,208,31,208,30,208,29,172,31,172,30,200,31,14,31,110,31,110,30,110,29,156,31,156,30,65,31,241,31,214,31,88,31,88,30,3,31,62,31,242,31,26,31,91,31,19,31,72,31,72,30,72,29,158,31,194,31,77,31,179,31,217,31,27,31,244,31,192,31,103,31,155,31,234,31,187,31,187,30,245,31,124,31,203,31,158,31,158,30,44,31,44,30,249,31,66,31,106,31,170,31,82,31,76,31,5,31,5,30,205,31,100,31,177,31,122,31,161,31,107,31,40,31,143,31,170,31,125,31,150,31,73,31,75,31,75,30,44,31,10,31,140,31,140,30,224,31,13,31,138,31,147,31,147,30,147,29,1,31,162,31,53,31,40,31,136,31,55,31,55,30,189,31,155,31,254,31,121,31,218,31,28,31,20,31,222,31,222,30,156,31,135,31,175,31,175,30,45,31,146,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
