-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_336 is
end project_tb_336;

architecture project_tb_arch_336 of project_tb_336 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 628;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,44,0,0,0,64,0,16,0,22,0,29,0,118,0,61,0,140,0,93,0,154,0,92,0,239,0,244,0,0,0,117,0,0,0,171,0,151,0,187,0,203,0,137,0,152,0,244,0,41,0,94,0,52,0,162,0,157,0,238,0,81,0,177,0,251,0,0,0,137,0,115,0,228,0,126,0,191,0,52,0,133,0,172,0,0,0,231,0,95,0,53,0,130,0,0,0,0,0,49,0,155,0,76,0,153,0,72,0,109,0,29,0,83,0,221,0,0,0,242,0,45,0,0,0,162,0,0,0,241,0,82,0,220,0,182,0,16,0,67,0,0,0,0,0,164,0,168,0,53,0,0,0,20,0,223,0,142,0,0,0,39,0,119,0,0,0,57,0,20,0,6,0,197,0,38,0,192,0,128,0,76,0,101,0,102,0,231,0,6,0,89,0,249,0,192,0,165,0,176,0,0,0,212,0,0,0,235,0,118,0,222,0,0,0,0,0,231,0,176,0,211,0,0,0,0,0,127,0,171,0,238,0,202,0,94,0,0,0,76,0,9,0,33,0,207,0,136,0,0,0,195,0,0,0,84,0,124,0,180,0,61,0,98,0,233,0,56,0,32,0,211,0,148,0,0,0,0,0,139,0,214,0,112,0,206,0,21,0,47,0,58,0,154,0,118,0,107,0,0,0,53,0,217,0,30,0,166,0,193,0,0,0,0,0,139,0,87,0,173,0,113,0,140,0,241,0,145,0,8,0,126,0,192,0,186,0,0,0,1,0,128,0,77,0,125,0,137,0,46,0,139,0,0,0,0,0,100,0,14,0,0,0,224,0,144,0,75,0,17,0,114,0,11,0,180,0,241,0,0,0,184,0,254,0,40,0,142,0,5,0,0,0,194,0,155,0,83,0,102,0,192,0,30,0,199,0,176,0,48,0,145,0,0,0,17,0,146,0,128,0,60,0,3,0,113,0,146,0,0,0,246,0,202,0,216,0,88,0,109,0,33,0,0,0,0,0,219,0,40,0,0,0,72,0,215,0,228,0,0,0,164,0,0,0,0,0,69,0,55,0,251,0,0,0,178,0,236,0,127,0,0,0,40,0,202,0,89,0,190,0,96,0,127,0,165,0,27,0,238,0,86,0,81,0,189,0,117,0,0,0,0,0,53,0,0,0,125,0,156,0,155,0,230,0,211,0,58,0,65,0,53,0,20,0,45,0,93,0,33,0,118,0,0,0,71,0,252,0,52,0,100,0,195,0,211,0,131,0,2,0,25,0,84,0,20,0,233,0,152,0,236,0,186,0,218,0,0,0,80,0,119,0,168,0,70,0,1,0,128,0,179,0,35,0,224,0,92,0,61,0,130,0,103,0,226,0,44,0,12,0,63,0,194,0,0,0,249,0,180,0,170,0,24,0,187,0,0,0,59,0,151,0,0,0,128,0,222,0,71,0,156,0,163,0,109,0,0,0,0,0,189,0,0,0,145,0,122,0,78,0,0,0,73,0,7,0,0,0,117,0,0,0,45,0,125,0,0,0,163,0,23,0,186,0,232,0,0,0,0,0,172,0,181,0,122,0,210,0,57,0,109,0,0,0,0,0,177,0,25,0,150,0,220,0,0,0,35,0,0,0,0,0,237,0,170,0,0,0,8,0,224,0,178,0,0,0,59,0,196,0,223,0,95,0,156,0,117,0,23,0,0,0,26,0,198,0,216,0,121,0,202,0,214,0,49,0,184,0,157,0,169,0,0,0,224,0,13,0,192,0,117,0,9,0,191,0,162,0,138,0,59,0,243,0,118,0,175,0,135,0,248,0,177,0,10,0,196,0,0,0,36,0,229,0,84,0,109,0,215,0,117,0,181,0,251,0,0,0,208,0,128,0,122,0,34,0,168,0,5,0,0,0,0,0,98,0,154,0,213,0,164,0,0,0,114,0,149,0,107,0,0,0,119,0,12,0,165,0,0,0,106,0,6,0,0,0,211,0,79,0,0,0,0,0,0,0,118,0,57,0,4,0,0,0,213,0,0,0,212,0,70,0,82,0,138,0,228,0,158,0,240,0,0,0,0,0,0,0,219,0,83,0,107,0,0,0,243,0,160,0,113,0,92,0,0,0,255,0,0,0,104,0,79,0,199,0,102,0,5,0,223,0,74,0,166,0,0,0,0,0,113,0,39,0,160,0,25,0,0,0,0,0,0,0,151,0,105,0,22,0,184,0,71,0,139,0,64,0,203,0,59,0,22,0,24,0,72,0,171,0,0,0,221,0,0,0,43,0,21,0,138,0,96,0,97,0,238,0,66,0,206,0,66,0,32,0,172,0,140,0,128,0,124,0,213,0,144,0,170,0,0,0,159,0,37,0,143,0,253,0,187,0,10,0,57,0,207,0,86,0,218,0,253,0,209,0,236,0,21,0,158,0,182,0,0,0,212,0,241,0,121,0,40,0,210,0,1,0,96,0,0,0,156,0,59,0,0,0,0,0,37,0,22,0,0,0,182,0,215,0,235,0,108,0,147,0,154,0,36,0,108,0,113,0,0,0,0,0,153,0,163,0,172,0,2,0,0,0,0,0,230,0,44,0,77,0,166,0,246,0,71,0,164,0,3,0,219,0,70,0,115,0,11,0,30,0,148,0,0,0,7,0,96,0,204,0,58,0,160,0,253,0,22,0,200,0,158,0,162,0,75,0,159,0,250,0,104,0,106,0,60,0,167,0,186,0,76,0,0,0,26,0,0,0,245,0,18,0,187,0,0,0,230,0,0,0,40,0,96,0,91,0,27,0,0,0,0,0,0,0,115,0,88,0,108,0,172,0,118,0,56,0,100,0);
signal scenario_full  : scenario_type := (83,31,44,31,44,30,64,31,16,31,22,31,29,31,118,31,61,31,140,31,93,31,154,31,92,31,239,31,244,31,244,30,117,31,117,30,171,31,151,31,187,31,203,31,137,31,152,31,244,31,41,31,94,31,52,31,162,31,157,31,238,31,81,31,177,31,251,31,251,30,137,31,115,31,228,31,126,31,191,31,52,31,133,31,172,31,172,30,231,31,95,31,53,31,130,31,130,30,130,29,49,31,155,31,76,31,153,31,72,31,109,31,29,31,83,31,221,31,221,30,242,31,45,31,45,30,162,31,162,30,241,31,82,31,220,31,182,31,16,31,67,31,67,30,67,29,164,31,168,31,53,31,53,30,20,31,223,31,142,31,142,30,39,31,119,31,119,30,57,31,20,31,6,31,197,31,38,31,192,31,128,31,76,31,101,31,102,31,231,31,6,31,89,31,249,31,192,31,165,31,176,31,176,30,212,31,212,30,235,31,118,31,222,31,222,30,222,29,231,31,176,31,211,31,211,30,211,29,127,31,171,31,238,31,202,31,94,31,94,30,76,31,9,31,33,31,207,31,136,31,136,30,195,31,195,30,84,31,124,31,180,31,61,31,98,31,233,31,56,31,32,31,211,31,148,31,148,30,148,29,139,31,214,31,112,31,206,31,21,31,47,31,58,31,154,31,118,31,107,31,107,30,53,31,217,31,30,31,166,31,193,31,193,30,193,29,139,31,87,31,173,31,113,31,140,31,241,31,145,31,8,31,126,31,192,31,186,31,186,30,1,31,128,31,77,31,125,31,137,31,46,31,139,31,139,30,139,29,100,31,14,31,14,30,224,31,144,31,75,31,17,31,114,31,11,31,180,31,241,31,241,30,184,31,254,31,40,31,142,31,5,31,5,30,194,31,155,31,83,31,102,31,192,31,30,31,199,31,176,31,48,31,145,31,145,30,17,31,146,31,128,31,60,31,3,31,113,31,146,31,146,30,246,31,202,31,216,31,88,31,109,31,33,31,33,30,33,29,219,31,40,31,40,30,72,31,215,31,228,31,228,30,164,31,164,30,164,29,69,31,55,31,251,31,251,30,178,31,236,31,127,31,127,30,40,31,202,31,89,31,190,31,96,31,127,31,165,31,27,31,238,31,86,31,81,31,189,31,117,31,117,30,117,29,53,31,53,30,125,31,156,31,155,31,230,31,211,31,58,31,65,31,53,31,20,31,45,31,93,31,33,31,118,31,118,30,71,31,252,31,52,31,100,31,195,31,211,31,131,31,2,31,25,31,84,31,20,31,233,31,152,31,236,31,186,31,218,31,218,30,80,31,119,31,168,31,70,31,1,31,128,31,179,31,35,31,224,31,92,31,61,31,130,31,103,31,226,31,44,31,12,31,63,31,194,31,194,30,249,31,180,31,170,31,24,31,187,31,187,30,59,31,151,31,151,30,128,31,222,31,71,31,156,31,163,31,109,31,109,30,109,29,189,31,189,30,145,31,122,31,78,31,78,30,73,31,7,31,7,30,117,31,117,30,45,31,125,31,125,30,163,31,23,31,186,31,232,31,232,30,232,29,172,31,181,31,122,31,210,31,57,31,109,31,109,30,109,29,177,31,25,31,150,31,220,31,220,30,35,31,35,30,35,29,237,31,170,31,170,30,8,31,224,31,178,31,178,30,59,31,196,31,223,31,95,31,156,31,117,31,23,31,23,30,26,31,198,31,216,31,121,31,202,31,214,31,49,31,184,31,157,31,169,31,169,30,224,31,13,31,192,31,117,31,9,31,191,31,162,31,138,31,59,31,243,31,118,31,175,31,135,31,248,31,177,31,10,31,196,31,196,30,36,31,229,31,84,31,109,31,215,31,117,31,181,31,251,31,251,30,208,31,128,31,122,31,34,31,168,31,5,31,5,30,5,29,98,31,154,31,213,31,164,31,164,30,114,31,149,31,107,31,107,30,119,31,12,31,165,31,165,30,106,31,6,31,6,30,211,31,79,31,79,30,79,29,79,28,118,31,57,31,4,31,4,30,213,31,213,30,212,31,70,31,82,31,138,31,228,31,158,31,240,31,240,30,240,29,240,28,219,31,83,31,107,31,107,30,243,31,160,31,113,31,92,31,92,30,255,31,255,30,104,31,79,31,199,31,102,31,5,31,223,31,74,31,166,31,166,30,166,29,113,31,39,31,160,31,25,31,25,30,25,29,25,28,151,31,105,31,22,31,184,31,71,31,139,31,64,31,203,31,59,31,22,31,24,31,72,31,171,31,171,30,221,31,221,30,43,31,21,31,138,31,96,31,97,31,238,31,66,31,206,31,66,31,32,31,172,31,140,31,128,31,124,31,213,31,144,31,170,31,170,30,159,31,37,31,143,31,253,31,187,31,10,31,57,31,207,31,86,31,218,31,253,31,209,31,236,31,21,31,158,31,182,31,182,30,212,31,241,31,121,31,40,31,210,31,1,31,96,31,96,30,156,31,59,31,59,30,59,29,37,31,22,31,22,30,182,31,215,31,235,31,108,31,147,31,154,31,36,31,108,31,113,31,113,30,113,29,153,31,163,31,172,31,2,31,2,30,2,29,230,31,44,31,77,31,166,31,246,31,71,31,164,31,3,31,219,31,70,31,115,31,11,31,30,31,148,31,148,30,7,31,96,31,204,31,58,31,160,31,253,31,22,31,200,31,158,31,162,31,75,31,159,31,250,31,104,31,106,31,60,31,167,31,186,31,76,31,76,30,26,31,26,30,245,31,18,31,187,31,187,30,230,31,230,30,40,31,96,31,91,31,27,31,27,30,27,29,27,28,115,31,88,31,108,31,172,31,118,31,56,31,100,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
