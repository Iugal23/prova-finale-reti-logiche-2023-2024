-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 766;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (13,0,0,0,0,0,56,0,197,0,100,0,211,0,227,0,238,0,0,0,0,0,0,0,31,0,148,0,0,0,166,0,0,0,185,0,248,0,66,0,126,0,83,0,100,0,147,0,226,0,0,0,95,0,253,0,46,0,67,0,178,0,95,0,140,0,175,0,74,0,149,0,202,0,5,0,64,0,168,0,173,0,17,0,194,0,96,0,226,0,0,0,229,0,88,0,110,0,34,0,229,0,138,0,85,0,129,0,172,0,0,0,0,0,194,0,4,0,248,0,25,0,159,0,0,0,66,0,66,0,0,0,214,0,163,0,172,0,9,0,75,0,181,0,61,0,8,0,0,0,53,0,16,0,30,0,0,0,0,0,110,0,103,0,17,0,168,0,170,0,41,0,0,0,169,0,210,0,248,0,142,0,144,0,80,0,164,0,186,0,136,0,37,0,0,0,237,0,0,0,20,0,71,0,14,0,227,0,169,0,58,0,194,0,131,0,244,0,0,0,198,0,241,0,101,0,155,0,122,0,5,0,67,0,241,0,186,0,126,0,91,0,202,0,123,0,190,0,132,0,0,0,195,0,199,0,158,0,181,0,105,0,251,0,178,0,249,0,0,0,242,0,71,0,170,0,26,0,56,0,207,0,138,0,64,0,50,0,84,0,184,0,0,0,0,0,92,0,163,0,21,0,18,0,37,0,0,0,119,0,101,0,58,0,68,0,54,0,166,0,251,0,115,0,247,0,36,0,0,0,10,0,11,0,0,0,195,0,222,0,0,0,0,0,87,0,53,0,100,0,25,0,72,0,0,0,251,0,23,0,113,0,120,0,0,0,0,0,0,0,165,0,144,0,89,0,197,0,125,0,55,0,73,0,249,0,145,0,122,0,0,0,130,0,169,0,27,0,53,0,102,0,15,0,0,0,129,0,61,0,65,0,218,0,0,0,142,0,0,0,180,0,138,0,145,0,244,0,0,0,0,0,30,0,205,0,219,0,119,0,0,0,197,0,238,0,74,0,239,0,222,0,202,0,68,0,145,0,0,0,94,0,245,0,3,0,150,0,178,0,62,0,0,0,122,0,77,0,0,0,0,0,92,0,45,0,33,0,0,0,0,0,0,0,151,0,236,0,244,0,108,0,193,0,177,0,0,0,77,0,0,0,178,0,40,0,165,0,168,0,0,0,36,0,104,0,0,0,141,0,219,0,37,0,186,0,184,0,81,0,185,0,0,0,44,0,5,0,75,0,0,0,131,0,146,0,0,0,0,0,248,0,213,0,103,0,160,0,209,0,150,0,0,0,58,0,215,0,96,0,208,0,14,0,60,0,45,0,0,0,204,0,94,0,50,0,3,0,113,0,181,0,0,0,210,0,91,0,105,0,0,0,132,0,213,0,204,0,88,0,232,0,0,0,206,0,0,0,17,0,84,0,0,0,193,0,55,0,38,0,141,0,48,0,189,0,207,0,245,0,0,0,0,0,0,0,19,0,77,0,0,0,242,0,176,0,47,0,80,0,41,0,100,0,228,0,0,0,0,0,202,0,59,0,113,0,48,0,0,0,27,0,3,0,251,0,230,0,7,0,170,0,27,0,1,0,105,0,253,0,82,0,0,0,0,0,62,0,0,0,68,0,141,0,244,0,75,0,7,0,0,0,230,0,74,0,124,0,248,0,0,0,223,0,0,0,102,0,213,0,230,0,17,0,136,0,44,0,124,0,0,0,225,0,143,0,0,0,0,0,0,0,140,0,0,0,20,0,210,0,241,0,125,0,237,0,79,0,0,0,15,0,198,0,37,0,240,0,0,0,65,0,180,0,58,0,211,0,0,0,191,0,168,0,171,0,249,0,21,0,71,0,0,0,58,0,216,0,242,0,36,0,136,0,115,0,0,0,0,0,175,0,0,0,8,0,72,0,56,0,60,0,0,0,237,0,0,0,71,0,141,0,0,0,0,0,200,0,0,0,9,0,99,0,241,0,249,0,242,0,110,0,34,0,145,0,102,0,246,0,19,0,172,0,0,0,181,0,77,0,0,0,242,0,193,0,0,0,67,0,116,0,114,0,186,0,21,0,196,0,52,0,55,0,0,0,40,0,15,0,237,0,206,0,50,0,227,0,160,0,227,0,220,0,198,0,88,0,236,0,135,0,0,0,110,0,78,0,19,0,191,0,13,0,110,0,171,0,223,0,154,0,206,0,0,0,1,0,179,0,233,0,74,0,0,0,187,0,107,0,85,0,32,0,79,0,169,0,0,0,3,0,83,0,106,0,0,0,138,0,12,0,0,0,116,0,197,0,196,0,131,0,85,0,137,0,10,0,129,0,195,0,32,0,52,0,185,0,122,0,75,0,143,0,165,0,0,0,41,0,215,0,213,0,115,0,62,0,122,0,0,0,47,0,154,0,0,0,253,0,162,0,103,0,26,0,0,0,255,0,0,0,102,0,27,0,200,0,70,0,165,0,240,0,59,0,0,0,5,0,0,0,71,0,0,0,74,0,2,0,114,0,253,0,66,0,4,0,192,0,227,0,240,0,176,0,185,0,52,0,0,0,0,0,0,0,45,0,20,0,164,0,224,0,108,0,54,0,241,0,60,0,118,0,17,0,0,0,168,0,21,0,99,0,96,0,11,0,61,0,2,0,248,0,105,0,104,0,194,0,103,0,0,0,73,0,216,0,226,0,215,0,27,0,2,0,0,0,203,0,110,0,190,0,24,0,133,0,56,0,45,0,174,0,0,0,118,0,108,0,158,0,61,0,125,0,167,0,38,0,152,0,202,0,0,0,238,0,0,0,222,0,5,0,96,0,0,0,21,0,140,0,110,0,32,0,0,0,111,0,225,0,0,0,104,0,0,0,0,0,67,0,0,0,131,0,150,0,138,0,54,0,100,0,125,0,28,0,85,0,190,0,0,0,1,0,118,0,177,0,91,0,208,0,252,0,0,0,230,0,130,0,206,0,87,0,0,0,231,0,112,0,130,0,0,0,1,0,120,0,0,0,0,0,6,0,0,0,0,0,10,0,194,0,148,0,44,0,139,0,218,0,204,0,0,0,31,0,140,0,20,0,0,0,130,0,185,0,55,0,0,0,194,0,84,0,69,0,0,0,247,0,189,0,230,0,219,0,142,0,197,0,153,0,239,0,151,0,159,0,214,0,133,0,68,0,138,0,0,0,135,0,0,0,239,0,146,0,250,0,79,0,0,0,120,0,57,0,22,0,242,0,0,0,224,0,20,0,58,0,148,0,93,0,180,0,218,0,109,0,0,0,15,0,0,0,45,0,0,0,249,0,16,0,248,0,125,0,136,0,38,0,55,0,190,0,45,0,0,0,174,0,24,0,104,0,143,0,173,0,18,0,0,0,0,0,0,0,248,0,168,0,255,0,203,0,113,0,222,0,98,0,43,0,247,0,0,0,0,0,98,0,64,0,249,0,95,0,0,0,46,0);
signal scenario_full  : scenario_type := (13,31,13,30,13,29,56,31,197,31,100,31,211,31,227,31,238,31,238,30,238,29,238,28,31,31,148,31,148,30,166,31,166,30,185,31,248,31,66,31,126,31,83,31,100,31,147,31,226,31,226,30,95,31,253,31,46,31,67,31,178,31,95,31,140,31,175,31,74,31,149,31,202,31,5,31,64,31,168,31,173,31,17,31,194,31,96,31,226,31,226,30,229,31,88,31,110,31,34,31,229,31,138,31,85,31,129,31,172,31,172,30,172,29,194,31,4,31,248,31,25,31,159,31,159,30,66,31,66,31,66,30,214,31,163,31,172,31,9,31,75,31,181,31,61,31,8,31,8,30,53,31,16,31,30,31,30,30,30,29,110,31,103,31,17,31,168,31,170,31,41,31,41,30,169,31,210,31,248,31,142,31,144,31,80,31,164,31,186,31,136,31,37,31,37,30,237,31,237,30,20,31,71,31,14,31,227,31,169,31,58,31,194,31,131,31,244,31,244,30,198,31,241,31,101,31,155,31,122,31,5,31,67,31,241,31,186,31,126,31,91,31,202,31,123,31,190,31,132,31,132,30,195,31,199,31,158,31,181,31,105,31,251,31,178,31,249,31,249,30,242,31,71,31,170,31,26,31,56,31,207,31,138,31,64,31,50,31,84,31,184,31,184,30,184,29,92,31,163,31,21,31,18,31,37,31,37,30,119,31,101,31,58,31,68,31,54,31,166,31,251,31,115,31,247,31,36,31,36,30,10,31,11,31,11,30,195,31,222,31,222,30,222,29,87,31,53,31,100,31,25,31,72,31,72,30,251,31,23,31,113,31,120,31,120,30,120,29,120,28,165,31,144,31,89,31,197,31,125,31,55,31,73,31,249,31,145,31,122,31,122,30,130,31,169,31,27,31,53,31,102,31,15,31,15,30,129,31,61,31,65,31,218,31,218,30,142,31,142,30,180,31,138,31,145,31,244,31,244,30,244,29,30,31,205,31,219,31,119,31,119,30,197,31,238,31,74,31,239,31,222,31,202,31,68,31,145,31,145,30,94,31,245,31,3,31,150,31,178,31,62,31,62,30,122,31,77,31,77,30,77,29,92,31,45,31,33,31,33,30,33,29,33,28,151,31,236,31,244,31,108,31,193,31,177,31,177,30,77,31,77,30,178,31,40,31,165,31,168,31,168,30,36,31,104,31,104,30,141,31,219,31,37,31,186,31,184,31,81,31,185,31,185,30,44,31,5,31,75,31,75,30,131,31,146,31,146,30,146,29,248,31,213,31,103,31,160,31,209,31,150,31,150,30,58,31,215,31,96,31,208,31,14,31,60,31,45,31,45,30,204,31,94,31,50,31,3,31,113,31,181,31,181,30,210,31,91,31,105,31,105,30,132,31,213,31,204,31,88,31,232,31,232,30,206,31,206,30,17,31,84,31,84,30,193,31,55,31,38,31,141,31,48,31,189,31,207,31,245,31,245,30,245,29,245,28,19,31,77,31,77,30,242,31,176,31,47,31,80,31,41,31,100,31,228,31,228,30,228,29,202,31,59,31,113,31,48,31,48,30,27,31,3,31,251,31,230,31,7,31,170,31,27,31,1,31,105,31,253,31,82,31,82,30,82,29,62,31,62,30,68,31,141,31,244,31,75,31,7,31,7,30,230,31,74,31,124,31,248,31,248,30,223,31,223,30,102,31,213,31,230,31,17,31,136,31,44,31,124,31,124,30,225,31,143,31,143,30,143,29,143,28,140,31,140,30,20,31,210,31,241,31,125,31,237,31,79,31,79,30,15,31,198,31,37,31,240,31,240,30,65,31,180,31,58,31,211,31,211,30,191,31,168,31,171,31,249,31,21,31,71,31,71,30,58,31,216,31,242,31,36,31,136,31,115,31,115,30,115,29,175,31,175,30,8,31,72,31,56,31,60,31,60,30,237,31,237,30,71,31,141,31,141,30,141,29,200,31,200,30,9,31,99,31,241,31,249,31,242,31,110,31,34,31,145,31,102,31,246,31,19,31,172,31,172,30,181,31,77,31,77,30,242,31,193,31,193,30,67,31,116,31,114,31,186,31,21,31,196,31,52,31,55,31,55,30,40,31,15,31,237,31,206,31,50,31,227,31,160,31,227,31,220,31,198,31,88,31,236,31,135,31,135,30,110,31,78,31,19,31,191,31,13,31,110,31,171,31,223,31,154,31,206,31,206,30,1,31,179,31,233,31,74,31,74,30,187,31,107,31,85,31,32,31,79,31,169,31,169,30,3,31,83,31,106,31,106,30,138,31,12,31,12,30,116,31,197,31,196,31,131,31,85,31,137,31,10,31,129,31,195,31,32,31,52,31,185,31,122,31,75,31,143,31,165,31,165,30,41,31,215,31,213,31,115,31,62,31,122,31,122,30,47,31,154,31,154,30,253,31,162,31,103,31,26,31,26,30,255,31,255,30,102,31,27,31,200,31,70,31,165,31,240,31,59,31,59,30,5,31,5,30,71,31,71,30,74,31,2,31,114,31,253,31,66,31,4,31,192,31,227,31,240,31,176,31,185,31,52,31,52,30,52,29,52,28,45,31,20,31,164,31,224,31,108,31,54,31,241,31,60,31,118,31,17,31,17,30,168,31,21,31,99,31,96,31,11,31,61,31,2,31,248,31,105,31,104,31,194,31,103,31,103,30,73,31,216,31,226,31,215,31,27,31,2,31,2,30,203,31,110,31,190,31,24,31,133,31,56,31,45,31,174,31,174,30,118,31,108,31,158,31,61,31,125,31,167,31,38,31,152,31,202,31,202,30,238,31,238,30,222,31,5,31,96,31,96,30,21,31,140,31,110,31,32,31,32,30,111,31,225,31,225,30,104,31,104,30,104,29,67,31,67,30,131,31,150,31,138,31,54,31,100,31,125,31,28,31,85,31,190,31,190,30,1,31,118,31,177,31,91,31,208,31,252,31,252,30,230,31,130,31,206,31,87,31,87,30,231,31,112,31,130,31,130,30,1,31,120,31,120,30,120,29,6,31,6,30,6,29,10,31,194,31,148,31,44,31,139,31,218,31,204,31,204,30,31,31,140,31,20,31,20,30,130,31,185,31,55,31,55,30,194,31,84,31,69,31,69,30,247,31,189,31,230,31,219,31,142,31,197,31,153,31,239,31,151,31,159,31,214,31,133,31,68,31,138,31,138,30,135,31,135,30,239,31,146,31,250,31,79,31,79,30,120,31,57,31,22,31,242,31,242,30,224,31,20,31,58,31,148,31,93,31,180,31,218,31,109,31,109,30,15,31,15,30,45,31,45,30,249,31,16,31,248,31,125,31,136,31,38,31,55,31,190,31,45,31,45,30,174,31,24,31,104,31,143,31,173,31,18,31,18,30,18,29,18,28,248,31,168,31,255,31,203,31,113,31,222,31,98,31,43,31,247,31,247,30,247,29,98,31,64,31,249,31,95,31,95,30,46,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
