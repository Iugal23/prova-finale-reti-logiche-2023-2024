-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 679;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (55,0,0,0,0,0,70,0,145,0,157,0,182,0,247,0,207,0,105,0,51,0,236,0,0,0,191,0,241,0,120,0,70,0,225,0,0,0,203,0,31,0,0,0,0,0,202,0,240,0,0,0,0,0,168,0,206,0,0,0,34,0,0,0,248,0,61,0,139,0,220,0,205,0,123,0,247,0,82,0,0,0,32,0,168,0,222,0,89,0,27,0,0,0,0,0,73,0,91,0,0,0,197,0,25,0,128,0,252,0,139,0,0,0,0,0,189,0,0,0,0,0,154,0,0,0,52,0,235,0,171,0,240,0,236,0,209,0,142,0,208,0,18,0,15,0,0,0,146,0,113,0,218,0,0,0,0,0,0,0,226,0,182,0,234,0,104,0,206,0,68,0,117,0,58,0,245,0,0,0,0,0,75,0,0,0,178,0,234,0,176,0,244,0,160,0,95,0,172,0,72,0,146,0,81,0,248,0,178,0,0,0,111,0,50,0,0,0,210,0,208,0,24,0,151,0,0,0,0,0,0,0,140,0,243,0,0,0,105,0,169,0,0,0,0,0,178,0,0,0,61,0,132,0,52,0,164,0,0,0,78,0,215,0,253,0,4,0,160,0,196,0,166,0,251,0,184,0,82,0,0,0,246,0,0,0,56,0,24,0,0,0,238,0,0,0,76,0,95,0,206,0,223,0,26,0,136,0,116,0,176,0,0,0,196,0,49,0,54,0,142,0,167,0,183,0,15,0,43,0,0,0,129,0,26,0,0,0,0,0,92,0,0,0,31,0,107,0,124,0,0,0,0,0,233,0,151,0,29,0,118,0,251,0,95,0,155,0,47,0,0,0,101,0,167,0,50,0,73,0,245,0,178,0,69,0,1,0,217,0,56,0,152,0,202,0,0,0,140,0,17,0,28,0,111,0,85,0,34,0,233,0,246,0,56,0,185,0,120,0,211,0,0,0,0,0,129,0,251,0,0,0,182,0,69,0,53,0,0,0,25,0,158,0,203,0,0,0,235,0,101,0,134,0,12,0,91,0,177,0,0,0,109,0,46,0,0,0,152,0,0,0,70,0,240,0,98,0,120,0,0,0,101,0,54,0,191,0,89,0,12,0,0,0,0,0,8,0,0,0,0,0,0,0,130,0,3,0,0,0,151,0,0,0,60,0,86,0,206,0,164,0,0,0,72,0,103,0,253,0,194,0,169,0,58,0,0,0,37,0,176,0,211,0,164,0,88,0,40,0,86,0,116,0,0,0,145,0,3,0,120,0,107,0,120,0,39,0,185,0,216,0,242,0,223,0,183,0,36,0,189,0,71,0,65,0,198,0,193,0,7,0,137,0,78,0,120,0,112,0,140,0,0,0,202,0,2,0,0,0,148,0,53,0,0,0,0,0,6,0,178,0,154,0,207,0,133,0,113,0,209,0,254,0,25,0,146,0,31,0,99,0,212,0,0,0,120,0,46,0,152,0,185,0,219,0,246,0,212,0,0,0,164,0,19,0,72,0,214,0,0,0,0,0,0,0,58,0,150,0,170,0,137,0,0,0,247,0,16,0,0,0,0,0,234,0,107,0,249,0,54,0,45,0,188,0,165,0,57,0,219,0,0,0,154,0,0,0,166,0,36,0,209,0,16,0,0,0,22,0,60,0,0,0,96,0,97,0,210,0,235,0,225,0,171,0,214,0,244,0,234,0,248,0,118,0,60,0,176,0,0,0,45,0,236,0,204,0,85,0,45,0,0,0,139,0,138,0,0,0,0,0,0,0,203,0,120,0,161,0,183,0,6,0,57,0,121,0,100,0,0,0,184,0,204,0,169,0,0,0,162,0,166,0,252,0,0,0,218,0,110,0,116,0,0,0,64,0,0,0,134,0,182,0,254,0,152,0,56,0,113,0,191,0,205,0,162,0,20,0,199,0,135,0,47,0,228,0,19,0,166,0,78,0,161,0,131,0,0,0,171,0,127,0,0,0,182,0,58,0,121,0,39,0,14,0,75,0,170,0,94,0,79,0,79,0,164,0,108,0,137,0,41,0,45,0,65,0,191,0,59,0,58,0,48,0,188,0,0,0,36,0,0,0,41,0,100,0,60,0,143,0,98,0,203,0,60,0,156,0,219,0,0,0,0,0,42,0,0,0,126,0,41,0,158,0,78,0,240,0,215,0,132,0,65,0,59,0,93,0,0,0,167,0,198,0,53,0,49,0,156,0,176,0,174,0,2,0,0,0,54,0,0,0,177,0,160,0,215,0,0,0,0,0,173,0,1,0,243,0,0,0,237,0,252,0,59,0,148,0,143,0,188,0,107,0,84,0,169,0,9,0,128,0,105,0,27,0,0,0,0,0,116,0,12,0,0,0,0,0,0,0,148,0,177,0,7,0,5,0,125,0,175,0,174,0,215,0,103,0,179,0,231,0,247,0,0,0,103,0,0,0,231,0,198,0,29,0,62,0,20,0,144,0,0,0,241,0,0,0,253,0,179,0,0,0,247,0,170,0,237,0,82,0,188,0,165,0,139,0,152,0,109,0,60,0,0,0,217,0,162,0,41,0,173,0,211,0,0,0,0,0,150,0,0,0,0,0,224,0,36,0,149,0,68,0,8,0,0,0,114,0,32,0,3,0,216,0,203,0,43,0,66,0,248,0,12,0,0,0,112,0,118,0,111,0,163,0,58,0,65,0,185,0,0,0,106,0,0,0,252,0,1,0,250,0,44,0,182,0,16,0,157,0,0,0,0,0,0,0,108,0,208,0,224,0,0,0,141,0,126,0,0,0,202,0,0,0,157,0,124,0,197,0,240,0,172,0,15,0,127,0,0,0,0,0,103,0,97,0,99,0,0,0,165,0,1,0,65,0,0,0,17,0,0,0,176,0,239,0,0,0,64,0,252,0,0,0,245,0,138,0,106,0,195,0,237,0,244,0,93,0,0,0,106,0,0,0,54,0,76,0,42,0,0,0,0,0,113,0,40,0,0,0,0,0,171,0,26,0,162,0,242,0,0,0,24,0,41,0,166,0,115,0,214,0,0,0,215,0,156,0,0,0,0,0,174,0);
signal scenario_full  : scenario_type := (55,31,55,30,55,29,70,31,145,31,157,31,182,31,247,31,207,31,105,31,51,31,236,31,236,30,191,31,241,31,120,31,70,31,225,31,225,30,203,31,31,31,31,30,31,29,202,31,240,31,240,30,240,29,168,31,206,31,206,30,34,31,34,30,248,31,61,31,139,31,220,31,205,31,123,31,247,31,82,31,82,30,32,31,168,31,222,31,89,31,27,31,27,30,27,29,73,31,91,31,91,30,197,31,25,31,128,31,252,31,139,31,139,30,139,29,189,31,189,30,189,29,154,31,154,30,52,31,235,31,171,31,240,31,236,31,209,31,142,31,208,31,18,31,15,31,15,30,146,31,113,31,218,31,218,30,218,29,218,28,226,31,182,31,234,31,104,31,206,31,68,31,117,31,58,31,245,31,245,30,245,29,75,31,75,30,178,31,234,31,176,31,244,31,160,31,95,31,172,31,72,31,146,31,81,31,248,31,178,31,178,30,111,31,50,31,50,30,210,31,208,31,24,31,151,31,151,30,151,29,151,28,140,31,243,31,243,30,105,31,169,31,169,30,169,29,178,31,178,30,61,31,132,31,52,31,164,31,164,30,78,31,215,31,253,31,4,31,160,31,196,31,166,31,251,31,184,31,82,31,82,30,246,31,246,30,56,31,24,31,24,30,238,31,238,30,76,31,95,31,206,31,223,31,26,31,136,31,116,31,176,31,176,30,196,31,49,31,54,31,142,31,167,31,183,31,15,31,43,31,43,30,129,31,26,31,26,30,26,29,92,31,92,30,31,31,107,31,124,31,124,30,124,29,233,31,151,31,29,31,118,31,251,31,95,31,155,31,47,31,47,30,101,31,167,31,50,31,73,31,245,31,178,31,69,31,1,31,217,31,56,31,152,31,202,31,202,30,140,31,17,31,28,31,111,31,85,31,34,31,233,31,246,31,56,31,185,31,120,31,211,31,211,30,211,29,129,31,251,31,251,30,182,31,69,31,53,31,53,30,25,31,158,31,203,31,203,30,235,31,101,31,134,31,12,31,91,31,177,31,177,30,109,31,46,31,46,30,152,31,152,30,70,31,240,31,98,31,120,31,120,30,101,31,54,31,191,31,89,31,12,31,12,30,12,29,8,31,8,30,8,29,8,28,130,31,3,31,3,30,151,31,151,30,60,31,86,31,206,31,164,31,164,30,72,31,103,31,253,31,194,31,169,31,58,31,58,30,37,31,176,31,211,31,164,31,88,31,40,31,86,31,116,31,116,30,145,31,3,31,120,31,107,31,120,31,39,31,185,31,216,31,242,31,223,31,183,31,36,31,189,31,71,31,65,31,198,31,193,31,7,31,137,31,78,31,120,31,112,31,140,31,140,30,202,31,2,31,2,30,148,31,53,31,53,30,53,29,6,31,178,31,154,31,207,31,133,31,113,31,209,31,254,31,25,31,146,31,31,31,99,31,212,31,212,30,120,31,46,31,152,31,185,31,219,31,246,31,212,31,212,30,164,31,19,31,72,31,214,31,214,30,214,29,214,28,58,31,150,31,170,31,137,31,137,30,247,31,16,31,16,30,16,29,234,31,107,31,249,31,54,31,45,31,188,31,165,31,57,31,219,31,219,30,154,31,154,30,166,31,36,31,209,31,16,31,16,30,22,31,60,31,60,30,96,31,97,31,210,31,235,31,225,31,171,31,214,31,244,31,234,31,248,31,118,31,60,31,176,31,176,30,45,31,236,31,204,31,85,31,45,31,45,30,139,31,138,31,138,30,138,29,138,28,203,31,120,31,161,31,183,31,6,31,57,31,121,31,100,31,100,30,184,31,204,31,169,31,169,30,162,31,166,31,252,31,252,30,218,31,110,31,116,31,116,30,64,31,64,30,134,31,182,31,254,31,152,31,56,31,113,31,191,31,205,31,162,31,20,31,199,31,135,31,47,31,228,31,19,31,166,31,78,31,161,31,131,31,131,30,171,31,127,31,127,30,182,31,58,31,121,31,39,31,14,31,75,31,170,31,94,31,79,31,79,31,164,31,108,31,137,31,41,31,45,31,65,31,191,31,59,31,58,31,48,31,188,31,188,30,36,31,36,30,41,31,100,31,60,31,143,31,98,31,203,31,60,31,156,31,219,31,219,30,219,29,42,31,42,30,126,31,41,31,158,31,78,31,240,31,215,31,132,31,65,31,59,31,93,31,93,30,167,31,198,31,53,31,49,31,156,31,176,31,174,31,2,31,2,30,54,31,54,30,177,31,160,31,215,31,215,30,215,29,173,31,1,31,243,31,243,30,237,31,252,31,59,31,148,31,143,31,188,31,107,31,84,31,169,31,9,31,128,31,105,31,27,31,27,30,27,29,116,31,12,31,12,30,12,29,12,28,148,31,177,31,7,31,5,31,125,31,175,31,174,31,215,31,103,31,179,31,231,31,247,31,247,30,103,31,103,30,231,31,198,31,29,31,62,31,20,31,144,31,144,30,241,31,241,30,253,31,179,31,179,30,247,31,170,31,237,31,82,31,188,31,165,31,139,31,152,31,109,31,60,31,60,30,217,31,162,31,41,31,173,31,211,31,211,30,211,29,150,31,150,30,150,29,224,31,36,31,149,31,68,31,8,31,8,30,114,31,32,31,3,31,216,31,203,31,43,31,66,31,248,31,12,31,12,30,112,31,118,31,111,31,163,31,58,31,65,31,185,31,185,30,106,31,106,30,252,31,1,31,250,31,44,31,182,31,16,31,157,31,157,30,157,29,157,28,108,31,208,31,224,31,224,30,141,31,126,31,126,30,202,31,202,30,157,31,124,31,197,31,240,31,172,31,15,31,127,31,127,30,127,29,103,31,97,31,99,31,99,30,165,31,1,31,65,31,65,30,17,31,17,30,176,31,239,31,239,30,64,31,252,31,252,30,245,31,138,31,106,31,195,31,237,31,244,31,93,31,93,30,106,31,106,30,54,31,76,31,42,31,42,30,42,29,113,31,40,31,40,30,40,29,171,31,26,31,162,31,242,31,242,30,24,31,41,31,166,31,115,31,214,31,214,30,215,31,156,31,156,30,156,29,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
