-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 592;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,174,0,32,0,44,0,121,0,169,0,66,0,61,0,187,0,148,0,92,0,0,0,0,0,182,0,0,0,233,0,96,0,209,0,206,0,0,0,237,0,0,0,0,0,0,0,93,0,133,0,147,0,67,0,146,0,110,0,137,0,98,0,216,0,20,0,76,0,153,0,88,0,204,0,172,0,248,0,176,0,226,0,83,0,182,0,59,0,231,0,210,0,197,0,187,0,128,0,0,0,182,0,35,0,50,0,164,0,127,0,15,0,130,0,237,0,0,0,0,0,149,0,117,0,138,0,0,0,8,0,32,0,115,0,185,0,158,0,0,0,135,0,169,0,156,0,186,0,110,0,0,0,101,0,222,0,185,0,0,0,254,0,0,0,189,0,220,0,205,0,128,0,104,0,90,0,163,0,72,0,0,0,36,0,63,0,0,0,0,0,50,0,150,0,220,0,134,0,30,0,7,0,46,0,62,0,206,0,1,0,215,0,78,0,187,0,144,0,124,0,128,0,213,0,36,0,127,0,0,0,0,0,22,0,218,0,252,0,83,0,0,0,95,0,0,0,0,0,0,0,110,0,89,0,176,0,47,0,114,0,219,0,39,0,151,0,6,0,0,0,5,0,7,0,0,0,226,0,84,0,41,0,159,0,0,0,213,0,242,0,194,0,127,0,104,0,199,0,23,0,0,0,112,0,175,0,121,0,155,0,42,0,107,0,177,0,177,0,245,0,0,0,112,0,61,0,0,0,61,0,0,0,0,0,79,0,95,0,0,0,216,0,9,0,161,0,204,0,79,0,68,0,0,0,0,0,189,0,0,0,211,0,59,0,170,0,157,0,153,0,61,0,169,0,0,0,33,0,203,0,145,0,213,0,243,0,175,0,24,0,143,0,91,0,46,0,64,0,210,0,4,0,177,0,0,0,0,0,169,0,0,0,140,0,95,0,227,0,0,0,69,0,0,0,168,0,23,0,26,0,160,0,35,0,5,0,164,0,0,0,152,0,43,0,1,0,80,0,0,0,0,0,67,0,0,0,160,0,253,0,205,0,24,0,78,0,33,0,20,0,2,0,217,0,221,0,117,0,0,0,0,0,138,0,162,0,37,0,0,0,47,0,103,0,59,0,0,0,105,0,202,0,97,0,70,0,107,0,0,0,62,0,197,0,60,0,196,0,0,0,0,0,0,0,179,0,233,0,214,0,106,0,156,0,0,0,0,0,249,0,135,0,101,0,201,0,242,0,91,0,0,0,0,0,0,0,136,0,0,0,24,0,0,0,114,0,64,0,226,0,0,0,0,0,177,0,15,0,158,0,68,0,0,0,0,0,136,0,115,0,185,0,0,0,216,0,59,0,0,0,109,0,9,0,229,0,206,0,62,0,6,0,163,0,116,0,0,0,45,0,41,0,100,0,24,0,13,0,0,0,217,0,54,0,212,0,1,0,131,0,0,0,216,0,249,0,107,0,180,0,108,0,126,0,108,0,167,0,127,0,9,0,85,0,223,0,187,0,225,0,232,0,38,0,202,0,39,0,91,0,157,0,0,0,165,0,140,0,231,0,103,0,0,0,39,0,172,0,77,0,0,0,0,0,127,0,93,0,0,0,134,0,106,0,194,0,52,0,163,0,160,0,13,0,191,0,102,0,178,0,152,0,100,0,99,0,0,0,232,0,0,0,209,0,145,0,167,0,247,0,243,0,14,0,0,0,180,0,0,0,119,0,201,0,133,0,62,0,227,0,76,0,125,0,0,0,184,0,136,0,84,0,194,0,152,0,184,0,231,0,159,0,196,0,125,0,191,0,0,0,136,0,151,0,0,0,173,0,206,0,9,0,68,0,83,0,58,0,254,0,196,0,0,0,54,0,129,0,173,0,116,0,42,0,0,0,173,0,194,0,146,0,187,0,0,0,120,0,28,0,255,0,110,0,134,0,0,0,6,0,0,0,0,0,249,0,0,0,103,0,23,0,132,0,199,0,212,0,222,0,253,0,16,0,226,0,0,0,97,0,0,0,7,0,24,0,45,0,96,0,0,0,130,0,0,0,219,0,116,0,178,0,0,0,180,0,80,0,236,0,187,0,233,0,217,0,223,0,218,0,141,0,162,0,34,0,93,0,176,0,202,0,210,0,91,0,50,0,101,0,169,0,0,0,235,0,1,0,19,0,21,0,84,0,36,0,21,0,3,0,0,0,254,0,99,0,41,0,79,0,118,0,133,0,160,0,192,0,242,0,150,0,156,0,0,0,4,0,51,0,51,0,159,0,82,0,197,0,161,0,124,0,239,0,155,0,227,0,25,0,34,0,64,0,99,0,246,0,0,0,203,0,57,0,187,0,0,0,148,0,103,0,50,0,189,0,0,0,103,0,72,0,22,0,250,0,0,0,0,0,9,0,232,0,0,0,0,0,141,0,102,0,74,0,0,0,226,0,239,0,166,0,0,0,28,0,53,0,127,0,103,0,65,0,56,0,0,0,225,0,195,0,97,0,0,0,128,0,0,0,106,0,0,0,0,0,0,0,0,0,33,0,111,0,36,0,194,0,0,0,83,0,86,0,220,0,47,0,182,0,164,0,16,0,123,0,244,0,0,0,169,0,98,0,71,0,247,0,0,0,160,0,8,0,98,0,121,0,6,0,239,0,0,0,0,0,0,0,192,0,3,0);
signal scenario_full  : scenario_type := (154,31,174,31,32,31,44,31,121,31,169,31,66,31,61,31,187,31,148,31,92,31,92,30,92,29,182,31,182,30,233,31,96,31,209,31,206,31,206,30,237,31,237,30,237,29,237,28,93,31,133,31,147,31,67,31,146,31,110,31,137,31,98,31,216,31,20,31,76,31,153,31,88,31,204,31,172,31,248,31,176,31,226,31,83,31,182,31,59,31,231,31,210,31,197,31,187,31,128,31,128,30,182,31,35,31,50,31,164,31,127,31,15,31,130,31,237,31,237,30,237,29,149,31,117,31,138,31,138,30,8,31,32,31,115,31,185,31,158,31,158,30,135,31,169,31,156,31,186,31,110,31,110,30,101,31,222,31,185,31,185,30,254,31,254,30,189,31,220,31,205,31,128,31,104,31,90,31,163,31,72,31,72,30,36,31,63,31,63,30,63,29,50,31,150,31,220,31,134,31,30,31,7,31,46,31,62,31,206,31,1,31,215,31,78,31,187,31,144,31,124,31,128,31,213,31,36,31,127,31,127,30,127,29,22,31,218,31,252,31,83,31,83,30,95,31,95,30,95,29,95,28,110,31,89,31,176,31,47,31,114,31,219,31,39,31,151,31,6,31,6,30,5,31,7,31,7,30,226,31,84,31,41,31,159,31,159,30,213,31,242,31,194,31,127,31,104,31,199,31,23,31,23,30,112,31,175,31,121,31,155,31,42,31,107,31,177,31,177,31,245,31,245,30,112,31,61,31,61,30,61,31,61,30,61,29,79,31,95,31,95,30,216,31,9,31,161,31,204,31,79,31,68,31,68,30,68,29,189,31,189,30,211,31,59,31,170,31,157,31,153,31,61,31,169,31,169,30,33,31,203,31,145,31,213,31,243,31,175,31,24,31,143,31,91,31,46,31,64,31,210,31,4,31,177,31,177,30,177,29,169,31,169,30,140,31,95,31,227,31,227,30,69,31,69,30,168,31,23,31,26,31,160,31,35,31,5,31,164,31,164,30,152,31,43,31,1,31,80,31,80,30,80,29,67,31,67,30,160,31,253,31,205,31,24,31,78,31,33,31,20,31,2,31,217,31,221,31,117,31,117,30,117,29,138,31,162,31,37,31,37,30,47,31,103,31,59,31,59,30,105,31,202,31,97,31,70,31,107,31,107,30,62,31,197,31,60,31,196,31,196,30,196,29,196,28,179,31,233,31,214,31,106,31,156,31,156,30,156,29,249,31,135,31,101,31,201,31,242,31,91,31,91,30,91,29,91,28,136,31,136,30,24,31,24,30,114,31,64,31,226,31,226,30,226,29,177,31,15,31,158,31,68,31,68,30,68,29,136,31,115,31,185,31,185,30,216,31,59,31,59,30,109,31,9,31,229,31,206,31,62,31,6,31,163,31,116,31,116,30,45,31,41,31,100,31,24,31,13,31,13,30,217,31,54,31,212,31,1,31,131,31,131,30,216,31,249,31,107,31,180,31,108,31,126,31,108,31,167,31,127,31,9,31,85,31,223,31,187,31,225,31,232,31,38,31,202,31,39,31,91,31,157,31,157,30,165,31,140,31,231,31,103,31,103,30,39,31,172,31,77,31,77,30,77,29,127,31,93,31,93,30,134,31,106,31,194,31,52,31,163,31,160,31,13,31,191,31,102,31,178,31,152,31,100,31,99,31,99,30,232,31,232,30,209,31,145,31,167,31,247,31,243,31,14,31,14,30,180,31,180,30,119,31,201,31,133,31,62,31,227,31,76,31,125,31,125,30,184,31,136,31,84,31,194,31,152,31,184,31,231,31,159,31,196,31,125,31,191,31,191,30,136,31,151,31,151,30,173,31,206,31,9,31,68,31,83,31,58,31,254,31,196,31,196,30,54,31,129,31,173,31,116,31,42,31,42,30,173,31,194,31,146,31,187,31,187,30,120,31,28,31,255,31,110,31,134,31,134,30,6,31,6,30,6,29,249,31,249,30,103,31,23,31,132,31,199,31,212,31,222,31,253,31,16,31,226,31,226,30,97,31,97,30,7,31,24,31,45,31,96,31,96,30,130,31,130,30,219,31,116,31,178,31,178,30,180,31,80,31,236,31,187,31,233,31,217,31,223,31,218,31,141,31,162,31,34,31,93,31,176,31,202,31,210,31,91,31,50,31,101,31,169,31,169,30,235,31,1,31,19,31,21,31,84,31,36,31,21,31,3,31,3,30,254,31,99,31,41,31,79,31,118,31,133,31,160,31,192,31,242,31,150,31,156,31,156,30,4,31,51,31,51,31,159,31,82,31,197,31,161,31,124,31,239,31,155,31,227,31,25,31,34,31,64,31,99,31,246,31,246,30,203,31,57,31,187,31,187,30,148,31,103,31,50,31,189,31,189,30,103,31,72,31,22,31,250,31,250,30,250,29,9,31,232,31,232,30,232,29,141,31,102,31,74,31,74,30,226,31,239,31,166,31,166,30,28,31,53,31,127,31,103,31,65,31,56,31,56,30,225,31,195,31,97,31,97,30,128,31,128,30,106,31,106,30,106,29,106,28,106,27,33,31,111,31,36,31,194,31,194,30,83,31,86,31,220,31,47,31,182,31,164,31,16,31,123,31,244,31,244,30,169,31,98,31,71,31,247,31,247,30,160,31,8,31,98,31,121,31,6,31,239,31,239,30,239,29,239,28,192,31,3,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
