-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 827;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (58,0,72,0,181,0,222,0,0,0,160,0,135,0,30,0,181,0,65,0,0,0,182,0,0,0,0,0,117,0,209,0,251,0,101,0,70,0,63,0,110,0,0,0,97,0,177,0,0,0,175,0,240,0,86,0,0,0,0,0,4,0,79,0,30,0,63,0,96,0,153,0,88,0,238,0,0,0,46,0,227,0,191,0,140,0,133,0,158,0,89,0,108,0,35,0,159,0,247,0,125,0,205,0,0,0,104,0,202,0,156,0,0,0,233,0,89,0,157,0,97,0,16,0,0,0,144,0,227,0,2,0,105,0,132,0,0,0,198,0,76,0,121,0,184,0,247,0,133,0,73,0,63,0,0,0,0,0,21,0,143,0,0,0,65,0,171,0,126,0,0,0,0,0,171,0,15,0,4,0,163,0,0,0,146,0,0,0,55,0,192,0,13,0,104,0,85,0,152,0,186,0,168,0,0,0,204,0,207,0,212,0,246,0,100,0,253,0,0,0,23,0,37,0,173,0,165,0,107,0,0,0,0,0,97,0,203,0,0,0,195,0,125,0,34,0,228,0,0,0,52,0,73,0,56,0,64,0,243,0,173,0,228,0,0,0,248,0,237,0,160,0,0,0,79,0,212,0,131,0,0,0,55,0,8,0,32,0,0,0,39,0,93,0,184,0,100,0,0,0,237,0,106,0,145,0,137,0,26,0,0,0,39,0,238,0,88,0,72,0,107,0,162,0,0,0,0,0,0,0,0,0,237,0,42,0,0,0,96,0,0,0,242,0,78,0,69,0,0,0,217,0,0,0,2,0,145,0,36,0,119,0,185,0,3,0,60,0,199,0,232,0,74,0,79,0,0,0,152,0,86,0,244,0,0,0,32,0,249,0,237,0,123,0,0,0,247,0,184,0,0,0,240,0,125,0,37,0,145,0,190,0,239,0,135,0,239,0,1,0,150,0,81,0,115,0,93,0,121,0,122,0,177,0,27,0,105,0,153,0,0,0,0,0,211,0,209,0,11,0,199,0,95,0,208,0,104,0,0,0,4,0,68,0,0,0,165,0,79,0,115,0,27,0,187,0,65,0,0,0,100,0,232,0,90,0,0,0,77,0,250,0,218,0,235,0,204,0,248,0,94,0,89,0,151,0,148,0,7,0,234,0,39,0,243,0,28,0,129,0,199,0,238,0,133,0,37,0,132,0,143,0,99,0,44,0,0,0,174,0,16,0,116,0,0,0,0,0,163,0,17,0,136,0,238,0,186,0,143,0,128,0,0,0,52,0,212,0,94,0,0,0,0,0,216,0,77,0,12,0,0,0,94,0,203,0,193,0,143,0,172,0,18,0,104,0,32,0,165,0,0,0,80,0,37,0,0,0,186,0,138,0,83,0,114,0,163,0,205,0,209,0,250,0,0,0,75,0,0,0,49,0,39,0,24,0,117,0,83,0,181,0,135,0,215,0,0,0,74,0,252,0,111,0,80,0,50,0,114,0,127,0,0,0,185,0,51,0,90,0,210,0,41,0,72,0,122,0,166,0,10,0,0,0,133,0,18,0,144,0,239,0,99,0,59,0,0,0,0,0,98,0,0,0,166,0,57,0,177,0,165,0,42,0,32,0,0,0,115,0,0,0,162,0,158,0,0,0,185,0,209,0,184,0,31,0,105,0,61,0,0,0,214,0,140,0,6,0,185,0,112,0,249,0,0,0,95,0,120,0,212,0,101,0,26,0,226,0,215,0,117,0,133,0,112,0,0,0,231,0,212,0,159,0,0,0,112,0,0,0,188,0,0,0,177,0,179,0,0,0,179,0,238,0,156,0,96,0,166,0,160,0,254,0,154,0,13,0,199,0,46,0,0,0,220,0,198,0,126,0,0,0,62,0,174,0,189,0,187,0,44,0,140,0,42,0,0,0,174,0,105,0,0,0,16,0,46,0,0,0,110,0,212,0,217,0,171,0,87,0,90,0,201,0,0,0,41,0,0,0,212,0,162,0,5,0,145,0,33,0,0,0,186,0,92,0,116,0,136,0,153,0,54,0,0,0,168,0,0,0,217,0,10,0,242,0,205,0,17,0,95,0,180,0,0,0,224,0,0,0,0,0,0,0,180,0,164,0,123,0,206,0,40,0,0,0,203,0,19,0,75,0,0,0,121,0,124,0,48,0,205,0,249,0,0,0,1,0,236,0,0,0,62,0,91,0,118,0,71,0,180,0,0,0,60,0,0,0,69,0,0,0,0,0,73,0,0,0,0,0,0,0,155,0,237,0,110,0,17,0,18,0,171,0,240,0,138,0,122,0,0,0,14,0,172,0,2,0,234,0,147,0,160,0,51,0,238,0,0,0,0,0,196,0,0,0,208,0,0,0,0,0,246,0,68,0,202,0,0,0,200,0,39,0,181,0,125,0,0,0,36,0,59,0,23,0,137,0,50,0,15,0,121,0,79,0,61,0,0,0,96,0,250,0,225,0,0,0,173,0,236,0,207,0,207,0,42,0,32,0,182,0,135,0,2,0,175,0,217,0,229,0,0,0,202,0,61,0,0,0,189,0,0,0,0,0,52,0,97,0,0,0,198,0,42,0,177,0,0,0,251,0,111,0,0,0,243,0,233,0,159,0,176,0,0,0,121,0,0,0,89,0,0,0,90,0,0,0,182,0,175,0,172,0,92,0,139,0,15,0,0,0,158,0,111,0,186,0,0,0,229,0,209,0,215,0,250,0,47,0,200,0,143,0,95,0,37,0,221,0,199,0,144,0,116,0,114,0,138,0,0,0,8,0,31,0,107,0,69,0,159,0,52,0,206,0,220,0,136,0,229,0,0,0,141,0,0,0,224,0,208,0,49,0,171,0,148,0,179,0,150,0,44,0,0,0,148,0,45,0,0,0,209,0,213,0,74,0,123,0,179,0,62,0,227,0,0,0,139,0,128,0,198,0,67,0,14,0,96,0,1,0,59,0,0,0,246,0,0,0,151,0,49,0,223,0,199,0,0,0,181,0,53,0,9,0,247,0,0,0,217,0,212,0,14,0,212,0,130,0,206,0,0,0,4,0,35,0,142,0,149,0,53,0,174,0,79,0,0,0,0,0,0,0,68,0,0,0,213,0,139,0,209,0,183,0,0,0,77,0,1,0,0,0,33,0,22,0,40,0,0,0,4,0,32,0,229,0,97,0,0,0,0,0,90,0,0,0,191,0,93,0,27,0,241,0,93,0,0,0,0,0,237,0,0,0,189,0,196,0,0,0,206,0,204,0,223,0,189,0,0,0,175,0,173,0,230,0,0,0,169,0,104,0,0,0,189,0,233,0,0,0,0,0,249,0,183,0,87,0,169,0,84,0,245,0,96,0,208,0,9,0,191,0,141,0,0,0,217,0,56,0,103,0,218,0,172,0,0,0,212,0,1,0,199,0,195,0,205,0,0,0,0,0,203,0,184,0,0,0,209,0,0,0,0,0,218,0,124,0,71,0,0,0,239,0,26,0,230,0,147,0,254,0,84,0,237,0,215,0,150,0,220,0,236,0,69,0,0,0,59,0,88,0,132,0,49,0,179,0,200,0,83,0,146,0,142,0,197,0,247,0,252,0,234,0,112,0,71,0,51,0,0,0,151,0,0,0,144,0,75,0,192,0,0,0,172,0,0,0,157,0,152,0,96,0,35,0,221,0,0,0,19,0,209,0,0,0,5,0,180,0,102,0,0,0,167,0,0,0,239,0,65,0);
signal scenario_full  : scenario_type := (58,31,72,31,181,31,222,31,222,30,160,31,135,31,30,31,181,31,65,31,65,30,182,31,182,30,182,29,117,31,209,31,251,31,101,31,70,31,63,31,110,31,110,30,97,31,177,31,177,30,175,31,240,31,86,31,86,30,86,29,4,31,79,31,30,31,63,31,96,31,153,31,88,31,238,31,238,30,46,31,227,31,191,31,140,31,133,31,158,31,89,31,108,31,35,31,159,31,247,31,125,31,205,31,205,30,104,31,202,31,156,31,156,30,233,31,89,31,157,31,97,31,16,31,16,30,144,31,227,31,2,31,105,31,132,31,132,30,198,31,76,31,121,31,184,31,247,31,133,31,73,31,63,31,63,30,63,29,21,31,143,31,143,30,65,31,171,31,126,31,126,30,126,29,171,31,15,31,4,31,163,31,163,30,146,31,146,30,55,31,192,31,13,31,104,31,85,31,152,31,186,31,168,31,168,30,204,31,207,31,212,31,246,31,100,31,253,31,253,30,23,31,37,31,173,31,165,31,107,31,107,30,107,29,97,31,203,31,203,30,195,31,125,31,34,31,228,31,228,30,52,31,73,31,56,31,64,31,243,31,173,31,228,31,228,30,248,31,237,31,160,31,160,30,79,31,212,31,131,31,131,30,55,31,8,31,32,31,32,30,39,31,93,31,184,31,100,31,100,30,237,31,106,31,145,31,137,31,26,31,26,30,39,31,238,31,88,31,72,31,107,31,162,31,162,30,162,29,162,28,162,27,237,31,42,31,42,30,96,31,96,30,242,31,78,31,69,31,69,30,217,31,217,30,2,31,145,31,36,31,119,31,185,31,3,31,60,31,199,31,232,31,74,31,79,31,79,30,152,31,86,31,244,31,244,30,32,31,249,31,237,31,123,31,123,30,247,31,184,31,184,30,240,31,125,31,37,31,145,31,190,31,239,31,135,31,239,31,1,31,150,31,81,31,115,31,93,31,121,31,122,31,177,31,27,31,105,31,153,31,153,30,153,29,211,31,209,31,11,31,199,31,95,31,208,31,104,31,104,30,4,31,68,31,68,30,165,31,79,31,115,31,27,31,187,31,65,31,65,30,100,31,232,31,90,31,90,30,77,31,250,31,218,31,235,31,204,31,248,31,94,31,89,31,151,31,148,31,7,31,234,31,39,31,243,31,28,31,129,31,199,31,238,31,133,31,37,31,132,31,143,31,99,31,44,31,44,30,174,31,16,31,116,31,116,30,116,29,163,31,17,31,136,31,238,31,186,31,143,31,128,31,128,30,52,31,212,31,94,31,94,30,94,29,216,31,77,31,12,31,12,30,94,31,203,31,193,31,143,31,172,31,18,31,104,31,32,31,165,31,165,30,80,31,37,31,37,30,186,31,138,31,83,31,114,31,163,31,205,31,209,31,250,31,250,30,75,31,75,30,49,31,39,31,24,31,117,31,83,31,181,31,135,31,215,31,215,30,74,31,252,31,111,31,80,31,50,31,114,31,127,31,127,30,185,31,51,31,90,31,210,31,41,31,72,31,122,31,166,31,10,31,10,30,133,31,18,31,144,31,239,31,99,31,59,31,59,30,59,29,98,31,98,30,166,31,57,31,177,31,165,31,42,31,32,31,32,30,115,31,115,30,162,31,158,31,158,30,185,31,209,31,184,31,31,31,105,31,61,31,61,30,214,31,140,31,6,31,185,31,112,31,249,31,249,30,95,31,120,31,212,31,101,31,26,31,226,31,215,31,117,31,133,31,112,31,112,30,231,31,212,31,159,31,159,30,112,31,112,30,188,31,188,30,177,31,179,31,179,30,179,31,238,31,156,31,96,31,166,31,160,31,254,31,154,31,13,31,199,31,46,31,46,30,220,31,198,31,126,31,126,30,62,31,174,31,189,31,187,31,44,31,140,31,42,31,42,30,174,31,105,31,105,30,16,31,46,31,46,30,110,31,212,31,217,31,171,31,87,31,90,31,201,31,201,30,41,31,41,30,212,31,162,31,5,31,145,31,33,31,33,30,186,31,92,31,116,31,136,31,153,31,54,31,54,30,168,31,168,30,217,31,10,31,242,31,205,31,17,31,95,31,180,31,180,30,224,31,224,30,224,29,224,28,180,31,164,31,123,31,206,31,40,31,40,30,203,31,19,31,75,31,75,30,121,31,124,31,48,31,205,31,249,31,249,30,1,31,236,31,236,30,62,31,91,31,118,31,71,31,180,31,180,30,60,31,60,30,69,31,69,30,69,29,73,31,73,30,73,29,73,28,155,31,237,31,110,31,17,31,18,31,171,31,240,31,138,31,122,31,122,30,14,31,172,31,2,31,234,31,147,31,160,31,51,31,238,31,238,30,238,29,196,31,196,30,208,31,208,30,208,29,246,31,68,31,202,31,202,30,200,31,39,31,181,31,125,31,125,30,36,31,59,31,23,31,137,31,50,31,15,31,121,31,79,31,61,31,61,30,96,31,250,31,225,31,225,30,173,31,236,31,207,31,207,31,42,31,32,31,182,31,135,31,2,31,175,31,217,31,229,31,229,30,202,31,61,31,61,30,189,31,189,30,189,29,52,31,97,31,97,30,198,31,42,31,177,31,177,30,251,31,111,31,111,30,243,31,233,31,159,31,176,31,176,30,121,31,121,30,89,31,89,30,90,31,90,30,182,31,175,31,172,31,92,31,139,31,15,31,15,30,158,31,111,31,186,31,186,30,229,31,209,31,215,31,250,31,47,31,200,31,143,31,95,31,37,31,221,31,199,31,144,31,116,31,114,31,138,31,138,30,8,31,31,31,107,31,69,31,159,31,52,31,206,31,220,31,136,31,229,31,229,30,141,31,141,30,224,31,208,31,49,31,171,31,148,31,179,31,150,31,44,31,44,30,148,31,45,31,45,30,209,31,213,31,74,31,123,31,179,31,62,31,227,31,227,30,139,31,128,31,198,31,67,31,14,31,96,31,1,31,59,31,59,30,246,31,246,30,151,31,49,31,223,31,199,31,199,30,181,31,53,31,9,31,247,31,247,30,217,31,212,31,14,31,212,31,130,31,206,31,206,30,4,31,35,31,142,31,149,31,53,31,174,31,79,31,79,30,79,29,79,28,68,31,68,30,213,31,139,31,209,31,183,31,183,30,77,31,1,31,1,30,33,31,22,31,40,31,40,30,4,31,32,31,229,31,97,31,97,30,97,29,90,31,90,30,191,31,93,31,27,31,241,31,93,31,93,30,93,29,237,31,237,30,189,31,196,31,196,30,206,31,204,31,223,31,189,31,189,30,175,31,173,31,230,31,230,30,169,31,104,31,104,30,189,31,233,31,233,30,233,29,249,31,183,31,87,31,169,31,84,31,245,31,96,31,208,31,9,31,191,31,141,31,141,30,217,31,56,31,103,31,218,31,172,31,172,30,212,31,1,31,199,31,195,31,205,31,205,30,205,29,203,31,184,31,184,30,209,31,209,30,209,29,218,31,124,31,71,31,71,30,239,31,26,31,230,31,147,31,254,31,84,31,237,31,215,31,150,31,220,31,236,31,69,31,69,30,59,31,88,31,132,31,49,31,179,31,200,31,83,31,146,31,142,31,197,31,247,31,252,31,234,31,112,31,71,31,51,31,51,30,151,31,151,30,144,31,75,31,192,31,192,30,172,31,172,30,157,31,152,31,96,31,35,31,221,31,221,30,19,31,209,31,209,30,5,31,180,31,102,31,102,30,167,31,167,30,239,31,65,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
