-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_979 is
end project_tb_979;

architecture project_tb_arch_979 of project_tb_979 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 815;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (57,0,154,0,16,0,211,0,155,0,51,0,96,0,192,0,167,0,66,0,222,0,33,0,240,0,0,0,210,0,54,0,163,0,253,0,112,0,133,0,0,0,54,0,63,0,84,0,89,0,23,0,13,0,108,0,220,0,90,0,201,0,44,0,67,0,18,0,140,0,143,0,54,0,184,0,100,0,171,0,118,0,123,0,251,0,142,0,118,0,17,0,0,0,202,0,2,0,195,0,151,0,0,0,193,0,179,0,103,0,156,0,107,0,222,0,0,0,49,0,106,0,0,0,211,0,127,0,231,0,171,0,143,0,246,0,6,0,0,0,148,0,209,0,42,0,210,0,91,0,108,0,131,0,78,0,105,0,245,0,143,0,100,0,0,0,15,0,73,0,0,0,157,0,0,0,0,0,230,0,41,0,62,0,143,0,181,0,114,0,0,0,194,0,148,0,227,0,19,0,0,0,216,0,15,0,0,0,0,0,232,0,174,0,41,0,56,0,85,0,237,0,0,0,197,0,47,0,0,0,3,0,87,0,183,0,0,0,0,0,99,0,0,0,118,0,225,0,222,0,121,0,236,0,242,0,176,0,58,0,38,0,125,0,101,0,113,0,85,0,156,0,52,0,89,0,123,0,0,0,14,0,0,0,24,0,152,0,238,0,230,0,35,0,51,0,0,0,15,0,244,0,0,0,85,0,142,0,42,0,176,0,35,0,108,0,0,0,0,0,83,0,189,0,137,0,156,0,0,0,102,0,238,0,35,0,202,0,81,0,89,0,138,0,39,0,236,0,0,0,186,0,199,0,25,0,0,0,199,0,100,0,57,0,104,0,101,0,102,0,193,0,0,0,0,0,60,0,50,0,97,0,15,0,0,0,0,0,0,0,127,0,136,0,177,0,148,0,0,0,114,0,251,0,8,0,0,0,43,0,154,0,146,0,40,0,52,0,130,0,0,0,198,0,107,0,84,0,98,0,90,0,146,0,73,0,0,0,119,0,27,0,5,0,203,0,121,0,218,0,66,0,165,0,54,0,186,0,235,0,61,0,112,0,62,0,217,0,10,0,214,0,189,0,129,0,166,0,60,0,237,0,0,0,0,0,0,0,24,0,180,0,35,0,36,0,113,0,0,0,242,0,85,0,1,0,228,0,51,0,160,0,114,0,0,0,66,0,131,0,54,0,122,0,204,0,116,0,96,0,75,0,91,0,0,0,25,0,121,0,40,0,211,0,0,0,183,0,41,0,101,0,131,0,0,0,147,0,162,0,0,0,58,0,52,0,139,0,15,0,117,0,250,0,64,0,192,0,55,0,0,0,150,0,77,0,1,0,35,0,143,0,0,0,127,0,0,0,0,0,74,0,11,0,98,0,114,0,133,0,133,0,151,0,0,0,119,0,30,0,167,0,173,0,79,0,187,0,12,0,9,0,247,0,0,0,196,0,0,0,242,0,135,0,0,0,37,0,0,0,74,0,104,0,128,0,153,0,250,0,0,0,0,0,121,0,0,0,205,0,183,0,0,0,17,0,0,0,10,0,33,0,11,0,71,0,71,0,115,0,227,0,198,0,86,0,19,0,0,0,225,0,134,0,154,0,37,0,253,0,0,0,0,0,121,0,229,0,0,0,108,0,1,0,0,0,0,0,0,0,70,0,0,0,0,0,0,0,33,0,0,0,212,0,49,0,0,0,154,0,0,0,42,0,217,0,133,0,119,0,187,0,237,0,49,0,35,0,249,0,94,0,0,0,168,0,28,0,27,0,83,0,0,0,234,0,5,0,223,0,0,0,79,0,73,0,0,0,240,0,0,0,0,0,0,0,0,0,54,0,12,0,10,0,86,0,210,0,158,0,193,0,137,0,71,0,54,0,155,0,222,0,217,0,0,0,13,0,118,0,199,0,186,0,172,0,216,0,51,0,236,0,0,0,209,0,2,0,4,0,48,0,129,0,0,0,172,0,171,0,69,0,0,0,255,0,44,0,0,0,0,0,0,0,47,0,0,0,193,0,198,0,82,0,188,0,114,0,159,0,210,0,100,0,8,0,56,0,240,0,183,0,162,0,180,0,205,0,53,0,131,0,0,0,119,0,0,0,0,0,80,0,1,0,238,0,81,0,3,0,247,0,25,0,0,0,0,0,21,0,156,0,22,0,117,0,172,0,0,0,157,0,106,0,231,0,122,0,211,0,252,0,237,0,0,0,38,0,54,0,37,0,160,0,24,0,4,0,11,0,169,0,146,0,229,0,124,0,124,0,45,0,144,0,48,0,0,0,119,0,24,0,124,0,165,0,0,0,0,0,204,0,135,0,0,0,133,0,38,0,0,0,214,0,97,0,231,0,205,0,109,0,14,0,82,0,171,0,168,0,176,0,171,0,136,0,37,0,0,0,139,0,144,0,82,0,223,0,43,0,1,0,0,0,226,0,0,0,125,0,6,0,35,0,128,0,172,0,46,0,183,0,125,0,231,0,0,0,143,0,54,0,0,0,189,0,140,0,119,0,122,0,131,0,186,0,75,0,15,0,0,0,0,0,174,0,60,0,0,0,185,0,0,0,208,0,45,0,234,0,209,0,217,0,70,0,195,0,142,0,47,0,0,0,242,0,0,0,232,0,122,0,134,0,92,0,0,0,189,0,9,0,28,0,165,0,0,0,35,0,99,0,2,0,0,0,142,0,120,0,39,0,230,0,45,0,195,0,202,0,255,0,71,0,204,0,249,0,0,0,245,0,0,0,146,0,227,0,183,0,69,0,0,0,195,0,99,0,188,0,246,0,164,0,244,0,0,0,0,0,23,0,183,0,227,0,0,0,77,0,97,0,85,0,171,0,61,0,0,0,25,0,147,0,25,0,253,0,127,0,179,0,248,0,1,0,89,0,123,0,200,0,222,0,106,0,25,0,161,0,1,0,62,0,146,0,0,0,117,0,99,0,8,0,126,0,79,0,100,0,185,0,105,0,183,0,0,0,0,0,0,0,171,0,253,0,206,0,183,0,230,0,64,0,224,0,217,0,0,0,154,0,0,0,87,0,0,0,232,0,118,0,0,0,198,0,33,0,58,0,10,0,0,0,0,0,188,0,0,0,235,0,102,0,29,0,167,0,195,0,214,0,127,0,0,0,236,0,181,0,129,0,148,0,195,0,112,0,0,0,34,0,196,0,146,0,49,0,90,0,216,0,168,0,225,0,34,0,0,0,106,0,0,0,73,0,0,0,0,0,237,0,174,0,190,0,61,0,172,0,168,0,212,0,117,0,0,0,0,0,160,0,188,0,1,0,0,0,133,0,164,0,0,0,196,0,0,0,240,0,211,0,129,0,160,0,214,0,33,0,128,0,176,0,161,0,53,0,251,0,0,0,231,0,94,0,99,0,211,0,6,0,0,0,155,0,227,0,208,0,155,0,35,0,45,0,98,0,159,0,190,0,172,0,89,0,30,0,0,0,125,0,173,0,225,0,0,0,90,0,242,0,48,0,0,0,113,0,218,0,53,0,179,0,0,0,39,0,165,0,54,0,169,0,0,0,160,0,0,0,235,0,0,0,169,0,0,0,0,0,173,0,206,0,85,0,234,0,117,0,0,0,0,0,0,0,254,0,199,0,207,0,212,0,172,0,231,0,162,0,14,0,75,0,0,0,149,0,3,0,254,0,110,0,0,0,91,0,76,0);
signal scenario_full  : scenario_type := (57,31,154,31,16,31,211,31,155,31,51,31,96,31,192,31,167,31,66,31,222,31,33,31,240,31,240,30,210,31,54,31,163,31,253,31,112,31,133,31,133,30,54,31,63,31,84,31,89,31,23,31,13,31,108,31,220,31,90,31,201,31,44,31,67,31,18,31,140,31,143,31,54,31,184,31,100,31,171,31,118,31,123,31,251,31,142,31,118,31,17,31,17,30,202,31,2,31,195,31,151,31,151,30,193,31,179,31,103,31,156,31,107,31,222,31,222,30,49,31,106,31,106,30,211,31,127,31,231,31,171,31,143,31,246,31,6,31,6,30,148,31,209,31,42,31,210,31,91,31,108,31,131,31,78,31,105,31,245,31,143,31,100,31,100,30,15,31,73,31,73,30,157,31,157,30,157,29,230,31,41,31,62,31,143,31,181,31,114,31,114,30,194,31,148,31,227,31,19,31,19,30,216,31,15,31,15,30,15,29,232,31,174,31,41,31,56,31,85,31,237,31,237,30,197,31,47,31,47,30,3,31,87,31,183,31,183,30,183,29,99,31,99,30,118,31,225,31,222,31,121,31,236,31,242,31,176,31,58,31,38,31,125,31,101,31,113,31,85,31,156,31,52,31,89,31,123,31,123,30,14,31,14,30,24,31,152,31,238,31,230,31,35,31,51,31,51,30,15,31,244,31,244,30,85,31,142,31,42,31,176,31,35,31,108,31,108,30,108,29,83,31,189,31,137,31,156,31,156,30,102,31,238,31,35,31,202,31,81,31,89,31,138,31,39,31,236,31,236,30,186,31,199,31,25,31,25,30,199,31,100,31,57,31,104,31,101,31,102,31,193,31,193,30,193,29,60,31,50,31,97,31,15,31,15,30,15,29,15,28,127,31,136,31,177,31,148,31,148,30,114,31,251,31,8,31,8,30,43,31,154,31,146,31,40,31,52,31,130,31,130,30,198,31,107,31,84,31,98,31,90,31,146,31,73,31,73,30,119,31,27,31,5,31,203,31,121,31,218,31,66,31,165,31,54,31,186,31,235,31,61,31,112,31,62,31,217,31,10,31,214,31,189,31,129,31,166,31,60,31,237,31,237,30,237,29,237,28,24,31,180,31,35,31,36,31,113,31,113,30,242,31,85,31,1,31,228,31,51,31,160,31,114,31,114,30,66,31,131,31,54,31,122,31,204,31,116,31,96,31,75,31,91,31,91,30,25,31,121,31,40,31,211,31,211,30,183,31,41,31,101,31,131,31,131,30,147,31,162,31,162,30,58,31,52,31,139,31,15,31,117,31,250,31,64,31,192,31,55,31,55,30,150,31,77,31,1,31,35,31,143,31,143,30,127,31,127,30,127,29,74,31,11,31,98,31,114,31,133,31,133,31,151,31,151,30,119,31,30,31,167,31,173,31,79,31,187,31,12,31,9,31,247,31,247,30,196,31,196,30,242,31,135,31,135,30,37,31,37,30,74,31,104,31,128,31,153,31,250,31,250,30,250,29,121,31,121,30,205,31,183,31,183,30,17,31,17,30,10,31,33,31,11,31,71,31,71,31,115,31,227,31,198,31,86,31,19,31,19,30,225,31,134,31,154,31,37,31,253,31,253,30,253,29,121,31,229,31,229,30,108,31,1,31,1,30,1,29,1,28,70,31,70,30,70,29,70,28,33,31,33,30,212,31,49,31,49,30,154,31,154,30,42,31,217,31,133,31,119,31,187,31,237,31,49,31,35,31,249,31,94,31,94,30,168,31,28,31,27,31,83,31,83,30,234,31,5,31,223,31,223,30,79,31,73,31,73,30,240,31,240,30,240,29,240,28,240,27,54,31,12,31,10,31,86,31,210,31,158,31,193,31,137,31,71,31,54,31,155,31,222,31,217,31,217,30,13,31,118,31,199,31,186,31,172,31,216,31,51,31,236,31,236,30,209,31,2,31,4,31,48,31,129,31,129,30,172,31,171,31,69,31,69,30,255,31,44,31,44,30,44,29,44,28,47,31,47,30,193,31,198,31,82,31,188,31,114,31,159,31,210,31,100,31,8,31,56,31,240,31,183,31,162,31,180,31,205,31,53,31,131,31,131,30,119,31,119,30,119,29,80,31,1,31,238,31,81,31,3,31,247,31,25,31,25,30,25,29,21,31,156,31,22,31,117,31,172,31,172,30,157,31,106,31,231,31,122,31,211,31,252,31,237,31,237,30,38,31,54,31,37,31,160,31,24,31,4,31,11,31,169,31,146,31,229,31,124,31,124,31,45,31,144,31,48,31,48,30,119,31,24,31,124,31,165,31,165,30,165,29,204,31,135,31,135,30,133,31,38,31,38,30,214,31,97,31,231,31,205,31,109,31,14,31,82,31,171,31,168,31,176,31,171,31,136,31,37,31,37,30,139,31,144,31,82,31,223,31,43,31,1,31,1,30,226,31,226,30,125,31,6,31,35,31,128,31,172,31,46,31,183,31,125,31,231,31,231,30,143,31,54,31,54,30,189,31,140,31,119,31,122,31,131,31,186,31,75,31,15,31,15,30,15,29,174,31,60,31,60,30,185,31,185,30,208,31,45,31,234,31,209,31,217,31,70,31,195,31,142,31,47,31,47,30,242,31,242,30,232,31,122,31,134,31,92,31,92,30,189,31,9,31,28,31,165,31,165,30,35,31,99,31,2,31,2,30,142,31,120,31,39,31,230,31,45,31,195,31,202,31,255,31,71,31,204,31,249,31,249,30,245,31,245,30,146,31,227,31,183,31,69,31,69,30,195,31,99,31,188,31,246,31,164,31,244,31,244,30,244,29,23,31,183,31,227,31,227,30,77,31,97,31,85,31,171,31,61,31,61,30,25,31,147,31,25,31,253,31,127,31,179,31,248,31,1,31,89,31,123,31,200,31,222,31,106,31,25,31,161,31,1,31,62,31,146,31,146,30,117,31,99,31,8,31,126,31,79,31,100,31,185,31,105,31,183,31,183,30,183,29,183,28,171,31,253,31,206,31,183,31,230,31,64,31,224,31,217,31,217,30,154,31,154,30,87,31,87,30,232,31,118,31,118,30,198,31,33,31,58,31,10,31,10,30,10,29,188,31,188,30,235,31,102,31,29,31,167,31,195,31,214,31,127,31,127,30,236,31,181,31,129,31,148,31,195,31,112,31,112,30,34,31,196,31,146,31,49,31,90,31,216,31,168,31,225,31,34,31,34,30,106,31,106,30,73,31,73,30,73,29,237,31,174,31,190,31,61,31,172,31,168,31,212,31,117,31,117,30,117,29,160,31,188,31,1,31,1,30,133,31,164,31,164,30,196,31,196,30,240,31,211,31,129,31,160,31,214,31,33,31,128,31,176,31,161,31,53,31,251,31,251,30,231,31,94,31,99,31,211,31,6,31,6,30,155,31,227,31,208,31,155,31,35,31,45,31,98,31,159,31,190,31,172,31,89,31,30,31,30,30,125,31,173,31,225,31,225,30,90,31,242,31,48,31,48,30,113,31,218,31,53,31,179,31,179,30,39,31,165,31,54,31,169,31,169,30,160,31,160,30,235,31,235,30,169,31,169,30,169,29,173,31,206,31,85,31,234,31,117,31,117,30,117,29,117,28,254,31,199,31,207,31,212,31,172,31,231,31,162,31,14,31,75,31,75,30,149,31,3,31,254,31,110,31,110,30,91,31,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
