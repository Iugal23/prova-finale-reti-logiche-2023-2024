-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_163 is
end project_tb_163;

architecture project_tb_arch_163 of project_tb_163 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 887;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (183,0,0,0,155,0,0,0,0,0,0,0,113,0,132,0,0,0,0,0,148,0,150,0,117,0,104,0,219,0,0,0,0,0,147,0,0,0,248,0,0,0,7,0,58,0,25,0,205,0,240,0,106,0,194,0,135,0,70,0,103,0,99,0,23,0,0,0,0,0,124,0,247,0,58,0,233,0,136,0,147,0,0,0,96,0,70,0,171,0,140,0,210,0,122,0,138,0,0,0,8,0,112,0,0,0,65,0,0,0,57,0,138,0,144,0,0,0,185,0,110,0,0,0,240,0,229,0,133,0,118,0,33,0,0,0,255,0,237,0,53,0,140,0,142,0,243,0,169,0,240,0,69,0,0,0,87,0,229,0,0,0,182,0,123,0,234,0,0,0,192,0,0,0,132,0,0,0,122,0,184,0,245,0,229,0,110,0,0,0,63,0,138,0,183,0,0,0,138,0,187,0,125,0,199,0,62,0,50,0,0,0,117,0,102,0,153,0,90,0,131,0,82,0,0,0,154,0,124,0,232,0,7,0,153,0,65,0,233,0,135,0,203,0,210,0,131,0,0,0,195,0,41,0,46,0,96,0,96,0,0,0,0,0,154,0,191,0,87,0,111,0,255,0,231,0,17,0,253,0,198,0,120,0,63,0,23,0,126,0,99,0,0,0,0,0,65,0,198,0,140,0,223,0,0,0,0,0,118,0,81,0,87,0,56,0,174,0,0,0,0,0,205,0,0,0,224,0,235,0,0,0,209,0,175,0,1,0,186,0,64,0,58,0,218,0,0,0,47,0,117,0,97,0,86,0,132,0,0,0,238,0,102,0,4,0,245,0,0,0,249,0,0,0,179,0,148,0,194,0,0,0,69,0,232,0,11,0,148,0,12,0,198,0,166,0,152,0,248,0,4,0,77,0,213,0,61,0,133,0,214,0,7,0,22,0,167,0,0,0,30,0,0,0,0,0,0,0,100,0,52,0,0,0,117,0,0,0,0,0,35,0,231,0,12,0,0,0,0,0,226,0,194,0,0,0,218,0,41,0,196,0,168,0,115,0,180,0,56,0,60,0,205,0,46,0,96,0,100,0,198,0,18,0,92,0,82,0,121,0,77,0,210,0,67,0,101,0,28,0,203,0,111,0,200,0,0,0,36,0,228,0,246,0,200,0,0,0,87,0,45,0,127,0,255,0,128,0,217,0,201,0,225,0,0,0,102,0,2,0,94,0,153,0,183,0,0,0,0,0,68,0,242,0,113,0,0,0,137,0,204,0,246,0,89,0,203,0,203,0,152,0,25,0,254,0,11,0,28,0,0,0,0,0,0,0,15,0,221,0,0,0,246,0,118,0,245,0,66,0,24,0,0,0,116,0,196,0,211,0,219,0,108,0,177,0,227,0,110,0,5,0,53,0,196,0,169,0,40,0,214,0,103,0,183,0,240,0,74,0,0,0,67,0,210,0,0,0,164,0,108,0,0,0,92,0,60,0,215,0,255,0,14,0,233,0,0,0,0,0,235,0,226,0,203,0,131,0,0,0,0,0,0,0,150,0,194,0,173,0,138,0,127,0,151,0,105,0,0,0,241,0,220,0,0,0,236,0,0,0,250,0,0,0,66,0,185,0,0,0,211,0,0,0,61,0,57,0,52,0,0,0,0,0,97,0,194,0,140,0,140,0,164,0,59,0,214,0,102,0,11,0,236,0,27,0,222,0,0,0,206,0,201,0,116,0,90,0,159,0,0,0,61,0,0,0,114,0,181,0,240,0,56,0,86,0,217,0,0,0,37,0,164,0,250,0,249,0,100,0,90,0,166,0,237,0,73,0,74,0,238,0,0,0,206,0,159,0,0,0,225,0,89,0,73,0,17,0,153,0,173,0,217,0,0,0,211,0,117,0,106,0,188,0,131,0,0,0,254,0,243,0,0,0,0,0,74,0,34,0,184,0,68,0,182,0,177,0,189,0,180,0,0,0,212,0,11,0,223,0,118,0,253,0,183,0,125,0,82,0,177,0,74,0,227,0,252,0,189,0,70,0,39,0,174,0,240,0,53,0,131,0,214,0,50,0,0,0,208,0,6,0,200,0,68,0,67,0,157,0,246,0,38,0,59,0,55,0,0,0,131,0,64,0,0,0,25,0,214,0,28,0,92,0,18,0,77,0,5,0,30,0,248,0,8,0,0,0,94,0,152,0,246,0,183,0,0,0,50,0,151,0,157,0,254,0,0,0,155,0,0,0,0,0,0,0,60,0,164,0,237,0,143,0,124,0,244,0,0,0,246,0,0,0,58,0,167,0,93,0,108,0,0,0,0,0,116,0,35,0,242,0,236,0,99,0,236,0,66,0,239,0,232,0,55,0,137,0,176,0,69,0,15,0,0,0,0,0,182,0,146,0,213,0,150,0,187,0,241,0,68,0,207,0,89,0,109,0,70,0,0,0,68,0,0,0,138,0,111,0,25,0,190,0,0,0,72,0,217,0,220,0,8,0,159,0,0,0,0,0,191,0,216,0,221,0,0,0,196,0,0,0,0,0,73,0,61,0,39,0,0,0,34,0,83,0,0,0,0,0,52,0,33,0,220,0,104,0,152,0,179,0,187,0,7,0,148,0,154,0,0,0,5,0,112,0,12,0,0,0,206,0,195,0,0,0,48,0,145,0,139,0,22,0,64,0,0,0,192,0,0,0,196,0,159,0,0,0,146,0,187,0,85,0,161,0,0,0,68,0,111,0,57,0,214,0,174,0,239,0,147,0,6,0,178,0,117,0,24,0,29,0,0,0,184,0,0,0,139,0,0,0,0,0,248,0,83,0,30,0,91,0,183,0,70,0,0,0,80,0,80,0,0,0,232,0,137,0,0,0,106,0,0,0,0,0,164,0,0,0,56,0,0,0,220,0,0,0,64,0,0,0,204,0,53,0,129,0,13,0,248,0,0,0,0,0,222,0,104,0,141,0,25,0,50,0,114,0,123,0,0,0,234,0,202,0,119,0,135,0,58,0,131,0,211,0,49,0,0,0,0,0,0,0,0,0,249,0,0,0,131,0,187,0,78,0,0,0,19,0,182,0,254,0,0,0,0,0,0,0,227,0,0,0,0,0,132,0,246,0,38,0,116,0,17,0,168,0,228,0,0,0,46,0,0,0,194,0,151,0,109,0,0,0,94,0,0,0,84,0,124,0,39,0,182,0,213,0,228,0,152,0,0,0,0,0,236,0,0,0,0,0,196,0,41,0,40,0,71,0,63,0,154,0,156,0,0,0,0,0,125,0,226,0,165,0,0,0,29,0,49,0,0,0,0,0,164,0,22,0,77,0,0,0,0,0,160,0,0,0,20,0,0,0,130,0,173,0,217,0,98,0,63,0,97,0,237,0,48,0,18,0,210,0,244,0,179,0,68,0,101,0,72,0,8,0,145,0,208,0,0,0,106,0,232,0,0,0,18,0,164,0,0,0,112,0,12,0,114,0,48,0,148,0,226,0,255,0,70,0,2,0,205,0,222,0,203,0,107,0,96,0,61,0,0,0,0,0,233,0,98,0,0,0,62,0,0,0,197,0,107,0,150,0,95,0,184,0,194,0,36,0,243,0,107,0,206,0,81,0,0,0,21,0,23,0,205,0,0,0,0,0,42,0,22,0,12,0,47,0,234,0,254,0,216,0,0,0,23,0,52,0,12,0,233,0,126,0,179,0,112,0,144,0,100,0,224,0,9,0,50,0,99,0,0,0,109,0,0,0,64,0,75,0,180,0,93,0,160,0,17,0,228,0,56,0,234,0,0,0,0,0,57,0,0,0,0,0,0,0,195,0,46,0,63,0,42,0,234,0,251,0,22,0,0,0,132,0,173,0,144,0,246,0,204,0,158,0,57,0,65,0,122,0,243,0,94,0,38,0,234,0,246,0,0,0,98,0,252,0,165,0,143,0,0,0,103,0,35,0,134,0,59,0,67,0,96,0,191,0,219,0,103,0,0,0,106,0,183,0,0,0,0,0);
signal scenario_full  : scenario_type := (183,31,183,30,155,31,155,30,155,29,155,28,113,31,132,31,132,30,132,29,148,31,150,31,117,31,104,31,219,31,219,30,219,29,147,31,147,30,248,31,248,30,7,31,58,31,25,31,205,31,240,31,106,31,194,31,135,31,70,31,103,31,99,31,23,31,23,30,23,29,124,31,247,31,58,31,233,31,136,31,147,31,147,30,96,31,70,31,171,31,140,31,210,31,122,31,138,31,138,30,8,31,112,31,112,30,65,31,65,30,57,31,138,31,144,31,144,30,185,31,110,31,110,30,240,31,229,31,133,31,118,31,33,31,33,30,255,31,237,31,53,31,140,31,142,31,243,31,169,31,240,31,69,31,69,30,87,31,229,31,229,30,182,31,123,31,234,31,234,30,192,31,192,30,132,31,132,30,122,31,184,31,245,31,229,31,110,31,110,30,63,31,138,31,183,31,183,30,138,31,187,31,125,31,199,31,62,31,50,31,50,30,117,31,102,31,153,31,90,31,131,31,82,31,82,30,154,31,124,31,232,31,7,31,153,31,65,31,233,31,135,31,203,31,210,31,131,31,131,30,195,31,41,31,46,31,96,31,96,31,96,30,96,29,154,31,191,31,87,31,111,31,255,31,231,31,17,31,253,31,198,31,120,31,63,31,23,31,126,31,99,31,99,30,99,29,65,31,198,31,140,31,223,31,223,30,223,29,118,31,81,31,87,31,56,31,174,31,174,30,174,29,205,31,205,30,224,31,235,31,235,30,209,31,175,31,1,31,186,31,64,31,58,31,218,31,218,30,47,31,117,31,97,31,86,31,132,31,132,30,238,31,102,31,4,31,245,31,245,30,249,31,249,30,179,31,148,31,194,31,194,30,69,31,232,31,11,31,148,31,12,31,198,31,166,31,152,31,248,31,4,31,77,31,213,31,61,31,133,31,214,31,7,31,22,31,167,31,167,30,30,31,30,30,30,29,30,28,100,31,52,31,52,30,117,31,117,30,117,29,35,31,231,31,12,31,12,30,12,29,226,31,194,31,194,30,218,31,41,31,196,31,168,31,115,31,180,31,56,31,60,31,205,31,46,31,96,31,100,31,198,31,18,31,92,31,82,31,121,31,77,31,210,31,67,31,101,31,28,31,203,31,111,31,200,31,200,30,36,31,228,31,246,31,200,31,200,30,87,31,45,31,127,31,255,31,128,31,217,31,201,31,225,31,225,30,102,31,2,31,94,31,153,31,183,31,183,30,183,29,68,31,242,31,113,31,113,30,137,31,204,31,246,31,89,31,203,31,203,31,152,31,25,31,254,31,11,31,28,31,28,30,28,29,28,28,15,31,221,31,221,30,246,31,118,31,245,31,66,31,24,31,24,30,116,31,196,31,211,31,219,31,108,31,177,31,227,31,110,31,5,31,53,31,196,31,169,31,40,31,214,31,103,31,183,31,240,31,74,31,74,30,67,31,210,31,210,30,164,31,108,31,108,30,92,31,60,31,215,31,255,31,14,31,233,31,233,30,233,29,235,31,226,31,203,31,131,31,131,30,131,29,131,28,150,31,194,31,173,31,138,31,127,31,151,31,105,31,105,30,241,31,220,31,220,30,236,31,236,30,250,31,250,30,66,31,185,31,185,30,211,31,211,30,61,31,57,31,52,31,52,30,52,29,97,31,194,31,140,31,140,31,164,31,59,31,214,31,102,31,11,31,236,31,27,31,222,31,222,30,206,31,201,31,116,31,90,31,159,31,159,30,61,31,61,30,114,31,181,31,240,31,56,31,86,31,217,31,217,30,37,31,164,31,250,31,249,31,100,31,90,31,166,31,237,31,73,31,74,31,238,31,238,30,206,31,159,31,159,30,225,31,89,31,73,31,17,31,153,31,173,31,217,31,217,30,211,31,117,31,106,31,188,31,131,31,131,30,254,31,243,31,243,30,243,29,74,31,34,31,184,31,68,31,182,31,177,31,189,31,180,31,180,30,212,31,11,31,223,31,118,31,253,31,183,31,125,31,82,31,177,31,74,31,227,31,252,31,189,31,70,31,39,31,174,31,240,31,53,31,131,31,214,31,50,31,50,30,208,31,6,31,200,31,68,31,67,31,157,31,246,31,38,31,59,31,55,31,55,30,131,31,64,31,64,30,25,31,214,31,28,31,92,31,18,31,77,31,5,31,30,31,248,31,8,31,8,30,94,31,152,31,246,31,183,31,183,30,50,31,151,31,157,31,254,31,254,30,155,31,155,30,155,29,155,28,60,31,164,31,237,31,143,31,124,31,244,31,244,30,246,31,246,30,58,31,167,31,93,31,108,31,108,30,108,29,116,31,35,31,242,31,236,31,99,31,236,31,66,31,239,31,232,31,55,31,137,31,176,31,69,31,15,31,15,30,15,29,182,31,146,31,213,31,150,31,187,31,241,31,68,31,207,31,89,31,109,31,70,31,70,30,68,31,68,30,138,31,111,31,25,31,190,31,190,30,72,31,217,31,220,31,8,31,159,31,159,30,159,29,191,31,216,31,221,31,221,30,196,31,196,30,196,29,73,31,61,31,39,31,39,30,34,31,83,31,83,30,83,29,52,31,33,31,220,31,104,31,152,31,179,31,187,31,7,31,148,31,154,31,154,30,5,31,112,31,12,31,12,30,206,31,195,31,195,30,48,31,145,31,139,31,22,31,64,31,64,30,192,31,192,30,196,31,159,31,159,30,146,31,187,31,85,31,161,31,161,30,68,31,111,31,57,31,214,31,174,31,239,31,147,31,6,31,178,31,117,31,24,31,29,31,29,30,184,31,184,30,139,31,139,30,139,29,248,31,83,31,30,31,91,31,183,31,70,31,70,30,80,31,80,31,80,30,232,31,137,31,137,30,106,31,106,30,106,29,164,31,164,30,56,31,56,30,220,31,220,30,64,31,64,30,204,31,53,31,129,31,13,31,248,31,248,30,248,29,222,31,104,31,141,31,25,31,50,31,114,31,123,31,123,30,234,31,202,31,119,31,135,31,58,31,131,31,211,31,49,31,49,30,49,29,49,28,49,27,249,31,249,30,131,31,187,31,78,31,78,30,19,31,182,31,254,31,254,30,254,29,254,28,227,31,227,30,227,29,132,31,246,31,38,31,116,31,17,31,168,31,228,31,228,30,46,31,46,30,194,31,151,31,109,31,109,30,94,31,94,30,84,31,124,31,39,31,182,31,213,31,228,31,152,31,152,30,152,29,236,31,236,30,236,29,196,31,41,31,40,31,71,31,63,31,154,31,156,31,156,30,156,29,125,31,226,31,165,31,165,30,29,31,49,31,49,30,49,29,164,31,22,31,77,31,77,30,77,29,160,31,160,30,20,31,20,30,130,31,173,31,217,31,98,31,63,31,97,31,237,31,48,31,18,31,210,31,244,31,179,31,68,31,101,31,72,31,8,31,145,31,208,31,208,30,106,31,232,31,232,30,18,31,164,31,164,30,112,31,12,31,114,31,48,31,148,31,226,31,255,31,70,31,2,31,205,31,222,31,203,31,107,31,96,31,61,31,61,30,61,29,233,31,98,31,98,30,62,31,62,30,197,31,107,31,150,31,95,31,184,31,194,31,36,31,243,31,107,31,206,31,81,31,81,30,21,31,23,31,205,31,205,30,205,29,42,31,22,31,12,31,47,31,234,31,254,31,216,31,216,30,23,31,52,31,12,31,233,31,126,31,179,31,112,31,144,31,100,31,224,31,9,31,50,31,99,31,99,30,109,31,109,30,64,31,75,31,180,31,93,31,160,31,17,31,228,31,56,31,234,31,234,30,234,29,57,31,57,30,57,29,57,28,195,31,46,31,63,31,42,31,234,31,251,31,22,31,22,30,132,31,173,31,144,31,246,31,204,31,158,31,57,31,65,31,122,31,243,31,94,31,38,31,234,31,246,31,246,30,98,31,252,31,165,31,143,31,143,30,103,31,35,31,134,31,59,31,67,31,96,31,191,31,219,31,103,31,103,30,106,31,183,31,183,30,183,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
