-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_714 is
end project_tb_714;

architecture project_tb_arch_714 of project_tb_714 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 613;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (222,0,169,0,239,0,227,0,0,0,21,0,205,0,0,0,33,0,0,0,152,0,158,0,206,0,202,0,112,0,112,0,0,0,216,0,37,0,0,0,77,0,197,0,117,0,77,0,0,0,16,0,225,0,243,0,79,0,0,0,110,0,211,0,44,0,208,0,21,0,123,0,163,0,15,0,156,0,135,0,213,0,0,0,115,0,26,0,79,0,194,0,164,0,163,0,67,0,224,0,0,0,132,0,167,0,78,0,211,0,232,0,0,0,38,0,103,0,63,0,0,0,161,0,42,0,68,0,65,0,48,0,181,0,120,0,174,0,0,0,0,0,106,0,0,0,0,0,0,0,84,0,223,0,0,0,56,0,0,0,16,0,37,0,0,0,119,0,183,0,201,0,0,0,31,0,50,0,171,0,92,0,73,0,215,0,0,0,253,0,150,0,138,0,62,0,8,0,200,0,38,0,1,0,54,0,243,0,208,0,0,0,113,0,36,0,235,0,155,0,0,0,143,0,166,0,148,0,221,0,254,0,226,0,180,0,18,0,254,0,0,0,141,0,120,0,0,0,69,0,240,0,0,0,249,0,110,0,39,0,0,0,102,0,122,0,35,0,0,0,60,0,99,0,23,0,170,0,11,0,65,0,167,0,0,0,0,0,157,0,90,0,167,0,61,0,202,0,120,0,204,0,151,0,93,0,68,0,126,0,34,0,177,0,83,0,0,0,209,0,255,0,93,0,84,0,167,0,169,0,82,0,22,0,28,0,94,0,120,0,9,0,69,0,112,0,0,0,0,0,239,0,168,0,187,0,124,0,41,0,213,0,0,0,54,0,0,0,78,0,93,0,200,0,104,0,0,0,41,0,208,0,83,0,1,0,0,0,71,0,0,0,117,0,15,0,72,0,209,0,0,0,151,0,247,0,190,0,0,0,0,0,57,0,74,0,240,0,55,0,89,0,72,0,245,0,86,0,0,0,59,0,210,0,59,0,152,0,6,0,245,0,251,0,101,0,124,0,0,0,201,0,187,0,9,0,125,0,253,0,0,0,175,0,0,0,24,0,71,0,158,0,86,0,251,0,0,0,236,0,158,0,45,0,163,0,0,0,80,0,184,0,12,0,36,0,127,0,155,0,220,0,222,0,119,0,44,0,0,0,0,0,99,0,229,0,163,0,114,0,21,0,98,0,35,0,0,0,41,0,0,0,12,0,183,0,76,0,16,0,55,0,245,0,139,0,198,0,240,0,93,0,27,0,0,0,0,0,70,0,240,0,182,0,0,0,0,0,45,0,104,0,24,0,78,0,0,0,84,0,165,0,153,0,140,0,89,0,123,0,0,0,10,0,25,0,16,0,83,0,140,0,191,0,220,0,255,0,0,0,0,0,57,0,210,0,245,0,0,0,62,0,192,0,110,0,168,0,176,0,0,0,181,0,212,0,0,0,0,0,184,0,194,0,181,0,197,0,126,0,92,0,0,0,0,0,5,0,19,0,60,0,111,0,25,0,236,0,167,0,220,0,0,0,97,0,0,0,0,0,70,0,95,0,76,0,244,0,0,0,29,0,0,0,158,0,161,0,32,0,228,0,10,0,89,0,235,0,83,0,177,0,17,0,163,0,232,0,136,0,69,0,35,0,0,0,159,0,228,0,38,0,106,0,162,0,129,0,0,0,0,0,228,0,159,0,3,0,11,0,12,0,10,0,0,0,46,0,206,0,0,0,0,0,32,0,90,0,26,0,109,0,178,0,20,0,44,0,0,0,34,0,0,0,173,0,180,0,142,0,195,0,87,0,0,0,27,0,150,0,255,0,253,0,110,0,133,0,0,0,17,0,89,0,227,0,210,0,198,0,9,0,85,0,83,0,47,0,21,0,11,0,0,0,138,0,122,0,244,0,147,0,252,0,0,0,85,0,0,0,0,0,179,0,106,0,0,0,144,0,31,0,207,0,63,0,217,0,239,0,127,0,239,0,45,0,242,0,7,0,151,0,0,0,12,0,57,0,229,0,173,0,95,0,185,0,27,0,194,0,77,0,92,0,206,0,156,0,111,0,179,0,0,0,0,0,13,0,79,0,85,0,0,0,253,0,0,0,161,0,201,0,131,0,156,0,165,0,0,0,120,0,58,0,50,0,69,0,254,0,244,0,81,0,35,0,217,0,232,0,76,0,67,0,0,0,160,0,47,0,63,0,44,0,0,0,23,0,142,0,0,0,0,0,0,0,0,0,133,0,51,0,246,0,234,0,184,0,34,0,89,0,40,0,0,0,59,0,123,0,200,0,0,0,0,0,133,0,69,0,0,0,127,0,46,0,113,0,10,0,163,0,134,0,42,0,0,0,47,0,241,0,92,0,163,0,0,0,122,0,0,0,94,0,78,0,67,0,86,0,200,0,208,0,76,0,11,0,121,0,203,0,71,0,224,0,0,0,187,0,0,0,170,0,0,0,88,0,175,0,125,0,38,0,84,0,126,0,91,0,0,0,95,0,181,0,69,0,126,0,159,0,183,0,208,0,0,0,35,0,226,0,67,0,79,0,73,0,218,0,0,0,0,0,0,0,242,0,154,0,31,0,0,0,0,0,49,0,135,0,44,0,0,0,136,0,181,0,74,0,61,0,61,0,144,0,228,0,210,0,225,0,251,0,133,0,202,0,225,0,212,0,0,0,13,0,53,0,68,0,0,0,50,0,60,0,62,0,187,0,16,0,34,0,34,0,143,0,200,0,93,0,0,0,0,0,14,0,56,0,137,0,21,0,122,0);
signal scenario_full  : scenario_type := (222,31,169,31,239,31,227,31,227,30,21,31,205,31,205,30,33,31,33,30,152,31,158,31,206,31,202,31,112,31,112,31,112,30,216,31,37,31,37,30,77,31,197,31,117,31,77,31,77,30,16,31,225,31,243,31,79,31,79,30,110,31,211,31,44,31,208,31,21,31,123,31,163,31,15,31,156,31,135,31,213,31,213,30,115,31,26,31,79,31,194,31,164,31,163,31,67,31,224,31,224,30,132,31,167,31,78,31,211,31,232,31,232,30,38,31,103,31,63,31,63,30,161,31,42,31,68,31,65,31,48,31,181,31,120,31,174,31,174,30,174,29,106,31,106,30,106,29,106,28,84,31,223,31,223,30,56,31,56,30,16,31,37,31,37,30,119,31,183,31,201,31,201,30,31,31,50,31,171,31,92,31,73,31,215,31,215,30,253,31,150,31,138,31,62,31,8,31,200,31,38,31,1,31,54,31,243,31,208,31,208,30,113,31,36,31,235,31,155,31,155,30,143,31,166,31,148,31,221,31,254,31,226,31,180,31,18,31,254,31,254,30,141,31,120,31,120,30,69,31,240,31,240,30,249,31,110,31,39,31,39,30,102,31,122,31,35,31,35,30,60,31,99,31,23,31,170,31,11,31,65,31,167,31,167,30,167,29,157,31,90,31,167,31,61,31,202,31,120,31,204,31,151,31,93,31,68,31,126,31,34,31,177,31,83,31,83,30,209,31,255,31,93,31,84,31,167,31,169,31,82,31,22,31,28,31,94,31,120,31,9,31,69,31,112,31,112,30,112,29,239,31,168,31,187,31,124,31,41,31,213,31,213,30,54,31,54,30,78,31,93,31,200,31,104,31,104,30,41,31,208,31,83,31,1,31,1,30,71,31,71,30,117,31,15,31,72,31,209,31,209,30,151,31,247,31,190,31,190,30,190,29,57,31,74,31,240,31,55,31,89,31,72,31,245,31,86,31,86,30,59,31,210,31,59,31,152,31,6,31,245,31,251,31,101,31,124,31,124,30,201,31,187,31,9,31,125,31,253,31,253,30,175,31,175,30,24,31,71,31,158,31,86,31,251,31,251,30,236,31,158,31,45,31,163,31,163,30,80,31,184,31,12,31,36,31,127,31,155,31,220,31,222,31,119,31,44,31,44,30,44,29,99,31,229,31,163,31,114,31,21,31,98,31,35,31,35,30,41,31,41,30,12,31,183,31,76,31,16,31,55,31,245,31,139,31,198,31,240,31,93,31,27,31,27,30,27,29,70,31,240,31,182,31,182,30,182,29,45,31,104,31,24,31,78,31,78,30,84,31,165,31,153,31,140,31,89,31,123,31,123,30,10,31,25,31,16,31,83,31,140,31,191,31,220,31,255,31,255,30,255,29,57,31,210,31,245,31,245,30,62,31,192,31,110,31,168,31,176,31,176,30,181,31,212,31,212,30,212,29,184,31,194,31,181,31,197,31,126,31,92,31,92,30,92,29,5,31,19,31,60,31,111,31,25,31,236,31,167,31,220,31,220,30,97,31,97,30,97,29,70,31,95,31,76,31,244,31,244,30,29,31,29,30,158,31,161,31,32,31,228,31,10,31,89,31,235,31,83,31,177,31,17,31,163,31,232,31,136,31,69,31,35,31,35,30,159,31,228,31,38,31,106,31,162,31,129,31,129,30,129,29,228,31,159,31,3,31,11,31,12,31,10,31,10,30,46,31,206,31,206,30,206,29,32,31,90,31,26,31,109,31,178,31,20,31,44,31,44,30,34,31,34,30,173,31,180,31,142,31,195,31,87,31,87,30,27,31,150,31,255,31,253,31,110,31,133,31,133,30,17,31,89,31,227,31,210,31,198,31,9,31,85,31,83,31,47,31,21,31,11,31,11,30,138,31,122,31,244,31,147,31,252,31,252,30,85,31,85,30,85,29,179,31,106,31,106,30,144,31,31,31,207,31,63,31,217,31,239,31,127,31,239,31,45,31,242,31,7,31,151,31,151,30,12,31,57,31,229,31,173,31,95,31,185,31,27,31,194,31,77,31,92,31,206,31,156,31,111,31,179,31,179,30,179,29,13,31,79,31,85,31,85,30,253,31,253,30,161,31,201,31,131,31,156,31,165,31,165,30,120,31,58,31,50,31,69,31,254,31,244,31,81,31,35,31,217,31,232,31,76,31,67,31,67,30,160,31,47,31,63,31,44,31,44,30,23,31,142,31,142,30,142,29,142,28,142,27,133,31,51,31,246,31,234,31,184,31,34,31,89,31,40,31,40,30,59,31,123,31,200,31,200,30,200,29,133,31,69,31,69,30,127,31,46,31,113,31,10,31,163,31,134,31,42,31,42,30,47,31,241,31,92,31,163,31,163,30,122,31,122,30,94,31,78,31,67,31,86,31,200,31,208,31,76,31,11,31,121,31,203,31,71,31,224,31,224,30,187,31,187,30,170,31,170,30,88,31,175,31,125,31,38,31,84,31,126,31,91,31,91,30,95,31,181,31,69,31,126,31,159,31,183,31,208,31,208,30,35,31,226,31,67,31,79,31,73,31,218,31,218,30,218,29,218,28,242,31,154,31,31,31,31,30,31,29,49,31,135,31,44,31,44,30,136,31,181,31,74,31,61,31,61,31,144,31,228,31,210,31,225,31,251,31,133,31,202,31,225,31,212,31,212,30,13,31,53,31,68,31,68,30,50,31,60,31,62,31,187,31,16,31,34,31,34,31,143,31,200,31,93,31,93,30,93,29,14,31,56,31,137,31,21,31,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
