-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_592 is
end project_tb_592;

architecture project_tb_arch_592 of project_tb_592 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 509;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (131,0,122,0,0,0,0,0,41,0,168,0,7,0,0,0,142,0,249,0,0,0,119,0,122,0,112,0,157,0,0,0,135,0,132,0,0,0,29,0,143,0,0,0,117,0,110,0,217,0,114,0,202,0,181,0,28,0,0,0,53,0,218,0,142,0,169,0,90,0,52,0,30,0,0,0,95,0,4,0,207,0,0,0,109,0,95,0,85,0,245,0,161,0,251,0,151,0,252,0,0,0,221,0,150,0,213,0,11,0,0,0,0,0,141,0,104,0,65,0,144,0,0,0,68,0,82,0,175,0,0,0,144,0,175,0,125,0,31,0,0,0,0,0,0,0,173,0,18,0,0,0,65,0,254,0,0,0,169,0,0,0,0,0,146,0,0,0,17,0,234,0,69,0,235,0,105,0,0,0,67,0,144,0,94,0,49,0,81,0,37,0,206,0,0,0,130,0,107,0,154,0,196,0,197,0,201,0,143,0,144,0,0,0,0,0,83,0,189,0,18,0,4,0,199,0,86,0,0,0,29,0,120,0,47,0,30,0,8,0,16,0,112,0,0,0,151,0,0,0,52,0,155,0,139,0,157,0,151,0,121,0,204,0,94,0,161,0,30,0,31,0,42,0,41,0,0,0,182,0,25,0,240,0,114,0,121,0,0,0,197,0,29,0,244,0,0,0,0,0,0,0,144,0,16,0,42,0,0,0,139,0,47,0,205,0,246,0,175,0,113,0,209,0,0,0,20,0,45,0,70,0,14,0,80,0,220,0,205,0,174,0,58,0,0,0,169,0,52,0,193,0,0,0,191,0,0,0,214,0,56,0,199,0,0,0,81,0,151,0,245,0,95,0,98,0,122,0,232,0,0,0,253,0,232,0,21,0,203,0,252,0,0,0,45,0,17,0,53,0,176,0,27,0,169,0,231,0,240,0,252,0,135,0,167,0,149,0,0,0,0,0,52,0,98,0,88,0,188,0,64,0,77,0,0,0,165,0,209,0,102,0,171,0,0,0,0,0,105,0,128,0,0,0,179,0,64,0,129,0,0,0,64,0,215,0,187,0,137,0,42,0,202,0,214,0,19,0,110,0,89,0,181,0,226,0,101,0,0,0,138,0,218,0,160,0,166,0,68,0,0,0,0,0,64,0,165,0,238,0,9,0,23,0,194,0,178,0,200,0,218,0,0,0,136,0,0,0,0,0,202,0,208,0,227,0,151,0,197,0,246,0,52,0,158,0,156,0,19,0,133,0,0,0,209,0,155,0,0,0,198,0,53,0,166,0,54,0,213,0,46,0,240,0,236,0,157,0,67,0,114,0,100,0,1,0,198,0,185,0,161,0,251,0,84,0,0,0,47,0,245,0,0,0,114,0,143,0,191,0,171,0,0,0,92,0,67,0,124,0,205,0,53,0,132,0,86,0,0,0,21,0,56,0,11,0,10,0,37,0,44,0,116,0,45,0,89,0,70,0,130,0,41,0,74,0,221,0,52,0,156,0,41,0,86,0,0,0,0,0,116,0,104,0,191,0,78,0,167,0,37,0,124,0,232,0,0,0,166,0,0,0,106,0,50,0,0,0,225,0,218,0,136,0,214,0,87,0,0,0,154,0,255,0,243,0,2,0,0,0,65,0,209,0,179,0,221,0,53,0,0,0,92,0,216,0,47,0,98,0,132,0,149,0,0,0,36,0,0,0,110,0,0,0,0,0,169,0,191,0,152,0,110,0,31,0,12,0,234,0,17,0,106,0,0,0,0,0,168,0,14,0,80,0,118,0,21,0,227,0,198,0,101,0,228,0,0,0,100,0,59,0,246,0,17,0,19,0,145,0,0,0,51,0,93,0,194,0,41,0,225,0,102,0,110,0,248,0,74,0,123,0,95,0,127,0,35,0,200,0,192,0,45,0,12,0,221,0,0,0,195,0,135,0,0,0,69,0,23,0,9,0,0,0,0,0,0,0,178,0,222,0,152,0,83,0,152,0,61,0,0,0,228,0,61,0,150,0,238,0,217,0,8,0,52,0,49,0,0,0,162,0,117,0,64,0,0,0,238,0,150,0,81,0,230,0,0,0,72,0,49,0,44,0,48,0,0,0,97,0,0,0,124,0,59,0,0,0,36,0,209,0,118,0,119,0,15,0,128,0,8,0,0,0,73,0,0,0,242,0,49,0,216,0,136,0,172,0,141,0,6,0,35,0,225,0,141,0,171,0,208,0,177,0,197,0,230,0,187,0,49,0,205,0,221,0,216,0,220,0,197,0,123,0,0,0,20,0,195,0,87,0,65,0,119,0,83,0);
signal scenario_full  : scenario_type := (131,31,122,31,122,30,122,29,41,31,168,31,7,31,7,30,142,31,249,31,249,30,119,31,122,31,112,31,157,31,157,30,135,31,132,31,132,30,29,31,143,31,143,30,117,31,110,31,217,31,114,31,202,31,181,31,28,31,28,30,53,31,218,31,142,31,169,31,90,31,52,31,30,31,30,30,95,31,4,31,207,31,207,30,109,31,95,31,85,31,245,31,161,31,251,31,151,31,252,31,252,30,221,31,150,31,213,31,11,31,11,30,11,29,141,31,104,31,65,31,144,31,144,30,68,31,82,31,175,31,175,30,144,31,175,31,125,31,31,31,31,30,31,29,31,28,173,31,18,31,18,30,65,31,254,31,254,30,169,31,169,30,169,29,146,31,146,30,17,31,234,31,69,31,235,31,105,31,105,30,67,31,144,31,94,31,49,31,81,31,37,31,206,31,206,30,130,31,107,31,154,31,196,31,197,31,201,31,143,31,144,31,144,30,144,29,83,31,189,31,18,31,4,31,199,31,86,31,86,30,29,31,120,31,47,31,30,31,8,31,16,31,112,31,112,30,151,31,151,30,52,31,155,31,139,31,157,31,151,31,121,31,204,31,94,31,161,31,30,31,31,31,42,31,41,31,41,30,182,31,25,31,240,31,114,31,121,31,121,30,197,31,29,31,244,31,244,30,244,29,244,28,144,31,16,31,42,31,42,30,139,31,47,31,205,31,246,31,175,31,113,31,209,31,209,30,20,31,45,31,70,31,14,31,80,31,220,31,205,31,174,31,58,31,58,30,169,31,52,31,193,31,193,30,191,31,191,30,214,31,56,31,199,31,199,30,81,31,151,31,245,31,95,31,98,31,122,31,232,31,232,30,253,31,232,31,21,31,203,31,252,31,252,30,45,31,17,31,53,31,176,31,27,31,169,31,231,31,240,31,252,31,135,31,167,31,149,31,149,30,149,29,52,31,98,31,88,31,188,31,64,31,77,31,77,30,165,31,209,31,102,31,171,31,171,30,171,29,105,31,128,31,128,30,179,31,64,31,129,31,129,30,64,31,215,31,187,31,137,31,42,31,202,31,214,31,19,31,110,31,89,31,181,31,226,31,101,31,101,30,138,31,218,31,160,31,166,31,68,31,68,30,68,29,64,31,165,31,238,31,9,31,23,31,194,31,178,31,200,31,218,31,218,30,136,31,136,30,136,29,202,31,208,31,227,31,151,31,197,31,246,31,52,31,158,31,156,31,19,31,133,31,133,30,209,31,155,31,155,30,198,31,53,31,166,31,54,31,213,31,46,31,240,31,236,31,157,31,67,31,114,31,100,31,1,31,198,31,185,31,161,31,251,31,84,31,84,30,47,31,245,31,245,30,114,31,143,31,191,31,171,31,171,30,92,31,67,31,124,31,205,31,53,31,132,31,86,31,86,30,21,31,56,31,11,31,10,31,37,31,44,31,116,31,45,31,89,31,70,31,130,31,41,31,74,31,221,31,52,31,156,31,41,31,86,31,86,30,86,29,116,31,104,31,191,31,78,31,167,31,37,31,124,31,232,31,232,30,166,31,166,30,106,31,50,31,50,30,225,31,218,31,136,31,214,31,87,31,87,30,154,31,255,31,243,31,2,31,2,30,65,31,209,31,179,31,221,31,53,31,53,30,92,31,216,31,47,31,98,31,132,31,149,31,149,30,36,31,36,30,110,31,110,30,110,29,169,31,191,31,152,31,110,31,31,31,12,31,234,31,17,31,106,31,106,30,106,29,168,31,14,31,80,31,118,31,21,31,227,31,198,31,101,31,228,31,228,30,100,31,59,31,246,31,17,31,19,31,145,31,145,30,51,31,93,31,194,31,41,31,225,31,102,31,110,31,248,31,74,31,123,31,95,31,127,31,35,31,200,31,192,31,45,31,12,31,221,31,221,30,195,31,135,31,135,30,69,31,23,31,9,31,9,30,9,29,9,28,178,31,222,31,152,31,83,31,152,31,61,31,61,30,228,31,61,31,150,31,238,31,217,31,8,31,52,31,49,31,49,30,162,31,117,31,64,31,64,30,238,31,150,31,81,31,230,31,230,30,72,31,49,31,44,31,48,31,48,30,97,31,97,30,124,31,59,31,59,30,36,31,209,31,118,31,119,31,15,31,128,31,8,31,8,30,73,31,73,30,242,31,49,31,216,31,136,31,172,31,141,31,6,31,35,31,225,31,141,31,171,31,208,31,177,31,197,31,230,31,187,31,49,31,205,31,221,31,216,31,220,31,197,31,123,31,123,30,20,31,195,31,87,31,65,31,119,31,83,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
