-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 341;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (5,0,254,0,157,0,4,0,61,0,11,0,129,0,49,0,255,0,234,0,0,0,190,0,0,0,95,0,170,0,137,0,199,0,98,0,86,0,25,0,0,0,0,0,244,0,242,0,55,0,0,0,205,0,226,0,183,0,218,0,0,0,78,0,120,0,194,0,236,0,0,0,0,0,0,0,130,0,241,0,215,0,177,0,135,0,242,0,91,0,218,0,192,0,153,0,0,0,243,0,199,0,21,0,162,0,16,0,0,0,0,0,166,0,0,0,0,0,228,0,40,0,89,0,105,0,92,0,216,0,222,0,130,0,0,0,246,0,21,0,138,0,155,0,0,0,92,0,90,0,185,0,183,0,104,0,13,0,3,0,115,0,255,0,189,0,117,0,180,0,13,0,30,0,39,0,203,0,229,0,212,0,0,0,253,0,96,0,0,0,236,0,0,0,0,0,57,0,120,0,53,0,39,0,33,0,0,0,251,0,192,0,118,0,0,0,127,0,179,0,96,0,177,0,40,0,16,0,164,0,126,0,9,0,94,0,108,0,0,0,0,0,7,0,0,0,55,0,58,0,0,0,0,0,75,0,243,0,74,0,0,0,7,0,14,0,112,0,8,0,0,0,0,0,129,0,13,0,113,0,0,0,0,0,22,0,0,0,127,0,40,0,225,0,0,0,79,0,107,0,239,0,38,0,169,0,0,0,18,0,0,0,4,0,0,0,24,0,24,0,94,0,100,0,49,0,161,0,0,0,174,0,44,0,0,0,0,0,211,0,0,0,222,0,149,0,177,0,213,0,41,0,65,0,0,0,114,0,250,0,70,0,88,0,195,0,0,0,45,0,0,0,193,0,0,0,39,0,0,0,201,0,0,0,66,0,34,0,5,0,238,0,119,0,101,0,78,0,125,0,98,0,74,0,187,0,101,0,0,0,42,0,42,0,169,0,0,0,136,0,249,0,206,0,0,0,240,0,15,0,0,0,0,0,236,0,239,0,23,0,0,0,187,0,0,0,200,0,146,0,172,0,65,0,110,0,0,0,80,0,0,0,128,0,248,0,0,0,89,0,109,0,95,0,107,0,0,0,105,0,100,0,49,0,123,0,97,0,75,0,0,0,249,0,0,0,174,0,0,0,113,0,67,0,0,0,253,0,220,0,41,0,31,0,235,0,0,0,218,0,0,0,254,0,244,0,176,0,209,0,0,0,206,0,91,0,237,0,0,0,59,0,251,0,129,0,254,0,146,0,0,0,140,0,95,0,0,0,215,0,165,0,214,0,138,0,184,0,29,0,214,0,243,0,139,0,196,0,157,0,216,0,18,0,127,0,40,0,205,0,71,0,0,0,215,0,180,0,70,0,244,0,162,0,81,0,193,0,48,0,44,0,19,0,216,0,203,0,106,0,154,0,165,0,188,0,71,0,212,0,159,0,62,0,0,0,18,0,247,0,126,0,6,0,0,0,212,0,0,0,0,0,0,0,86,0,202,0,63,0,106,0,178,0,126,0,63,0,102,0,0,0,135,0,175,0,219,0,61,0,2,0);
signal scenario_full  : scenario_type := (5,31,254,31,157,31,4,31,61,31,11,31,129,31,49,31,255,31,234,31,234,30,190,31,190,30,95,31,170,31,137,31,199,31,98,31,86,31,25,31,25,30,25,29,244,31,242,31,55,31,55,30,205,31,226,31,183,31,218,31,218,30,78,31,120,31,194,31,236,31,236,30,236,29,236,28,130,31,241,31,215,31,177,31,135,31,242,31,91,31,218,31,192,31,153,31,153,30,243,31,199,31,21,31,162,31,16,31,16,30,16,29,166,31,166,30,166,29,228,31,40,31,89,31,105,31,92,31,216,31,222,31,130,31,130,30,246,31,21,31,138,31,155,31,155,30,92,31,90,31,185,31,183,31,104,31,13,31,3,31,115,31,255,31,189,31,117,31,180,31,13,31,30,31,39,31,203,31,229,31,212,31,212,30,253,31,96,31,96,30,236,31,236,30,236,29,57,31,120,31,53,31,39,31,33,31,33,30,251,31,192,31,118,31,118,30,127,31,179,31,96,31,177,31,40,31,16,31,164,31,126,31,9,31,94,31,108,31,108,30,108,29,7,31,7,30,55,31,58,31,58,30,58,29,75,31,243,31,74,31,74,30,7,31,14,31,112,31,8,31,8,30,8,29,129,31,13,31,113,31,113,30,113,29,22,31,22,30,127,31,40,31,225,31,225,30,79,31,107,31,239,31,38,31,169,31,169,30,18,31,18,30,4,31,4,30,24,31,24,31,94,31,100,31,49,31,161,31,161,30,174,31,44,31,44,30,44,29,211,31,211,30,222,31,149,31,177,31,213,31,41,31,65,31,65,30,114,31,250,31,70,31,88,31,195,31,195,30,45,31,45,30,193,31,193,30,39,31,39,30,201,31,201,30,66,31,34,31,5,31,238,31,119,31,101,31,78,31,125,31,98,31,74,31,187,31,101,31,101,30,42,31,42,31,169,31,169,30,136,31,249,31,206,31,206,30,240,31,15,31,15,30,15,29,236,31,239,31,23,31,23,30,187,31,187,30,200,31,146,31,172,31,65,31,110,31,110,30,80,31,80,30,128,31,248,31,248,30,89,31,109,31,95,31,107,31,107,30,105,31,100,31,49,31,123,31,97,31,75,31,75,30,249,31,249,30,174,31,174,30,113,31,67,31,67,30,253,31,220,31,41,31,31,31,235,31,235,30,218,31,218,30,254,31,244,31,176,31,209,31,209,30,206,31,91,31,237,31,237,30,59,31,251,31,129,31,254,31,146,31,146,30,140,31,95,31,95,30,215,31,165,31,214,31,138,31,184,31,29,31,214,31,243,31,139,31,196,31,157,31,216,31,18,31,127,31,40,31,205,31,71,31,71,30,215,31,180,31,70,31,244,31,162,31,81,31,193,31,48,31,44,31,19,31,216,31,203,31,106,31,154,31,165,31,188,31,71,31,212,31,159,31,62,31,62,30,18,31,247,31,126,31,6,31,6,30,212,31,212,30,212,29,212,28,86,31,202,31,63,31,106,31,178,31,126,31,63,31,102,31,102,30,135,31,175,31,219,31,61,31,2,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
