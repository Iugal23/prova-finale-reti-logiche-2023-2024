-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_697 is
end project_tb_697;

architecture project_tb_arch_697 of project_tb_697 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 290;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,55,0,229,0,214,0,0,0,81,0,16,0,30,0,153,0,18,0,38,0,221,0,225,0,206,0,11,0,0,0,192,0,131,0,205,0,63,0,204,0,69,0,202,0,240,0,224,0,223,0,66,0,65,0,0,0,0,0,248,0,0,0,243,0,0,0,7,0,0,0,92,0,238,0,126,0,136,0,16,0,0,0,149,0,212,0,74,0,84,0,161,0,75,0,83,0,137,0,29,0,156,0,143,0,100,0,0,0,0,0,238,0,201,0,0,0,36,0,93,0,0,0,226,0,0,0,212,0,51,0,143,0,41,0,5,0,130,0,253,0,0,0,254,0,0,0,170,0,64,0,186,0,122,0,135,0,215,0,240,0,95,0,60,0,255,0,41,0,0,0,0,0,227,0,19,0,75,0,247,0,0,0,18,0,0,0,64,0,0,0,0,0,0,0,4,0,129,0,34,0,0,0,105,0,191,0,37,0,78,0,58,0,0,0,13,0,62,0,242,0,104,0,0,0,108,0,231,0,114,0,143,0,0,0,201,0,89,0,73,0,29,0,142,0,41,0,44,0,0,0,0,0,184,0,14,0,201,0,0,0,138,0,144,0,0,0,0,0,193,0,41,0,139,0,190,0,52,0,96,0,222,0,28,0,0,0,231,0,44,0,53,0,29,0,112,0,0,0,137,0,15,0,139,0,0,0,227,0,190,0,124,0,252,0,115,0,227,0,0,0,11,0,255,0,60,0,70,0,122,0,70,0,0,0,0,0,72,0,204,0,20,0,236,0,225,0,61,0,37,0,138,0,0,0,153,0,0,0,114,0,139,0,175,0,224,0,63,0,17,0,0,0,37,0,39,0,150,0,92,0,2,0,0,0,10,0,196,0,218,0,0,0,24,0,27,0,191,0,76,0,161,0,36,0,199,0,137,0,0,0,0,0,229,0,218,0,144,0,0,0,35,0,95,0,0,0,0,0,50,0,167,0,234,0,133,0,163,0,188,0,191,0,0,0,145,0,122,0,101,0,100,0,211,0,10,0,121,0,228,0,80,0,136,0,130,0,0,0,0,0,30,0,23,0,19,0,0,0,160,0,255,0,95,0,29,0,0,0,143,0,124,0,147,0,216,0,0,0,95,0,0,0,230,0,30,0,243,0,0,0,240,0,120,0,26,0,0,0,117,0,233,0,95,0,0,0,2,0,192,0,0,0,240,0,36,0,109,0,0,0,0,0,204,0,0,0,172,0,0,0,0,0,0,0,167,0,205,0,94,0,0,0,158,0,166,0,0,0,28,0,165,0,0,0,151,0,38,0);
signal scenario_full  : scenario_type := (201,31,55,31,229,31,214,31,214,30,81,31,16,31,30,31,153,31,18,31,38,31,221,31,225,31,206,31,11,31,11,30,192,31,131,31,205,31,63,31,204,31,69,31,202,31,240,31,224,31,223,31,66,31,65,31,65,30,65,29,248,31,248,30,243,31,243,30,7,31,7,30,92,31,238,31,126,31,136,31,16,31,16,30,149,31,212,31,74,31,84,31,161,31,75,31,83,31,137,31,29,31,156,31,143,31,100,31,100,30,100,29,238,31,201,31,201,30,36,31,93,31,93,30,226,31,226,30,212,31,51,31,143,31,41,31,5,31,130,31,253,31,253,30,254,31,254,30,170,31,64,31,186,31,122,31,135,31,215,31,240,31,95,31,60,31,255,31,41,31,41,30,41,29,227,31,19,31,75,31,247,31,247,30,18,31,18,30,64,31,64,30,64,29,64,28,4,31,129,31,34,31,34,30,105,31,191,31,37,31,78,31,58,31,58,30,13,31,62,31,242,31,104,31,104,30,108,31,231,31,114,31,143,31,143,30,201,31,89,31,73,31,29,31,142,31,41,31,44,31,44,30,44,29,184,31,14,31,201,31,201,30,138,31,144,31,144,30,144,29,193,31,41,31,139,31,190,31,52,31,96,31,222,31,28,31,28,30,231,31,44,31,53,31,29,31,112,31,112,30,137,31,15,31,139,31,139,30,227,31,190,31,124,31,252,31,115,31,227,31,227,30,11,31,255,31,60,31,70,31,122,31,70,31,70,30,70,29,72,31,204,31,20,31,236,31,225,31,61,31,37,31,138,31,138,30,153,31,153,30,114,31,139,31,175,31,224,31,63,31,17,31,17,30,37,31,39,31,150,31,92,31,2,31,2,30,10,31,196,31,218,31,218,30,24,31,27,31,191,31,76,31,161,31,36,31,199,31,137,31,137,30,137,29,229,31,218,31,144,31,144,30,35,31,95,31,95,30,95,29,50,31,167,31,234,31,133,31,163,31,188,31,191,31,191,30,145,31,122,31,101,31,100,31,211,31,10,31,121,31,228,31,80,31,136,31,130,31,130,30,130,29,30,31,23,31,19,31,19,30,160,31,255,31,95,31,29,31,29,30,143,31,124,31,147,31,216,31,216,30,95,31,95,30,230,31,30,31,243,31,243,30,240,31,120,31,26,31,26,30,117,31,233,31,95,31,95,30,2,31,192,31,192,30,240,31,36,31,109,31,109,30,109,29,204,31,204,30,172,31,172,30,172,29,172,28,167,31,205,31,94,31,94,30,158,31,166,31,166,30,28,31,165,31,165,30,151,31,38,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
