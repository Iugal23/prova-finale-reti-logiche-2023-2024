-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 326;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (160,0,83,0,150,0,166,0,126,0,116,0,252,0,0,0,144,0,217,0,0,0,2,0,115,0,189,0,244,0,79,0,0,0,0,0,13,0,31,0,73,0,0,0,0,0,0,0,0,0,0,0,36,0,0,0,81,0,48,0,74,0,0,0,78,0,135,0,0,0,149,0,104,0,205,0,0,0,130,0,100,0,0,0,99,0,0,0,61,0,74,0,0,0,56,0,0,0,0,0,87,0,13,0,0,0,253,0,70,0,0,0,111,0,116,0,0,0,59,0,194,0,67,0,30,0,225,0,118,0,87,0,0,0,0,0,0,0,108,0,85,0,36,0,178,0,10,0,0,0,17,0,187,0,70,0,0,0,64,0,0,0,0,0,162,0,96,0,0,0,94,0,0,0,188,0,66,0,118,0,247,0,0,0,6,0,51,0,0,0,0,0,190,0,155,0,155,0,77,0,146,0,141,0,32,0,65,0,56,0,75,0,0,0,16,0,136,0,179,0,0,0,0,0,72,0,206,0,3,0,133,0,52,0,0,0,52,0,138,0,0,0,0,0,131,0,58,0,0,0,230,0,21,0,0,0,104,0,77,0,251,0,36,0,96,0,153,0,19,0,4,0,95,0,203,0,27,0,70,0,55,0,239,0,221,0,0,0,76,0,163,0,97,0,140,0,176,0,0,0,176,0,0,0,217,0,86,0,0,0,152,0,0,0,176,0,158,0,99,0,223,0,181,0,72,0,105,0,154,0,237,0,0,0,20,0,226,0,89,0,211,0,171,0,107,0,95,0,188,0,33,0,127,0,0,0,159,0,227,0,0,0,37,0,91,0,0,0,100,0,242,0,194,0,76,0,105,0,237,0,95,0,79,0,246,0,155,0,8,0,69,0,41,0,0,0,89,0,247,0,126,0,0,0,0,0,0,0,129,0,217,0,63,0,228,0,217,0,73,0,5,0,0,0,106,0,18,0,105,0,253,0,181,0,75,0,0,0,170,0,0,0,156,0,47,0,58,0,83,0,160,0,115,0,192,0,219,0,81,0,221,0,0,0,24,0,80,0,0,0,161,0,232,0,6,0,216,0,35,0,57,0,0,0,54,0,23,0,0,0,170,0,0,0,200,0,99,0,185,0,187,0,39,0,142,0,249,0,215,0,157,0,241,0,103,0,0,0,196,0,218,0,127,0,0,0,115,0,0,0,126,0,0,0,93,0,1,0,232,0,190,0,252,0,0,0,0,0,105,0,172,0,190,0,122,0,152,0,13,0,219,0,80,0,0,0,135,0,227,0,15,0,184,0,96,0,5,0,84,0,0,0,58,0,129,0,131,0,191,0,149,0,76,0,105,0,0,0,0,0,246,0,0,0,181,0,245,0,0,0,159,0,116,0,150,0,0,0,107,0,14,0,97,0,117,0,176,0,233,0,0,0,0,0,0,0,26,0,64,0,29,0,0,0,212,0,209,0,11,0,68,0);
signal scenario_full  : scenario_type := (160,31,83,31,150,31,166,31,126,31,116,31,252,31,252,30,144,31,217,31,217,30,2,31,115,31,189,31,244,31,79,31,79,30,79,29,13,31,31,31,73,31,73,30,73,29,73,28,73,27,73,26,36,31,36,30,81,31,48,31,74,31,74,30,78,31,135,31,135,30,149,31,104,31,205,31,205,30,130,31,100,31,100,30,99,31,99,30,61,31,74,31,74,30,56,31,56,30,56,29,87,31,13,31,13,30,253,31,70,31,70,30,111,31,116,31,116,30,59,31,194,31,67,31,30,31,225,31,118,31,87,31,87,30,87,29,87,28,108,31,85,31,36,31,178,31,10,31,10,30,17,31,187,31,70,31,70,30,64,31,64,30,64,29,162,31,96,31,96,30,94,31,94,30,188,31,66,31,118,31,247,31,247,30,6,31,51,31,51,30,51,29,190,31,155,31,155,31,77,31,146,31,141,31,32,31,65,31,56,31,75,31,75,30,16,31,136,31,179,31,179,30,179,29,72,31,206,31,3,31,133,31,52,31,52,30,52,31,138,31,138,30,138,29,131,31,58,31,58,30,230,31,21,31,21,30,104,31,77,31,251,31,36,31,96,31,153,31,19,31,4,31,95,31,203,31,27,31,70,31,55,31,239,31,221,31,221,30,76,31,163,31,97,31,140,31,176,31,176,30,176,31,176,30,217,31,86,31,86,30,152,31,152,30,176,31,158,31,99,31,223,31,181,31,72,31,105,31,154,31,237,31,237,30,20,31,226,31,89,31,211,31,171,31,107,31,95,31,188,31,33,31,127,31,127,30,159,31,227,31,227,30,37,31,91,31,91,30,100,31,242,31,194,31,76,31,105,31,237,31,95,31,79,31,246,31,155,31,8,31,69,31,41,31,41,30,89,31,247,31,126,31,126,30,126,29,126,28,129,31,217,31,63,31,228,31,217,31,73,31,5,31,5,30,106,31,18,31,105,31,253,31,181,31,75,31,75,30,170,31,170,30,156,31,47,31,58,31,83,31,160,31,115,31,192,31,219,31,81,31,221,31,221,30,24,31,80,31,80,30,161,31,232,31,6,31,216,31,35,31,57,31,57,30,54,31,23,31,23,30,170,31,170,30,200,31,99,31,185,31,187,31,39,31,142,31,249,31,215,31,157,31,241,31,103,31,103,30,196,31,218,31,127,31,127,30,115,31,115,30,126,31,126,30,93,31,1,31,232,31,190,31,252,31,252,30,252,29,105,31,172,31,190,31,122,31,152,31,13,31,219,31,80,31,80,30,135,31,227,31,15,31,184,31,96,31,5,31,84,31,84,30,58,31,129,31,131,31,191,31,149,31,76,31,105,31,105,30,105,29,246,31,246,30,181,31,245,31,245,30,159,31,116,31,150,31,150,30,107,31,14,31,97,31,117,31,176,31,233,31,233,30,233,29,233,28,26,31,64,31,29,31,29,30,212,31,209,31,11,31,68,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
