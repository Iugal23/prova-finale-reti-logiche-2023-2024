-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_723 is
end project_tb_723;

architecture project_tb_arch_723 of project_tb_723 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 812;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,157,0,40,0,92,0,7,0,0,0,79,0,34,0,0,0,191,0,64,0,74,0,47,0,0,0,0,0,156,0,46,0,0,0,154,0,109,0,197,0,18,0,215,0,7,0,129,0,120,0,226,0,14,0,158,0,170,0,0,0,165,0,253,0,90,0,0,0,143,0,0,0,199,0,250,0,100,0,186,0,34,0,162,0,143,0,0,0,4,0,56,0,0,0,215,0,247,0,187,0,24,0,224,0,206,0,0,0,87,0,63,0,64,0,73,0,0,0,214,0,45,0,0,0,113,0,146,0,218,0,0,0,170,0,0,0,0,0,85,0,51,0,159,0,17,0,167,0,230,0,135,0,0,0,45,0,239,0,135,0,0,0,48,0,0,0,196,0,0,0,0,0,173,0,222,0,37,0,87,0,39,0,220,0,0,0,230,0,131,0,130,0,242,0,176,0,0,0,98,0,112,0,15,0,0,0,120,0,16,0,17,0,26,0,246,0,64,0,132,0,188,0,244,0,227,0,226,0,231,0,0,0,154,0,0,0,216,0,162,0,114,0,114,0,222,0,247,0,189,0,97,0,220,0,0,0,139,0,87,0,0,0,125,0,0,0,53,0,2,0,189,0,61,0,0,0,28,0,133,0,232,0,0,0,11,0,192,0,199,0,0,0,10,0,60,0,137,0,61,0,113,0,58,0,152,0,92,0,47,0,0,0,0,0,127,0,30,0,214,0,108,0,243,0,10,0,14,0,129,0,6,0,142,0,52,0,199,0,69,0,53,0,135,0,0,0,0,0,227,0,150,0,0,0,93,0,116,0,95,0,92,0,37,0,0,0,191,0,40,0,238,0,177,0,196,0,242,0,211,0,240,0,103,0,252,0,83,0,176,0,128,0,0,0,66,0,20,0,27,0,158,0,30,0,146,0,175,0,90,0,233,0,98,0,142,0,125,0,69,0,153,0,11,0,247,0,249,0,15,0,94,0,28,0,177,0,230,0,53,0,131,0,108,0,248,0,16,0,184,0,191,0,147,0,239,0,148,0,199,0,144,0,208,0,114,0,19,0,130,0,239,0,157,0,156,0,0,0,69,0,198,0,166,0,17,0,0,0,143,0,0,0,132,0,164,0,117,0,0,0,6,0,29,0,177,0,0,0,45,0,11,0,158,0,59,0,138,0,106,0,0,0,24,0,239,0,0,0,0,0,50,0,0,0,160,0,242,0,137,0,37,0,159,0,0,0,63,0,128,0,187,0,0,0,144,0,0,0,196,0,191,0,212,0,148,0,0,0,0,0,96,0,197,0,0,0,0,0,124,0,24,0,19,0,169,0,174,0,246,0,171,0,0,0,145,0,5,0,122,0,120,0,73,0,148,0,121,0,251,0,169,0,0,0,199,0,106,0,9,0,186,0,252,0,118,0,165,0,62,0,211,0,101,0,44,0,187,0,0,0,78,0,0,0,0,0,60,0,141,0,239,0,232,0,142,0,175,0,0,0,165,0,5,0,114,0,140,0,145,0,201,0,241,0,90,0,203,0,206,0,133,0,187,0,0,0,0,0,47,0,200,0,111,0,168,0,61,0,89,0,231,0,165,0,161,0,145,0,99,0,248,0,195,0,71,0,141,0,224,0,105,0,208,0,44,0,192,0,25,0,137,0,34,0,90,0,51,0,17,0,3,0,140,0,13,0,0,0,0,0,48,0,142,0,230,0,157,0,0,0,0,0,15,0,144,0,60,0,16,0,84,0,207,0,193,0,0,0,87,0,153,0,5,0,0,0,0,0,31,0,224,0,177,0,144,0,255,0,138,0,95,0,10,0,0,0,76,0,77,0,201,0,62,0,167,0,76,0,249,0,0,0,138,0,193,0,0,0,146,0,143,0,107,0,25,0,166,0,25,0,169,0,240,0,148,0,0,0,0,0,0,0,226,0,141,0,0,0,103,0,186,0,0,0,120,0,0,0,105,0,0,0,0,0,49,0,62,0,0,0,72,0,0,0,0,0,234,0,0,0,191,0,0,0,218,0,135,0,249,0,80,0,74,0,0,0,138,0,0,0,21,0,0,0,0,0,97,0,0,0,98,0,56,0,105,0,0,0,161,0,131,0,58,0,121,0,7,0,96,0,28,0,97,0,0,0,36,0,26,0,163,0,157,0,29,0,211,0,233,0,165,0,150,0,0,0,5,0,162,0,0,0,19,0,18,0,40,0,174,0,0,0,217,0,239,0,52,0,0,0,92,0,29,0,160,0,1,0,132,0,234,0,60,0,184,0,182,0,106,0,224,0,201,0,84,0,73,0,169,0,180,0,209,0,179,0,207,0,138,0,228,0,192,0,247,0,94,0,180,0,14,0,0,0,115,0,104,0,193,0,176,0,0,0,218,0,115,0,25,0,0,0,227,0,0,0,226,0,0,0,41,0,0,0,231,0,101,0,150,0,0,0,74,0,8,0,0,0,20,0,0,0,155,0,156,0,248,0,53,0,80,0,24,0,172,0,61,0,0,0,204,0,198,0,49,0,0,0,0,0,101,0,16,0,57,0,104,0,0,0,0,0,61,0,59,0,45,0,115,0,0,0,143,0,119,0,227,0,153,0,160,0,172,0,28,0,176,0,211,0,210,0,71,0,31,0,10,0,0,0,98,0,110,0,142,0,233,0,204,0,0,0,0,0,191,0,108,0,223,0,148,0,203,0,95,0,0,0,0,0,100,0,222,0,0,0,0,0,64,0,81,0,127,0,237,0,152,0,193,0,0,0,10,0,87,0,75,0,0,0,0,0,6,0,0,0,160,0,128,0,112,0,88,0,0,0,96,0,50,0,126,0,0,0,0,0,105,0,28,0,244,0,50,0,176,0,220,0,65,0,215,0,126,0,0,0,143,0,0,0,61,0,0,0,0,0,0,0,162,0,152,0,197,0,0,0,75,0,0,0,181,0,61,0,211,0,29,0,19,0,96,0,0,0,78,0,0,0,112,0,176,0,233,0,39,0,47,0,2,0,198,0,178,0,38,0,36,0,0,0,168,0,2,0,205,0,177,0,145,0,175,0,0,0,231,0,173,0,0,0,0,0,86,0,0,0,207,0,235,0,31,0,227,0,159,0,94,0,0,0,0,0,103,0,0,0,238,0,132,0,0,0,0,0,204,0,16,0,228,0,202,0,143,0,150,0,244,0,0,0,122,0,193,0,200,0,41,0,31,0,0,0,216,0,127,0,127,0,0,0,0,0,228,0,0,0,0,0,121,0,58,0,127,0,39,0,176,0,97,0,0,0,68,0,231,0,84,0,116,0,22,0,84,0,17,0,53,0,126,0,145,0,38,0,0,0,0,0,0,0,101,0,128,0,150,0,83,0,0,0,0,0,39,0,175,0,0,0,0,0,211,0,145,0,160,0,0,0,179,0,0,0,118,0,161,0,0,0,226,0,193,0,56,0,233,0,255,0,0,0,245,0,160,0,108,0,179,0,165,0,90,0,130,0,35,0,56,0,110,0,150,0,0,0,247,0,28,0,127,0,189,0,43,0,210,0,31,0,0,0,0,0,139,0,235,0,0,0,210,0,33,0,0,0,174,0,0,0,248,0,23,0,0,0,30,0,101,0,253,0,60,0,206,0,11,0,5,0,0,0,0,0,0,0,148,0,213,0,23,0,243,0);
signal scenario_full  : scenario_type := (0,0,157,31,40,31,92,31,7,31,7,30,79,31,34,31,34,30,191,31,64,31,74,31,47,31,47,30,47,29,156,31,46,31,46,30,154,31,109,31,197,31,18,31,215,31,7,31,129,31,120,31,226,31,14,31,158,31,170,31,170,30,165,31,253,31,90,31,90,30,143,31,143,30,199,31,250,31,100,31,186,31,34,31,162,31,143,31,143,30,4,31,56,31,56,30,215,31,247,31,187,31,24,31,224,31,206,31,206,30,87,31,63,31,64,31,73,31,73,30,214,31,45,31,45,30,113,31,146,31,218,31,218,30,170,31,170,30,170,29,85,31,51,31,159,31,17,31,167,31,230,31,135,31,135,30,45,31,239,31,135,31,135,30,48,31,48,30,196,31,196,30,196,29,173,31,222,31,37,31,87,31,39,31,220,31,220,30,230,31,131,31,130,31,242,31,176,31,176,30,98,31,112,31,15,31,15,30,120,31,16,31,17,31,26,31,246,31,64,31,132,31,188,31,244,31,227,31,226,31,231,31,231,30,154,31,154,30,216,31,162,31,114,31,114,31,222,31,247,31,189,31,97,31,220,31,220,30,139,31,87,31,87,30,125,31,125,30,53,31,2,31,189,31,61,31,61,30,28,31,133,31,232,31,232,30,11,31,192,31,199,31,199,30,10,31,60,31,137,31,61,31,113,31,58,31,152,31,92,31,47,31,47,30,47,29,127,31,30,31,214,31,108,31,243,31,10,31,14,31,129,31,6,31,142,31,52,31,199,31,69,31,53,31,135,31,135,30,135,29,227,31,150,31,150,30,93,31,116,31,95,31,92,31,37,31,37,30,191,31,40,31,238,31,177,31,196,31,242,31,211,31,240,31,103,31,252,31,83,31,176,31,128,31,128,30,66,31,20,31,27,31,158,31,30,31,146,31,175,31,90,31,233,31,98,31,142,31,125,31,69,31,153,31,11,31,247,31,249,31,15,31,94,31,28,31,177,31,230,31,53,31,131,31,108,31,248,31,16,31,184,31,191,31,147,31,239,31,148,31,199,31,144,31,208,31,114,31,19,31,130,31,239,31,157,31,156,31,156,30,69,31,198,31,166,31,17,31,17,30,143,31,143,30,132,31,164,31,117,31,117,30,6,31,29,31,177,31,177,30,45,31,11,31,158,31,59,31,138,31,106,31,106,30,24,31,239,31,239,30,239,29,50,31,50,30,160,31,242,31,137,31,37,31,159,31,159,30,63,31,128,31,187,31,187,30,144,31,144,30,196,31,191,31,212,31,148,31,148,30,148,29,96,31,197,31,197,30,197,29,124,31,24,31,19,31,169,31,174,31,246,31,171,31,171,30,145,31,5,31,122,31,120,31,73,31,148,31,121,31,251,31,169,31,169,30,199,31,106,31,9,31,186,31,252,31,118,31,165,31,62,31,211,31,101,31,44,31,187,31,187,30,78,31,78,30,78,29,60,31,141,31,239,31,232,31,142,31,175,31,175,30,165,31,5,31,114,31,140,31,145,31,201,31,241,31,90,31,203,31,206,31,133,31,187,31,187,30,187,29,47,31,200,31,111,31,168,31,61,31,89,31,231,31,165,31,161,31,145,31,99,31,248,31,195,31,71,31,141,31,224,31,105,31,208,31,44,31,192,31,25,31,137,31,34,31,90,31,51,31,17,31,3,31,140,31,13,31,13,30,13,29,48,31,142,31,230,31,157,31,157,30,157,29,15,31,144,31,60,31,16,31,84,31,207,31,193,31,193,30,87,31,153,31,5,31,5,30,5,29,31,31,224,31,177,31,144,31,255,31,138,31,95,31,10,31,10,30,76,31,77,31,201,31,62,31,167,31,76,31,249,31,249,30,138,31,193,31,193,30,146,31,143,31,107,31,25,31,166,31,25,31,169,31,240,31,148,31,148,30,148,29,148,28,226,31,141,31,141,30,103,31,186,31,186,30,120,31,120,30,105,31,105,30,105,29,49,31,62,31,62,30,72,31,72,30,72,29,234,31,234,30,191,31,191,30,218,31,135,31,249,31,80,31,74,31,74,30,138,31,138,30,21,31,21,30,21,29,97,31,97,30,98,31,56,31,105,31,105,30,161,31,131,31,58,31,121,31,7,31,96,31,28,31,97,31,97,30,36,31,26,31,163,31,157,31,29,31,211,31,233,31,165,31,150,31,150,30,5,31,162,31,162,30,19,31,18,31,40,31,174,31,174,30,217,31,239,31,52,31,52,30,92,31,29,31,160,31,1,31,132,31,234,31,60,31,184,31,182,31,106,31,224,31,201,31,84,31,73,31,169,31,180,31,209,31,179,31,207,31,138,31,228,31,192,31,247,31,94,31,180,31,14,31,14,30,115,31,104,31,193,31,176,31,176,30,218,31,115,31,25,31,25,30,227,31,227,30,226,31,226,30,41,31,41,30,231,31,101,31,150,31,150,30,74,31,8,31,8,30,20,31,20,30,155,31,156,31,248,31,53,31,80,31,24,31,172,31,61,31,61,30,204,31,198,31,49,31,49,30,49,29,101,31,16,31,57,31,104,31,104,30,104,29,61,31,59,31,45,31,115,31,115,30,143,31,119,31,227,31,153,31,160,31,172,31,28,31,176,31,211,31,210,31,71,31,31,31,10,31,10,30,98,31,110,31,142,31,233,31,204,31,204,30,204,29,191,31,108,31,223,31,148,31,203,31,95,31,95,30,95,29,100,31,222,31,222,30,222,29,64,31,81,31,127,31,237,31,152,31,193,31,193,30,10,31,87,31,75,31,75,30,75,29,6,31,6,30,160,31,128,31,112,31,88,31,88,30,96,31,50,31,126,31,126,30,126,29,105,31,28,31,244,31,50,31,176,31,220,31,65,31,215,31,126,31,126,30,143,31,143,30,61,31,61,30,61,29,61,28,162,31,152,31,197,31,197,30,75,31,75,30,181,31,61,31,211,31,29,31,19,31,96,31,96,30,78,31,78,30,112,31,176,31,233,31,39,31,47,31,2,31,198,31,178,31,38,31,36,31,36,30,168,31,2,31,205,31,177,31,145,31,175,31,175,30,231,31,173,31,173,30,173,29,86,31,86,30,207,31,235,31,31,31,227,31,159,31,94,31,94,30,94,29,103,31,103,30,238,31,132,31,132,30,132,29,204,31,16,31,228,31,202,31,143,31,150,31,244,31,244,30,122,31,193,31,200,31,41,31,31,31,31,30,216,31,127,31,127,31,127,30,127,29,228,31,228,30,228,29,121,31,58,31,127,31,39,31,176,31,97,31,97,30,68,31,231,31,84,31,116,31,22,31,84,31,17,31,53,31,126,31,145,31,38,31,38,30,38,29,38,28,101,31,128,31,150,31,83,31,83,30,83,29,39,31,175,31,175,30,175,29,211,31,145,31,160,31,160,30,179,31,179,30,118,31,161,31,161,30,226,31,193,31,56,31,233,31,255,31,255,30,245,31,160,31,108,31,179,31,165,31,90,31,130,31,35,31,56,31,110,31,150,31,150,30,247,31,28,31,127,31,189,31,43,31,210,31,31,31,31,30,31,29,139,31,235,31,235,30,210,31,33,31,33,30,174,31,174,30,248,31,23,31,23,30,30,31,101,31,253,31,60,31,206,31,11,31,5,31,5,30,5,29,5,28,148,31,213,31,23,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
