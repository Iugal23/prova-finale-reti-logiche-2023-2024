-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1003;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,110,0,209,0,47,0,100,0,240,0,236,0,156,0,255,0,100,0,63,0,246,0,81,0,204,0,0,0,95,0,245,0,15,0,187,0,71,0,27,0,0,0,0,0,0,0,14,0,229,0,104,0,36,0,221,0,179,0,0,0,60,0,167,0,0,0,3,0,0,0,131,0,98,0,229,0,139,0,210,0,169,0,177,0,76,0,0,0,237,0,123,0,68,0,224,0,46,0,76,0,55,0,172,0,247,0,0,0,113,0,0,0,1,0,78,0,66,0,170,0,56,0,90,0,0,0,89,0,70,0,210,0,32,0,253,0,175,0,2,0,204,0,17,0,81,0,12,0,60,0,63,0,32,0,125,0,202,0,117,0,92,0,182,0,230,0,174,0,72,0,152,0,82,0,198,0,71,0,137,0,75,0,0,0,0,0,124,0,12,0,146,0,0,0,0,0,223,0,143,0,0,0,187,0,253,0,0,0,175,0,0,0,187,0,218,0,0,0,0,0,139,0,162,0,228,0,238,0,158,0,197,0,0,0,30,0,255,0,250,0,139,0,154,0,36,0,74,0,51,0,0,0,0,0,205,0,119,0,97,0,185,0,50,0,114,0,174,0,102,0,245,0,54,0,47,0,62,0,29,0,79,0,25,0,189,0,52,0,46,0,233,0,193,0,0,0,0,0,180,0,1,0,46,0,244,0,126,0,237,0,0,0,159,0,227,0,142,0,0,0,32,0,240,0,112,0,241,0,0,0,138,0,175,0,187,0,35,0,254,0,12,0,30,0,187,0,216,0,12,0,0,0,83,0,0,0,97,0,90,0,199,0,79,0,0,0,185,0,0,0,6,0,56,0,0,0,0,0,243,0,81,0,43,0,0,0,87,0,155,0,86,0,222,0,158,0,0,0,0,0,219,0,64,0,0,0,0,0,0,0,199,0,193,0,147,0,155,0,168,0,54,0,53,0,88,0,0,0,252,0,103,0,116,0,0,0,0,0,92,0,82,0,0,0,87,0,38,0,196,0,167,0,29,0,120,0,138,0,44,0,58,0,191,0,240,0,160,0,17,0,250,0,252,0,144,0,192,0,33,0,201,0,19,0,51,0,189,0,231,0,0,0,63,0,41,0,24,0,243,0,0,0,146,0,0,0,179,0,4,0,196,0,99,0,70,0,134,0,74,0,133,0,172,0,93,0,39,0,158,0,0,0,96,0,135,0,80,0,100,0,251,0,21,0,82,0,234,0,65,0,0,0,243,0,138,0,232,0,15,0,171,0,34,0,247,0,169,0,13,0,23,0,202,0,242,0,58,0,241,0,83,0,170,0,0,0,0,0,98,0,0,0,114,0,232,0,67,0,0,0,103,0,223,0,249,0,122,0,0,0,133,0,0,0,22,0,84,0,202,0,164,0,49,0,47,0,91,0,183,0,0,0,156,0,9,0,0,0,0,0,14,0,0,0,0,0,104,0,101,0,113,0,27,0,200,0,174,0,0,0,225,0,5,0,0,0,181,0,0,0,46,0,37,0,130,0,241,0,0,0,187,0,0,0,123,0,34,0,0,0,161,0,106,0,109,0,131,0,0,0,194,0,247,0,204,0,0,0,52,0,167,0,174,0,17,0,125,0,109,0,203,0,132,0,0,0,44,0,69,0,14,0,0,0,42,0,0,0,0,0,213,0,119,0,119,0,6,0,169,0,0,0,158,0,195,0,38,0,167,0,239,0,64,0,238,0,169,0,0,0,0,0,106,0,252,0,154,0,117,0,163,0,190,0,131,0,88,0,162,0,166,0,147,0,200,0,68,0,196,0,245,0,0,0,11,0,107,0,88,0,116,0,219,0,152,0,253,0,237,0,5,0,194,0,42,0,0,0,10,0,159,0,62,0,188,0,0,0,78,0,187,0,89,0,0,0,94,0,190,0,31,0,0,0,75,0,43,0,0,0,39,0,69,0,94,0,0,0,0,0,103,0,161,0,191,0,0,0,0,0,137,0,1,0,255,0,0,0,0,0,40,0,21,0,136,0,120,0,160,0,177,0,117,0,67,0,0,0,0,0,54,0,241,0,201,0,253,0,0,0,86,0,10,0,0,0,228,0,36,0,244,0,228,0,0,0,0,0,45,0,198,0,229,0,237,0,69,0,28,0,29,0,156,0,213,0,24,0,175,0,156,0,233,0,91,0,139,0,171,0,178,0,79,0,0,0,139,0,0,0,227,0,35,0,77,0,30,0,162,0,20,0,0,0,250,0,103,0,43,0,45,0,0,0,237,0,76,0,236,0,185,0,128,0,226,0,248,0,83,0,74,0,241,0,47,0,8,0,26,0,148,0,43,0,219,0,215,0,232,0,72,0,193,0,40,0,229,0,60,0,0,0,152,0,187,0,0,0,29,0,0,0,11,0,113,0,0,0,70,0,5,0,240,0,63,0,96,0,202,0,162,0,0,0,27,0,166,0,192,0,0,0,38,0,44,0,218,0,171,0,63,0,11,0,206,0,115,0,116,0,144,0,151,0,115,0,201,0,138,0,196,0,0,0,0,0,0,0,251,0,75,0,210,0,191,0,188,0,77,0,137,0,0,0,115,0,83,0,198,0,155,0,100,0,240,0,18,0,0,0,133,0,235,0,0,0,0,0,185,0,14,0,13,0,74,0,224,0,0,0,86,0,69,0,0,0,67,0,194,0,0,0,0,0,162,0,212,0,183,0,17,0,255,0,0,0,185,0,0,0,77,0,71,0,3,0,130,0,130,0,219,0,25,0,137,0,0,0,222,0,239,0,34,0,192,0,0,0,15,0,60,0,33,0,0,0,0,0,241,0,0,0,238,0,59,0,17,0,252,0,196,0,0,0,189,0,0,0,121,0,180,0,117,0,0,0,0,0,0,0,0,0,205,0,0,0,194,0,39,0,48,0,44,0,33,0,247,0,81,0,145,0,9,0,42,0,0,0,178,0,40,0,204,0,0,0,51,0,53,0,158,0,56,0,0,0,164,0,218,0,102,0,0,0,128,0,220,0,204,0,236,0,158,0,0,0,219,0,0,0,28,0,166,0,113,0,56,0,246,0,169,0,43,0,44,0,39,0,253,0,240,0,84,0,183,0,34,0,0,0,108,0,232,0,238,0,173,0,0,0,154,0,112,0,184,0,0,0,25,0,44,0,92,0,195,0,247,0,38,0,0,0,39,0,240,0,25,0,129,0,9,0,98,0,41,0,211,0,48,0,233,0,48,0,177,0,166,0,4,0,167,0,242,0,235,0,48,0,251,0,215,0,16,0,93,0,148,0,213,0,153,0,59,0,86,0,112,0,207,0,173,0,117,0,169,0,245,0,137,0,201,0,84,0,116,0,250,0,0,0,64,0,255,0,163,0,102,0,185,0,254,0,44,0,0,0,0,0,68,0,91,0,228,0,15,0,92,0,80,0,98,0,108,0,96,0,42,0,183,0,0,0,0,0,0,0,181,0,112,0,16,0,84,0,217,0,0,0,40,0,36,0,212,0,116,0,147,0,0,0,196,0,25,0,0,0,0,0,163,0,60,0,76,0,139,0,0,0,0,0,210,0,0,0,40,0,216,0,30,0,236,0,190,0,180,0,138,0,91,0,144,0,0,0,0,0,249,0,216,0,169,0,159,0,72,0,244,0,148,0,64,0,129,0,0,0,148,0,0,0,77,0,202,0,99,0,0,0,165,0,122,0,122,0,0,0,0,0,250,0,81,0,21,0,63,0,252,0,188,0,42,0,0,0,254,0,206,0,88,0,62,0,49,0,156,0,0,0,126,0,204,0,118,0,38,0,65,0,0,0,0,0,23,0,31,0,215,0,206,0,172,0,186,0,160,0,15,0,133,0,122,0,160,0,79,0,82,0,0,0,123,0,33,0,49,0,131,0,0,0,178,0,83,0,37,0,246,0,196,0,0,0,0,0,41,0,32,0,72,0,227,0,183,0,48,0,117,0,215,0,200,0,57,0,244,0,130,0,19,0,253,0,107,0,109,0,0,0,152,0,118,0,29,0,218,0,195,0,0,0,65,0,154,0,58,0,66,0,31,0,0,0,160,0,0,0,198,0,81,0,238,0,46,0,101,0,0,0,0,0,175,0,135,0,72,0,56,0,157,0,0,0,0,0,0,0,135,0,0,0,251,0,239,0,205,0,0,0,148,0,166,0,20,0,80,0,25,0,82,0,183,0,187,0,10,0,168,0,0,0,237,0,143,0,21,0,0,0,64,0,230,0,16,0,105,0,104,0,93,0,216,0,0,0,136,0,7,0,85,0,151,0,0,0,3,0,92,0,196,0,83,0,0,0,237,0,172,0,205,0,243,0,145,0,168,0,223,0,134,0,171,0,31,0,52,0,133,0,67,0,0,0,134,0,241,0,26,0,50,0,0,0,0,0,86,0,187,0,40,0,213,0,0,0,103,0,61,0,198,0,253,0,0,0,0,0,174,0,192,0,0,0,0,0,194,0,207,0,0,0,0,0,179,0,0,0,51,0,0,0,18,0,165,0);
signal scenario_full  : scenario_type := (0,0,110,31,209,31,47,31,100,31,240,31,236,31,156,31,255,31,100,31,63,31,246,31,81,31,204,31,204,30,95,31,245,31,15,31,187,31,71,31,27,31,27,30,27,29,27,28,14,31,229,31,104,31,36,31,221,31,179,31,179,30,60,31,167,31,167,30,3,31,3,30,131,31,98,31,229,31,139,31,210,31,169,31,177,31,76,31,76,30,237,31,123,31,68,31,224,31,46,31,76,31,55,31,172,31,247,31,247,30,113,31,113,30,1,31,78,31,66,31,170,31,56,31,90,31,90,30,89,31,70,31,210,31,32,31,253,31,175,31,2,31,204,31,17,31,81,31,12,31,60,31,63,31,32,31,125,31,202,31,117,31,92,31,182,31,230,31,174,31,72,31,152,31,82,31,198,31,71,31,137,31,75,31,75,30,75,29,124,31,12,31,146,31,146,30,146,29,223,31,143,31,143,30,187,31,253,31,253,30,175,31,175,30,187,31,218,31,218,30,218,29,139,31,162,31,228,31,238,31,158,31,197,31,197,30,30,31,255,31,250,31,139,31,154,31,36,31,74,31,51,31,51,30,51,29,205,31,119,31,97,31,185,31,50,31,114,31,174,31,102,31,245,31,54,31,47,31,62,31,29,31,79,31,25,31,189,31,52,31,46,31,233,31,193,31,193,30,193,29,180,31,1,31,46,31,244,31,126,31,237,31,237,30,159,31,227,31,142,31,142,30,32,31,240,31,112,31,241,31,241,30,138,31,175,31,187,31,35,31,254,31,12,31,30,31,187,31,216,31,12,31,12,30,83,31,83,30,97,31,90,31,199,31,79,31,79,30,185,31,185,30,6,31,56,31,56,30,56,29,243,31,81,31,43,31,43,30,87,31,155,31,86,31,222,31,158,31,158,30,158,29,219,31,64,31,64,30,64,29,64,28,199,31,193,31,147,31,155,31,168,31,54,31,53,31,88,31,88,30,252,31,103,31,116,31,116,30,116,29,92,31,82,31,82,30,87,31,38,31,196,31,167,31,29,31,120,31,138,31,44,31,58,31,191,31,240,31,160,31,17,31,250,31,252,31,144,31,192,31,33,31,201,31,19,31,51,31,189,31,231,31,231,30,63,31,41,31,24,31,243,31,243,30,146,31,146,30,179,31,4,31,196,31,99,31,70,31,134,31,74,31,133,31,172,31,93,31,39,31,158,31,158,30,96,31,135,31,80,31,100,31,251,31,21,31,82,31,234,31,65,31,65,30,243,31,138,31,232,31,15,31,171,31,34,31,247,31,169,31,13,31,23,31,202,31,242,31,58,31,241,31,83,31,170,31,170,30,170,29,98,31,98,30,114,31,232,31,67,31,67,30,103,31,223,31,249,31,122,31,122,30,133,31,133,30,22,31,84,31,202,31,164,31,49,31,47,31,91,31,183,31,183,30,156,31,9,31,9,30,9,29,14,31,14,30,14,29,104,31,101,31,113,31,27,31,200,31,174,31,174,30,225,31,5,31,5,30,181,31,181,30,46,31,37,31,130,31,241,31,241,30,187,31,187,30,123,31,34,31,34,30,161,31,106,31,109,31,131,31,131,30,194,31,247,31,204,31,204,30,52,31,167,31,174,31,17,31,125,31,109,31,203,31,132,31,132,30,44,31,69,31,14,31,14,30,42,31,42,30,42,29,213,31,119,31,119,31,6,31,169,31,169,30,158,31,195,31,38,31,167,31,239,31,64,31,238,31,169,31,169,30,169,29,106,31,252,31,154,31,117,31,163,31,190,31,131,31,88,31,162,31,166,31,147,31,200,31,68,31,196,31,245,31,245,30,11,31,107,31,88,31,116,31,219,31,152,31,253,31,237,31,5,31,194,31,42,31,42,30,10,31,159,31,62,31,188,31,188,30,78,31,187,31,89,31,89,30,94,31,190,31,31,31,31,30,75,31,43,31,43,30,39,31,69,31,94,31,94,30,94,29,103,31,161,31,191,31,191,30,191,29,137,31,1,31,255,31,255,30,255,29,40,31,21,31,136,31,120,31,160,31,177,31,117,31,67,31,67,30,67,29,54,31,241,31,201,31,253,31,253,30,86,31,10,31,10,30,228,31,36,31,244,31,228,31,228,30,228,29,45,31,198,31,229,31,237,31,69,31,28,31,29,31,156,31,213,31,24,31,175,31,156,31,233,31,91,31,139,31,171,31,178,31,79,31,79,30,139,31,139,30,227,31,35,31,77,31,30,31,162,31,20,31,20,30,250,31,103,31,43,31,45,31,45,30,237,31,76,31,236,31,185,31,128,31,226,31,248,31,83,31,74,31,241,31,47,31,8,31,26,31,148,31,43,31,219,31,215,31,232,31,72,31,193,31,40,31,229,31,60,31,60,30,152,31,187,31,187,30,29,31,29,30,11,31,113,31,113,30,70,31,5,31,240,31,63,31,96,31,202,31,162,31,162,30,27,31,166,31,192,31,192,30,38,31,44,31,218,31,171,31,63,31,11,31,206,31,115,31,116,31,144,31,151,31,115,31,201,31,138,31,196,31,196,30,196,29,196,28,251,31,75,31,210,31,191,31,188,31,77,31,137,31,137,30,115,31,83,31,198,31,155,31,100,31,240,31,18,31,18,30,133,31,235,31,235,30,235,29,185,31,14,31,13,31,74,31,224,31,224,30,86,31,69,31,69,30,67,31,194,31,194,30,194,29,162,31,212,31,183,31,17,31,255,31,255,30,185,31,185,30,77,31,71,31,3,31,130,31,130,31,219,31,25,31,137,31,137,30,222,31,239,31,34,31,192,31,192,30,15,31,60,31,33,31,33,30,33,29,241,31,241,30,238,31,59,31,17,31,252,31,196,31,196,30,189,31,189,30,121,31,180,31,117,31,117,30,117,29,117,28,117,27,205,31,205,30,194,31,39,31,48,31,44,31,33,31,247,31,81,31,145,31,9,31,42,31,42,30,178,31,40,31,204,31,204,30,51,31,53,31,158,31,56,31,56,30,164,31,218,31,102,31,102,30,128,31,220,31,204,31,236,31,158,31,158,30,219,31,219,30,28,31,166,31,113,31,56,31,246,31,169,31,43,31,44,31,39,31,253,31,240,31,84,31,183,31,34,31,34,30,108,31,232,31,238,31,173,31,173,30,154,31,112,31,184,31,184,30,25,31,44,31,92,31,195,31,247,31,38,31,38,30,39,31,240,31,25,31,129,31,9,31,98,31,41,31,211,31,48,31,233,31,48,31,177,31,166,31,4,31,167,31,242,31,235,31,48,31,251,31,215,31,16,31,93,31,148,31,213,31,153,31,59,31,86,31,112,31,207,31,173,31,117,31,169,31,245,31,137,31,201,31,84,31,116,31,250,31,250,30,64,31,255,31,163,31,102,31,185,31,254,31,44,31,44,30,44,29,68,31,91,31,228,31,15,31,92,31,80,31,98,31,108,31,96,31,42,31,183,31,183,30,183,29,183,28,181,31,112,31,16,31,84,31,217,31,217,30,40,31,36,31,212,31,116,31,147,31,147,30,196,31,25,31,25,30,25,29,163,31,60,31,76,31,139,31,139,30,139,29,210,31,210,30,40,31,216,31,30,31,236,31,190,31,180,31,138,31,91,31,144,31,144,30,144,29,249,31,216,31,169,31,159,31,72,31,244,31,148,31,64,31,129,31,129,30,148,31,148,30,77,31,202,31,99,31,99,30,165,31,122,31,122,31,122,30,122,29,250,31,81,31,21,31,63,31,252,31,188,31,42,31,42,30,254,31,206,31,88,31,62,31,49,31,156,31,156,30,126,31,204,31,118,31,38,31,65,31,65,30,65,29,23,31,31,31,215,31,206,31,172,31,186,31,160,31,15,31,133,31,122,31,160,31,79,31,82,31,82,30,123,31,33,31,49,31,131,31,131,30,178,31,83,31,37,31,246,31,196,31,196,30,196,29,41,31,32,31,72,31,227,31,183,31,48,31,117,31,215,31,200,31,57,31,244,31,130,31,19,31,253,31,107,31,109,31,109,30,152,31,118,31,29,31,218,31,195,31,195,30,65,31,154,31,58,31,66,31,31,31,31,30,160,31,160,30,198,31,81,31,238,31,46,31,101,31,101,30,101,29,175,31,135,31,72,31,56,31,157,31,157,30,157,29,157,28,135,31,135,30,251,31,239,31,205,31,205,30,148,31,166,31,20,31,80,31,25,31,82,31,183,31,187,31,10,31,168,31,168,30,237,31,143,31,21,31,21,30,64,31,230,31,16,31,105,31,104,31,93,31,216,31,216,30,136,31,7,31,85,31,151,31,151,30,3,31,92,31,196,31,83,31,83,30,237,31,172,31,205,31,243,31,145,31,168,31,223,31,134,31,171,31,31,31,52,31,133,31,67,31,67,30,134,31,241,31,26,31,50,31,50,30,50,29,86,31,187,31,40,31,213,31,213,30,103,31,61,31,198,31,253,31,253,30,253,29,174,31,192,31,192,30,192,29,194,31,207,31,207,30,207,29,179,31,179,30,51,31,51,30,18,31,165,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
