-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 368;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,169,0,81,0,55,0,191,0,32,0,136,0,58,0,228,0,146,0,109,0,14,0,95,0,213,0,192,0,42,0,0,0,146,0,145,0,123,0,61,0,50,0,43,0,90,0,0,0,4,0,124,0,182,0,0,0,122,0,176,0,0,0,62,0,69,0,248,0,187,0,25,0,225,0,0,0,83,0,105,0,71,0,80,0,144,0,160,0,0,0,241,0,53,0,158,0,13,0,247,0,176,0,65,0,243,0,198,0,221,0,245,0,234,0,152,0,155,0,190,0,94,0,230,0,19,0,140,0,1,0,81,0,166,0,0,0,78,0,0,0,0,0,248,0,189,0,73,0,206,0,73,0,0,0,0,0,22,0,82,0,49,0,64,0,235,0,0,0,93,0,0,0,2,0,121,0,46,0,174,0,0,0,0,0,0,0,124,0,99,0,246,0,64,0,127,0,206,0,198,0,126,0,49,0,211,0,197,0,90,0,80,0,197,0,94,0,145,0,29,0,242,0,137,0,157,0,174,0,123,0,219,0,200,0,238,0,35,0,120,0,179,0,0,0,27,0,36,0,68,0,95,0,80,0,130,0,189,0,55,0,8,0,0,0,181,0,0,0,243,0,81,0,0,0,168,0,11,0,175,0,176,0,144,0,131,0,95,0,193,0,244,0,114,0,52,0,60,0,0,0,157,0,169,0,70,0,0,0,159,0,73,0,77,0,0,0,146,0,143,0,170,0,27,0,130,0,48,0,72,0,0,0,0,0,210,0,37,0,85,0,0,0,143,0,235,0,196,0,173,0,163,0,0,0,197,0,191,0,170,0,169,0,105,0,132,0,66,0,106,0,92,0,250,0,187,0,38,0,254,0,247,0,130,0,1,0,0,0,107,0,159,0,24,0,157,0,236,0,218,0,224,0,242,0,167,0,109,0,254,0,0,0,18,0,13,0,0,0,211,0,46,0,0,0,20,0,145,0,0,0,190,0,67,0,121,0,0,0,68,0,0,0,35,0,113,0,153,0,0,0,198,0,65,0,64,0,0,0,180,0,228,0,126,0,0,0,89,0,0,0,54,0,9,0,40,0,180,0,81,0,43,0,121,0,0,0,142,0,0,0,64,0,0,0,0,0,187,0,0,0,12,0,174,0,0,0,0,0,161,0,210,0,91,0,164,0,248,0,40,0,47,0,1,0,0,0,251,0,244,0,102,0,130,0,0,0,67,0,0,0,207,0,235,0,33,0,0,0,0,0,228,0,194,0,184,0,225,0,97,0,134,0,126,0,194,0,61,0,204,0,58,0,29,0,20,0,129,0,173,0,24,0,151,0,226,0,184,0,34,0,128,0,232,0,0,0,106,0,30,0,12,0,131,0,101,0,104,0,33,0,235,0,158,0,0,0,174,0,174,0,175,0,0,0,13,0,0,0,205,0,3,0,231,0,139,0,249,0,0,0,24,0,137,0,43,0,231,0,241,0,233,0,20,0,243,0,137,0,44,0,0,0,0,0,121,0,0,0,252,0,101,0,52,0,165,0,129,0,252,0,95,0,75,0,0,0,0,0,30,0,247,0,233,0,0,0,202,0,29,0,250,0,205,0,12,0,0,0,72,0,195,0,0,0,147,0,152,0,245,0,110,0,61,0,169,0,33,0,81,0,0,0,174,0);
signal scenario_full  : scenario_type := (0,0,169,31,81,31,55,31,191,31,32,31,136,31,58,31,228,31,146,31,109,31,14,31,95,31,213,31,192,31,42,31,42,30,146,31,145,31,123,31,61,31,50,31,43,31,90,31,90,30,4,31,124,31,182,31,182,30,122,31,176,31,176,30,62,31,69,31,248,31,187,31,25,31,225,31,225,30,83,31,105,31,71,31,80,31,144,31,160,31,160,30,241,31,53,31,158,31,13,31,247,31,176,31,65,31,243,31,198,31,221,31,245,31,234,31,152,31,155,31,190,31,94,31,230,31,19,31,140,31,1,31,81,31,166,31,166,30,78,31,78,30,78,29,248,31,189,31,73,31,206,31,73,31,73,30,73,29,22,31,82,31,49,31,64,31,235,31,235,30,93,31,93,30,2,31,121,31,46,31,174,31,174,30,174,29,174,28,124,31,99,31,246,31,64,31,127,31,206,31,198,31,126,31,49,31,211,31,197,31,90,31,80,31,197,31,94,31,145,31,29,31,242,31,137,31,157,31,174,31,123,31,219,31,200,31,238,31,35,31,120,31,179,31,179,30,27,31,36,31,68,31,95,31,80,31,130,31,189,31,55,31,8,31,8,30,181,31,181,30,243,31,81,31,81,30,168,31,11,31,175,31,176,31,144,31,131,31,95,31,193,31,244,31,114,31,52,31,60,31,60,30,157,31,169,31,70,31,70,30,159,31,73,31,77,31,77,30,146,31,143,31,170,31,27,31,130,31,48,31,72,31,72,30,72,29,210,31,37,31,85,31,85,30,143,31,235,31,196,31,173,31,163,31,163,30,197,31,191,31,170,31,169,31,105,31,132,31,66,31,106,31,92,31,250,31,187,31,38,31,254,31,247,31,130,31,1,31,1,30,107,31,159,31,24,31,157,31,236,31,218,31,224,31,242,31,167,31,109,31,254,31,254,30,18,31,13,31,13,30,211,31,46,31,46,30,20,31,145,31,145,30,190,31,67,31,121,31,121,30,68,31,68,30,35,31,113,31,153,31,153,30,198,31,65,31,64,31,64,30,180,31,228,31,126,31,126,30,89,31,89,30,54,31,9,31,40,31,180,31,81,31,43,31,121,31,121,30,142,31,142,30,64,31,64,30,64,29,187,31,187,30,12,31,174,31,174,30,174,29,161,31,210,31,91,31,164,31,248,31,40,31,47,31,1,31,1,30,251,31,244,31,102,31,130,31,130,30,67,31,67,30,207,31,235,31,33,31,33,30,33,29,228,31,194,31,184,31,225,31,97,31,134,31,126,31,194,31,61,31,204,31,58,31,29,31,20,31,129,31,173,31,24,31,151,31,226,31,184,31,34,31,128,31,232,31,232,30,106,31,30,31,12,31,131,31,101,31,104,31,33,31,235,31,158,31,158,30,174,31,174,31,175,31,175,30,13,31,13,30,205,31,3,31,231,31,139,31,249,31,249,30,24,31,137,31,43,31,231,31,241,31,233,31,20,31,243,31,137,31,44,31,44,30,44,29,121,31,121,30,252,31,101,31,52,31,165,31,129,31,252,31,95,31,75,31,75,30,75,29,30,31,247,31,233,31,233,30,202,31,29,31,250,31,205,31,12,31,12,30,72,31,195,31,195,30,147,31,152,31,245,31,110,31,61,31,169,31,33,31,81,31,81,30,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
