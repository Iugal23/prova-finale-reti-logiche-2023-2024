-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 726;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (156,0,241,0,65,0,166,0,212,0,251,0,225,0,97,0,68,0,203,0,172,0,63,0,0,0,0,0,169,0,0,0,0,0,28,0,84,0,194,0,190,0,183,0,0,0,49,0,13,0,0,0,120,0,156,0,0,0,110,0,36,0,148,0,83,0,107,0,48,0,109,0,46,0,22,0,0,0,172,0,119,0,0,0,0,0,0,0,97,0,117,0,244,0,0,0,0,0,144,0,252,0,204,0,208,0,237,0,122,0,77,0,31,0,0,0,232,0,168,0,145,0,135,0,172,0,112,0,0,0,78,0,233,0,227,0,68,0,242,0,173,0,164,0,118,0,50,0,243,0,0,0,151,0,162,0,55,0,17,0,53,0,159,0,118,0,65,0,86,0,84,0,77,0,227,0,205,0,211,0,0,0,66,0,111,0,225,0,145,0,0,0,88,0,99,0,147,0,34,0,53,0,172,0,0,0,0,0,0,0,134,0,150,0,0,0,100,0,207,0,14,0,156,0,0,0,0,0,176,0,31,0,90,0,91,0,35,0,57,0,218,0,79,0,16,0,84,0,132,0,144,0,0,0,36,0,0,0,0,0,243,0,0,0,7,0,98,0,207,0,0,0,106,0,0,0,227,0,186,0,137,0,239,0,1,0,0,0,10,0,96,0,0,0,65,0,0,0,253,0,41,0,0,0,37,0,164,0,71,0,33,0,142,0,209,0,0,0,138,0,157,0,6,0,40,0,70,0,150,0,249,0,26,0,223,0,0,0,0,0,167,0,177,0,53,0,255,0,52,0,0,0,0,0,87,0,80,0,246,0,60,0,175,0,126,0,196,0,0,0,0,0,11,0,244,0,184,0,47,0,109,0,135,0,0,0,0,0,119,0,0,0,129,0,117,0,52,0,191,0,181,0,186,0,86,0,241,0,15,0,153,0,108,0,0,0,50,0,177,0,0,0,139,0,42,0,0,0,174,0,72,0,251,0,121,0,71,0,253,0,221,0,55,0,186,0,15,0,14,0,190,0,66,0,43,0,97,0,53,0,0,0,144,0,48,0,180,0,0,0,119,0,168,0,7,0,81,0,232,0,114,0,0,0,51,0,217,0,200,0,216,0,93,0,100,0,0,0,205,0,29,0,213,0,0,0,88,0,41,0,177,0,27,0,121,0,0,0,57,0,223,0,95,0,20,0,72,0,69,0,128,0,131,0,0,0,108,0,201,0,136,0,153,0,0,0,152,0,199,0,0,0,130,0,157,0,95,0,72,0,174,0,0,0,165,0,0,0,68,0,85,0,100,0,40,0,153,0,130,0,236,0,186,0,13,0,212,0,13,0,0,0,0,0,112,0,104,0,50,0,179,0,197,0,0,0,96,0,108,0,0,0,71,0,57,0,228,0,80,0,94,0,0,0,0,0,9,0,5,0,17,0,63,0,60,0,225,0,147,0,104,0,197,0,0,0,9,0,31,0,0,0,192,0,200,0,254,0,36,0,248,0,165,0,24,0,69,0,171,0,84,0,158,0,0,0,35,0,176,0,171,0,133,0,185,0,223,0,185,0,60,0,212,0,93,0,18,0,70,0,120,0,227,0,109,0,133,0,203,0,169,0,187,0,40,0,249,0,188,0,198,0,168,0,21,0,175,0,212,0,173,0,246,0,115,0,0,0,207,0,14,0,138,0,0,0,147,0,30,0,178,0,5,0,0,0,114,0,161,0,217,0,196,0,118,0,236,0,0,0,163,0,154,0,182,0,213,0,191,0,180,0,161,0,14,0,237,0,200,0,44,0,125,0,2,0,161,0,164,0,115,0,160,0,0,0,0,0,0,0,103,0,214,0,188,0,71,0,0,0,0,0,176,0,239,0,153,0,94,0,11,0,33,0,255,0,79,0,103,0,33,0,42,0,218,0,213,0,146,0,63,0,199,0,67,0,57,0,173,0,80,0,212,0,196,0,176,0,0,0,238,0,194,0,236,0,0,0,0,0,38,0,0,0,196,0,0,0,0,0,57,0,20,0,76,0,246,0,226,0,0,0,103,0,164,0,207,0,0,0,233,0,69,0,253,0,176,0,176,0,49,0,124,0,184,0,205,0,0,0,112,0,42,0,0,0,250,0,78,0,202,0,222,0,7,0,187,0,205,0,45,0,0,0,0,0,159,0,211,0,253,0,48,0,173,0,205,0,130,0,242,0,151,0,128,0,122,0,108,0,244,0,108,0,114,0,15,0,91,0,201,0,10,0,37,0,160,0,163,0,57,0,165,0,60,0,128,0,241,0,209,0,27,0,0,0,0,0,250,0,0,0,213,0,199,0,0,0,4,0,214,0,173,0,224,0,35,0,48,0,56,0,0,0,98,0,181,0,184,0,248,0,0,0,37,0,200,0,160,0,0,0,5,0,61,0,71,0,114,0,96,0,117,0,204,0,149,0,0,0,0,0,255,0,202,0,47,0,0,0,200,0,109,0,7,0,36,0,226,0,175,0,73,0,229,0,210,0,76,0,0,0,184,0,0,0,232,0,214,0,0,0,30,0,158,0,235,0,243,0,120,0,44,0,0,0,53,0,182,0,15,0,0,0,0,0,160,0,79,0,42,0,0,0,50,0,124,0,22,0,242,0,41,0,181,0,218,0,30,0,0,0,21,0,70,0,243,0,0,0,0,0,60,0,0,0,217,0,18,0,241,0,62,0,73,0,228,0,181,0,94,0,0,0,232,0,0,0,131,0,214,0,122,0,249,0,0,0,0,0,239,0,0,0,158,0,162,0,0,0,22,0,188,0,180,0,0,0,213,0,62,0,193,0,47,0,254,0,107,0,127,0,87,0,97,0,108,0,147,0,92,0,102,0,105,0,0,0,143,0,6,0,254,0,176,0,2,0,31,0,0,0,211,0,84,0,112,0,135,0,181,0,0,0,218,0,67,0,197,0,0,0,176,0,95,0,26,0,76,0,99,0,44,0,245,0,62,0,12,0,159,0,0,0,37,0,172,0,238,0,232,0,0,0,120,0,11,0,225,0,71,0,229,0,87,0,0,0,115,0,0,0,8,0,21,0,174,0,109,0,0,0,188,0,0,0,0,0,250,0,205,0,208,0,25,0,105,0,59,0,90,0,225,0,233,0,104,0,0,0,4,0,0,0,151,0,60,0,47,0,26,0,239,0,184,0,0,0,223,0,151,0,215,0,37,0,0,0,0,0,174,0,0,0,0,0,252,0,225,0,102,0,32,0,0,0,131,0,48,0,0,0,229,0,41,0,217,0,201,0,96,0);
signal scenario_full  : scenario_type := (156,31,241,31,65,31,166,31,212,31,251,31,225,31,97,31,68,31,203,31,172,31,63,31,63,30,63,29,169,31,169,30,169,29,28,31,84,31,194,31,190,31,183,31,183,30,49,31,13,31,13,30,120,31,156,31,156,30,110,31,36,31,148,31,83,31,107,31,48,31,109,31,46,31,22,31,22,30,172,31,119,31,119,30,119,29,119,28,97,31,117,31,244,31,244,30,244,29,144,31,252,31,204,31,208,31,237,31,122,31,77,31,31,31,31,30,232,31,168,31,145,31,135,31,172,31,112,31,112,30,78,31,233,31,227,31,68,31,242,31,173,31,164,31,118,31,50,31,243,31,243,30,151,31,162,31,55,31,17,31,53,31,159,31,118,31,65,31,86,31,84,31,77,31,227,31,205,31,211,31,211,30,66,31,111,31,225,31,145,31,145,30,88,31,99,31,147,31,34,31,53,31,172,31,172,30,172,29,172,28,134,31,150,31,150,30,100,31,207,31,14,31,156,31,156,30,156,29,176,31,31,31,90,31,91,31,35,31,57,31,218,31,79,31,16,31,84,31,132,31,144,31,144,30,36,31,36,30,36,29,243,31,243,30,7,31,98,31,207,31,207,30,106,31,106,30,227,31,186,31,137,31,239,31,1,31,1,30,10,31,96,31,96,30,65,31,65,30,253,31,41,31,41,30,37,31,164,31,71,31,33,31,142,31,209,31,209,30,138,31,157,31,6,31,40,31,70,31,150,31,249,31,26,31,223,31,223,30,223,29,167,31,177,31,53,31,255,31,52,31,52,30,52,29,87,31,80,31,246,31,60,31,175,31,126,31,196,31,196,30,196,29,11,31,244,31,184,31,47,31,109,31,135,31,135,30,135,29,119,31,119,30,129,31,117,31,52,31,191,31,181,31,186,31,86,31,241,31,15,31,153,31,108,31,108,30,50,31,177,31,177,30,139,31,42,31,42,30,174,31,72,31,251,31,121,31,71,31,253,31,221,31,55,31,186,31,15,31,14,31,190,31,66,31,43,31,97,31,53,31,53,30,144,31,48,31,180,31,180,30,119,31,168,31,7,31,81,31,232,31,114,31,114,30,51,31,217,31,200,31,216,31,93,31,100,31,100,30,205,31,29,31,213,31,213,30,88,31,41,31,177,31,27,31,121,31,121,30,57,31,223,31,95,31,20,31,72,31,69,31,128,31,131,31,131,30,108,31,201,31,136,31,153,31,153,30,152,31,199,31,199,30,130,31,157,31,95,31,72,31,174,31,174,30,165,31,165,30,68,31,85,31,100,31,40,31,153,31,130,31,236,31,186,31,13,31,212,31,13,31,13,30,13,29,112,31,104,31,50,31,179,31,197,31,197,30,96,31,108,31,108,30,71,31,57,31,228,31,80,31,94,31,94,30,94,29,9,31,5,31,17,31,63,31,60,31,225,31,147,31,104,31,197,31,197,30,9,31,31,31,31,30,192,31,200,31,254,31,36,31,248,31,165,31,24,31,69,31,171,31,84,31,158,31,158,30,35,31,176,31,171,31,133,31,185,31,223,31,185,31,60,31,212,31,93,31,18,31,70,31,120,31,227,31,109,31,133,31,203,31,169,31,187,31,40,31,249,31,188,31,198,31,168,31,21,31,175,31,212,31,173,31,246,31,115,31,115,30,207,31,14,31,138,31,138,30,147,31,30,31,178,31,5,31,5,30,114,31,161,31,217,31,196,31,118,31,236,31,236,30,163,31,154,31,182,31,213,31,191,31,180,31,161,31,14,31,237,31,200,31,44,31,125,31,2,31,161,31,164,31,115,31,160,31,160,30,160,29,160,28,103,31,214,31,188,31,71,31,71,30,71,29,176,31,239,31,153,31,94,31,11,31,33,31,255,31,79,31,103,31,33,31,42,31,218,31,213,31,146,31,63,31,199,31,67,31,57,31,173,31,80,31,212,31,196,31,176,31,176,30,238,31,194,31,236,31,236,30,236,29,38,31,38,30,196,31,196,30,196,29,57,31,20,31,76,31,246,31,226,31,226,30,103,31,164,31,207,31,207,30,233,31,69,31,253,31,176,31,176,31,49,31,124,31,184,31,205,31,205,30,112,31,42,31,42,30,250,31,78,31,202,31,222,31,7,31,187,31,205,31,45,31,45,30,45,29,159,31,211,31,253,31,48,31,173,31,205,31,130,31,242,31,151,31,128,31,122,31,108,31,244,31,108,31,114,31,15,31,91,31,201,31,10,31,37,31,160,31,163,31,57,31,165,31,60,31,128,31,241,31,209,31,27,31,27,30,27,29,250,31,250,30,213,31,199,31,199,30,4,31,214,31,173,31,224,31,35,31,48,31,56,31,56,30,98,31,181,31,184,31,248,31,248,30,37,31,200,31,160,31,160,30,5,31,61,31,71,31,114,31,96,31,117,31,204,31,149,31,149,30,149,29,255,31,202,31,47,31,47,30,200,31,109,31,7,31,36,31,226,31,175,31,73,31,229,31,210,31,76,31,76,30,184,31,184,30,232,31,214,31,214,30,30,31,158,31,235,31,243,31,120,31,44,31,44,30,53,31,182,31,15,31,15,30,15,29,160,31,79,31,42,31,42,30,50,31,124,31,22,31,242,31,41,31,181,31,218,31,30,31,30,30,21,31,70,31,243,31,243,30,243,29,60,31,60,30,217,31,18,31,241,31,62,31,73,31,228,31,181,31,94,31,94,30,232,31,232,30,131,31,214,31,122,31,249,31,249,30,249,29,239,31,239,30,158,31,162,31,162,30,22,31,188,31,180,31,180,30,213,31,62,31,193,31,47,31,254,31,107,31,127,31,87,31,97,31,108,31,147,31,92,31,102,31,105,31,105,30,143,31,6,31,254,31,176,31,2,31,31,31,31,30,211,31,84,31,112,31,135,31,181,31,181,30,218,31,67,31,197,31,197,30,176,31,95,31,26,31,76,31,99,31,44,31,245,31,62,31,12,31,159,31,159,30,37,31,172,31,238,31,232,31,232,30,120,31,11,31,225,31,71,31,229,31,87,31,87,30,115,31,115,30,8,31,21,31,174,31,109,31,109,30,188,31,188,30,188,29,250,31,205,31,208,31,25,31,105,31,59,31,90,31,225,31,233,31,104,31,104,30,4,31,4,30,151,31,60,31,47,31,26,31,239,31,184,31,184,30,223,31,151,31,215,31,37,31,37,30,37,29,174,31,174,30,174,29,252,31,225,31,102,31,32,31,32,30,131,31,48,31,48,30,229,31,41,31,217,31,201,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
