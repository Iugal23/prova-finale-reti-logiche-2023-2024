-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 797;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,249,0,88,0,137,0,130,0,103,0,30,0,125,0,167,0,117,0,223,0,116,0,37,0,209,0,0,0,64,0,229,0,0,0,0,0,206,0,148,0,27,0,240,0,76,0,0,0,0,0,20,0,83,0,84,0,131,0,194,0,211,0,0,0,222,0,187,0,171,0,253,0,161,0,0,0,202,0,172,0,0,0,0,0,241,0,149,0,174,0,0,0,93,0,81,0,197,0,23,0,0,0,48,0,191,0,48,0,34,0,0,0,24,0,0,0,0,0,210,0,0,0,181,0,0,0,245,0,80,0,165,0,158,0,233,0,159,0,209,0,151,0,158,0,238,0,214,0,189,0,132,0,61,0,18,0,158,0,0,0,0,0,203,0,0,0,0,0,169,0,143,0,90,0,178,0,26,0,212,0,240,0,235,0,66,0,132,0,36,0,71,0,191,0,193,0,178,0,218,0,218,0,63,0,143,0,0,0,0,0,145,0,47,0,55,0,234,0,116,0,0,0,41,0,190,0,0,0,238,0,0,0,0,0,134,0,0,0,91,0,174,0,220,0,152,0,154,0,0,0,109,0,0,0,88,0,171,0,143,0,25,0,156,0,42,0,50,0,204,0,0,0,98,0,71,0,212,0,94,0,156,0,79,0,0,0,9,0,175,0,110,0,0,0,53,0,149,0,0,0,24,0,44,0,137,0,179,0,49,0,43,0,55,0,171,0,50,0,0,0,207,0,0,0,0,0,115,0,0,0,205,0,34,0,24,0,173,0,0,0,93,0,209,0,182,0,250,0,117,0,24,0,0,0,213,0,20,0,148,0,133,0,243,0,178,0,241,0,27,0,0,0,104,0,56,0,74,0,189,0,51,0,150,0,45,0,63,0,247,0,0,0,27,0,57,0,85,0,0,0,222,0,148,0,233,0,211,0,185,0,62,0,67,0,253,0,141,0,106,0,0,0,211,0,13,0,213,0,247,0,78,0,0,0,155,0,82,0,182,0,129,0,31,0,84,0,143,0,248,0,122,0,108,0,91,0,127,0,250,0,145,0,186,0,196,0,0,0,143,0,0,0,0,0,181,0,26,0,0,0,88,0,254,0,25,0,0,0,129,0,229,0,204,0,0,0,87,0,147,0,65,0,101,0,254,0,19,0,77,0,241,0,0,0,215,0,63,0,64,0,120,0,209,0,151,0,202,0,146,0,72,0,114,0,0,0,0,0,203,0,224,0,22,0,176,0,173,0,0,0,185,0,0,0,0,0,61,0,88,0,150,0,21,0,188,0,241,0,0,0,5,0,77,0,126,0,137,0,60,0,64,0,74,0,231,0,35,0,202,0,0,0,96,0,27,0,253,0,194,0,183,0,145,0,178,0,222,0,0,0,155,0,167,0,22,0,116,0,148,0,159,0,174,0,216,0,115,0,105,0,107,0,26,0,149,0,252,0,69,0,54,0,198,0,0,0,84,0,254,0,201,0,124,0,253,0,241,0,27,0,0,0,209,0,213,0,174,0,7,0,247,0,129,0,246,0,104,0,182,0,87,0,98,0,139,0,224,0,97,0,251,0,224,0,81,0,110,0,129,0,75,0,145,0,203,0,0,0,94,0,32,0,211,0,124,0,61,0,203,0,70,0,241,0,13,0,50,0,56,0,90,0,0,0,175,0,44,0,214,0,144,0,119,0,220,0,18,0,155,0,63,0,119,0,148,0,0,0,0,0,158,0,0,0,108,0,121,0,0,0,87,0,171,0,144,0,12,0,186,0,3,0,39,0,241,0,112,0,0,0,104,0,0,0,135,0,161,0,148,0,216,0,152,0,67,0,16,0,55,0,243,0,0,0,44,0,194,0,0,0,68,0,128,0,104,0,0,0,18,0,69,0,72,0,91,0,168,0,130,0,154,0,132,0,0,0,92,0,224,0,128,0,41,0,0,0,0,0,12,0,0,0,25,0,0,0,192,0,103,0,10,0,173,0,0,0,0,0,109,0,23,0,154,0,89,0,74,0,161,0,92,0,61,0,211,0,58,0,199,0,230,0,99,0,0,0,138,0,194,0,0,0,130,0,55,0,58,0,137,0,103,0,128,0,201,0,17,0,0,0,234,0,179,0,85,0,0,0,11,0,95,0,19,0,213,0,195,0,127,0,0,0,0,0,37,0,135,0,207,0,228,0,231,0,65,0,92,0,228,0,0,0,204,0,164,0,132,0,65,0,0,0,61,0,160,0,0,0,175,0,0,0,0,0,138,0,191,0,138,0,150,0,82,0,214,0,179,0,20,0,127,0,123,0,195,0,166,0,0,0,250,0,69,0,205,0,229,0,31,0,50,0,255,0,213,0,0,0,230,0,7,0,0,0,150,0,193,0,184,0,0,0,206,0,183,0,218,0,26,0,160,0,235,0,161,0,0,0,105,0,0,0,0,0,202,0,24,0,215,0,202,0,201,0,201,0,34,0,0,0,43,0,89,0,136,0,209,0,28,0,41,0,215,0,26,0,161,0,26,0,244,0,118,0,0,0,31,0,157,0,37,0,176,0,51,0,0,0,133,0,231,0,219,0,100,0,86,0,212,0,49,0,0,0,234,0,150,0,100,0,148,0,138,0,248,0,102,0,110,0,134,0,73,0,170,0,106,0,241,0,150,0,178,0,193,0,19,0,63,0,49,0,247,0,0,0,27,0,131,0,158,0,148,0,50,0,247,0,0,0,23,0,207,0,68,0,102,0,191,0,185,0,70,0,34,0,103,0,196,0,59,0,0,0,107,0,210,0,88,0,132,0,19,0,22,0,14,0,238,0,197,0,113,0,176,0,105,0,152,0,0,0,83,0,72,0,175,0,87,0,96,0,12,0,173,0,103,0,0,0,91,0,0,0,0,0,106,0,7,0,129,0,22,0,209,0,152,0,0,0,124,0,33,0,0,0,93,0,107,0,221,0,102,0,36,0,129,0,229,0,250,0,70,0,89,0,172,0,22,0,0,0,138,0,207,0,81,0,160,0,243,0,29,0,45,0,153,0,3,0,0,0,249,0,0,0,60,0,0,0,102,0,49,0,239,0,40,0,231,0,0,0,0,0,214,0,149,0,213,0,99,0,0,0,180,0,67,0,0,0,230,0,0,0,0,0,0,0,118,0,26,0,147,0,231,0,0,0,237,0,108,0,224,0,244,0,2,0,0,0,121,0,87,0,0,0,116,0,0,0,28,0,65,0,134,0,208,0,182,0,221,0,68,0,8,0,230,0,32,0,164,0,63,0,29,0,88,0,84,0,60,0,39,0,0,0,109,0,0,0,92,0,132,0,239,0,0,0,22,0,31,0,1,0,131,0,81,0,108,0,0,0,0,0,2,0,129,0,189,0,89,0,95,0,0,0,41,0,0,0,255,0,11,0,0,0,241,0,95,0,5,0,239,0,0,0,247,0,0,0,38,0,223,0,78,0,218,0,117,0,41,0,0,0,50,0,179,0,123,0,78,0,0,0,43,0,165,0,193,0,0,0,139,0,53,0,156,0,164,0,199,0,53,0,0,0,32,0,167,0,236,0,42,0,0,0,123,0,206,0,193,0,58,0,60,0,0,0,1,0,96,0);
signal scenario_full  : scenario_type := (16,31,249,31,88,31,137,31,130,31,103,31,30,31,125,31,167,31,117,31,223,31,116,31,37,31,209,31,209,30,64,31,229,31,229,30,229,29,206,31,148,31,27,31,240,31,76,31,76,30,76,29,20,31,83,31,84,31,131,31,194,31,211,31,211,30,222,31,187,31,171,31,253,31,161,31,161,30,202,31,172,31,172,30,172,29,241,31,149,31,174,31,174,30,93,31,81,31,197,31,23,31,23,30,48,31,191,31,48,31,34,31,34,30,24,31,24,30,24,29,210,31,210,30,181,31,181,30,245,31,80,31,165,31,158,31,233,31,159,31,209,31,151,31,158,31,238,31,214,31,189,31,132,31,61,31,18,31,158,31,158,30,158,29,203,31,203,30,203,29,169,31,143,31,90,31,178,31,26,31,212,31,240,31,235,31,66,31,132,31,36,31,71,31,191,31,193,31,178,31,218,31,218,31,63,31,143,31,143,30,143,29,145,31,47,31,55,31,234,31,116,31,116,30,41,31,190,31,190,30,238,31,238,30,238,29,134,31,134,30,91,31,174,31,220,31,152,31,154,31,154,30,109,31,109,30,88,31,171,31,143,31,25,31,156,31,42,31,50,31,204,31,204,30,98,31,71,31,212,31,94,31,156,31,79,31,79,30,9,31,175,31,110,31,110,30,53,31,149,31,149,30,24,31,44,31,137,31,179,31,49,31,43,31,55,31,171,31,50,31,50,30,207,31,207,30,207,29,115,31,115,30,205,31,34,31,24,31,173,31,173,30,93,31,209,31,182,31,250,31,117,31,24,31,24,30,213,31,20,31,148,31,133,31,243,31,178,31,241,31,27,31,27,30,104,31,56,31,74,31,189,31,51,31,150,31,45,31,63,31,247,31,247,30,27,31,57,31,85,31,85,30,222,31,148,31,233,31,211,31,185,31,62,31,67,31,253,31,141,31,106,31,106,30,211,31,13,31,213,31,247,31,78,31,78,30,155,31,82,31,182,31,129,31,31,31,84,31,143,31,248,31,122,31,108,31,91,31,127,31,250,31,145,31,186,31,196,31,196,30,143,31,143,30,143,29,181,31,26,31,26,30,88,31,254,31,25,31,25,30,129,31,229,31,204,31,204,30,87,31,147,31,65,31,101,31,254,31,19,31,77,31,241,31,241,30,215,31,63,31,64,31,120,31,209,31,151,31,202,31,146,31,72,31,114,31,114,30,114,29,203,31,224,31,22,31,176,31,173,31,173,30,185,31,185,30,185,29,61,31,88,31,150,31,21,31,188,31,241,31,241,30,5,31,77,31,126,31,137,31,60,31,64,31,74,31,231,31,35,31,202,31,202,30,96,31,27,31,253,31,194,31,183,31,145,31,178,31,222,31,222,30,155,31,167,31,22,31,116,31,148,31,159,31,174,31,216,31,115,31,105,31,107,31,26,31,149,31,252,31,69,31,54,31,198,31,198,30,84,31,254,31,201,31,124,31,253,31,241,31,27,31,27,30,209,31,213,31,174,31,7,31,247,31,129,31,246,31,104,31,182,31,87,31,98,31,139,31,224,31,97,31,251,31,224,31,81,31,110,31,129,31,75,31,145,31,203,31,203,30,94,31,32,31,211,31,124,31,61,31,203,31,70,31,241,31,13,31,50,31,56,31,90,31,90,30,175,31,44,31,214,31,144,31,119,31,220,31,18,31,155,31,63,31,119,31,148,31,148,30,148,29,158,31,158,30,108,31,121,31,121,30,87,31,171,31,144,31,12,31,186,31,3,31,39,31,241,31,112,31,112,30,104,31,104,30,135,31,161,31,148,31,216,31,152,31,67,31,16,31,55,31,243,31,243,30,44,31,194,31,194,30,68,31,128,31,104,31,104,30,18,31,69,31,72,31,91,31,168,31,130,31,154,31,132,31,132,30,92,31,224,31,128,31,41,31,41,30,41,29,12,31,12,30,25,31,25,30,192,31,103,31,10,31,173,31,173,30,173,29,109,31,23,31,154,31,89,31,74,31,161,31,92,31,61,31,211,31,58,31,199,31,230,31,99,31,99,30,138,31,194,31,194,30,130,31,55,31,58,31,137,31,103,31,128,31,201,31,17,31,17,30,234,31,179,31,85,31,85,30,11,31,95,31,19,31,213,31,195,31,127,31,127,30,127,29,37,31,135,31,207,31,228,31,231,31,65,31,92,31,228,31,228,30,204,31,164,31,132,31,65,31,65,30,61,31,160,31,160,30,175,31,175,30,175,29,138,31,191,31,138,31,150,31,82,31,214,31,179,31,20,31,127,31,123,31,195,31,166,31,166,30,250,31,69,31,205,31,229,31,31,31,50,31,255,31,213,31,213,30,230,31,7,31,7,30,150,31,193,31,184,31,184,30,206,31,183,31,218,31,26,31,160,31,235,31,161,31,161,30,105,31,105,30,105,29,202,31,24,31,215,31,202,31,201,31,201,31,34,31,34,30,43,31,89,31,136,31,209,31,28,31,41,31,215,31,26,31,161,31,26,31,244,31,118,31,118,30,31,31,157,31,37,31,176,31,51,31,51,30,133,31,231,31,219,31,100,31,86,31,212,31,49,31,49,30,234,31,150,31,100,31,148,31,138,31,248,31,102,31,110,31,134,31,73,31,170,31,106,31,241,31,150,31,178,31,193,31,19,31,63,31,49,31,247,31,247,30,27,31,131,31,158,31,148,31,50,31,247,31,247,30,23,31,207,31,68,31,102,31,191,31,185,31,70,31,34,31,103,31,196,31,59,31,59,30,107,31,210,31,88,31,132,31,19,31,22,31,14,31,238,31,197,31,113,31,176,31,105,31,152,31,152,30,83,31,72,31,175,31,87,31,96,31,12,31,173,31,103,31,103,30,91,31,91,30,91,29,106,31,7,31,129,31,22,31,209,31,152,31,152,30,124,31,33,31,33,30,93,31,107,31,221,31,102,31,36,31,129,31,229,31,250,31,70,31,89,31,172,31,22,31,22,30,138,31,207,31,81,31,160,31,243,31,29,31,45,31,153,31,3,31,3,30,249,31,249,30,60,31,60,30,102,31,49,31,239,31,40,31,231,31,231,30,231,29,214,31,149,31,213,31,99,31,99,30,180,31,67,31,67,30,230,31,230,30,230,29,230,28,118,31,26,31,147,31,231,31,231,30,237,31,108,31,224,31,244,31,2,31,2,30,121,31,87,31,87,30,116,31,116,30,28,31,65,31,134,31,208,31,182,31,221,31,68,31,8,31,230,31,32,31,164,31,63,31,29,31,88,31,84,31,60,31,39,31,39,30,109,31,109,30,92,31,132,31,239,31,239,30,22,31,31,31,1,31,131,31,81,31,108,31,108,30,108,29,2,31,129,31,189,31,89,31,95,31,95,30,41,31,41,30,255,31,11,31,11,30,241,31,95,31,5,31,239,31,239,30,247,31,247,30,38,31,223,31,78,31,218,31,117,31,41,31,41,30,50,31,179,31,123,31,78,31,78,30,43,31,165,31,193,31,193,30,139,31,53,31,156,31,164,31,199,31,53,31,53,30,32,31,167,31,236,31,42,31,42,30,123,31,206,31,193,31,58,31,60,31,60,30,1,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
