-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_471 is
end project_tb_471;

architecture project_tb_arch_471 of project_tb_471 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 453;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,0,0,0,0,222,0,96,0,227,0,58,0,85,0,0,0,0,0,250,0,63,0,133,0,255,0,0,0,58,0,172,0,0,0,4,0,163,0,229,0,146,0,204,0,145,0,201,0,53,0,19,0,232,0,0,0,208,0,44,0,117,0,72,0,167,0,167,0,248,0,203,0,63,0,0,0,247,0,68,0,115,0,199,0,0,0,46,0,27,0,240,0,96,0,0,0,191,0,85,0,225,0,16,0,163,0,5,0,70,0,50,0,0,0,0,0,61,0,29,0,47,0,37,0,34,0,159,0,162,0,136,0,46,0,3,0,1,0,135,0,245,0,204,0,175,0,207,0,142,0,99,0,151,0,213,0,28,0,157,0,229,0,211,0,0,0,0,0,229,0,230,0,44,0,234,0,88,0,0,0,172,0,0,0,3,0,0,0,132,0,51,0,0,0,146,0,45,0,18,0,227,0,97,0,132,0,87,0,0,0,22,0,190,0,110,0,0,0,0,0,242,0,107,0,167,0,239,0,136,0,51,0,218,0,218,0,229,0,140,0,195,0,207,0,0,0,240,0,160,0,147,0,146,0,21,0,237,0,214,0,0,0,64,0,223,0,144,0,0,0,0,0,140,0,244,0,43,0,4,0,196,0,34,0,0,0,80,0,12,0,93,0,216,0,115,0,245,0,15,0,31,0,55,0,44,0,0,0,6,0,0,0,39,0,247,0,0,0,98,0,212,0,237,0,109,0,0,0,112,0,0,0,112,0,218,0,59,0,0,0,203,0,48,0,0,0,102,0,146,0,161,0,176,0,117,0,89,0,93,0,102,0,111,0,1,0,219,0,162,0,127,0,227,0,169,0,176,0,108,0,131,0,27,0,164,0,202,0,47,0,0,0,143,0,108,0,195,0,60,0,0,0,9,0,0,0,63,0,11,0,0,0,113,0,114,0,187,0,61,0,181,0,159,0,50,0,0,0,0,0,34,0,16,0,0,0,178,0,104,0,36,0,156,0,0,0,172,0,0,0,3,0,53,0,228,0,176,0,0,0,47,0,59,0,142,0,114,0,51,0,0,0,31,0,154,0,234,0,117,0,0,0,101,0,211,0,123,0,166,0,142,0,75,0,0,0,68,0,140,0,36,0,169,0,31,0,0,0,110,0,251,0,80,0,35,0,0,0,82,0,137,0,0,0,211,0,52,0,35,0,0,0,152,0,97,0,59,0,0,0,179,0,0,0,127,0,224,0,219,0,203,0,193,0,152,0,0,0,10,0,237,0,54,0,255,0,72,0,216,0,0,0,28,0,104,0,60,0,102,0,2,0,215,0,69,0,36,0,33,0,0,0,206,0,11,0,0,0,220,0,0,0,57,0,0,0,0,0,52,0,198,0,128,0,162,0,0,0,4,0,211,0,251,0,197,0,174,0,57,0,0,0,208,0,34,0,164,0,61,0,107,0,239,0,0,0,240,0,185,0,251,0,177,0,213,0,75,0,248,0,96,0,0,0,101,0,130,0,79,0,0,0,0,0,78,0,88,0,127,0,132,0,59,0,93,0,82,0,135,0,34,0,163,0,21,0,233,0,45,0,232,0,0,0,229,0,6,0,0,0,0,0,192,0,0,0,140,0,103,0,136,0,176,0,169,0,246,0,0,0,15,0,1,0,0,0,25,0,248,0,33,0,93,0,0,0,0,0,170,0,0,0,26,0,249,0,88,0,208,0,129,0,154,0,34,0,253,0,90,0,107,0,53,0,0,0,184,0,195,0,67,0,54,0,229,0,54,0,84,0,0,0,63,0,253,0,218,0,171,0,163,0,128,0,0,0,76,0,157,0,217,0,252,0,25,0,94,0,0,0,243,0,123,0,252,0,98,0,155,0,185,0,100,0,239,0,109,0,167,0,184,0,0,0,229,0,229,0,0,0,143,0,9,0,26,0,0,0,69,0,35,0,36,0,201,0,7,0,218,0,89,0,203,0,29,0,179,0,20,0,118,0,110,0,11,0,143,0,14,0,25,0,240,0,198,0,0,0,64,0,128,0,104,0);
signal scenario_full  : scenario_type := (245,31,245,30,245,29,222,31,96,31,227,31,58,31,85,31,85,30,85,29,250,31,63,31,133,31,255,31,255,30,58,31,172,31,172,30,4,31,163,31,229,31,146,31,204,31,145,31,201,31,53,31,19,31,232,31,232,30,208,31,44,31,117,31,72,31,167,31,167,31,248,31,203,31,63,31,63,30,247,31,68,31,115,31,199,31,199,30,46,31,27,31,240,31,96,31,96,30,191,31,85,31,225,31,16,31,163,31,5,31,70,31,50,31,50,30,50,29,61,31,29,31,47,31,37,31,34,31,159,31,162,31,136,31,46,31,3,31,1,31,135,31,245,31,204,31,175,31,207,31,142,31,99,31,151,31,213,31,28,31,157,31,229,31,211,31,211,30,211,29,229,31,230,31,44,31,234,31,88,31,88,30,172,31,172,30,3,31,3,30,132,31,51,31,51,30,146,31,45,31,18,31,227,31,97,31,132,31,87,31,87,30,22,31,190,31,110,31,110,30,110,29,242,31,107,31,167,31,239,31,136,31,51,31,218,31,218,31,229,31,140,31,195,31,207,31,207,30,240,31,160,31,147,31,146,31,21,31,237,31,214,31,214,30,64,31,223,31,144,31,144,30,144,29,140,31,244,31,43,31,4,31,196,31,34,31,34,30,80,31,12,31,93,31,216,31,115,31,245,31,15,31,31,31,55,31,44,31,44,30,6,31,6,30,39,31,247,31,247,30,98,31,212,31,237,31,109,31,109,30,112,31,112,30,112,31,218,31,59,31,59,30,203,31,48,31,48,30,102,31,146,31,161,31,176,31,117,31,89,31,93,31,102,31,111,31,1,31,219,31,162,31,127,31,227,31,169,31,176,31,108,31,131,31,27,31,164,31,202,31,47,31,47,30,143,31,108,31,195,31,60,31,60,30,9,31,9,30,63,31,11,31,11,30,113,31,114,31,187,31,61,31,181,31,159,31,50,31,50,30,50,29,34,31,16,31,16,30,178,31,104,31,36,31,156,31,156,30,172,31,172,30,3,31,53,31,228,31,176,31,176,30,47,31,59,31,142,31,114,31,51,31,51,30,31,31,154,31,234,31,117,31,117,30,101,31,211,31,123,31,166,31,142,31,75,31,75,30,68,31,140,31,36,31,169,31,31,31,31,30,110,31,251,31,80,31,35,31,35,30,82,31,137,31,137,30,211,31,52,31,35,31,35,30,152,31,97,31,59,31,59,30,179,31,179,30,127,31,224,31,219,31,203,31,193,31,152,31,152,30,10,31,237,31,54,31,255,31,72,31,216,31,216,30,28,31,104,31,60,31,102,31,2,31,215,31,69,31,36,31,33,31,33,30,206,31,11,31,11,30,220,31,220,30,57,31,57,30,57,29,52,31,198,31,128,31,162,31,162,30,4,31,211,31,251,31,197,31,174,31,57,31,57,30,208,31,34,31,164,31,61,31,107,31,239,31,239,30,240,31,185,31,251,31,177,31,213,31,75,31,248,31,96,31,96,30,101,31,130,31,79,31,79,30,79,29,78,31,88,31,127,31,132,31,59,31,93,31,82,31,135,31,34,31,163,31,21,31,233,31,45,31,232,31,232,30,229,31,6,31,6,30,6,29,192,31,192,30,140,31,103,31,136,31,176,31,169,31,246,31,246,30,15,31,1,31,1,30,25,31,248,31,33,31,93,31,93,30,93,29,170,31,170,30,26,31,249,31,88,31,208,31,129,31,154,31,34,31,253,31,90,31,107,31,53,31,53,30,184,31,195,31,67,31,54,31,229,31,54,31,84,31,84,30,63,31,253,31,218,31,171,31,163,31,128,31,128,30,76,31,157,31,217,31,252,31,25,31,94,31,94,30,243,31,123,31,252,31,98,31,155,31,185,31,100,31,239,31,109,31,167,31,184,31,184,30,229,31,229,31,229,30,143,31,9,31,26,31,26,30,69,31,35,31,36,31,201,31,7,31,218,31,89,31,203,31,29,31,179,31,20,31,118,31,110,31,11,31,143,31,14,31,25,31,240,31,198,31,198,30,64,31,128,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
