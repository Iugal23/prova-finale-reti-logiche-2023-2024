-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_783 is
end project_tb_783;

architecture project_tb_arch_783 of project_tb_783 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,0,0,152,0,144,0,75,0,181,0,110,0,239,0,61,0,115,0,0,0,39,0,68,0,161,0,217,0,226,0,146,0,0,0,235,0,116,0,238,0,80,0,37,0,0,0,0,0,21,0,171,0,1,0,18,0,237,0,200,0,249,0,0,0,61,0,149,0,242,0,0,0,0,0,233,0,0,0,207,0,106,0,31,0,217,0,151,0,99,0,129,0,183,0,56,0,229,0,188,0,129,0,99,0,108,0,65,0,78,0,101,0,190,0,6,0,102,0,6,0,19,0,122,0,14,0,0,0,220,0,80,0,168,0,146,0,0,0,52,0,0,0,0,0,0,0,222,0,188,0,0,0,112,0,74,0,115,0,0,0,187,0,51,0,96,0,46,0,10,0,68,0,99,0,155,0,239,0,147,0,222,0,33,0,2,0,0,0,128,0,140,0,240,0,37,0,153,0,0,0,152,0,0,0,234,0,214,0,181,0,89,0,0,0,32,0,161,0,5,0,0,0,0,0,131,0,16,0,74,0,236,0,0,0,64,0,153,0,76,0,89,0,23,0,0,0,8,0,174,0,102,0,0,0,169,0,64,0,0,0,31,0,249,0,0,0,239,0,220,0,0,0,84,0,232,0,116,0,253,0,96,0,19,0,167,0,66,0,15,0,0,0,17,0,76,0,14,0,0,0,47,0,241,0,183,0,128,0,5,0,57,0,20,0,49,0,0,0,218,0,48,0,24,0,94,0,176,0,174,0,51,0,199,0,14,0,138,0,0,0,0,0,247,0,95,0,241,0,177,0,188,0,217,0,25,0,243,0,126,0,196,0,51,0,236,0,106,0,107,0,0,0,140,0,167,0,0,0,0,0,249,0,162,0,123,0,0,0,66,0,0,0,226,0,27,0,84,0,210,0,134,0,165,0,57,0,207,0,57,0,0,0,75,0,52,0,245,0,179,0,168,0,0,0,235,0,87,0,207,0,75,0,0,0,180,0,20,0,201,0,133,0,97,0,242,0,221,0,136,0,115,0,255,0,249,0,244,0,17,0,53,0,200,0,100,0,203,0,156,0,134,0,163,0,0,0,249,0,0,0,92,0,186,0,0,0,0,0,0,0,0,0,224,0,0,0,219,0,93,0,202,0,0,0,70,0,176,0,64,0,119,0,0,0,95,0,134,0,74,0,178,0,139,0,235,0,45,0,168,0,125,0,161,0,42,0,151,0,228,0,0,0,170,0,45,0,180,0,225,0,10,0,23,0,0,0,0,0,0,0,129,0,176,0,209,0,73,0,0,0,198,0,94,0,125,0,66,0,26,0,203,0,3,0,116,0,115,0,143,0,0,0,23,0,76,0,73,0,30,0,184,0,59,0,236,0,240,0,100,0,155,0,172,0,24,0,105,0,213,0,245,0,120,0,0,0,227,0,178,0,126,0,3,0,0,0,58,0,57,0,213,0,0,0,67,0,0,0,158,0,0,0,251,0,192,0,250,0,108,0,168,0,153,0,189,0,0,0,79,0,42,0,218,0,120,0,136,0,0,0,0,0,167,0,184,0,12,0,165,0,187,0,188,0,140,0,0,0,204,0,55,0,71,0,188,0,197,0,53,0,62,0,2,0,7,0,9,0,128,0,63,0,137,0,87,0,252,0,126,0,50,0,0,0,194,0,149,0,196,0,109,0,122,0,174,0,0,0,191,0,218,0,6,0,254,0,0,0,87,0,19,0,0,0,111,0,99,0,145,0,0,0,222,0,212,0,197,0,196,0,76,0,216,0,172,0,143,0,28,0,1,0,79,0,62,0,238,0,49,0,31,0,1,0,28,0,49,0,224,0,225,0,0,0,250,0,0,0,4,0,0,0,23,0,181,0,0,0,68,0,41,0,198,0,173,0,85,0,0,0,106,0,30,0,132,0,230,0,77,0,0,0,0,0,0,0,0,0,0,0,129,0,35,0,228,0,188,0,0,0,3,0,143,0,0,0,76,0,226,0,121,0,42,0,0,0,164,0,218,0,95,0,9,0,113,0,53,0,0,0,148,0,11,0,69,0,158,0,40,0,199,0,17,0,63,0,234,0,29,0,6,0,41,0,0,0,136,0,24,0,181,0,0,0,0,0,171,0,27,0,239,0,81,0,3,0,219,0,0,0,87,0,111,0,2,0,220,0,227,0,79,0,0,0,0,0,229,0,56,0,70,0,0,0,45,0,199,0,0,0,177,0,185,0,146,0,58,0,123,0,94,0,41,0,0,0,252,0,0,0,0,0,227,0,171,0,179,0,221,0,48,0,65,0,171,0,21,0,132,0,0,0,105,0,130,0,128,0,20,0,95,0,138,0,0,0,164,0,27,0,0,0,31,0,36,0,224,0,25,0,219,0,63,0,23,0,252,0,0,0,63,0,244,0,187,0,98,0,129,0,177,0,0,0,142,0,84,0,102,0,76,0,253,0,0,0,34,0,252,0,149,0,0,0,23,0,0,0,231,0,12,0,0,0,233,0,28,0,114,0,83,0,172,0,51,0,57,0,63,0,0,0,18,0,0,0,58,0,0,0,106,0,101,0,0,0,0,0,96,0,206,0,0,0,64,0,129,0,0,0,214,0,159,0,228,0,120,0,18,0,33,0,0,0,240,0,238,0,145,0,232,0,25,0,1,0,168,0,253,0,109,0,124,0,21,0,174,0,37,0,255,0,205,0,47,0,214,0,0,0,0,0,167,0,111,0,0,0,113,0,83,0,79,0,180,0,0,0,14,0,222,0,195,0,220,0,236,0,200,0,0,0,0,0,12,0,0,0,28,0,78,0,89,0,16,0,222,0,181,0,229,0,85,0,121,0,253,0,122,0,100,0,181,0,99,0,62,0,180,0,12,0,117,0,185,0,239,0,155,0,56,0,122,0,230,0,0,0,132,0);
signal scenario_full  : scenario_type := (195,31,195,30,152,31,144,31,75,31,181,31,110,31,239,31,61,31,115,31,115,30,39,31,68,31,161,31,217,31,226,31,146,31,146,30,235,31,116,31,238,31,80,31,37,31,37,30,37,29,21,31,171,31,1,31,18,31,237,31,200,31,249,31,249,30,61,31,149,31,242,31,242,30,242,29,233,31,233,30,207,31,106,31,31,31,217,31,151,31,99,31,129,31,183,31,56,31,229,31,188,31,129,31,99,31,108,31,65,31,78,31,101,31,190,31,6,31,102,31,6,31,19,31,122,31,14,31,14,30,220,31,80,31,168,31,146,31,146,30,52,31,52,30,52,29,52,28,222,31,188,31,188,30,112,31,74,31,115,31,115,30,187,31,51,31,96,31,46,31,10,31,68,31,99,31,155,31,239,31,147,31,222,31,33,31,2,31,2,30,128,31,140,31,240,31,37,31,153,31,153,30,152,31,152,30,234,31,214,31,181,31,89,31,89,30,32,31,161,31,5,31,5,30,5,29,131,31,16,31,74,31,236,31,236,30,64,31,153,31,76,31,89,31,23,31,23,30,8,31,174,31,102,31,102,30,169,31,64,31,64,30,31,31,249,31,249,30,239,31,220,31,220,30,84,31,232,31,116,31,253,31,96,31,19,31,167,31,66,31,15,31,15,30,17,31,76,31,14,31,14,30,47,31,241,31,183,31,128,31,5,31,57,31,20,31,49,31,49,30,218,31,48,31,24,31,94,31,176,31,174,31,51,31,199,31,14,31,138,31,138,30,138,29,247,31,95,31,241,31,177,31,188,31,217,31,25,31,243,31,126,31,196,31,51,31,236,31,106,31,107,31,107,30,140,31,167,31,167,30,167,29,249,31,162,31,123,31,123,30,66,31,66,30,226,31,27,31,84,31,210,31,134,31,165,31,57,31,207,31,57,31,57,30,75,31,52,31,245,31,179,31,168,31,168,30,235,31,87,31,207,31,75,31,75,30,180,31,20,31,201,31,133,31,97,31,242,31,221,31,136,31,115,31,255,31,249,31,244,31,17,31,53,31,200,31,100,31,203,31,156,31,134,31,163,31,163,30,249,31,249,30,92,31,186,31,186,30,186,29,186,28,186,27,224,31,224,30,219,31,93,31,202,31,202,30,70,31,176,31,64,31,119,31,119,30,95,31,134,31,74,31,178,31,139,31,235,31,45,31,168,31,125,31,161,31,42,31,151,31,228,31,228,30,170,31,45,31,180,31,225,31,10,31,23,31,23,30,23,29,23,28,129,31,176,31,209,31,73,31,73,30,198,31,94,31,125,31,66,31,26,31,203,31,3,31,116,31,115,31,143,31,143,30,23,31,76,31,73,31,30,31,184,31,59,31,236,31,240,31,100,31,155,31,172,31,24,31,105,31,213,31,245,31,120,31,120,30,227,31,178,31,126,31,3,31,3,30,58,31,57,31,213,31,213,30,67,31,67,30,158,31,158,30,251,31,192,31,250,31,108,31,168,31,153,31,189,31,189,30,79,31,42,31,218,31,120,31,136,31,136,30,136,29,167,31,184,31,12,31,165,31,187,31,188,31,140,31,140,30,204,31,55,31,71,31,188,31,197,31,53,31,62,31,2,31,7,31,9,31,128,31,63,31,137,31,87,31,252,31,126,31,50,31,50,30,194,31,149,31,196,31,109,31,122,31,174,31,174,30,191,31,218,31,6,31,254,31,254,30,87,31,19,31,19,30,111,31,99,31,145,31,145,30,222,31,212,31,197,31,196,31,76,31,216,31,172,31,143,31,28,31,1,31,79,31,62,31,238,31,49,31,31,31,1,31,28,31,49,31,224,31,225,31,225,30,250,31,250,30,4,31,4,30,23,31,181,31,181,30,68,31,41,31,198,31,173,31,85,31,85,30,106,31,30,31,132,31,230,31,77,31,77,30,77,29,77,28,77,27,77,26,129,31,35,31,228,31,188,31,188,30,3,31,143,31,143,30,76,31,226,31,121,31,42,31,42,30,164,31,218,31,95,31,9,31,113,31,53,31,53,30,148,31,11,31,69,31,158,31,40,31,199,31,17,31,63,31,234,31,29,31,6,31,41,31,41,30,136,31,24,31,181,31,181,30,181,29,171,31,27,31,239,31,81,31,3,31,219,31,219,30,87,31,111,31,2,31,220,31,227,31,79,31,79,30,79,29,229,31,56,31,70,31,70,30,45,31,199,31,199,30,177,31,185,31,146,31,58,31,123,31,94,31,41,31,41,30,252,31,252,30,252,29,227,31,171,31,179,31,221,31,48,31,65,31,171,31,21,31,132,31,132,30,105,31,130,31,128,31,20,31,95,31,138,31,138,30,164,31,27,31,27,30,31,31,36,31,224,31,25,31,219,31,63,31,23,31,252,31,252,30,63,31,244,31,187,31,98,31,129,31,177,31,177,30,142,31,84,31,102,31,76,31,253,31,253,30,34,31,252,31,149,31,149,30,23,31,23,30,231,31,12,31,12,30,233,31,28,31,114,31,83,31,172,31,51,31,57,31,63,31,63,30,18,31,18,30,58,31,58,30,106,31,101,31,101,30,101,29,96,31,206,31,206,30,64,31,129,31,129,30,214,31,159,31,228,31,120,31,18,31,33,31,33,30,240,31,238,31,145,31,232,31,25,31,1,31,168,31,253,31,109,31,124,31,21,31,174,31,37,31,255,31,205,31,47,31,214,31,214,30,214,29,167,31,111,31,111,30,113,31,83,31,79,31,180,31,180,30,14,31,222,31,195,31,220,31,236,31,200,31,200,30,200,29,12,31,12,30,28,31,78,31,89,31,16,31,222,31,181,31,229,31,85,31,121,31,253,31,122,31,100,31,181,31,99,31,62,31,180,31,12,31,117,31,185,31,239,31,155,31,56,31,122,31,230,31,230,30,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
