-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 840;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,200,0,231,0,0,0,145,0,108,0,213,0,0,0,158,0,2,0,178,0,81,0,217,0,108,0,195,0,62,0,210,0,5,0,99,0,3,0,0,0,10,0,15,0,140,0,136,0,0,0,205,0,151,0,77,0,0,0,72,0,50,0,167,0,0,0,0,0,0,0,90,0,0,0,0,0,184,0,107,0,108,0,0,0,136,0,31,0,216,0,220,0,130,0,127,0,0,0,69,0,184,0,11,0,124,0,75,0,247,0,92,0,64,0,131,0,83,0,223,0,236,0,143,0,59,0,185,0,187,0,139,0,188,0,78,0,189,0,0,0,20,0,170,0,216,0,182,0,103,0,240,0,30,0,160,0,222,0,47,0,0,0,85,0,100,0,102,0,0,0,0,0,192,0,117,0,0,0,72,0,254,0,1,0,131,0,111,0,201,0,62,0,4,0,255,0,182,0,192,0,0,0,34,0,13,0,116,0,41,0,57,0,231,0,38,0,223,0,43,0,213,0,246,0,20,0,208,0,0,0,131,0,123,0,160,0,146,0,223,0,89,0,133,0,235,0,175,0,223,0,253,0,132,0,57,0,0,0,115,0,182,0,166,0,98,0,56,0,214,0,0,0,246,0,70,0,99,0,228,0,207,0,0,0,182,0,210,0,169,0,225,0,41,0,134,0,141,0,0,0,105,0,83,0,221,0,25,0,13,0,0,0,118,0,44,0,214,0,174,0,98,0,169,0,211,0,47,0,90,0,241,0,26,0,0,0,62,0,0,0,217,0,164,0,0,0,104,0,39,0,55,0,0,0,190,0,122,0,0,0,149,0,0,0,227,0,0,0,62,0,117,0,0,0,34,0,165,0,244,0,11,0,125,0,7,0,72,0,204,0,0,0,0,0,11,0,0,0,163,0,52,0,0,0,181,0,170,0,149,0,16,0,73,0,114,0,47,0,0,0,89,0,249,0,170,0,179,0,231,0,193,0,202,0,26,0,57,0,178,0,175,0,172,0,93,0,209,0,0,0,220,0,0,0,79,0,0,0,28,0,170,0,76,0,158,0,0,0,7,0,196,0,0,0,13,0,153,0,211,0,0,0,133,0,86,0,74,0,0,0,0,0,121,0,61,0,0,0,87,0,0,0,80,0,0,0,230,0,0,0,97,0,120,0,237,0,2,0,239,0,19,0,0,0,163,0,26,0,233,0,134,0,74,0,54,0,229,0,7,0,31,0,40,0,127,0,141,0,120,0,34,0,0,0,225,0,146,0,119,0,0,0,213,0,219,0,27,0,81,0,0,0,35,0,120,0,8,0,57,0,0,0,251,0,0,0,223,0,230,0,0,0,184,0,183,0,81,0,103,0,44,0,109,0,0,0,145,0,0,0,69,0,233,0,54,0,242,0,160,0,244,0,0,0,0,0,194,0,0,0,152,0,209,0,211,0,138,0,170,0,138,0,42,0,11,0,17,0,185,0,180,0,79,0,98,0,232,0,221,0,246,0,134,0,21,0,68,0,0,0,26,0,98,0,167,0,240,0,71,0,75,0,142,0,221,0,0,0,197,0,252,0,18,0,249,0,0,0,105,0,198,0,0,0,243,0,176,0,55,0,255,0,64,0,0,0,108,0,70,0,6,0,154,0,23,0,66,0,214,0,125,0,75,0,23,0,0,0,105,0,109,0,248,0,143,0,9,0,147,0,255,0,0,0,12,0,0,0,0,0,252,0,0,0,114,0,0,0,107,0,0,0,214,0,211,0,99,0,232,0,1,0,224,0,19,0,102,0,179,0,184,0,253,0,213,0,104,0,100,0,177,0,97,0,227,0,8,0,41,0,160,0,216,0,39,0,186,0,190,0,95,0,31,0,160,0,215,0,0,0,20,0,131,0,0,0,216,0,195,0,208,0,184,0,220,0,0,0,86,0,115,0,127,0,141,0,214,0,37,0,8,0,176,0,0,0,201,0,237,0,0,0,149,0,250,0,80,0,15,0,162,0,252,0,42,0,0,0,0,0,0,0,117,0,189,0,210,0,26,0,207,0,85,0,0,0,162,0,0,0,143,0,39,0,0,0,187,0,0,0,123,0,202,0,215,0,69,0,201,0,189,0,71,0,0,0,177,0,242,0,29,0,146,0,107,0,3,0,0,0,36,0,0,0,70,0,122,0,48,0,200,0,175,0,119,0,162,0,202,0,111,0,211,0,157,0,27,0,56,0,155,0,0,0,171,0,79,0,15,0,54,0,227,0,85,0,14,0,227,0,64,0,40,0,243,0,227,0,67,0,30,0,159,0,0,0,106,0,11,0,248,0,163,0,214,0,60,0,153,0,210,0,0,0,205,0,246,0,69,0,217,0,0,0,184,0,113,0,198,0,0,0,192,0,117,0,0,0,114,0,205,0,0,0,146,0,29,0,0,0,53,0,241,0,68,0,160,0,0,0,33,0,243,0,0,0,0,0,116,0,183,0,0,0,240,0,230,0,0,0,148,0,0,0,94,0,89,0,113,0,196,0,29,0,214,0,83,0,146,0,0,0,186,0,19,0,87,0,220,0,73,0,161,0,0,0,15,0,249,0,0,0,123,0,0,0,224,0,211,0,246,0,0,0,78,0,0,0,236,0,0,0,167,0,0,0,22,0,230,0,0,0,23,0,238,0,152,0,33,0,0,0,93,0,171,0,135,0,77,0,49,0,160,0,0,0,214,0,0,0,104,0,112,0,0,0,199,0,0,0,190,0,34,0,99,0,19,0,0,0,0,0,244,0,197,0,145,0,22,0,0,0,39,0,192,0,59,0,67,0,203,0,137,0,223,0,0,0,0,0,218,0,210,0,209,0,88,0,23,0,63,0,55,0,0,0,0,0,81,0,194,0,0,0,120,0,0,0,172,0,68,0,128,0,198,0,0,0,230,0,245,0,82,0,59,0,246,0,204,0,246,0,53,0,31,0,83,0,237,0,206,0,95,0,179,0,202,0,151,0,50,0,180,0,153,0,132,0,84,0,0,0,105,0,142,0,149,0,153,0,57,0,2,0,106,0,36,0,34,0,0,0,0,0,0,0,32,0,53,0,142,0,105,0,139,0,217,0,197,0,235,0,137,0,201,0,166,0,109,0,200,0,193,0,120,0,0,0,152,0,136,0,201,0,222,0,123,0,142,0,91,0,0,0,173,0,130,0,218,0,100,0,139,0,147,0,229,0,82,0,247,0,140,0,53,0,0,0,91,0,0,0,53,0,14,0,222,0,77,0,122,0,22,0,182,0,194,0,43,0,237,0,134,0,0,0,80,0,186,0,1,0,0,0,244,0,148,0,150,0,1,0,0,0,0,0,0,0,105,0,75,0,57,0,1,0,235,0,96,0,0,0,0,0,153,0,2,0,0,0,142,0,133,0,108,0,230,0,143,0,65,0,120,0,49,0,133,0,0,0,134,0,216,0,188,0,206,0,71,0,49,0,190,0,240,0,133,0,225,0,0,0,248,0,43,0,29,0,71,0,0,0,130,0,179,0,109,0,0,0,12,0,0,0,162,0,31,0,190,0,230,0,0,0,1,0,33,0,154,0,152,0,247,0,0,0,19,0,120,0,0,0,79,0,251,0,119,0,160,0,209,0,0,0,180,0,0,0,61,0,241,0,7,0,255,0,205,0,0,0,52,0,138,0,26,0,0,0,217,0,0,0,97,0,88,0,9,0,241,0,98,0,40,0,226,0,233,0,228,0,0,0,1,0,251,0,85,0,0,0,0,0,71,0,208,0,86,0,252,0,109,0,240,0,234,0,53,0);
signal scenario_full  : scenario_type := (0,0,200,31,231,31,231,30,145,31,108,31,213,31,213,30,158,31,2,31,178,31,81,31,217,31,108,31,195,31,62,31,210,31,5,31,99,31,3,31,3,30,10,31,15,31,140,31,136,31,136,30,205,31,151,31,77,31,77,30,72,31,50,31,167,31,167,30,167,29,167,28,90,31,90,30,90,29,184,31,107,31,108,31,108,30,136,31,31,31,216,31,220,31,130,31,127,31,127,30,69,31,184,31,11,31,124,31,75,31,247,31,92,31,64,31,131,31,83,31,223,31,236,31,143,31,59,31,185,31,187,31,139,31,188,31,78,31,189,31,189,30,20,31,170,31,216,31,182,31,103,31,240,31,30,31,160,31,222,31,47,31,47,30,85,31,100,31,102,31,102,30,102,29,192,31,117,31,117,30,72,31,254,31,1,31,131,31,111,31,201,31,62,31,4,31,255,31,182,31,192,31,192,30,34,31,13,31,116,31,41,31,57,31,231,31,38,31,223,31,43,31,213,31,246,31,20,31,208,31,208,30,131,31,123,31,160,31,146,31,223,31,89,31,133,31,235,31,175,31,223,31,253,31,132,31,57,31,57,30,115,31,182,31,166,31,98,31,56,31,214,31,214,30,246,31,70,31,99,31,228,31,207,31,207,30,182,31,210,31,169,31,225,31,41,31,134,31,141,31,141,30,105,31,83,31,221,31,25,31,13,31,13,30,118,31,44,31,214,31,174,31,98,31,169,31,211,31,47,31,90,31,241,31,26,31,26,30,62,31,62,30,217,31,164,31,164,30,104,31,39,31,55,31,55,30,190,31,122,31,122,30,149,31,149,30,227,31,227,30,62,31,117,31,117,30,34,31,165,31,244,31,11,31,125,31,7,31,72,31,204,31,204,30,204,29,11,31,11,30,163,31,52,31,52,30,181,31,170,31,149,31,16,31,73,31,114,31,47,31,47,30,89,31,249,31,170,31,179,31,231,31,193,31,202,31,26,31,57,31,178,31,175,31,172,31,93,31,209,31,209,30,220,31,220,30,79,31,79,30,28,31,170,31,76,31,158,31,158,30,7,31,196,31,196,30,13,31,153,31,211,31,211,30,133,31,86,31,74,31,74,30,74,29,121,31,61,31,61,30,87,31,87,30,80,31,80,30,230,31,230,30,97,31,120,31,237,31,2,31,239,31,19,31,19,30,163,31,26,31,233,31,134,31,74,31,54,31,229,31,7,31,31,31,40,31,127,31,141,31,120,31,34,31,34,30,225,31,146,31,119,31,119,30,213,31,219,31,27,31,81,31,81,30,35,31,120,31,8,31,57,31,57,30,251,31,251,30,223,31,230,31,230,30,184,31,183,31,81,31,103,31,44,31,109,31,109,30,145,31,145,30,69,31,233,31,54,31,242,31,160,31,244,31,244,30,244,29,194,31,194,30,152,31,209,31,211,31,138,31,170,31,138,31,42,31,11,31,17,31,185,31,180,31,79,31,98,31,232,31,221,31,246,31,134,31,21,31,68,31,68,30,26,31,98,31,167,31,240,31,71,31,75,31,142,31,221,31,221,30,197,31,252,31,18,31,249,31,249,30,105,31,198,31,198,30,243,31,176,31,55,31,255,31,64,31,64,30,108,31,70,31,6,31,154,31,23,31,66,31,214,31,125,31,75,31,23,31,23,30,105,31,109,31,248,31,143,31,9,31,147,31,255,31,255,30,12,31,12,30,12,29,252,31,252,30,114,31,114,30,107,31,107,30,214,31,211,31,99,31,232,31,1,31,224,31,19,31,102,31,179,31,184,31,253,31,213,31,104,31,100,31,177,31,97,31,227,31,8,31,41,31,160,31,216,31,39,31,186,31,190,31,95,31,31,31,160,31,215,31,215,30,20,31,131,31,131,30,216,31,195,31,208,31,184,31,220,31,220,30,86,31,115,31,127,31,141,31,214,31,37,31,8,31,176,31,176,30,201,31,237,31,237,30,149,31,250,31,80,31,15,31,162,31,252,31,42,31,42,30,42,29,42,28,117,31,189,31,210,31,26,31,207,31,85,31,85,30,162,31,162,30,143,31,39,31,39,30,187,31,187,30,123,31,202,31,215,31,69,31,201,31,189,31,71,31,71,30,177,31,242,31,29,31,146,31,107,31,3,31,3,30,36,31,36,30,70,31,122,31,48,31,200,31,175,31,119,31,162,31,202,31,111,31,211,31,157,31,27,31,56,31,155,31,155,30,171,31,79,31,15,31,54,31,227,31,85,31,14,31,227,31,64,31,40,31,243,31,227,31,67,31,30,31,159,31,159,30,106,31,11,31,248,31,163,31,214,31,60,31,153,31,210,31,210,30,205,31,246,31,69,31,217,31,217,30,184,31,113,31,198,31,198,30,192,31,117,31,117,30,114,31,205,31,205,30,146,31,29,31,29,30,53,31,241,31,68,31,160,31,160,30,33,31,243,31,243,30,243,29,116,31,183,31,183,30,240,31,230,31,230,30,148,31,148,30,94,31,89,31,113,31,196,31,29,31,214,31,83,31,146,31,146,30,186,31,19,31,87,31,220,31,73,31,161,31,161,30,15,31,249,31,249,30,123,31,123,30,224,31,211,31,246,31,246,30,78,31,78,30,236,31,236,30,167,31,167,30,22,31,230,31,230,30,23,31,238,31,152,31,33,31,33,30,93,31,171,31,135,31,77,31,49,31,160,31,160,30,214,31,214,30,104,31,112,31,112,30,199,31,199,30,190,31,34,31,99,31,19,31,19,30,19,29,244,31,197,31,145,31,22,31,22,30,39,31,192,31,59,31,67,31,203,31,137,31,223,31,223,30,223,29,218,31,210,31,209,31,88,31,23,31,63,31,55,31,55,30,55,29,81,31,194,31,194,30,120,31,120,30,172,31,68,31,128,31,198,31,198,30,230,31,245,31,82,31,59,31,246,31,204,31,246,31,53,31,31,31,83,31,237,31,206,31,95,31,179,31,202,31,151,31,50,31,180,31,153,31,132,31,84,31,84,30,105,31,142,31,149,31,153,31,57,31,2,31,106,31,36,31,34,31,34,30,34,29,34,28,32,31,53,31,142,31,105,31,139,31,217,31,197,31,235,31,137,31,201,31,166,31,109,31,200,31,193,31,120,31,120,30,152,31,136,31,201,31,222,31,123,31,142,31,91,31,91,30,173,31,130,31,218,31,100,31,139,31,147,31,229,31,82,31,247,31,140,31,53,31,53,30,91,31,91,30,53,31,14,31,222,31,77,31,122,31,22,31,182,31,194,31,43,31,237,31,134,31,134,30,80,31,186,31,1,31,1,30,244,31,148,31,150,31,1,31,1,30,1,29,1,28,105,31,75,31,57,31,1,31,235,31,96,31,96,30,96,29,153,31,2,31,2,30,142,31,133,31,108,31,230,31,143,31,65,31,120,31,49,31,133,31,133,30,134,31,216,31,188,31,206,31,71,31,49,31,190,31,240,31,133,31,225,31,225,30,248,31,43,31,29,31,71,31,71,30,130,31,179,31,109,31,109,30,12,31,12,30,162,31,31,31,190,31,230,31,230,30,1,31,33,31,154,31,152,31,247,31,247,30,19,31,120,31,120,30,79,31,251,31,119,31,160,31,209,31,209,30,180,31,180,30,61,31,241,31,7,31,255,31,205,31,205,30,52,31,138,31,26,31,26,30,217,31,217,30,97,31,88,31,9,31,241,31,98,31,40,31,226,31,233,31,228,31,228,30,1,31,251,31,85,31,85,30,85,29,71,31,208,31,86,31,252,31,109,31,240,31,234,31,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
