-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_559 is
end project_tb_559;

architecture project_tb_arch_559 of project_tb_559 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 700;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (46,0,246,0,36,0,0,0,103,0,70,0,128,0,0,0,246,0,124,0,169,0,91,0,122,0,136,0,69,0,172,0,144,0,103,0,175,0,119,0,0,0,229,0,60,0,78,0,0,0,0,0,102,0,0,0,7,0,210,0,0,0,159,0,163,0,247,0,56,0,173,0,9,0,167,0,246,0,62,0,106,0,0,0,112,0,1,0,97,0,61,0,9,0,143,0,0,0,202,0,126,0,201,0,0,0,244,0,93,0,0,0,27,0,0,0,0,0,5,0,140,0,117,0,56,0,0,0,0,0,112,0,101,0,154,0,0,0,229,0,212,0,118,0,0,0,103,0,0,0,187,0,218,0,56,0,56,0,105,0,133,0,185,0,172,0,163,0,118,0,36,0,2,0,44,0,148,0,209,0,136,0,194,0,249,0,144,0,170,0,154,0,166,0,184,0,81,0,163,0,122,0,170,0,255,0,225,0,160,0,56,0,0,0,0,0,112,0,0,0,235,0,53,0,38,0,53,0,151,0,197,0,38,0,0,0,0,0,51,0,153,0,51,0,119,0,129,0,215,0,141,0,80,0,0,0,238,0,37,0,185,0,146,0,0,0,50,0,0,0,199,0,0,0,156,0,0,0,6,0,238,0,173,0,12,0,146,0,231,0,56,0,226,0,73,0,0,0,100,0,45,0,152,0,99,0,80,0,237,0,48,0,242,0,204,0,74,0,119,0,53,0,167,0,89,0,0,0,76,0,45,0,170,0,0,0,136,0,214,0,179,0,211,0,162,0,101,0,80,0,0,0,161,0,144,0,126,0,1,0,0,0,50,0,133,0,234,0,189,0,236,0,4,0,0,0,245,0,195,0,203,0,107,0,33,0,0,0,0,0,232,0,139,0,111,0,45,0,247,0,176,0,46,0,15,0,213,0,0,0,211,0,101,0,15,0,4,0,53,0,74,0,2,0,237,0,117,0,10,0,0,0,176,0,0,0,192,0,0,0,190,0,0,0,153,0,4,0,0,0,215,0,78,0,36,0,243,0,0,0,0,0,0,0,105,0,201,0,30,0,71,0,235,0,34,0,0,0,0,0,161,0,250,0,15,0,17,0,119,0,242,0,122,0,21,0,48,0,109,0,253,0,95,0,193,0,133,0,191,0,0,0,148,0,173,0,115,0,218,0,70,0,101,0,0,0,21,0,0,0,243,0,161,0,36,0,137,0,30,0,0,0,129,0,136,0,244,0,159,0,75,0,208,0,43,0,209,0,107,0,37,0,0,0,138,0,163,0,250,0,193,0,241,0,230,0,78,0,152,0,104,0,0,0,4,0,82,0,11,0,145,0,51,0,248,0,198,0,0,0,0,0,0,0,128,0,113,0,206,0,20,0,9,0,95,0,62,0,183,0,63,0,53,0,234,0,79,0,52,0,66,0,94,0,196,0,79,0,89,0,68,0,0,0,220,0,125,0,246,0,144,0,182,0,213,0,0,0,200,0,0,0,0,0,25,0,55,0,153,0,226,0,233,0,0,0,92,0,200,0,98,0,210,0,112,0,48,0,21,0,81,0,159,0,95,0,95,0,216,0,0,0,0,0,207,0,159,0,196,0,15,0,120,0,219,0,26,0,216,0,96,0,88,0,195,0,129,0,0,0,94,0,39,0,79,0,91,0,26,0,0,0,126,0,71,0,37,0,0,0,4,0,0,0,228,0,118,0,18,0,142,0,38,0,208,0,117,0,255,0,238,0,0,0,254,0,184,0,167,0,0,0,150,0,89,0,192,0,34,0,247,0,0,0,0,0,157,0,0,0,203,0,81,0,0,0,146,0,0,0,61,0,208,0,53,0,0,0,0,0,141,0,229,0,239,0,89,0,0,0,150,0,0,0,0,0,182,0,64,0,205,0,142,0,123,0,173,0,220,0,0,0,200,0,9,0,208,0,127,0,174,0,0,0,0,0,81,0,156,0,63,0,0,0,180,0,8,0,92,0,20,0,90,0,216,0,148,0,76,0,85,0,100,0,82,0,241,0,9,0,0,0,40,0,155,0,65,0,220,0,100,0,240,0,16,0,200,0,32,0,179,0,66,0,128,0,180,0,0,0,218,0,199,0,0,0,11,0,103,0,133,0,0,0,105,0,0,0,167,0,192,0,129,0,131,0,200,0,83,0,0,0,48,0,227,0,87,0,108,0,252,0,127,0,212,0,0,0,82,0,81,0,0,0,79,0,0,0,0,0,29,0,18,0,0,0,114,0,0,0,84,0,41,0,158,0,0,0,0,0,183,0,170,0,69,0,0,0,12,0,110,0,189,0,179,0,0,0,0,0,0,0,150,0,40,0,172,0,83,0,0,0,160,0,164,0,0,0,0,0,149,0,232,0,30,0,141,0,205,0,0,0,188,0,199,0,34,0,75,0,44,0,152,0,107,0,78,0,80,0,31,0,228,0,73,0,60,0,0,0,237,0,28,0,24,0,245,0,242,0,3,0,4,0,247,0,207,0,44,0,0,0,98,0,192,0,101,0,0,0,142,0,186,0,0,0,84,0,195,0,95,0,103,0,236,0,21,0,225,0,140,0,0,0,129,0,210,0,207,0,6,0,96,0,0,0,86,0,187,0,0,0,33,0,226,0,90,0,186,0,11,0,0,0,0,0,0,0,130,0,0,0,0,0,209,0,129,0,15,0,0,0,202,0,13,0,19,0,129,0,0,0,107,0,0,0,145,0,251,0,255,0,83,0,0,0,69,0,65,0,180,0,218,0,7,0,116,0,123,0,34,0,42,0,96,0,244,0,0,0,70,0,44,0,0,0,0,0,243,0,117,0,128,0,214,0,66,0,116,0,224,0,138,0,152,0,0,0,243,0,229,0,157,0,155,0,38,0,227,0,0,0,0,0,0,0,121,0,40,0,239,0,0,0,48,0,45,0,135,0,0,0,145,0,0,0,56,0,0,0,119,0,47,0,212,0,222,0,97,0,122,0,63,0,9,0,183,0,0,0,82,0,30,0,254,0,0,0,157,0,0,0,100,0,245,0,217,0,66,0,180,0,175,0,34,0,146,0,124,0,0,0,108,0,0,0,237,0,247,0,137,0,227,0,41,0,221,0,0,0,59,0,48,0,68,0,96,0,129,0,80,0,70,0,79,0,23,0,205,0);
signal scenario_full  : scenario_type := (46,31,246,31,36,31,36,30,103,31,70,31,128,31,128,30,246,31,124,31,169,31,91,31,122,31,136,31,69,31,172,31,144,31,103,31,175,31,119,31,119,30,229,31,60,31,78,31,78,30,78,29,102,31,102,30,7,31,210,31,210,30,159,31,163,31,247,31,56,31,173,31,9,31,167,31,246,31,62,31,106,31,106,30,112,31,1,31,97,31,61,31,9,31,143,31,143,30,202,31,126,31,201,31,201,30,244,31,93,31,93,30,27,31,27,30,27,29,5,31,140,31,117,31,56,31,56,30,56,29,112,31,101,31,154,31,154,30,229,31,212,31,118,31,118,30,103,31,103,30,187,31,218,31,56,31,56,31,105,31,133,31,185,31,172,31,163,31,118,31,36,31,2,31,44,31,148,31,209,31,136,31,194,31,249,31,144,31,170,31,154,31,166,31,184,31,81,31,163,31,122,31,170,31,255,31,225,31,160,31,56,31,56,30,56,29,112,31,112,30,235,31,53,31,38,31,53,31,151,31,197,31,38,31,38,30,38,29,51,31,153,31,51,31,119,31,129,31,215,31,141,31,80,31,80,30,238,31,37,31,185,31,146,31,146,30,50,31,50,30,199,31,199,30,156,31,156,30,6,31,238,31,173,31,12,31,146,31,231,31,56,31,226,31,73,31,73,30,100,31,45,31,152,31,99,31,80,31,237,31,48,31,242,31,204,31,74,31,119,31,53,31,167,31,89,31,89,30,76,31,45,31,170,31,170,30,136,31,214,31,179,31,211,31,162,31,101,31,80,31,80,30,161,31,144,31,126,31,1,31,1,30,50,31,133,31,234,31,189,31,236,31,4,31,4,30,245,31,195,31,203,31,107,31,33,31,33,30,33,29,232,31,139,31,111,31,45,31,247,31,176,31,46,31,15,31,213,31,213,30,211,31,101,31,15,31,4,31,53,31,74,31,2,31,237,31,117,31,10,31,10,30,176,31,176,30,192,31,192,30,190,31,190,30,153,31,4,31,4,30,215,31,78,31,36,31,243,31,243,30,243,29,243,28,105,31,201,31,30,31,71,31,235,31,34,31,34,30,34,29,161,31,250,31,15,31,17,31,119,31,242,31,122,31,21,31,48,31,109,31,253,31,95,31,193,31,133,31,191,31,191,30,148,31,173,31,115,31,218,31,70,31,101,31,101,30,21,31,21,30,243,31,161,31,36,31,137,31,30,31,30,30,129,31,136,31,244,31,159,31,75,31,208,31,43,31,209,31,107,31,37,31,37,30,138,31,163,31,250,31,193,31,241,31,230,31,78,31,152,31,104,31,104,30,4,31,82,31,11,31,145,31,51,31,248,31,198,31,198,30,198,29,198,28,128,31,113,31,206,31,20,31,9,31,95,31,62,31,183,31,63,31,53,31,234,31,79,31,52,31,66,31,94,31,196,31,79,31,89,31,68,31,68,30,220,31,125,31,246,31,144,31,182,31,213,31,213,30,200,31,200,30,200,29,25,31,55,31,153,31,226,31,233,31,233,30,92,31,200,31,98,31,210,31,112,31,48,31,21,31,81,31,159,31,95,31,95,31,216,31,216,30,216,29,207,31,159,31,196,31,15,31,120,31,219,31,26,31,216,31,96,31,88,31,195,31,129,31,129,30,94,31,39,31,79,31,91,31,26,31,26,30,126,31,71,31,37,31,37,30,4,31,4,30,228,31,118,31,18,31,142,31,38,31,208,31,117,31,255,31,238,31,238,30,254,31,184,31,167,31,167,30,150,31,89,31,192,31,34,31,247,31,247,30,247,29,157,31,157,30,203,31,81,31,81,30,146,31,146,30,61,31,208,31,53,31,53,30,53,29,141,31,229,31,239,31,89,31,89,30,150,31,150,30,150,29,182,31,64,31,205,31,142,31,123,31,173,31,220,31,220,30,200,31,9,31,208,31,127,31,174,31,174,30,174,29,81,31,156,31,63,31,63,30,180,31,8,31,92,31,20,31,90,31,216,31,148,31,76,31,85,31,100,31,82,31,241,31,9,31,9,30,40,31,155,31,65,31,220,31,100,31,240,31,16,31,200,31,32,31,179,31,66,31,128,31,180,31,180,30,218,31,199,31,199,30,11,31,103,31,133,31,133,30,105,31,105,30,167,31,192,31,129,31,131,31,200,31,83,31,83,30,48,31,227,31,87,31,108,31,252,31,127,31,212,31,212,30,82,31,81,31,81,30,79,31,79,30,79,29,29,31,18,31,18,30,114,31,114,30,84,31,41,31,158,31,158,30,158,29,183,31,170,31,69,31,69,30,12,31,110,31,189,31,179,31,179,30,179,29,179,28,150,31,40,31,172,31,83,31,83,30,160,31,164,31,164,30,164,29,149,31,232,31,30,31,141,31,205,31,205,30,188,31,199,31,34,31,75,31,44,31,152,31,107,31,78,31,80,31,31,31,228,31,73,31,60,31,60,30,237,31,28,31,24,31,245,31,242,31,3,31,4,31,247,31,207,31,44,31,44,30,98,31,192,31,101,31,101,30,142,31,186,31,186,30,84,31,195,31,95,31,103,31,236,31,21,31,225,31,140,31,140,30,129,31,210,31,207,31,6,31,96,31,96,30,86,31,187,31,187,30,33,31,226,31,90,31,186,31,11,31,11,30,11,29,11,28,130,31,130,30,130,29,209,31,129,31,15,31,15,30,202,31,13,31,19,31,129,31,129,30,107,31,107,30,145,31,251,31,255,31,83,31,83,30,69,31,65,31,180,31,218,31,7,31,116,31,123,31,34,31,42,31,96,31,244,31,244,30,70,31,44,31,44,30,44,29,243,31,117,31,128,31,214,31,66,31,116,31,224,31,138,31,152,31,152,30,243,31,229,31,157,31,155,31,38,31,227,31,227,30,227,29,227,28,121,31,40,31,239,31,239,30,48,31,45,31,135,31,135,30,145,31,145,30,56,31,56,30,119,31,47,31,212,31,222,31,97,31,122,31,63,31,9,31,183,31,183,30,82,31,30,31,254,31,254,30,157,31,157,30,100,31,245,31,217,31,66,31,180,31,175,31,34,31,146,31,124,31,124,30,108,31,108,30,237,31,247,31,137,31,227,31,41,31,221,31,221,30,59,31,48,31,68,31,96,31,129,31,80,31,70,31,79,31,23,31,205,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
