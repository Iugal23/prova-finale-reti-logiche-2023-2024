-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_387 is
end project_tb_387;

architecture project_tb_arch_387 of project_tb_387 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 787;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,221,0,46,0,173,0,0,0,247,0,244,0,8,0,138,0,0,0,167,0,172,0,0,0,84,0,156,0,61,0,243,0,0,0,174,0,96,0,0,0,214,0,91,0,4,0,11,0,8,0,223,0,216,0,40,0,58,0,0,0,187,0,181,0,226,0,172,0,75,0,244,0,95,0,231,0,0,0,157,0,116,0,105,0,46,0,209,0,148,0,148,0,129,0,12,0,147,0,73,0,65,0,82,0,164,0,55,0,51,0,186,0,189,0,104,0,0,0,231,0,247,0,118,0,0,0,84,0,246,0,121,0,122,0,0,0,28,0,241,0,0,0,4,0,159,0,66,0,242,0,243,0,76,0,30,0,0,0,161,0,85,0,82,0,0,0,56,0,49,0,12,0,188,0,0,0,0,0,52,0,94,0,0,0,7,0,0,0,188,0,58,0,237,0,50,0,0,0,0,0,0,0,100,0,231,0,110,0,80,0,0,0,74,0,168,0,181,0,51,0,98,0,160,0,0,0,216,0,185,0,247,0,214,0,0,0,249,0,28,0,180,0,116,0,169,0,141,0,0,0,164,0,138,0,175,0,113,0,55,0,42,0,0,0,139,0,95,0,175,0,219,0,155,0,52,0,30,0,0,0,0,0,0,0,174,0,1,0,0,0,0,0,0,0,74,0,145,0,0,0,6,0,0,0,61,0,69,0,189,0,0,0,65,0,150,0,183,0,209,0,0,0,230,0,104,0,95,0,0,0,0,0,191,0,49,0,133,0,25,0,89,0,52,0,102,0,135,0,0,0,208,0,110,0,66,0,157,0,99,0,102,0,48,0,21,0,216,0,218,0,87,0,56,0,216,0,20,0,193,0,253,0,252,0,81,0,40,0,145,0,73,0,90,0,0,0,0,0,133,0,30,0,35,0,210,0,247,0,84,0,251,0,134,0,252,0,0,0,158,0,0,0,0,0,142,0,0,0,239,0,11,0,152,0,0,0,0,0,0,0,0,0,200,0,61,0,28,0,18,0,78,0,0,0,119,0,160,0,230,0,48,0,64,0,0,0,247,0,45,0,197,0,221,0,0,0,237,0,0,0,238,0,0,0,35,0,203,0,7,0,86,0,0,0,255,0,72,0,0,0,0,0,169,0,77,0,205,0,204,0,163,0,145,0,115,0,87,0,33,0,167,0,11,0,229,0,0,0,99,0,71,0,243,0,215,0,232,0,26,0,141,0,155,0,164,0,82,0,188,0,62,0,120,0,109,0,128,0,100,0,216,0,0,0,153,0,82,0,10,0,0,0,249,0,6,0,0,0,11,0,155,0,59,0,223,0,0,0,136,0,0,0,0,0,76,0,16,0,43,0,204,0,6,0,237,0,110,0,0,0,179,0,0,0,249,0,75,0,180,0,71,0,26,0,28,0,76,0,0,0,75,0,102,0,51,0,249,0,238,0,197,0,43,0,185,0,0,0,0,0,119,0,0,0,229,0,0,0,84,0,0,0,0,0,41,0,79,0,0,0,0,0,77,0,0,0,163,0,227,0,235,0,33,0,216,0,15,0,225,0,68,0,0,0,255,0,49,0,95,0,153,0,0,0,198,0,72,0,68,0,175,0,36,0,0,0,38,0,140,0,205,0,0,0,239,0,254,0,136,0,24,0,156,0,141,0,108,0,130,0,196,0,10,0,243,0,200,0,83,0,0,0,0,0,51,0,155,0,23,0,88,0,150,0,0,0,223,0,200,0,228,0,25,0,0,0,149,0,5,0,181,0,220,0,11,0,40,0,245,0,174,0,176,0,163,0,163,0,234,0,211,0,174,0,188,0,250,0,95,0,144,0,0,0,85,0,156,0,0,0,41,0,164,0,0,0,59,0,147,0,195,0,0,0,31,0,0,0,211,0,186,0,131,0,130,0,228,0,167,0,0,0,94,0,24,0,0,0,0,0,19,0,0,0,214,0,0,0,87,0,7,0,124,0,42,0,0,0,62,0,6,0,114,0,130,0,208,0,34,0,0,0,36,0,32,0,240,0,0,0,204,0,137,0,0,0,0,0,181,0,242,0,0,0,116,0,0,0,159,0,53,0,0,0,229,0,96,0,212,0,118,0,35,0,206,0,150,0,182,0,236,0,79,0,0,0,119,0,0,0,0,0,21,0,43,0,108,0,44,0,0,0,99,0,117,0,252,0,131,0,219,0,120,0,0,0,54,0,243,0,188,0,0,0,0,0,148,0,229,0,26,0,175,0,255,0,133,0,219,0,0,0,171,0,0,0,21,0,79,0,31,0,98,0,0,0,70,0,94,0,77,0,179,0,164,0,66,0,71,0,156,0,185,0,89,0,0,0,255,0,74,0,105,0,107,0,16,0,61,0,0,0,34,0,209,0,250,0,0,0,134,0,252,0,0,0,0,0,53,0,244,0,249,0,175,0,238,0,1,0,85,0,137,0,217,0,200,0,195,0,0,0,224,0,147,0,132,0,0,0,191,0,62,0,196,0,68,0,160,0,60,0,143,0,167,0,162,0,185,0,94,0,0,0,251,0,120,0,0,0,23,0,0,0,249,0,179,0,93,0,31,0,42,0,0,0,224,0,88,0,52,0,134,0,43,0,83,0,25,0,0,0,105,0,0,0,197,0,79,0,65,0,124,0,0,0,171,0,153,0,122,0,176,0,0,0,233,0,0,0,31,0,54,0,117,0,228,0,216,0,240,0,225,0,252,0,159,0,219,0,37,0,204,0,14,0,138,0,181,0,164,0,187,0,249,0,21,0,105,0,111,0,209,0,140,0,210,0,190,0,59,0,43,0,213,0,178,0,244,0,64,0,122,0,0,0,253,0,66,0,0,0,105,0,249,0,24,0,0,0,169,0,159,0,0,0,114,0,187,0,160,0,0,0,50,0,0,0,130,0,207,0,255,0,219,0,181,0,186,0,78,0,134,0,69,0,249,0,46,0,0,0,159,0,230,0,209,0,0,0,164,0,228,0,0,0,149,0,201,0,228,0,177,0,0,0,66,0,134,0,160,0,0,0,122,0,220,0,0,0,0,0,237,0,77,0,81,0,0,0,26,0,40,0,188,0,0,0,130,0,45,0,41,0,45,0,16,0,154,0,42,0,253,0,0,0,53,0,64,0,79,0,0,0,232,0,249,0,4,0,241,0,0,0,13,0,0,0,25,0,214,0,251,0,219,0,221,0,124,0,0,0,137,0,0,0,84,0,77,0,0,0,238,0,0,0,95,0,134,0,38,0,135,0,242,0,118,0,0,0,138,0,68,0,0,0,0,0,78,0,76,0,186,0,130,0,157,0,10,0,0,0,5,0,126,0,218,0,169,0,225,0,125,0,182,0,0,0,157,0,175,0,170,0,254,0,0,0,224,0,13,0,0,0,77,0,0,0,0,0,0,0,151,0,0,0,0,0,185,0,116,0,0,0,9,0,225,0,0,0,0,0,172,0,112,0,222,0,0,0,19,0,192,0,0,0,46,0,133,0,158,0,146,0,100,0,0,0,0,0,0,0,155,0,202,0,93,0,252,0,193,0);
signal scenario_full  : scenario_type := (0,0,221,31,46,31,173,31,173,30,247,31,244,31,8,31,138,31,138,30,167,31,172,31,172,30,84,31,156,31,61,31,243,31,243,30,174,31,96,31,96,30,214,31,91,31,4,31,11,31,8,31,223,31,216,31,40,31,58,31,58,30,187,31,181,31,226,31,172,31,75,31,244,31,95,31,231,31,231,30,157,31,116,31,105,31,46,31,209,31,148,31,148,31,129,31,12,31,147,31,73,31,65,31,82,31,164,31,55,31,51,31,186,31,189,31,104,31,104,30,231,31,247,31,118,31,118,30,84,31,246,31,121,31,122,31,122,30,28,31,241,31,241,30,4,31,159,31,66,31,242,31,243,31,76,31,30,31,30,30,161,31,85,31,82,31,82,30,56,31,49,31,12,31,188,31,188,30,188,29,52,31,94,31,94,30,7,31,7,30,188,31,58,31,237,31,50,31,50,30,50,29,50,28,100,31,231,31,110,31,80,31,80,30,74,31,168,31,181,31,51,31,98,31,160,31,160,30,216,31,185,31,247,31,214,31,214,30,249,31,28,31,180,31,116,31,169,31,141,31,141,30,164,31,138,31,175,31,113,31,55,31,42,31,42,30,139,31,95,31,175,31,219,31,155,31,52,31,30,31,30,30,30,29,30,28,174,31,1,31,1,30,1,29,1,28,74,31,145,31,145,30,6,31,6,30,61,31,69,31,189,31,189,30,65,31,150,31,183,31,209,31,209,30,230,31,104,31,95,31,95,30,95,29,191,31,49,31,133,31,25,31,89,31,52,31,102,31,135,31,135,30,208,31,110,31,66,31,157,31,99,31,102,31,48,31,21,31,216,31,218,31,87,31,56,31,216,31,20,31,193,31,253,31,252,31,81,31,40,31,145,31,73,31,90,31,90,30,90,29,133,31,30,31,35,31,210,31,247,31,84,31,251,31,134,31,252,31,252,30,158,31,158,30,158,29,142,31,142,30,239,31,11,31,152,31,152,30,152,29,152,28,152,27,200,31,61,31,28,31,18,31,78,31,78,30,119,31,160,31,230,31,48,31,64,31,64,30,247,31,45,31,197,31,221,31,221,30,237,31,237,30,238,31,238,30,35,31,203,31,7,31,86,31,86,30,255,31,72,31,72,30,72,29,169,31,77,31,205,31,204,31,163,31,145,31,115,31,87,31,33,31,167,31,11,31,229,31,229,30,99,31,71,31,243,31,215,31,232,31,26,31,141,31,155,31,164,31,82,31,188,31,62,31,120,31,109,31,128,31,100,31,216,31,216,30,153,31,82,31,10,31,10,30,249,31,6,31,6,30,11,31,155,31,59,31,223,31,223,30,136,31,136,30,136,29,76,31,16,31,43,31,204,31,6,31,237,31,110,31,110,30,179,31,179,30,249,31,75,31,180,31,71,31,26,31,28,31,76,31,76,30,75,31,102,31,51,31,249,31,238,31,197,31,43,31,185,31,185,30,185,29,119,31,119,30,229,31,229,30,84,31,84,30,84,29,41,31,79,31,79,30,79,29,77,31,77,30,163,31,227,31,235,31,33,31,216,31,15,31,225,31,68,31,68,30,255,31,49,31,95,31,153,31,153,30,198,31,72,31,68,31,175,31,36,31,36,30,38,31,140,31,205,31,205,30,239,31,254,31,136,31,24,31,156,31,141,31,108,31,130,31,196,31,10,31,243,31,200,31,83,31,83,30,83,29,51,31,155,31,23,31,88,31,150,31,150,30,223,31,200,31,228,31,25,31,25,30,149,31,5,31,181,31,220,31,11,31,40,31,245,31,174,31,176,31,163,31,163,31,234,31,211,31,174,31,188,31,250,31,95,31,144,31,144,30,85,31,156,31,156,30,41,31,164,31,164,30,59,31,147,31,195,31,195,30,31,31,31,30,211,31,186,31,131,31,130,31,228,31,167,31,167,30,94,31,24,31,24,30,24,29,19,31,19,30,214,31,214,30,87,31,7,31,124,31,42,31,42,30,62,31,6,31,114,31,130,31,208,31,34,31,34,30,36,31,32,31,240,31,240,30,204,31,137,31,137,30,137,29,181,31,242,31,242,30,116,31,116,30,159,31,53,31,53,30,229,31,96,31,212,31,118,31,35,31,206,31,150,31,182,31,236,31,79,31,79,30,119,31,119,30,119,29,21,31,43,31,108,31,44,31,44,30,99,31,117,31,252,31,131,31,219,31,120,31,120,30,54,31,243,31,188,31,188,30,188,29,148,31,229,31,26,31,175,31,255,31,133,31,219,31,219,30,171,31,171,30,21,31,79,31,31,31,98,31,98,30,70,31,94,31,77,31,179,31,164,31,66,31,71,31,156,31,185,31,89,31,89,30,255,31,74,31,105,31,107,31,16,31,61,31,61,30,34,31,209,31,250,31,250,30,134,31,252,31,252,30,252,29,53,31,244,31,249,31,175,31,238,31,1,31,85,31,137,31,217,31,200,31,195,31,195,30,224,31,147,31,132,31,132,30,191,31,62,31,196,31,68,31,160,31,60,31,143,31,167,31,162,31,185,31,94,31,94,30,251,31,120,31,120,30,23,31,23,30,249,31,179,31,93,31,31,31,42,31,42,30,224,31,88,31,52,31,134,31,43,31,83,31,25,31,25,30,105,31,105,30,197,31,79,31,65,31,124,31,124,30,171,31,153,31,122,31,176,31,176,30,233,31,233,30,31,31,54,31,117,31,228,31,216,31,240,31,225,31,252,31,159,31,219,31,37,31,204,31,14,31,138,31,181,31,164,31,187,31,249,31,21,31,105,31,111,31,209,31,140,31,210,31,190,31,59,31,43,31,213,31,178,31,244,31,64,31,122,31,122,30,253,31,66,31,66,30,105,31,249,31,24,31,24,30,169,31,159,31,159,30,114,31,187,31,160,31,160,30,50,31,50,30,130,31,207,31,255,31,219,31,181,31,186,31,78,31,134,31,69,31,249,31,46,31,46,30,159,31,230,31,209,31,209,30,164,31,228,31,228,30,149,31,201,31,228,31,177,31,177,30,66,31,134,31,160,31,160,30,122,31,220,31,220,30,220,29,237,31,77,31,81,31,81,30,26,31,40,31,188,31,188,30,130,31,45,31,41,31,45,31,16,31,154,31,42,31,253,31,253,30,53,31,64,31,79,31,79,30,232,31,249,31,4,31,241,31,241,30,13,31,13,30,25,31,214,31,251,31,219,31,221,31,124,31,124,30,137,31,137,30,84,31,77,31,77,30,238,31,238,30,95,31,134,31,38,31,135,31,242,31,118,31,118,30,138,31,68,31,68,30,68,29,78,31,76,31,186,31,130,31,157,31,10,31,10,30,5,31,126,31,218,31,169,31,225,31,125,31,182,31,182,30,157,31,175,31,170,31,254,31,254,30,224,31,13,31,13,30,77,31,77,30,77,29,77,28,151,31,151,30,151,29,185,31,116,31,116,30,9,31,225,31,225,30,225,29,172,31,112,31,222,31,222,30,19,31,192,31,192,30,46,31,133,31,158,31,146,31,100,31,100,30,100,29,100,28,155,31,202,31,93,31,252,31,193,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
