-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_749 is
end project_tb_749;

architecture project_tb_arch_749 of project_tb_749 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 480;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (12,0,85,0,173,0,43,0,182,0,40,0,170,0,253,0,246,0,159,0,121,0,0,0,121,0,233,0,11,0,26,0,0,0,162,0,0,0,79,0,245,0,175,0,16,0,155,0,0,0,0,0,9,0,83,0,22,0,106,0,0,0,0,0,197,0,87,0,9,0,235,0,7,0,0,0,254,0,62,0,129,0,223,0,196,0,66,0,35,0,140,0,141,0,10,0,62,0,29,0,176,0,120,0,45,0,160,0,253,0,104,0,232,0,69,0,26,0,240,0,197,0,88,0,114,0,0,0,84,0,0,0,123,0,6,0,173,0,163,0,239,0,214,0,40,0,171,0,52,0,0,0,226,0,218,0,12,0,0,0,12,0,170,0,79,0,14,0,177,0,232,0,184,0,147,0,198,0,0,0,58,0,235,0,167,0,197,0,107,0,60,0,133,0,121,0,60,0,195,0,76,0,0,0,77,0,220,0,108,0,177,0,0,0,98,0,187,0,87,0,184,0,0,0,182,0,25,0,86,0,190,0,35,0,27,0,199,0,13,0,210,0,32,0,72,0,244,0,158,0,173,0,67,0,149,0,182,0,124,0,144,0,194,0,5,0,247,0,194,0,0,0,187,0,172,0,18,0,38,0,0,0,41,0,45,0,0,0,99,0,0,0,152,0,183,0,146,0,48,0,77,0,0,0,232,0,16,0,0,0,158,0,83,0,2,0,109,0,195,0,248,0,0,0,0,0,162,0,0,0,211,0,52,0,0,0,203,0,0,0,204,0,0,0,239,0,17,0,0,0,223,0,133,0,190,0,167,0,189,0,212,0,0,0,159,0,169,0,0,0,240,0,84,0,33,0,187,0,242,0,0,0,42,0,186,0,0,0,106,0,9,0,187,0,167,0,14,0,174,0,0,0,24,0,58,0,0,0,0,0,247,0,229,0,178,0,248,0,0,0,25,0,86,0,0,0,0,0,0,0,134,0,0,0,0,0,25,0,61,0,136,0,104,0,63,0,157,0,0,0,0,0,0,0,98,0,12,0,175,0,69,0,157,0,145,0,187,0,0,0,0,0,246,0,41,0,0,0,233,0,42,0,213,0,60,0,0,0,86,0,142,0,150,0,113,0,51,0,0,0,152,0,191,0,173,0,165,0,55,0,21,0,243,0,0,0,213,0,236,0,0,0,0,0,109,0,41,0,105,0,110,0,144,0,221,0,118,0,184,0,23,0,88,0,0,0,184,0,31,0,157,0,100,0,0,0,176,0,0,0,51,0,192,0,240,0,0,0,209,0,82,0,53,0,207,0,0,0,7,0,209,0,0,0,247,0,94,0,143,0,47,0,42,0,183,0,210,0,9,0,247,0,250,0,163,0,205,0,0,0,35,0,165,0,154,0,25,0,172,0,16,0,0,0,8,0,69,0,0,0,172,0,0,0,26,0,0,0,0,0,82,0,74,0,212,0,168,0,0,0,0,0,219,0,59,0,175,0,245,0,0,0,146,0,193,0,252,0,35,0,204,0,26,0,0,0,119,0,177,0,116,0,250,0,28,0,10,0,22,0,109,0,68,0,77,0,124,0,186,0,165,0,39,0,69,0,7,0,210,0,62,0,146,0,0,0,87,0,0,0,1,0,0,0,147,0,78,0,78,0,114,0,188,0,21,0,3,0,220,0,0,0,175,0,105,0,51,0,94,0,101,0,219,0,43,0,0,0,80,0,199,0,141,0,73,0,140,0,68,0,53,0,66,0,115,0,0,0,90,0,0,0,0,0,0,0,58,0,94,0,70,0,85,0,164,0,181,0,210,0,0,0,64,0,0,0,24,0,25,0,192,0,7,0,255,0,157,0,209,0,170,0,161,0,153,0,220,0,200,0,176,0,120,0,0,0,50,0,142,0,139,0,53,0,143,0,5,0,253,0,108,0,89,0,34,0,58,0,228,0,76,0,82,0,50,0,0,0,236,0,0,0,121,0,55,0,21,0,0,0,249,0,0,0,0,0,206,0,0,0,146,0,194,0,112,0,242,0,171,0,251,0,0,0,0,0,98,0,225,0,157,0,196,0,20,0,185,0,94,0,167,0,144,0,122,0,247,0,222,0,238,0,94,0,235,0,228,0,28,0,14,0,76,0,0,0,0,0,173,0,178,0,110,0,116,0,163,0,0,0);
signal scenario_full  : scenario_type := (12,31,85,31,173,31,43,31,182,31,40,31,170,31,253,31,246,31,159,31,121,31,121,30,121,31,233,31,11,31,26,31,26,30,162,31,162,30,79,31,245,31,175,31,16,31,155,31,155,30,155,29,9,31,83,31,22,31,106,31,106,30,106,29,197,31,87,31,9,31,235,31,7,31,7,30,254,31,62,31,129,31,223,31,196,31,66,31,35,31,140,31,141,31,10,31,62,31,29,31,176,31,120,31,45,31,160,31,253,31,104,31,232,31,69,31,26,31,240,31,197,31,88,31,114,31,114,30,84,31,84,30,123,31,6,31,173,31,163,31,239,31,214,31,40,31,171,31,52,31,52,30,226,31,218,31,12,31,12,30,12,31,170,31,79,31,14,31,177,31,232,31,184,31,147,31,198,31,198,30,58,31,235,31,167,31,197,31,107,31,60,31,133,31,121,31,60,31,195,31,76,31,76,30,77,31,220,31,108,31,177,31,177,30,98,31,187,31,87,31,184,31,184,30,182,31,25,31,86,31,190,31,35,31,27,31,199,31,13,31,210,31,32,31,72,31,244,31,158,31,173,31,67,31,149,31,182,31,124,31,144,31,194,31,5,31,247,31,194,31,194,30,187,31,172,31,18,31,38,31,38,30,41,31,45,31,45,30,99,31,99,30,152,31,183,31,146,31,48,31,77,31,77,30,232,31,16,31,16,30,158,31,83,31,2,31,109,31,195,31,248,31,248,30,248,29,162,31,162,30,211,31,52,31,52,30,203,31,203,30,204,31,204,30,239,31,17,31,17,30,223,31,133,31,190,31,167,31,189,31,212,31,212,30,159,31,169,31,169,30,240,31,84,31,33,31,187,31,242,31,242,30,42,31,186,31,186,30,106,31,9,31,187,31,167,31,14,31,174,31,174,30,24,31,58,31,58,30,58,29,247,31,229,31,178,31,248,31,248,30,25,31,86,31,86,30,86,29,86,28,134,31,134,30,134,29,25,31,61,31,136,31,104,31,63,31,157,31,157,30,157,29,157,28,98,31,12,31,175,31,69,31,157,31,145,31,187,31,187,30,187,29,246,31,41,31,41,30,233,31,42,31,213,31,60,31,60,30,86,31,142,31,150,31,113,31,51,31,51,30,152,31,191,31,173,31,165,31,55,31,21,31,243,31,243,30,213,31,236,31,236,30,236,29,109,31,41,31,105,31,110,31,144,31,221,31,118,31,184,31,23,31,88,31,88,30,184,31,31,31,157,31,100,31,100,30,176,31,176,30,51,31,192,31,240,31,240,30,209,31,82,31,53,31,207,31,207,30,7,31,209,31,209,30,247,31,94,31,143,31,47,31,42,31,183,31,210,31,9,31,247,31,250,31,163,31,205,31,205,30,35,31,165,31,154,31,25,31,172,31,16,31,16,30,8,31,69,31,69,30,172,31,172,30,26,31,26,30,26,29,82,31,74,31,212,31,168,31,168,30,168,29,219,31,59,31,175,31,245,31,245,30,146,31,193,31,252,31,35,31,204,31,26,31,26,30,119,31,177,31,116,31,250,31,28,31,10,31,22,31,109,31,68,31,77,31,124,31,186,31,165,31,39,31,69,31,7,31,210,31,62,31,146,31,146,30,87,31,87,30,1,31,1,30,147,31,78,31,78,31,114,31,188,31,21,31,3,31,220,31,220,30,175,31,105,31,51,31,94,31,101,31,219,31,43,31,43,30,80,31,199,31,141,31,73,31,140,31,68,31,53,31,66,31,115,31,115,30,90,31,90,30,90,29,90,28,58,31,94,31,70,31,85,31,164,31,181,31,210,31,210,30,64,31,64,30,24,31,25,31,192,31,7,31,255,31,157,31,209,31,170,31,161,31,153,31,220,31,200,31,176,31,120,31,120,30,50,31,142,31,139,31,53,31,143,31,5,31,253,31,108,31,89,31,34,31,58,31,228,31,76,31,82,31,50,31,50,30,236,31,236,30,121,31,55,31,21,31,21,30,249,31,249,30,249,29,206,31,206,30,146,31,194,31,112,31,242,31,171,31,251,31,251,30,251,29,98,31,225,31,157,31,196,31,20,31,185,31,94,31,167,31,144,31,122,31,247,31,222,31,238,31,94,31,235,31,228,31,28,31,14,31,76,31,76,30,76,29,173,31,178,31,110,31,116,31,163,31,163,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
