-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_546 is
end project_tb_546;

architecture project_tb_arch_546 of project_tb_546 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 771;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,182,0,125,0,162,0,187,0,0,0,18,0,0,0,100,0,232,0,61,0,173,0,85,0,250,0,0,0,0,0,0,0,145,0,127,0,0,0,210,0,0,0,231,0,98,0,140,0,163,0,203,0,0,0,132,0,17,0,155,0,9,0,59,0,18,0,0,0,38,0,15,0,0,0,239,0,126,0,156,0,71,0,0,0,0,0,96,0,37,0,86,0,9,0,248,0,15,0,184,0,0,0,204,0,143,0,236,0,78,0,196,0,178,0,44,0,194,0,161,0,236,0,236,0,57,0,112,0,226,0,206,0,0,0,128,0,191,0,142,0,44,0,29,0,210,0,241,0,143,0,0,0,0,0,154,0,0,0,144,0,96,0,0,0,0,0,203,0,0,0,171,0,0,0,55,0,0,0,0,0,114,0,77,0,0,0,182,0,171,0,3,0,199,0,76,0,220,0,68,0,235,0,61,0,0,0,176,0,219,0,70,0,0,0,0,0,0,0,112,0,0,0,124,0,159,0,249,0,118,0,147,0,67,0,55,0,151,0,251,0,60,0,83,0,65,0,168,0,153,0,210,0,7,0,44,0,141,0,0,0,69,0,76,0,213,0,212,0,107,0,181,0,0,0,229,0,61,0,8,0,178,0,174,0,255,0,105,0,0,0,168,0,136,0,0,0,138,0,0,0,77,0,136,0,26,0,0,0,115,0,42,0,249,0,83,0,8,0,0,0,121,0,14,0,103,0,120,0,14,0,247,0,0,0,252,0,0,0,168,0,150,0,176,0,253,0,0,0,0,0,42,0,51,0,193,0,171,0,97,0,156,0,36,0,33,0,211,0,193,0,25,0,0,0,112,0,78,0,131,0,165,0,140,0,180,0,0,0,237,0,0,0,229,0,144,0,24,0,188,0,73,0,157,0,44,0,206,0,200,0,62,0,154,0,173,0,86,0,7,0,0,0,201,0,0,0,0,0,232,0,246,0,42,0,0,0,41,0,57,0,65,0,244,0,136,0,161,0,0,0,131,0,239,0,132,0,3,0,0,0,135,0,145,0,232,0,207,0,0,0,15,0,167,0,228,0,190,0,220,0,28,0,106,0,49,0,199,0,226,0,0,0,0,0,0,0,127,0,19,0,214,0,12,0,179,0,199,0,151,0,0,0,60,0,96,0,134,0,73,0,116,0,167,0,1,0,249,0,40,0,218,0,65,0,173,0,222,0,233,0,227,0,95,0,221,0,0,0,30,0,21,0,72,0,0,0,125,0,48,0,0,0,0,0,249,0,0,0,0,0,0,0,65,0,0,0,0,0,0,0,9,0,187,0,136,0,122,0,247,0,138,0,161,0,242,0,0,0,202,0,239,0,33,0,58,0,72,0,9,0,187,0,159,0,30,0,186,0,125,0,109,0,234,0,17,0,0,0,253,0,13,0,237,0,238,0,45,0,159,0,160,0,22,0,200,0,235,0,78,0,163,0,219,0,52,0,182,0,0,0,84,0,2,0,118,0,245,0,0,0,154,0,137,0,197,0,229,0,200,0,54,0,154,0,98,0,216,0,0,0,102,0,218,0,51,0,0,0,242,0,67,0,0,0,98,0,141,0,177,0,247,0,115,0,8,0,120,0,77,0,22,0,141,0,39,0,72,0,213,0,95,0,74,0,56,0,182,0,34,0,243,0,252,0,84,0,197,0,60,0,59,0,110,0,9,0,185,0,160,0,193,0,0,0,140,0,19,0,107,0,108,0,164,0,145,0,0,0,37,0,0,0,205,0,149,0,5,0,0,0,22,0,0,0,0,0,187,0,209,0,0,0,0,0,82,0,0,0,17,0,3,0,151,0,0,0,194,0,254,0,0,0,254,0,47,0,177,0,156,0,217,0,151,0,245,0,213,0,153,0,61,0,0,0,159,0,162,0,80,0,5,0,40,0,123,0,143,0,169,0,15,0,0,0,225,0,170,0,20,0,248,0,252,0,188,0,31,0,205,0,0,0,0,0,147,0,255,0,192,0,5,0,230,0,179,0,162,0,104,0,0,0,138,0,137,0,0,0,143,0,147,0,189,0,18,0,114,0,167,0,179,0,75,0,209,0,158,0,165,0,0,0,73,0,73,0,0,0,30,0,76,0,0,0,33,0,0,0,201,0,192,0,10,0,74,0,0,0,25,0,113,0,34,0,146,0,30,0,187,0,202,0,58,0,101,0,53,0,146,0,17,0,230,0,83,0,66,0,196,0,189,0,113,0,50,0,26,0,138,0,52,0,49,0,116,0,119,0,52,0,52,0,0,0,86,0,200,0,0,0,0,0,152,0,42,0,193,0,28,0,172,0,0,0,98,0,150,0,105,0,131,0,200,0,0,0,11,0,182,0,112,0,190,0,217,0,64,0,24,0,207,0,22,0,195,0,37,0,0,0,246,0,0,0,0,0,205,0,198,0,0,0,210,0,57,0,76,0,0,0,45,0,119,0,138,0,0,0,255,0,94,0,170,0,164,0,39,0,123,0,14,0,242,0,86,0,242,0,51,0,0,0,65,0,0,0,23,0,11,0,0,0,201,0,0,0,149,0,95,0,32,0,230,0,134,0,10,0,0,0,8,0,36,0,211,0,151,0,54,0,135,0,0,0,192,0,184,0,141,0,0,0,149,0,112,0,55,0,239,0,220,0,0,0,81,0,212,0,253,0,26,0,236,0,169,0,74,0,0,0,224,0,255,0,152,0,33,0,0,0,201,0,86,0,101,0,102,0,137,0,169,0,61,0,51,0,0,0,59,0,0,0,84,0,164,0,61,0,37,0,40,0,165,0,129,0,0,0,115,0,29,0,62,0,105,0,25,0,204,0,180,0,87,0,204,0,56,0,4,0,0,0,76,0,196,0,234,0,215,0,67,0,0,0,96,0,0,0,183,0,18,0,0,0,47,0,79,0,251,0,79,0,255,0,0,0,132,0,67,0,179,0,220,0,110,0,25,0,0,0,133,0,234,0,150,0,227,0,137,0,152,0,0,0,0,0,48,0,117,0,177,0,70,0,95,0,119,0,181,0,192,0,99,0,250,0,56,0,22,0,199,0,0,0,201,0,46,0,132,0,171,0,37,0,114,0,20,0,36,0,0,0,30,0,230,0,168,0,0,0,162,0,42,0,158,0,130,0,0,0,0,0,0,0,0,0,192,0,79,0,74,0,131,0,72,0,0,0,204,0,122,0,0,0,0,0,237,0,185,0,214,0,190,0,15,0,0,0,172,0,200,0,21,0,215,0,8,0,154,0,21,0,86,0,97,0,0,0,0,0,205,0,86,0,130,0,17,0,5,0,176,0,247,0,244,0,92,0,73,0,52,0,124,0,0,0,0,0,140,0,128,0,166,0,27,0,133,0,0,0,6,0,54,0,145,0,234,0,0,0,251,0,162,0,251,0,179,0,75,0,9,0,24,0,239,0,0,0,0,0,215,0,190,0,0,0,219,0,208,0);
signal scenario_full  : scenario_type := (0,0,182,31,125,31,162,31,187,31,187,30,18,31,18,30,100,31,232,31,61,31,173,31,85,31,250,31,250,30,250,29,250,28,145,31,127,31,127,30,210,31,210,30,231,31,98,31,140,31,163,31,203,31,203,30,132,31,17,31,155,31,9,31,59,31,18,31,18,30,38,31,15,31,15,30,239,31,126,31,156,31,71,31,71,30,71,29,96,31,37,31,86,31,9,31,248,31,15,31,184,31,184,30,204,31,143,31,236,31,78,31,196,31,178,31,44,31,194,31,161,31,236,31,236,31,57,31,112,31,226,31,206,31,206,30,128,31,191,31,142,31,44,31,29,31,210,31,241,31,143,31,143,30,143,29,154,31,154,30,144,31,96,31,96,30,96,29,203,31,203,30,171,31,171,30,55,31,55,30,55,29,114,31,77,31,77,30,182,31,171,31,3,31,199,31,76,31,220,31,68,31,235,31,61,31,61,30,176,31,219,31,70,31,70,30,70,29,70,28,112,31,112,30,124,31,159,31,249,31,118,31,147,31,67,31,55,31,151,31,251,31,60,31,83,31,65,31,168,31,153,31,210,31,7,31,44,31,141,31,141,30,69,31,76,31,213,31,212,31,107,31,181,31,181,30,229,31,61,31,8,31,178,31,174,31,255,31,105,31,105,30,168,31,136,31,136,30,138,31,138,30,77,31,136,31,26,31,26,30,115,31,42,31,249,31,83,31,8,31,8,30,121,31,14,31,103,31,120,31,14,31,247,31,247,30,252,31,252,30,168,31,150,31,176,31,253,31,253,30,253,29,42,31,51,31,193,31,171,31,97,31,156,31,36,31,33,31,211,31,193,31,25,31,25,30,112,31,78,31,131,31,165,31,140,31,180,31,180,30,237,31,237,30,229,31,144,31,24,31,188,31,73,31,157,31,44,31,206,31,200,31,62,31,154,31,173,31,86,31,7,31,7,30,201,31,201,30,201,29,232,31,246,31,42,31,42,30,41,31,57,31,65,31,244,31,136,31,161,31,161,30,131,31,239,31,132,31,3,31,3,30,135,31,145,31,232,31,207,31,207,30,15,31,167,31,228,31,190,31,220,31,28,31,106,31,49,31,199,31,226,31,226,30,226,29,226,28,127,31,19,31,214,31,12,31,179,31,199,31,151,31,151,30,60,31,96,31,134,31,73,31,116,31,167,31,1,31,249,31,40,31,218,31,65,31,173,31,222,31,233,31,227,31,95,31,221,31,221,30,30,31,21,31,72,31,72,30,125,31,48,31,48,30,48,29,249,31,249,30,249,29,249,28,65,31,65,30,65,29,65,28,9,31,187,31,136,31,122,31,247,31,138,31,161,31,242,31,242,30,202,31,239,31,33,31,58,31,72,31,9,31,187,31,159,31,30,31,186,31,125,31,109,31,234,31,17,31,17,30,253,31,13,31,237,31,238,31,45,31,159,31,160,31,22,31,200,31,235,31,78,31,163,31,219,31,52,31,182,31,182,30,84,31,2,31,118,31,245,31,245,30,154,31,137,31,197,31,229,31,200,31,54,31,154,31,98,31,216,31,216,30,102,31,218,31,51,31,51,30,242,31,67,31,67,30,98,31,141,31,177,31,247,31,115,31,8,31,120,31,77,31,22,31,141,31,39,31,72,31,213,31,95,31,74,31,56,31,182,31,34,31,243,31,252,31,84,31,197,31,60,31,59,31,110,31,9,31,185,31,160,31,193,31,193,30,140,31,19,31,107,31,108,31,164,31,145,31,145,30,37,31,37,30,205,31,149,31,5,31,5,30,22,31,22,30,22,29,187,31,209,31,209,30,209,29,82,31,82,30,17,31,3,31,151,31,151,30,194,31,254,31,254,30,254,31,47,31,177,31,156,31,217,31,151,31,245,31,213,31,153,31,61,31,61,30,159,31,162,31,80,31,5,31,40,31,123,31,143,31,169,31,15,31,15,30,225,31,170,31,20,31,248,31,252,31,188,31,31,31,205,31,205,30,205,29,147,31,255,31,192,31,5,31,230,31,179,31,162,31,104,31,104,30,138,31,137,31,137,30,143,31,147,31,189,31,18,31,114,31,167,31,179,31,75,31,209,31,158,31,165,31,165,30,73,31,73,31,73,30,30,31,76,31,76,30,33,31,33,30,201,31,192,31,10,31,74,31,74,30,25,31,113,31,34,31,146,31,30,31,187,31,202,31,58,31,101,31,53,31,146,31,17,31,230,31,83,31,66,31,196,31,189,31,113,31,50,31,26,31,138,31,52,31,49,31,116,31,119,31,52,31,52,31,52,30,86,31,200,31,200,30,200,29,152,31,42,31,193,31,28,31,172,31,172,30,98,31,150,31,105,31,131,31,200,31,200,30,11,31,182,31,112,31,190,31,217,31,64,31,24,31,207,31,22,31,195,31,37,31,37,30,246,31,246,30,246,29,205,31,198,31,198,30,210,31,57,31,76,31,76,30,45,31,119,31,138,31,138,30,255,31,94,31,170,31,164,31,39,31,123,31,14,31,242,31,86,31,242,31,51,31,51,30,65,31,65,30,23,31,11,31,11,30,201,31,201,30,149,31,95,31,32,31,230,31,134,31,10,31,10,30,8,31,36,31,211,31,151,31,54,31,135,31,135,30,192,31,184,31,141,31,141,30,149,31,112,31,55,31,239,31,220,31,220,30,81,31,212,31,253,31,26,31,236,31,169,31,74,31,74,30,224,31,255,31,152,31,33,31,33,30,201,31,86,31,101,31,102,31,137,31,169,31,61,31,51,31,51,30,59,31,59,30,84,31,164,31,61,31,37,31,40,31,165,31,129,31,129,30,115,31,29,31,62,31,105,31,25,31,204,31,180,31,87,31,204,31,56,31,4,31,4,30,76,31,196,31,234,31,215,31,67,31,67,30,96,31,96,30,183,31,18,31,18,30,47,31,79,31,251,31,79,31,255,31,255,30,132,31,67,31,179,31,220,31,110,31,25,31,25,30,133,31,234,31,150,31,227,31,137,31,152,31,152,30,152,29,48,31,117,31,177,31,70,31,95,31,119,31,181,31,192,31,99,31,250,31,56,31,22,31,199,31,199,30,201,31,46,31,132,31,171,31,37,31,114,31,20,31,36,31,36,30,30,31,230,31,168,31,168,30,162,31,42,31,158,31,130,31,130,30,130,29,130,28,130,27,192,31,79,31,74,31,131,31,72,31,72,30,204,31,122,31,122,30,122,29,237,31,185,31,214,31,190,31,15,31,15,30,172,31,200,31,21,31,215,31,8,31,154,31,21,31,86,31,97,31,97,30,97,29,205,31,86,31,130,31,17,31,5,31,176,31,247,31,244,31,92,31,73,31,52,31,124,31,124,30,124,29,140,31,128,31,166,31,27,31,133,31,133,30,6,31,54,31,145,31,234,31,234,30,251,31,162,31,251,31,179,31,75,31,9,31,24,31,239,31,239,30,239,29,215,31,190,31,190,30,219,31,208,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
