-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_618 is
end project_tb_618;

architecture project_tb_arch_618 of project_tb_618 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 686;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (48,0,145,0,93,0,0,0,114,0,60,0,130,0,193,0,55,0,197,0,161,0,97,0,68,0,96,0,51,0,3,0,229,0,43,0,251,0,0,0,190,0,201,0,32,0,65,0,0,0,124,0,243,0,121,0,0,0,9,0,0,0,145,0,97,0,21,0,130,0,0,0,227,0,122,0,73,0,0,0,105,0,105,0,235,0,0,0,0,0,83,0,82,0,0,0,0,0,94,0,169,0,69,0,182,0,0,0,182,0,60,0,7,0,111,0,73,0,65,0,129,0,62,0,27,0,0,0,0,0,224,0,169,0,185,0,212,0,253,0,18,0,135,0,130,0,229,0,104,0,0,0,184,0,125,0,39,0,239,0,2,0,26,0,98,0,143,0,122,0,150,0,236,0,108,0,125,0,116,0,48,0,1,0,142,0,91,0,146,0,38,0,130,0,0,0,98,0,0,0,57,0,212,0,128,0,145,0,0,0,0,0,24,0,2,0,231,0,10,0,0,0,29,0,238,0,241,0,211,0,248,0,0,0,121,0,86,0,85,0,0,0,216,0,59,0,20,0,114,0,153,0,151,0,205,0,17,0,188,0,44,0,205,0,187,0,104,0,0,0,24,0,227,0,212,0,217,0,17,0,0,0,12,0,0,0,186,0,127,0,46,0,138,0,46,0,12,0,150,0,210,0,220,0,81,0,111,0,97,0,0,0,169,0,108,0,85,0,235,0,164,0,215,0,0,0,176,0,222,0,0,0,33,0,3,0,0,0,13,0,49,0,72,0,56,0,251,0,246,0,42,0,0,0,36,0,121,0,169,0,218,0,0,0,0,0,125,0,68,0,135,0,0,0,148,0,9,0,84,0,154,0,148,0,156,0,247,0,105,0,0,0,45,0,83,0,0,0,0,0,90,0,248,0,180,0,237,0,118,0,251,0,235,0,0,0,17,0,0,0,122,0,113,0,227,0,120,0,0,0,42,0,0,0,0,0,150,0,248,0,114,0,167,0,0,0,7,0,242,0,218,0,64,0,73,0,84,0,92,0,127,0,153,0,237,0,29,0,184,0,163,0,120,0,185,0,157,0,0,0,221,0,96,0,220,0,0,0,0,0,117,0,0,0,1,0,237,0,34,0,216,0,142,0,0,0,252,0,196,0,102,0,42,0,118,0,94,0,68,0,230,0,254,0,0,0,185,0,0,0,49,0,173,0,133,0,0,0,147,0,226,0,113,0,0,0,34,0,124,0,129,0,18,0,155,0,235,0,135,0,91,0,0,0,0,0,229,0,0,0,198,0,150,0,99,0,226,0,0,0,223,0,216,0,0,0,24,0,94,0,81,0,0,0,7,0,0,0,209,0,0,0,0,0,135,0,96,0,148,0,0,0,98,0,0,0,55,0,174,0,0,0,129,0,31,0,0,0,23,0,54,0,237,0,199,0,81,0,76,0,206,0,190,0,86,0,148,0,210,0,218,0,228,0,112,0,108,0,242,0,212,0,175,0,115,0,0,0,0,0,60,0,184,0,66,0,162,0,216,0,61,0,0,0,216,0,188,0,76,0,236,0,39,0,50,0,0,0,127,0,0,0,140,0,93,0,216,0,170,0,72,0,79,0,36,0,113,0,244,0,97,0,8,0,212,0,13,0,220,0,122,0,171,0,117,0,231,0,0,0,241,0,139,0,69,0,173,0,0,0,156,0,24,0,162,0,0,0,208,0,118,0,249,0,129,0,106,0,15,0,71,0,18,0,199,0,133,0,216,0,218,0,0,0,0,0,0,0,192,0,34,0,218,0,116,0,211,0,232,0,242,0,77,0,63,0,63,0,170,0,222,0,201,0,72,0,117,0,86,0,0,0,0,0,226,0,0,0,97,0,0,0,244,0,139,0,228,0,141,0,162,0,0,0,186,0,54,0,71,0,0,0,209,0,73,0,0,0,179,0,233,0,218,0,0,0,184,0,0,0,0,0,60,0,230,0,44,0,150,0,50,0,61,0,204,0,226,0,221,0,225,0,137,0,172,0,95,0,228,0,96,0,0,0,118,0,186,0,125,0,0,0,36,0,129,0,239,0,102,0,23,0,43,0,184,0,213,0,201,0,184,0,51,0,183,0,146,0,223,0,0,0,181,0,50,0,23,0,0,0,62,0,60,0,190,0,245,0,98,0,13,0,94,0,0,0,3,0,73,0,66,0,43,0,0,0,0,0,74,0,43,0,59,0,91,0,0,0,219,0,27,0,99,0,211,0,0,0,142,0,112,0,169,0,0,0,205,0,0,0,179,0,112,0,26,0,138,0,61,0,239,0,49,0,0,0,11,0,0,0,178,0,0,0,186,0,205,0,94,0,217,0,64,0,219,0,119,0,181,0,0,0,39,0,60,0,29,0,103,0,161,0,177,0,247,0,0,0,19,0,94,0,0,0,9,0,53,0,134,0,182,0,16,0,226,0,0,0,157,0,113,0,0,0,161,0,22,0,149,0,208,0,0,0,123,0,242,0,136,0,35,0,235,0,91,0,164,0,7,0,76,0,115,0,162,0,17,0,166,0,100,0,88,0,189,0,156,0,117,0,0,0,67,0,67,0,0,0,174,0,177,0,138,0,193,0,159,0,148,0,199,0,71,0,0,0,42,0,25,0,14,0,255,0,39,0,219,0,0,0,230,0,128,0,9,0,69,0,113,0,32,0,213,0,91,0,192,0,88,0,6,0,158,0,219,0,206,0,242,0,169,0,146,0,187,0,0,0,29,0,182,0,221,0,18,0,8,0,0,0,0,0,0,0,37,0,0,0,210,0,106,0,27,0,28,0,238,0,221,0,46,0,195,0,0,0,102,0,53,0,141,0,159,0,176,0,0,0,138,0,148,0,110,0,219,0,195,0,176,0,0,0,243,0,222,0,0,0,47,0,0,0,127,0,85,0,242,0,209,0,53,0,137,0,0,0,230,0,137,0,64,0,33,0,46,0,0,0,212,0,100,0,103,0,212,0,0,0,139,0,0,0,151,0,153,0,36,0,0,0,221,0,108,0,24,0,160,0,136,0,0,0,36,0,33,0,0,0,214,0,0,0,101,0,49,0,186,0,158,0,0,0);
signal scenario_full  : scenario_type := (48,31,145,31,93,31,93,30,114,31,60,31,130,31,193,31,55,31,197,31,161,31,97,31,68,31,96,31,51,31,3,31,229,31,43,31,251,31,251,30,190,31,201,31,32,31,65,31,65,30,124,31,243,31,121,31,121,30,9,31,9,30,145,31,97,31,21,31,130,31,130,30,227,31,122,31,73,31,73,30,105,31,105,31,235,31,235,30,235,29,83,31,82,31,82,30,82,29,94,31,169,31,69,31,182,31,182,30,182,31,60,31,7,31,111,31,73,31,65,31,129,31,62,31,27,31,27,30,27,29,224,31,169,31,185,31,212,31,253,31,18,31,135,31,130,31,229,31,104,31,104,30,184,31,125,31,39,31,239,31,2,31,26,31,98,31,143,31,122,31,150,31,236,31,108,31,125,31,116,31,48,31,1,31,142,31,91,31,146,31,38,31,130,31,130,30,98,31,98,30,57,31,212,31,128,31,145,31,145,30,145,29,24,31,2,31,231,31,10,31,10,30,29,31,238,31,241,31,211,31,248,31,248,30,121,31,86,31,85,31,85,30,216,31,59,31,20,31,114,31,153,31,151,31,205,31,17,31,188,31,44,31,205,31,187,31,104,31,104,30,24,31,227,31,212,31,217,31,17,31,17,30,12,31,12,30,186,31,127,31,46,31,138,31,46,31,12,31,150,31,210,31,220,31,81,31,111,31,97,31,97,30,169,31,108,31,85,31,235,31,164,31,215,31,215,30,176,31,222,31,222,30,33,31,3,31,3,30,13,31,49,31,72,31,56,31,251,31,246,31,42,31,42,30,36,31,121,31,169,31,218,31,218,30,218,29,125,31,68,31,135,31,135,30,148,31,9,31,84,31,154,31,148,31,156,31,247,31,105,31,105,30,45,31,83,31,83,30,83,29,90,31,248,31,180,31,237,31,118,31,251,31,235,31,235,30,17,31,17,30,122,31,113,31,227,31,120,31,120,30,42,31,42,30,42,29,150,31,248,31,114,31,167,31,167,30,7,31,242,31,218,31,64,31,73,31,84,31,92,31,127,31,153,31,237,31,29,31,184,31,163,31,120,31,185,31,157,31,157,30,221,31,96,31,220,31,220,30,220,29,117,31,117,30,1,31,237,31,34,31,216,31,142,31,142,30,252,31,196,31,102,31,42,31,118,31,94,31,68,31,230,31,254,31,254,30,185,31,185,30,49,31,173,31,133,31,133,30,147,31,226,31,113,31,113,30,34,31,124,31,129,31,18,31,155,31,235,31,135,31,91,31,91,30,91,29,229,31,229,30,198,31,150,31,99,31,226,31,226,30,223,31,216,31,216,30,24,31,94,31,81,31,81,30,7,31,7,30,209,31,209,30,209,29,135,31,96,31,148,31,148,30,98,31,98,30,55,31,174,31,174,30,129,31,31,31,31,30,23,31,54,31,237,31,199,31,81,31,76,31,206,31,190,31,86,31,148,31,210,31,218,31,228,31,112,31,108,31,242,31,212,31,175,31,115,31,115,30,115,29,60,31,184,31,66,31,162,31,216,31,61,31,61,30,216,31,188,31,76,31,236,31,39,31,50,31,50,30,127,31,127,30,140,31,93,31,216,31,170,31,72,31,79,31,36,31,113,31,244,31,97,31,8,31,212,31,13,31,220,31,122,31,171,31,117,31,231,31,231,30,241,31,139,31,69,31,173,31,173,30,156,31,24,31,162,31,162,30,208,31,118,31,249,31,129,31,106,31,15,31,71,31,18,31,199,31,133,31,216,31,218,31,218,30,218,29,218,28,192,31,34,31,218,31,116,31,211,31,232,31,242,31,77,31,63,31,63,31,170,31,222,31,201,31,72,31,117,31,86,31,86,30,86,29,226,31,226,30,97,31,97,30,244,31,139,31,228,31,141,31,162,31,162,30,186,31,54,31,71,31,71,30,209,31,73,31,73,30,179,31,233,31,218,31,218,30,184,31,184,30,184,29,60,31,230,31,44,31,150,31,50,31,61,31,204,31,226,31,221,31,225,31,137,31,172,31,95,31,228,31,96,31,96,30,118,31,186,31,125,31,125,30,36,31,129,31,239,31,102,31,23,31,43,31,184,31,213,31,201,31,184,31,51,31,183,31,146,31,223,31,223,30,181,31,50,31,23,31,23,30,62,31,60,31,190,31,245,31,98,31,13,31,94,31,94,30,3,31,73,31,66,31,43,31,43,30,43,29,74,31,43,31,59,31,91,31,91,30,219,31,27,31,99,31,211,31,211,30,142,31,112,31,169,31,169,30,205,31,205,30,179,31,112,31,26,31,138,31,61,31,239,31,49,31,49,30,11,31,11,30,178,31,178,30,186,31,205,31,94,31,217,31,64,31,219,31,119,31,181,31,181,30,39,31,60,31,29,31,103,31,161,31,177,31,247,31,247,30,19,31,94,31,94,30,9,31,53,31,134,31,182,31,16,31,226,31,226,30,157,31,113,31,113,30,161,31,22,31,149,31,208,31,208,30,123,31,242,31,136,31,35,31,235,31,91,31,164,31,7,31,76,31,115,31,162,31,17,31,166,31,100,31,88,31,189,31,156,31,117,31,117,30,67,31,67,31,67,30,174,31,177,31,138,31,193,31,159,31,148,31,199,31,71,31,71,30,42,31,25,31,14,31,255,31,39,31,219,31,219,30,230,31,128,31,9,31,69,31,113,31,32,31,213,31,91,31,192,31,88,31,6,31,158,31,219,31,206,31,242,31,169,31,146,31,187,31,187,30,29,31,182,31,221,31,18,31,8,31,8,30,8,29,8,28,37,31,37,30,210,31,106,31,27,31,28,31,238,31,221,31,46,31,195,31,195,30,102,31,53,31,141,31,159,31,176,31,176,30,138,31,148,31,110,31,219,31,195,31,176,31,176,30,243,31,222,31,222,30,47,31,47,30,127,31,85,31,242,31,209,31,53,31,137,31,137,30,230,31,137,31,64,31,33,31,46,31,46,30,212,31,100,31,103,31,212,31,212,30,139,31,139,30,151,31,153,31,36,31,36,30,221,31,108,31,24,31,160,31,136,31,136,30,36,31,33,31,33,30,214,31,214,30,101,31,49,31,186,31,158,31,158,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
