-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_704 is
end project_tb_704;

architecture project_tb_arch_704 of project_tb_704 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 629;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,0,0,94,0,143,0,0,0,98,0,0,0,0,0,247,0,95,0,10,0,0,0,70,0,155,0,0,0,218,0,0,0,60,0,95,0,35,0,250,0,0,0,148,0,129,0,133,0,119,0,131,0,94,0,103,0,0,0,0,0,33,0,22,0,116,0,53,0,183,0,0,0,102,0,80,0,182,0,245,0,247,0,226,0,218,0,223,0,64,0,118,0,181,0,24,0,0,0,224,0,136,0,189,0,195,0,165,0,253,0,214,0,8,0,0,0,69,0,78,0,61,0,76,0,0,0,145,0,1,0,190,0,240,0,70,0,248,0,195,0,28,0,97,0,106,0,132,0,163,0,91,0,0,0,204,0,167,0,0,0,110,0,0,0,177,0,0,0,248,0,0,0,243,0,192,0,235,0,79,0,202,0,5,0,77,0,182,0,40,0,118,0,156,0,13,0,194,0,0,0,0,0,85,0,0,0,139,0,35,0,82,0,158,0,49,0,67,0,240,0,61,0,9,0,227,0,176,0,0,0,46,0,0,0,0,0,103,0,123,0,0,0,201,0,0,0,219,0,118,0,35,0,0,0,0,0,193,0,117,0,51,0,34,0,9,0,0,0,128,0,103,0,135,0,195,0,190,0,0,0,2,0,85,0,141,0,86,0,0,0,0,0,0,0,18,0,23,0,146,0,190,0,0,0,215,0,70,0,223,0,0,0,155,0,226,0,120,0,238,0,0,0,215,0,173,0,49,0,0,0,183,0,148,0,86,0,74,0,0,0,157,0,213,0,46,0,21,0,17,0,210,0,91,0,0,0,0,0,235,0,69,0,36,0,0,0,231,0,66,0,0,0,154,0,109,0,213,0,252,0,119,0,0,0,82,0,187,0,0,0,253,0,114,0,167,0,0,0,0,0,133,0,0,0,66,0,0,0,149,0,163,0,158,0,0,0,169,0,152,0,114,0,97,0,92,0,0,0,0,0,0,0,41,0,240,0,0,0,75,0,50,0,137,0,223,0,8,0,0,0,134,0,61,0,50,0,0,0,126,0,196,0,28,0,121,0,127,0,145,0,151,0,65,0,152,0,49,0,55,0,36,0,128,0,161,0,237,0,58,0,170,0,8,0,41,0,108,0,235,0,80,0,154,0,98,0,140,0,198,0,0,0,236,0,254,0,48,0,117,0,176,0,128,0,0,0,208,0,114,0,78,0,187,0,245,0,231,0,25,0,0,0,127,0,135,0,0,0,60,0,0,0,1,0,144,0,122,0,0,0,213,0,0,0,25,0,204,0,202,0,71,0,0,0,163,0,226,0,129,0,62,0,109,0,225,0,116,0,121,0,132,0,164,0,168,0,161,0,0,0,19,0,244,0,222,0,0,0,103,0,159,0,175,0,196,0,20,0,80,0,0,0,51,0,32,0,202,0,178,0,251,0,93,0,98,0,122,0,24,0,0,0,0,0,0,0,112,0,64,0,0,0,161,0,190,0,82,0,0,0,0,0,16,0,27,0,73,0,250,0,1,0,21,0,0,0,78,0,28,0,66,0,1,0,0,0,33,0,30,0,25,0,100,0,60,0,130,0,0,0,113,0,195,0,0,0,223,0,160,0,194,0,236,0,61,0,215,0,0,0,0,0,163,0,102,0,159,0,224,0,181,0,51,0,0,0,20,0,199,0,87,0,37,0,23,0,250,0,165,0,0,0,0,0,173,0,250,0,0,0,80,0,0,0,218,0,108,0,7,0,0,0,240,0,88,0,0,0,200,0,27,0,219,0,190,0,24,0,4,0,0,0,2,0,201,0,0,0,212,0,179,0,0,0,0,0,0,0,213,0,10,0,88,0,16,0,96,0,0,0,241,0,178,0,197,0,167,0,45,0,68,0,181,0,147,0,94,0,0,0,207,0,0,0,147,0,0,0,14,0,204,0,149,0,129,0,206,0,180,0,195,0,0,0,99,0,0,0,210,0,214,0,41,0,0,0,109,0,243,0,0,0,253,0,238,0,0,0,52,0,87,0,226,0,0,0,71,0,198,0,162,0,0,0,174,0,138,0,202,0,23,0,121,0,100,0,6,0,203,0,0,0,0,0,83,0,0,0,46,0,168,0,72,0,160,0,218,0,0,0,24,0,31,0,0,0,102,0,0,0,7,0,40,0,0,0,42,0,221,0,137,0,180,0,166,0,220,0,71,0,0,0,184,0,9,0,93,0,0,0,69,0,92,0,158,0,0,0,193,0,70,0,0,0,113,0,90,0,69,0,0,0,0,0,139,0,56,0,2,0,0,0,19,0,93,0,249,0,165,0,233,0,0,0,222,0,188,0,0,0,0,0,5,0,152,0,119,0,0,0,83,0,28,0,48,0,133,0,0,0,255,0,245,0,212,0,140,0,0,0,0,0,222,0,0,0,101,0,142,0,163,0,140,0,0,0,82,0,221,0,249,0,185,0,25,0,32,0,0,0,0,0,41,0,255,0,179,0,0,0,87,0,68,0,165,0,106,0,184,0,127,0,0,0,253,0,103,0,10,0,57,0,226,0,102,0,60,0,0,0,46,0,13,0,19,0,0,0,243,0,0,0,51,0,0,0,177,0,0,0,71,0,189,0,17,0,108,0,253,0,72,0,0,0,217,0,130,0,204,0,11,0,76,0,0,0,20,0,0,0,233,0,106,0,173,0,128,0,220,0,128,0,202,0,136,0,0,0,87,0,0,0,135,0,38,0,9,0,86,0,4,0,118,0,220,0,47,0,208,0,246,0,211,0,246,0,99,0,74,0,52,0,114,0,0,0,0,0,133,0,126,0,0,0,27,0,104,0,0,0,97,0,111,0,106,0);
signal scenario_full  : scenario_type := (40,31,40,30,94,31,143,31,143,30,98,31,98,30,98,29,247,31,95,31,10,31,10,30,70,31,155,31,155,30,218,31,218,30,60,31,95,31,35,31,250,31,250,30,148,31,129,31,133,31,119,31,131,31,94,31,103,31,103,30,103,29,33,31,22,31,116,31,53,31,183,31,183,30,102,31,80,31,182,31,245,31,247,31,226,31,218,31,223,31,64,31,118,31,181,31,24,31,24,30,224,31,136,31,189,31,195,31,165,31,253,31,214,31,8,31,8,30,69,31,78,31,61,31,76,31,76,30,145,31,1,31,190,31,240,31,70,31,248,31,195,31,28,31,97,31,106,31,132,31,163,31,91,31,91,30,204,31,167,31,167,30,110,31,110,30,177,31,177,30,248,31,248,30,243,31,192,31,235,31,79,31,202,31,5,31,77,31,182,31,40,31,118,31,156,31,13,31,194,31,194,30,194,29,85,31,85,30,139,31,35,31,82,31,158,31,49,31,67,31,240,31,61,31,9,31,227,31,176,31,176,30,46,31,46,30,46,29,103,31,123,31,123,30,201,31,201,30,219,31,118,31,35,31,35,30,35,29,193,31,117,31,51,31,34,31,9,31,9,30,128,31,103,31,135,31,195,31,190,31,190,30,2,31,85,31,141,31,86,31,86,30,86,29,86,28,18,31,23,31,146,31,190,31,190,30,215,31,70,31,223,31,223,30,155,31,226,31,120,31,238,31,238,30,215,31,173,31,49,31,49,30,183,31,148,31,86,31,74,31,74,30,157,31,213,31,46,31,21,31,17,31,210,31,91,31,91,30,91,29,235,31,69,31,36,31,36,30,231,31,66,31,66,30,154,31,109,31,213,31,252,31,119,31,119,30,82,31,187,31,187,30,253,31,114,31,167,31,167,30,167,29,133,31,133,30,66,31,66,30,149,31,163,31,158,31,158,30,169,31,152,31,114,31,97,31,92,31,92,30,92,29,92,28,41,31,240,31,240,30,75,31,50,31,137,31,223,31,8,31,8,30,134,31,61,31,50,31,50,30,126,31,196,31,28,31,121,31,127,31,145,31,151,31,65,31,152,31,49,31,55,31,36,31,128,31,161,31,237,31,58,31,170,31,8,31,41,31,108,31,235,31,80,31,154,31,98,31,140,31,198,31,198,30,236,31,254,31,48,31,117,31,176,31,128,31,128,30,208,31,114,31,78,31,187,31,245,31,231,31,25,31,25,30,127,31,135,31,135,30,60,31,60,30,1,31,144,31,122,31,122,30,213,31,213,30,25,31,204,31,202,31,71,31,71,30,163,31,226,31,129,31,62,31,109,31,225,31,116,31,121,31,132,31,164,31,168,31,161,31,161,30,19,31,244,31,222,31,222,30,103,31,159,31,175,31,196,31,20,31,80,31,80,30,51,31,32,31,202,31,178,31,251,31,93,31,98,31,122,31,24,31,24,30,24,29,24,28,112,31,64,31,64,30,161,31,190,31,82,31,82,30,82,29,16,31,27,31,73,31,250,31,1,31,21,31,21,30,78,31,28,31,66,31,1,31,1,30,33,31,30,31,25,31,100,31,60,31,130,31,130,30,113,31,195,31,195,30,223,31,160,31,194,31,236,31,61,31,215,31,215,30,215,29,163,31,102,31,159,31,224,31,181,31,51,31,51,30,20,31,199,31,87,31,37,31,23,31,250,31,165,31,165,30,165,29,173,31,250,31,250,30,80,31,80,30,218,31,108,31,7,31,7,30,240,31,88,31,88,30,200,31,27,31,219,31,190,31,24,31,4,31,4,30,2,31,201,31,201,30,212,31,179,31,179,30,179,29,179,28,213,31,10,31,88,31,16,31,96,31,96,30,241,31,178,31,197,31,167,31,45,31,68,31,181,31,147,31,94,31,94,30,207,31,207,30,147,31,147,30,14,31,204,31,149,31,129,31,206,31,180,31,195,31,195,30,99,31,99,30,210,31,214,31,41,31,41,30,109,31,243,31,243,30,253,31,238,31,238,30,52,31,87,31,226,31,226,30,71,31,198,31,162,31,162,30,174,31,138,31,202,31,23,31,121,31,100,31,6,31,203,31,203,30,203,29,83,31,83,30,46,31,168,31,72,31,160,31,218,31,218,30,24,31,31,31,31,30,102,31,102,30,7,31,40,31,40,30,42,31,221,31,137,31,180,31,166,31,220,31,71,31,71,30,184,31,9,31,93,31,93,30,69,31,92,31,158,31,158,30,193,31,70,31,70,30,113,31,90,31,69,31,69,30,69,29,139,31,56,31,2,31,2,30,19,31,93,31,249,31,165,31,233,31,233,30,222,31,188,31,188,30,188,29,5,31,152,31,119,31,119,30,83,31,28,31,48,31,133,31,133,30,255,31,245,31,212,31,140,31,140,30,140,29,222,31,222,30,101,31,142,31,163,31,140,31,140,30,82,31,221,31,249,31,185,31,25,31,32,31,32,30,32,29,41,31,255,31,179,31,179,30,87,31,68,31,165,31,106,31,184,31,127,31,127,30,253,31,103,31,10,31,57,31,226,31,102,31,60,31,60,30,46,31,13,31,19,31,19,30,243,31,243,30,51,31,51,30,177,31,177,30,71,31,189,31,17,31,108,31,253,31,72,31,72,30,217,31,130,31,204,31,11,31,76,31,76,30,20,31,20,30,233,31,106,31,173,31,128,31,220,31,128,31,202,31,136,31,136,30,87,31,87,30,135,31,38,31,9,31,86,31,4,31,118,31,220,31,47,31,208,31,246,31,211,31,246,31,99,31,74,31,52,31,114,31,114,30,114,29,133,31,126,31,126,30,27,31,104,31,104,30,97,31,111,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
