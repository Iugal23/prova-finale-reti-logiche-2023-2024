-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_547 is
end project_tb_547;

architecture project_tb_arch_547 of project_tb_547 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 497;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (57,0,89,0,120,0,75,0,69,0,170,0,171,0,103,0,95,0,0,0,114,0,190,0,0,0,0,0,239,0,140,0,0,0,228,0,156,0,31,0,22,0,87,0,0,0,106,0,111,0,0,0,182,0,129,0,133,0,76,0,238,0,195,0,152,0,192,0,98,0,187,0,176,0,0,0,58,0,0,0,0,0,0,0,204,0,0,0,0,0,242,0,68,0,44,0,213,0,161,0,228,0,27,0,187,0,185,0,197,0,0,0,4,0,0,0,120,0,135,0,80,0,79,0,61,0,92,0,250,0,0,0,52,0,0,0,157,0,138,0,125,0,0,0,79,0,34,0,0,0,19,0,194,0,179,0,135,0,60,0,0,0,0,0,37,0,20,0,221,0,169,0,152,0,97,0,47,0,150,0,228,0,145,0,166,0,74,0,67,0,8,0,105,0,161,0,0,0,0,0,84,0,103,0,219,0,130,0,187,0,122,0,173,0,248,0,67,0,66,0,71,0,48,0,184,0,57,0,129,0,199,0,13,0,84,0,0,0,180,0,60,0,167,0,64,0,193,0,217,0,0,0,182,0,180,0,197,0,0,0,0,0,0,0,7,0,227,0,39,0,122,0,50,0,80,0,69,0,244,0,0,0,81,0,197,0,141,0,52,0,74,0,214,0,0,0,0,0,47,0,10,0,87,0,146,0,42,0,5,0,133,0,104,0,18,0,1,0,0,0,31,0,134,0,245,0,251,0,0,0,65,0,0,0,159,0,13,0,212,0,73,0,106,0,207,0,3,0,105,0,65,0,157,0,70,0,220,0,0,0,224,0,37,0,31,0,176,0,0,0,50,0,201,0,31,0,232,0,40,0,0,0,124,0,0,0,73,0,0,0,238,0,0,0,0,0,27,0,131,0,60,0,41,0,224,0,102,0,210,0,0,0,104,0,67,0,89,0,247,0,122,0,238,0,2,0,67,0,198,0,208,0,140,0,97,0,74,0,0,0,0,0,121,0,0,0,232,0,175,0,11,0,24,0,157,0,0,0,1,0,165,0,125,0,18,0,164,0,70,0,19,0,0,0,0,0,0,0,120,0,69,0,142,0,0,0,186,0,153,0,155,0,203,0,233,0,0,0,233,0,125,0,0,0,0,0,142,0,240,0,0,0,155,0,0,0,0,0,205,0,220,0,0,0,234,0,91,0,43,0,74,0,162,0,200,0,132,0,211,0,11,0,174,0,155,0,208,0,183,0,233,0,119,0,79,0,11,0,248,0,57,0,175,0,186,0,123,0,6,0,103,0,43,0,194,0,217,0,190,0,22,0,188,0,234,0,91,0,161,0,155,0,149,0,64,0,186,0,29,0,216,0,130,0,75,0,95,0,198,0,106,0,214,0,7,0,136,0,30,0,22,0,64,0,0,0,82,0,178,0,210,0,144,0,133,0,95,0,21,0,36,0,116,0,214,0,234,0,142,0,221,0,226,0,154,0,74,0,150,0,0,0,0,0,0,0,0,0,0,0,60,0,25,0,190,0,90,0,98,0,0,0,17,0,0,0,74,0,193,0,203,0,188,0,11,0,0,0,0,0,222,0,194,0,0,0,213,0,59,0,0,0,0,0,111,0,218,0,100,0,0,0,29,0,0,0,0,0,23,0,0,0,0,0,33,0,52,0,0,0,185,0,177,0,17,0,38,0,78,0,0,0,179,0,200,0,40,0,160,0,73,0,62,0,29,0,50,0,166,0,36,0,89,0,203,0,0,0,134,0,37,0,205,0,84,0,0,0,7,0,0,0,244,0,1,0,196,0,205,0,175,0,77,0,0,0,15,0,54,0,61,0,154,0,5,0,0,0,109,0,195,0,149,0,108,0,51,0,14,0,236,0,235,0,30,0,0,0,85,0,171,0,171,0,2,0,131,0,0,0,24,0,0,0,0,0,204,0,44,0,14,0,178,0,170,0,252,0,0,0,48,0,136,0,0,0,150,0,252,0,211,0,184,0,103,0,1,0,77,0,255,0,46,0,19,0,0,0,62,0,176,0,238,0,15,0,55,0,73,0,165,0,112,0,216,0,195,0,184,0,18,0,247,0,90,0,0,0,35,0,181,0,211,0,131,0,224,0,188,0,223,0,199,0,187,0,235,0,129,0,161,0,143,0,220,0,63,0,214,0,169,0,218,0,0,0,172,0,55,0,119,0,122,0,192,0,129,0,124,0,149,0,0,0,0,0,21,0,0,0,0,0,64,0);
signal scenario_full  : scenario_type := (57,31,89,31,120,31,75,31,69,31,170,31,171,31,103,31,95,31,95,30,114,31,190,31,190,30,190,29,239,31,140,31,140,30,228,31,156,31,31,31,22,31,87,31,87,30,106,31,111,31,111,30,182,31,129,31,133,31,76,31,238,31,195,31,152,31,192,31,98,31,187,31,176,31,176,30,58,31,58,30,58,29,58,28,204,31,204,30,204,29,242,31,68,31,44,31,213,31,161,31,228,31,27,31,187,31,185,31,197,31,197,30,4,31,4,30,120,31,135,31,80,31,79,31,61,31,92,31,250,31,250,30,52,31,52,30,157,31,138,31,125,31,125,30,79,31,34,31,34,30,19,31,194,31,179,31,135,31,60,31,60,30,60,29,37,31,20,31,221,31,169,31,152,31,97,31,47,31,150,31,228,31,145,31,166,31,74,31,67,31,8,31,105,31,161,31,161,30,161,29,84,31,103,31,219,31,130,31,187,31,122,31,173,31,248,31,67,31,66,31,71,31,48,31,184,31,57,31,129,31,199,31,13,31,84,31,84,30,180,31,60,31,167,31,64,31,193,31,217,31,217,30,182,31,180,31,197,31,197,30,197,29,197,28,7,31,227,31,39,31,122,31,50,31,80,31,69,31,244,31,244,30,81,31,197,31,141,31,52,31,74,31,214,31,214,30,214,29,47,31,10,31,87,31,146,31,42,31,5,31,133,31,104,31,18,31,1,31,1,30,31,31,134,31,245,31,251,31,251,30,65,31,65,30,159,31,13,31,212,31,73,31,106,31,207,31,3,31,105,31,65,31,157,31,70,31,220,31,220,30,224,31,37,31,31,31,176,31,176,30,50,31,201,31,31,31,232,31,40,31,40,30,124,31,124,30,73,31,73,30,238,31,238,30,238,29,27,31,131,31,60,31,41,31,224,31,102,31,210,31,210,30,104,31,67,31,89,31,247,31,122,31,238,31,2,31,67,31,198,31,208,31,140,31,97,31,74,31,74,30,74,29,121,31,121,30,232,31,175,31,11,31,24,31,157,31,157,30,1,31,165,31,125,31,18,31,164,31,70,31,19,31,19,30,19,29,19,28,120,31,69,31,142,31,142,30,186,31,153,31,155,31,203,31,233,31,233,30,233,31,125,31,125,30,125,29,142,31,240,31,240,30,155,31,155,30,155,29,205,31,220,31,220,30,234,31,91,31,43,31,74,31,162,31,200,31,132,31,211,31,11,31,174,31,155,31,208,31,183,31,233,31,119,31,79,31,11,31,248,31,57,31,175,31,186,31,123,31,6,31,103,31,43,31,194,31,217,31,190,31,22,31,188,31,234,31,91,31,161,31,155,31,149,31,64,31,186,31,29,31,216,31,130,31,75,31,95,31,198,31,106,31,214,31,7,31,136,31,30,31,22,31,64,31,64,30,82,31,178,31,210,31,144,31,133,31,95,31,21,31,36,31,116,31,214,31,234,31,142,31,221,31,226,31,154,31,74,31,150,31,150,30,150,29,150,28,150,27,150,26,60,31,25,31,190,31,90,31,98,31,98,30,17,31,17,30,74,31,193,31,203,31,188,31,11,31,11,30,11,29,222,31,194,31,194,30,213,31,59,31,59,30,59,29,111,31,218,31,100,31,100,30,29,31,29,30,29,29,23,31,23,30,23,29,33,31,52,31,52,30,185,31,177,31,17,31,38,31,78,31,78,30,179,31,200,31,40,31,160,31,73,31,62,31,29,31,50,31,166,31,36,31,89,31,203,31,203,30,134,31,37,31,205,31,84,31,84,30,7,31,7,30,244,31,1,31,196,31,205,31,175,31,77,31,77,30,15,31,54,31,61,31,154,31,5,31,5,30,109,31,195,31,149,31,108,31,51,31,14,31,236,31,235,31,30,31,30,30,85,31,171,31,171,31,2,31,131,31,131,30,24,31,24,30,24,29,204,31,44,31,14,31,178,31,170,31,252,31,252,30,48,31,136,31,136,30,150,31,252,31,211,31,184,31,103,31,1,31,77,31,255,31,46,31,19,31,19,30,62,31,176,31,238,31,15,31,55,31,73,31,165,31,112,31,216,31,195,31,184,31,18,31,247,31,90,31,90,30,35,31,181,31,211,31,131,31,224,31,188,31,223,31,199,31,187,31,235,31,129,31,161,31,143,31,220,31,63,31,214,31,169,31,218,31,218,30,172,31,55,31,119,31,122,31,192,31,129,31,124,31,149,31,149,30,149,29,21,31,21,30,21,29,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
