-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 225;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (207,0,0,0,35,0,28,0,197,0,247,0,235,0,16,0,174,0,135,0,0,0,0,0,238,0,107,0,0,0,85,0,248,0,42,0,178,0,31,0,231,0,0,0,32,0,229,0,56,0,58,0,89,0,71,0,0,0,136,0,0,0,167,0,0,0,174,0,43,0,133,0,0,0,0,0,40,0,205,0,88,0,127,0,81,0,0,0,154,0,51,0,121,0,199,0,187,0,0,0,252,0,233,0,178,0,148,0,65,0,195,0,0,0,66,0,189,0,60,0,0,0,16,0,186,0,33,0,99,0,0,0,179,0,17,0,0,0,5,0,187,0,0,0,96,0,0,0,21,0,179,0,151,0,0,0,93,0,0,0,112,0,0,0,0,0,224,0,229,0,184,0,197,0,171,0,238,0,58,0,112,0,176,0,75,0,0,0,221,0,156,0,27,0,46,0,0,0,243,0,219,0,34,0,158,0,71,0,0,0,253,0,0,0,84,0,0,0,64,0,43,0,88,0,235,0,232,0,154,0,121,0,48,0,0,0,76,0,159,0,233,0,15,0,0,0,157,0,191,0,0,0,0,0,9,0,0,0,138,0,0,0,253,0,163,0,28,0,198,0,100,0,249,0,200,0,44,0,247,0,14,0,209,0,73,0,148,0,93,0,57,0,69,0,157,0,32,0,0,0,226,0,212,0,137,0,0,0,233,0,252,0,27,0,0,0,243,0,12,0,144,0,183,0,227,0,7,0,67,0,152,0,49,0,25,0,160,0,192,0,0,0,77,0,0,0,212,0,0,0,226,0,0,0,174,0,107,0,176,0,53,0,181,0,247,0,0,0,95,0,41,0,92,0,176,0,70,0,12,0,235,0,62,0,0,0,99,0,0,0,90,0,118,0,0,0,0,0,35,0,0,0,0,0,0,0,33,0,190,0,104,0,218,0,0,0,177,0,0,0,0,0,210,0,94,0,146,0,9,0,37,0,0,0,5,0,120,0,243,0,177,0,221,0,114,0,0,0,73,0);
signal scenario_full  : scenario_type := (207,31,207,30,35,31,28,31,197,31,247,31,235,31,16,31,174,31,135,31,135,30,135,29,238,31,107,31,107,30,85,31,248,31,42,31,178,31,31,31,231,31,231,30,32,31,229,31,56,31,58,31,89,31,71,31,71,30,136,31,136,30,167,31,167,30,174,31,43,31,133,31,133,30,133,29,40,31,205,31,88,31,127,31,81,31,81,30,154,31,51,31,121,31,199,31,187,31,187,30,252,31,233,31,178,31,148,31,65,31,195,31,195,30,66,31,189,31,60,31,60,30,16,31,186,31,33,31,99,31,99,30,179,31,17,31,17,30,5,31,187,31,187,30,96,31,96,30,21,31,179,31,151,31,151,30,93,31,93,30,112,31,112,30,112,29,224,31,229,31,184,31,197,31,171,31,238,31,58,31,112,31,176,31,75,31,75,30,221,31,156,31,27,31,46,31,46,30,243,31,219,31,34,31,158,31,71,31,71,30,253,31,253,30,84,31,84,30,64,31,43,31,88,31,235,31,232,31,154,31,121,31,48,31,48,30,76,31,159,31,233,31,15,31,15,30,157,31,191,31,191,30,191,29,9,31,9,30,138,31,138,30,253,31,163,31,28,31,198,31,100,31,249,31,200,31,44,31,247,31,14,31,209,31,73,31,148,31,93,31,57,31,69,31,157,31,32,31,32,30,226,31,212,31,137,31,137,30,233,31,252,31,27,31,27,30,243,31,12,31,144,31,183,31,227,31,7,31,67,31,152,31,49,31,25,31,160,31,192,31,192,30,77,31,77,30,212,31,212,30,226,31,226,30,174,31,107,31,176,31,53,31,181,31,247,31,247,30,95,31,41,31,92,31,176,31,70,31,12,31,235,31,62,31,62,30,99,31,99,30,90,31,118,31,118,30,118,29,35,31,35,30,35,29,35,28,33,31,190,31,104,31,218,31,218,30,177,31,177,30,177,29,210,31,94,31,146,31,9,31,37,31,37,30,5,31,120,31,243,31,177,31,221,31,114,31,114,30,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
