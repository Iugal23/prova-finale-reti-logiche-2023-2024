-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_767 is
end project_tb_767;

architecture project_tb_arch_767 of project_tb_767 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 309;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,214,0,205,0,23,0,159,0,127,0,230,0,182,0,53,0,0,0,161,0,0,0,81,0,49,0,170,0,44,0,177,0,184,0,0,0,186,0,195,0,227,0,64,0,198,0,0,0,196,0,162,0,249,0,0,0,255,0,39,0,0,0,241,0,221,0,123,0,67,0,0,0,0,0,63,0,177,0,89,0,241,0,21,0,142,0,234,0,71,0,101,0,64,0,0,0,0,0,133,0,159,0,52,0,123,0,180,0,242,0,201,0,0,0,0,0,0,0,212,0,156,0,134,0,121,0,63,0,134,0,201,0,0,0,239,0,134,0,70,0,0,0,52,0,12,0,36,0,197,0,51,0,0,0,4,0,104,0,199,0,132,0,61,0,115,0,151,0,24,0,214,0,0,0,199,0,0,0,206,0,221,0,167,0,36,0,166,0,73,0,0,0,54,0,90,0,38,0,96,0,123,0,78,0,0,0,20,0,161,0,129,0,0,0,4,0,1,0,12,0,29,0,55,0,0,0,0,0,155,0,100,0,114,0,0,0,63,0,168,0,188,0,32,0,9,0,177,0,0,0,169,0,99,0,171,0,59,0,200,0,2,0,218,0,0,0,32,0,229,0,0,0,192,0,0,0,16,0,207,0,161,0,0,0,131,0,22,0,232,0,78,0,0,0,109,0,0,0,78,0,0,0,139,0,179,0,32,0,5,0,248,0,56,0,0,0,0,0,0,0,182,0,6,0,63,0,94,0,0,0,167,0,9,0,0,0,0,0,0,0,0,0,142,0,205,0,11,0,14,0,218,0,71,0,0,0,75,0,111,0,77,0,71,0,210,0,131,0,0,0,54,0,28,0,60,0,149,0,15,0,214,0,73,0,191,0,250,0,0,0,8,0,139,0,69,0,135,0,167,0,167,0,158,0,0,0,185,0,143,0,166,0,54,0,210,0,167,0,6,0,0,0,27,0,124,0,63,0,50,0,139,0,0,0,0,0,103,0,103,0,232,0,218,0,103,0,219,0,63,0,52,0,95,0,80,0,187,0,241,0,92,0,0,0,107,0,247,0,0,0,229,0,79,0,141,0,0,0,0,0,137,0,179,0,0,0,83,0,84,0,191,0,217,0,195,0,34,0,0,0,131,0,134,0,165,0,0,0,201,0,222,0,47,0,0,0,243,0,233,0,0,0,40,0,252,0,187,0,214,0,0,0,139,0,93,0,126,0,170,0,37,0,152,0,0,0,27,0,220,0,56,0,237,0,60,0,0,0,19,0,0,0,139,0,185,0,199,0,95,0,155,0,208,0,43,0,17,0,173,0,0,0,243,0,0,0,137,0,0,0,10,0,25,0,233,0,43,0,154,0,211,0,220,0,101,0,130,0,234,0,0,0,0,0,233,0);
signal scenario_full  : scenario_type := (9,31,214,31,205,31,23,31,159,31,127,31,230,31,182,31,53,31,53,30,161,31,161,30,81,31,49,31,170,31,44,31,177,31,184,31,184,30,186,31,195,31,227,31,64,31,198,31,198,30,196,31,162,31,249,31,249,30,255,31,39,31,39,30,241,31,221,31,123,31,67,31,67,30,67,29,63,31,177,31,89,31,241,31,21,31,142,31,234,31,71,31,101,31,64,31,64,30,64,29,133,31,159,31,52,31,123,31,180,31,242,31,201,31,201,30,201,29,201,28,212,31,156,31,134,31,121,31,63,31,134,31,201,31,201,30,239,31,134,31,70,31,70,30,52,31,12,31,36,31,197,31,51,31,51,30,4,31,104,31,199,31,132,31,61,31,115,31,151,31,24,31,214,31,214,30,199,31,199,30,206,31,221,31,167,31,36,31,166,31,73,31,73,30,54,31,90,31,38,31,96,31,123,31,78,31,78,30,20,31,161,31,129,31,129,30,4,31,1,31,12,31,29,31,55,31,55,30,55,29,155,31,100,31,114,31,114,30,63,31,168,31,188,31,32,31,9,31,177,31,177,30,169,31,99,31,171,31,59,31,200,31,2,31,218,31,218,30,32,31,229,31,229,30,192,31,192,30,16,31,207,31,161,31,161,30,131,31,22,31,232,31,78,31,78,30,109,31,109,30,78,31,78,30,139,31,179,31,32,31,5,31,248,31,56,31,56,30,56,29,56,28,182,31,6,31,63,31,94,31,94,30,167,31,9,31,9,30,9,29,9,28,9,27,142,31,205,31,11,31,14,31,218,31,71,31,71,30,75,31,111,31,77,31,71,31,210,31,131,31,131,30,54,31,28,31,60,31,149,31,15,31,214,31,73,31,191,31,250,31,250,30,8,31,139,31,69,31,135,31,167,31,167,31,158,31,158,30,185,31,143,31,166,31,54,31,210,31,167,31,6,31,6,30,27,31,124,31,63,31,50,31,139,31,139,30,139,29,103,31,103,31,232,31,218,31,103,31,219,31,63,31,52,31,95,31,80,31,187,31,241,31,92,31,92,30,107,31,247,31,247,30,229,31,79,31,141,31,141,30,141,29,137,31,179,31,179,30,83,31,84,31,191,31,217,31,195,31,34,31,34,30,131,31,134,31,165,31,165,30,201,31,222,31,47,31,47,30,243,31,233,31,233,30,40,31,252,31,187,31,214,31,214,30,139,31,93,31,126,31,170,31,37,31,152,31,152,30,27,31,220,31,56,31,237,31,60,31,60,30,19,31,19,30,139,31,185,31,199,31,95,31,155,31,208,31,43,31,17,31,173,31,173,30,243,31,243,30,137,31,137,30,10,31,25,31,233,31,43,31,154,31,211,31,220,31,101,31,130,31,234,31,234,30,234,29,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
