-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 688;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (143,0,45,0,110,0,0,0,0,0,0,0,120,0,0,0,114,0,0,0,51,0,241,0,252,0,125,0,211,0,150,0,3,0,0,0,0,0,156,0,122,0,53,0,125,0,231,0,142,0,0,0,81,0,209,0,242,0,0,0,223,0,136,0,141,0,126,0,150,0,0,0,3,0,0,0,220,0,1,0,38,0,126,0,121,0,177,0,228,0,21,0,211,0,50,0,0,0,7,0,111,0,181,0,54,0,71,0,0,0,0,0,248,0,175,0,203,0,165,0,172,0,188,0,35,0,39,0,45,0,116,0,83,0,50,0,0,0,184,0,101,0,0,0,51,0,71,0,205,0,180,0,10,0,89,0,134,0,202,0,139,0,205,0,152,0,200,0,92,0,229,0,176,0,22,0,202,0,0,0,68,0,123,0,229,0,0,0,205,0,0,0,0,0,14,0,0,0,197,0,52,0,247,0,172,0,18,0,85,0,30,0,24,0,17,0,0,0,14,0,102,0,254,0,0,0,85,0,170,0,19,0,239,0,0,0,161,0,0,0,218,0,21,0,0,0,0,0,117,0,27,0,0,0,202,0,28,0,53,0,0,0,231,0,115,0,0,0,199,0,0,0,0,0,29,0,245,0,82,0,204,0,0,0,0,0,155,0,207,0,0,0,0,0,28,0,215,0,86,0,163,0,140,0,135,0,84,0,60,0,0,0,0,0,216,0,0,0,99,0,248,0,115,0,198,0,191,0,106,0,121,0,175,0,119,0,187,0,220,0,96,0,220,0,225,0,216,0,71,0,20,0,233,0,209,0,4,0,118,0,0,0,70,0,88,0,48,0,0,0,237,0,72,0,124,0,175,0,0,0,0,0,117,0,35,0,175,0,42,0,129,0,115,0,49,0,251,0,0,0,93,0,238,0,174,0,87,0,58,0,43,0,75,0,223,0,147,0,110,0,0,0,89,0,225,0,218,0,15,0,211,0,0,0,18,0,0,0,130,0,232,0,105,0,49,0,67,0,113,0,123,0,0,0,64,0,51,0,154,0,2,0,171,0,89,0,117,0,127,0,0,0,223,0,89,0,83,0,253,0,29,0,106,0,16,0,7,0,40,0,103,0,203,0,11,0,7,0,0,0,158,0,75,0,27,0,211,0,51,0,57,0,171,0,46,0,128,0,2,0,60,0,0,0,9,0,138,0,82,0,136,0,154,0,244,0,0,0,15,0,196,0,66,0,89,0,230,0,33,0,230,0,113,0,0,0,0,0,164,0,189,0,135,0,84,0,107,0,19,0,86,0,117,0,0,0,178,0,0,0,120,0,243,0,8,0,0,0,103,0,115,0,87,0,222,0,0,0,5,0,80,0,141,0,89,0,216,0,203,0,47,0,187,0,36,0,99,0,54,0,235,0,30,0,158,0,10,0,99,0,241,0,28,0,252,0,0,0,48,0,252,0,23,0,34,0,14,0,236,0,0,0,226,0,105,0,65,0,27,0,244,0,0,0,40,0,44,0,0,0,186,0,0,0,51,0,0,0,184,0,56,0,98,0,0,0,145,0,69,0,0,0,128,0,185,0,254,0,251,0,94,0,0,0,61,0,110,0,58,0,169,0,108,0,127,0,76,0,244,0,88,0,0,0,50,0,73,0,216,0,62,0,97,0,16,0,222,0,132,0,81,0,116,0,246,0,44,0,142,0,64,0,200,0,74,0,43,0,0,0,238,0,41,0,182,0,167,0,137,0,243,0,0,0,227,0,206,0,0,0,126,0,167,0,152,0,226,0,41,0,39,0,114,0,154,0,52,0,218,0,168,0,0,0,167,0,0,0,52,0,112,0,200,0,202,0,56,0,0,0,137,0,79,0,190,0,93,0,48,0,99,0,125,0,161,0,63,0,145,0,220,0,227,0,234,0,109,0,8,0,0,0,32,0,0,0,189,0,0,0,178,0,0,0,208,0,0,0,138,0,0,0,0,0,6,0,14,0,213,0,0,0,245,0,60,0,0,0,254,0,74,0,16,0,84,0,0,0,189,0,115,0,0,0,175,0,103,0,31,0,60,0,152,0,0,0,157,0,214,0,42,0,76,0,163,0,166,0,165,0,0,0,39,0,243,0,79,0,0,0,34,0,159,0,131,0,189,0,37,0,107,0,159,0,68,0,39,0,221,0,94,0,53,0,230,0,0,0,221,0,123,0,1,0,38,0,81,0,166,0,106,0,205,0,0,0,0,0,155,0,0,0,30,0,53,0,48,0,57,0,82,0,36,0,202,0,119,0,136,0,10,0,0,0,133,0,246,0,200,0,10,0,244,0,0,0,180,0,156,0,2,0,217,0,72,0,206,0,196,0,113,0,0,0,165,0,138,0,7,0,125,0,95,0,141,0,224,0,252,0,130,0,19,0,0,0,0,0,0,0,112,0,0,0,195,0,242,0,196,0,213,0,215,0,216,0,164,0,105,0,34,0,195,0,141,0,18,0,103,0,0,0,19,0,90,0,101,0,136,0,188,0,0,0,202,0,136,0,207,0,0,0,0,0,0,0,35,0,101,0,194,0,151,0,167,0,157,0,0,0,196,0,142,0,148,0,0,0,128,0,0,0,9,0,0,0,112,0,205,0,0,0,184,0,253,0,121,0,238,0,0,0,29,0,0,0,60,0,191,0,0,0,77,0,0,0,69,0,178,0,176,0,212,0,0,0,0,0,5,0,222,0,0,0,0,0,197,0,31,0,0,0,0,0,108,0,130,0,90,0,129,0,159,0,76,0,0,0,50,0,5,0,0,0,252,0,0,0,0,0,213,0,121,0,13,0,51,0,118,0,204,0,219,0,0,0,40,0,0,0,49,0,5,0,150,0,147,0,172,0,107,0,188,0,60,0,0,0,0,0,0,0,189,0,0,0,80,0,227,0,27,0,140,0,134,0,0,0,0,0,0,0,0,0,193,0,0,0,246,0,51,0,224,0,6,0,26,0,0,0,38,0,241,0,0,0,199,0,129,0,245,0,105,0,129,0,177,0,197,0,201,0,0,0,188,0,71,0,0,0,0,0,244,0,10,0,52,0,238,0,15,0,8,0,228,0,124,0,79,0,112,0,197,0,8,0);
signal scenario_full  : scenario_type := (143,31,45,31,110,31,110,30,110,29,110,28,120,31,120,30,114,31,114,30,51,31,241,31,252,31,125,31,211,31,150,31,3,31,3,30,3,29,156,31,122,31,53,31,125,31,231,31,142,31,142,30,81,31,209,31,242,31,242,30,223,31,136,31,141,31,126,31,150,31,150,30,3,31,3,30,220,31,1,31,38,31,126,31,121,31,177,31,228,31,21,31,211,31,50,31,50,30,7,31,111,31,181,31,54,31,71,31,71,30,71,29,248,31,175,31,203,31,165,31,172,31,188,31,35,31,39,31,45,31,116,31,83,31,50,31,50,30,184,31,101,31,101,30,51,31,71,31,205,31,180,31,10,31,89,31,134,31,202,31,139,31,205,31,152,31,200,31,92,31,229,31,176,31,22,31,202,31,202,30,68,31,123,31,229,31,229,30,205,31,205,30,205,29,14,31,14,30,197,31,52,31,247,31,172,31,18,31,85,31,30,31,24,31,17,31,17,30,14,31,102,31,254,31,254,30,85,31,170,31,19,31,239,31,239,30,161,31,161,30,218,31,21,31,21,30,21,29,117,31,27,31,27,30,202,31,28,31,53,31,53,30,231,31,115,31,115,30,199,31,199,30,199,29,29,31,245,31,82,31,204,31,204,30,204,29,155,31,207,31,207,30,207,29,28,31,215,31,86,31,163,31,140,31,135,31,84,31,60,31,60,30,60,29,216,31,216,30,99,31,248,31,115,31,198,31,191,31,106,31,121,31,175,31,119,31,187,31,220,31,96,31,220,31,225,31,216,31,71,31,20,31,233,31,209,31,4,31,118,31,118,30,70,31,88,31,48,31,48,30,237,31,72,31,124,31,175,31,175,30,175,29,117,31,35,31,175,31,42,31,129,31,115,31,49,31,251,31,251,30,93,31,238,31,174,31,87,31,58,31,43,31,75,31,223,31,147,31,110,31,110,30,89,31,225,31,218,31,15,31,211,31,211,30,18,31,18,30,130,31,232,31,105,31,49,31,67,31,113,31,123,31,123,30,64,31,51,31,154,31,2,31,171,31,89,31,117,31,127,31,127,30,223,31,89,31,83,31,253,31,29,31,106,31,16,31,7,31,40,31,103,31,203,31,11,31,7,31,7,30,158,31,75,31,27,31,211,31,51,31,57,31,171,31,46,31,128,31,2,31,60,31,60,30,9,31,138,31,82,31,136,31,154,31,244,31,244,30,15,31,196,31,66,31,89,31,230,31,33,31,230,31,113,31,113,30,113,29,164,31,189,31,135,31,84,31,107,31,19,31,86,31,117,31,117,30,178,31,178,30,120,31,243,31,8,31,8,30,103,31,115,31,87,31,222,31,222,30,5,31,80,31,141,31,89,31,216,31,203,31,47,31,187,31,36,31,99,31,54,31,235,31,30,31,158,31,10,31,99,31,241,31,28,31,252,31,252,30,48,31,252,31,23,31,34,31,14,31,236,31,236,30,226,31,105,31,65,31,27,31,244,31,244,30,40,31,44,31,44,30,186,31,186,30,51,31,51,30,184,31,56,31,98,31,98,30,145,31,69,31,69,30,128,31,185,31,254,31,251,31,94,31,94,30,61,31,110,31,58,31,169,31,108,31,127,31,76,31,244,31,88,31,88,30,50,31,73,31,216,31,62,31,97,31,16,31,222,31,132,31,81,31,116,31,246,31,44,31,142,31,64,31,200,31,74,31,43,31,43,30,238,31,41,31,182,31,167,31,137,31,243,31,243,30,227,31,206,31,206,30,126,31,167,31,152,31,226,31,41,31,39,31,114,31,154,31,52,31,218,31,168,31,168,30,167,31,167,30,52,31,112,31,200,31,202,31,56,31,56,30,137,31,79,31,190,31,93,31,48,31,99,31,125,31,161,31,63,31,145,31,220,31,227,31,234,31,109,31,8,31,8,30,32,31,32,30,189,31,189,30,178,31,178,30,208,31,208,30,138,31,138,30,138,29,6,31,14,31,213,31,213,30,245,31,60,31,60,30,254,31,74,31,16,31,84,31,84,30,189,31,115,31,115,30,175,31,103,31,31,31,60,31,152,31,152,30,157,31,214,31,42,31,76,31,163,31,166,31,165,31,165,30,39,31,243,31,79,31,79,30,34,31,159,31,131,31,189,31,37,31,107,31,159,31,68,31,39,31,221,31,94,31,53,31,230,31,230,30,221,31,123,31,1,31,38,31,81,31,166,31,106,31,205,31,205,30,205,29,155,31,155,30,30,31,53,31,48,31,57,31,82,31,36,31,202,31,119,31,136,31,10,31,10,30,133,31,246,31,200,31,10,31,244,31,244,30,180,31,156,31,2,31,217,31,72,31,206,31,196,31,113,31,113,30,165,31,138,31,7,31,125,31,95,31,141,31,224,31,252,31,130,31,19,31,19,30,19,29,19,28,112,31,112,30,195,31,242,31,196,31,213,31,215,31,216,31,164,31,105,31,34,31,195,31,141,31,18,31,103,31,103,30,19,31,90,31,101,31,136,31,188,31,188,30,202,31,136,31,207,31,207,30,207,29,207,28,35,31,101,31,194,31,151,31,167,31,157,31,157,30,196,31,142,31,148,31,148,30,128,31,128,30,9,31,9,30,112,31,205,31,205,30,184,31,253,31,121,31,238,31,238,30,29,31,29,30,60,31,191,31,191,30,77,31,77,30,69,31,178,31,176,31,212,31,212,30,212,29,5,31,222,31,222,30,222,29,197,31,31,31,31,30,31,29,108,31,130,31,90,31,129,31,159,31,76,31,76,30,50,31,5,31,5,30,252,31,252,30,252,29,213,31,121,31,13,31,51,31,118,31,204,31,219,31,219,30,40,31,40,30,49,31,5,31,150,31,147,31,172,31,107,31,188,31,60,31,60,30,60,29,60,28,189,31,189,30,80,31,227,31,27,31,140,31,134,31,134,30,134,29,134,28,134,27,193,31,193,30,246,31,51,31,224,31,6,31,26,31,26,30,38,31,241,31,241,30,199,31,129,31,245,31,105,31,129,31,177,31,197,31,201,31,201,30,188,31,71,31,71,30,71,29,244,31,10,31,52,31,238,31,15,31,8,31,228,31,124,31,79,31,112,31,197,31,8,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
