-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1021;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,31,0,110,0,99,0,0,0,0,0,98,0,221,0,37,0,0,0,0,0,107,0,121,0,90,0,69,0,140,0,10,0,65,0,63,0,0,0,160,0,41,0,0,0,164,0,97,0,15,0,181,0,209,0,141,0,186,0,47,0,71,0,173,0,205,0,125,0,102,0,42,0,199,0,160,0,59,0,245,0,0,0,249,0,0,0,120,0,26,0,12,0,124,0,219,0,222,0,116,0,107,0,33,0,0,0,53,0,0,0,18,0,39,0,0,0,217,0,0,0,0,0,129,0,214,0,0,0,42,0,0,0,139,0,0,0,67,0,109,0,0,0,63,0,166,0,14,0,0,0,13,0,0,0,64,0,106,0,255,0,190,0,251,0,0,0,65,0,127,0,221,0,88,0,92,0,70,0,213,0,0,0,49,0,130,0,61,0,3,0,30,0,3,0,88,0,129,0,255,0,27,0,23,0,117,0,144,0,8,0,219,0,153,0,128,0,98,0,199,0,186,0,134,0,225,0,118,0,45,0,100,0,208,0,58,0,189,0,0,0,2,0,42,0,191,0,160,0,135,0,229,0,0,0,0,0,128,0,226,0,95,0,0,0,171,0,217,0,106,0,53,0,230,0,152,0,0,0,233,0,54,0,153,0,91,0,231,0,158,0,94,0,194,0,0,0,192,0,0,0,122,0,0,0,88,0,0,0,135,0,232,0,43,0,246,0,163,0,39,0,0,0,254,0,176,0,0,0,0,0,139,0,0,0,134,0,212,0,3,0,112,0,76,0,158,0,206,0,238,0,59,0,0,0,224,0,78,0,140,0,211,0,210,0,104,0,204,0,142,0,33,0,85,0,153,0,17,0,0,0,130,0,90,0,0,0,115,0,69,0,20,0,0,0,98,0,0,0,55,0,141,0,11,0,27,0,226,0,0,0,149,0,17,0,5,0,0,0,171,0,101,0,252,0,138,0,20,0,0,0,0,0,10,0,53,0,165,0,0,0,0,0,155,0,111,0,80,0,81,0,202,0,100,0,0,0,0,0,0,0,176,0,0,0,75,0,42,0,0,0,173,0,33,0,220,0,242,0,0,0,10,0,0,0,0,0,233,0,0,0,23,0,10,0,0,0,75,0,0,0,123,0,0,0,2,0,227,0,199,0,17,0,165,0,53,0,0,0,56,0,195,0,199,0,77,0,145,0,115,0,225,0,189,0,0,0,250,0,197,0,222,0,96,0,143,0,190,0,0,0,111,0,103,0,17,0,0,0,194,0,168,0,23,0,4,0,214,0,168,0,75,0,237,0,139,0,206,0,0,0,63,0,204,0,0,0,0,0,7,0,0,0,121,0,25,0,225,0,229,0,45,0,96,0,29,0,0,0,36,0,162,0,0,0,227,0,203,0,126,0,18,0,0,0,46,0,0,0,30,0,63,0,79,0,111,0,0,0,1,0,129,0,35,0,0,0,214,0,0,0,93,0,181,0,0,0,0,0,125,0,221,0,0,0,103,0,27,0,189,0,196,0,120,0,12,0,100,0,189,0,0,0,0,0,124,0,67,0,0,0,39,0,151,0,128,0,152,0,0,0,100,0,30,0,214,0,0,0,0,0,0,0,194,0,197,0,52,0,0,0,228,0,0,0,0,0,0,0,60,0,74,0,58,0,141,0,27,0,48,0,0,0,201,0,210,0,2,0,188,0,82,0,163,0,85,0,0,0,236,0,0,0,46,0,214,0,184,0,204,0,197,0,123,0,115,0,139,0,0,0,0,0,28,0,0,0,101,0,122,0,144,0,216,0,98,0,213,0,60,0,148,0,59,0,215,0,42,0,11,0,79,0,165,0,211,0,37,0,167,0,154,0,48,0,0,0,33,0,200,0,235,0,0,0,12,0,86,0,201,0,12,0,63,0,0,0,0,0,93,0,227,0,232,0,60,0,63,0,6,0,93,0,95,0,154,0,117,0,142,0,33,0,153,0,161,0,0,0,87,0,34,0,0,0,133,0,48,0,57,0,189,0,32,0,200,0,241,0,176,0,186,0,229,0,194,0,143,0,193,0,245,0,111,0,182,0,169,0,193,0,87,0,0,0,151,0,8,0,0,0,218,0,170,0,36,0,27,0,34,0,130,0,244,0,192,0,208,0,145,0,206,0,0,0,35,0,30,0,251,0,0,0,171,0,45,0,15,0,65,0,3,0,35,0,31,0,169,0,161,0,5,0,32,0,93,0,0,0,0,0,3,0,0,0,14,0,233,0,0,0,150,0,81,0,103,0,78,0,110,0,76,0,15,0,250,0,224,0,31,0,76,0,0,0,95,0,0,0,129,0,185,0,120,0,26,0,7,0,216,0,145,0,0,0,43,0,72,0,199,0,177,0,132,0,0,0,196,0,123,0,156,0,75,0,146,0,3,0,44,0,112,0,144,0,172,0,0,0,111,0,158,0,106,0,22,0,181,0,0,0,176,0,8,0,74,0,31,0,244,0,133,0,160,0,91,0,216,0,41,0,193,0,127,0,120,0,0,0,147,0,236,0,70,0,255,0,0,0,79,0,61,0,214,0,37,0,229,0,10,0,133,0,0,0,0,0,3,0,0,0,201,0,79,0,0,0,213,0,164,0,0,0,132,0,233,0,250,0,0,0,50,0,48,0,211,0,0,0,249,0,182,0,0,0,229,0,73,0,1,0,40,0,98,0,238,0,0,0,223,0,202,0,193,0,71,0,0,0,0,0,137,0,0,0,100,0,9,0,129,0,38,0,212,0,182,0,55,0,249,0,0,0,171,0,149,0,0,0,200,0,0,0,0,0,231,0,237,0,0,0,202,0,33,0,70,0,148,0,28,0,0,0,148,0,191,0,94,0,201,0,186,0,90,0,180,0,57,0,9,0,84,0,0,0,0,0,75,0,40,0,0,0,43,0,138,0,13,0,201,0,112,0,229,0,212,0,100,0,0,0,67,0,0,0,0,0,130,0,38,0,55,0,79,0,220,0,80,0,0,0,104,0,151,0,138,0,247,0,180,0,25,0,0,0,195,0,14,0,144,0,165,0,181,0,125,0,153,0,0,0,0,0,217,0,169,0,0,0,0,0,227,0,11,0,66,0,207,0,54,0,204,0,0,0,55,0,193,0,14,0,72,0,240,0,221,0,1,0,233,0,28,0,253,0,0,0,148,0,0,0,69,0,69,0,0,0,0,0,91,0,246,0,0,0,61,0,0,0,12,0,0,0,11,0,114,0,49,0,209,0,245,0,106,0,54,0,133,0,201,0,0,0,93,0,0,0,15,0,0,0,117,0,83,0,54,0,4,0,242,0,208,0,242,0,0,0,174,0,78,0,77,0,118,0,0,0,224,0,0,0,47,0,0,0,251,0,8,0,25,0,145,0,165,0,39,0,110,0,216,0,0,0,217,0,108,0,81,0,4,0,250,0,221,0,202,0,116,0,0,0,127,0,0,0,0,0,203,0,0,0,177,0,108,0,231,0,169,0,119,0,111,0,70,0,201,0,0,0,175,0,167,0,132,0,228,0,123,0,0,0,126,0,18,0,0,0,124,0,0,0,83,0,204,0,0,0,0,0,0,0,225,0,56,0,0,0,22,0,37,0,225,0,93,0,0,0,110,0,0,0,115,0,5,0,193,0,0,0,249,0,115,0,0,0,126,0,45,0,44,0,252,0,245,0,92,0,0,0,26,0,139,0,195,0,0,0,114,0,169,0,0,0,79,0,48,0,14,0,0,0,212,0,131,0,215,0,16,0,226,0,84,0,121,0,113,0,254,0,214,0,135,0,114,0,241,0,207,0,80,0,225,0,0,0,107,0,160,0,47,0,31,0,54,0,189,0,213,0,0,0,0,0,243,0,90,0,0,0,27,0,106,0,49,0,36,0,0,0,162,0,151,0,7,0,13,0,0,0,179,0,37,0,0,0,206,0,148,0,0,0,207,0,0,0,123,0,24,0,149,0,121,0,141,0,160,0,167,0,88,0,137,0,99,0,0,0,208,0,103,0,0,0,233,0,81,0,38,0,231,0,0,0,0,0,35,0,97,0,0,0,93,0,116,0,0,0,181,0,0,0,0,0,56,0,173,0,148,0,0,0,0,0,193,0,255,0,156,0,201,0,107,0,96,0,156,0,78,0,207,0,149,0,40,0,232,0,243,0,0,0,15,0,191,0,0,0,205,0,22,0,92,0,0,0,101,0,188,0,96,0,149,0,41,0,141,0,83,0,142,0,134,0,60,0,43,0,0,0,0,0,0,0,237,0,193,0,8,0,45,0,0,0,201,0,122,0,208,0,36,0,172,0,0,0,0,0,133,0,0,0,0,0,23,0,242,0,0,0,0,0,0,0,198,0,138,0,0,0,227,0,0,0,169,0,114,0,0,0,229,0,169,0,140,0,172,0,137,0,0,0,82,0,18,0,0,0,230,0,201,0,142,0,142,0,0,0,141,0,32,0,221,0,8,0,0,0,126,0,33,0,0,0,42,0,0,0,2,0,0,0,216,0,0,0,185,0,0,0,109,0,0,0,28,0,78,0,122,0,169,0,38,0,152,0,58,0,0,0,0,0,117,0,47,0,129,0,31,0,136,0);
signal scenario_full  : scenario_type := (69,31,31,31,110,31,99,31,99,30,99,29,98,31,221,31,37,31,37,30,37,29,107,31,121,31,90,31,69,31,140,31,10,31,65,31,63,31,63,30,160,31,41,31,41,30,164,31,97,31,15,31,181,31,209,31,141,31,186,31,47,31,71,31,173,31,205,31,125,31,102,31,42,31,199,31,160,31,59,31,245,31,245,30,249,31,249,30,120,31,26,31,12,31,124,31,219,31,222,31,116,31,107,31,33,31,33,30,53,31,53,30,18,31,39,31,39,30,217,31,217,30,217,29,129,31,214,31,214,30,42,31,42,30,139,31,139,30,67,31,109,31,109,30,63,31,166,31,14,31,14,30,13,31,13,30,64,31,106,31,255,31,190,31,251,31,251,30,65,31,127,31,221,31,88,31,92,31,70,31,213,31,213,30,49,31,130,31,61,31,3,31,30,31,3,31,88,31,129,31,255,31,27,31,23,31,117,31,144,31,8,31,219,31,153,31,128,31,98,31,199,31,186,31,134,31,225,31,118,31,45,31,100,31,208,31,58,31,189,31,189,30,2,31,42,31,191,31,160,31,135,31,229,31,229,30,229,29,128,31,226,31,95,31,95,30,171,31,217,31,106,31,53,31,230,31,152,31,152,30,233,31,54,31,153,31,91,31,231,31,158,31,94,31,194,31,194,30,192,31,192,30,122,31,122,30,88,31,88,30,135,31,232,31,43,31,246,31,163,31,39,31,39,30,254,31,176,31,176,30,176,29,139,31,139,30,134,31,212,31,3,31,112,31,76,31,158,31,206,31,238,31,59,31,59,30,224,31,78,31,140,31,211,31,210,31,104,31,204,31,142,31,33,31,85,31,153,31,17,31,17,30,130,31,90,31,90,30,115,31,69,31,20,31,20,30,98,31,98,30,55,31,141,31,11,31,27,31,226,31,226,30,149,31,17,31,5,31,5,30,171,31,101,31,252,31,138,31,20,31,20,30,20,29,10,31,53,31,165,31,165,30,165,29,155,31,111,31,80,31,81,31,202,31,100,31,100,30,100,29,100,28,176,31,176,30,75,31,42,31,42,30,173,31,33,31,220,31,242,31,242,30,10,31,10,30,10,29,233,31,233,30,23,31,10,31,10,30,75,31,75,30,123,31,123,30,2,31,227,31,199,31,17,31,165,31,53,31,53,30,56,31,195,31,199,31,77,31,145,31,115,31,225,31,189,31,189,30,250,31,197,31,222,31,96,31,143,31,190,31,190,30,111,31,103,31,17,31,17,30,194,31,168,31,23,31,4,31,214,31,168,31,75,31,237,31,139,31,206,31,206,30,63,31,204,31,204,30,204,29,7,31,7,30,121,31,25,31,225,31,229,31,45,31,96,31,29,31,29,30,36,31,162,31,162,30,227,31,203,31,126,31,18,31,18,30,46,31,46,30,30,31,63,31,79,31,111,31,111,30,1,31,129,31,35,31,35,30,214,31,214,30,93,31,181,31,181,30,181,29,125,31,221,31,221,30,103,31,27,31,189,31,196,31,120,31,12,31,100,31,189,31,189,30,189,29,124,31,67,31,67,30,39,31,151,31,128,31,152,31,152,30,100,31,30,31,214,31,214,30,214,29,214,28,194,31,197,31,52,31,52,30,228,31,228,30,228,29,228,28,60,31,74,31,58,31,141,31,27,31,48,31,48,30,201,31,210,31,2,31,188,31,82,31,163,31,85,31,85,30,236,31,236,30,46,31,214,31,184,31,204,31,197,31,123,31,115,31,139,31,139,30,139,29,28,31,28,30,101,31,122,31,144,31,216,31,98,31,213,31,60,31,148,31,59,31,215,31,42,31,11,31,79,31,165,31,211,31,37,31,167,31,154,31,48,31,48,30,33,31,200,31,235,31,235,30,12,31,86,31,201,31,12,31,63,31,63,30,63,29,93,31,227,31,232,31,60,31,63,31,6,31,93,31,95,31,154,31,117,31,142,31,33,31,153,31,161,31,161,30,87,31,34,31,34,30,133,31,48,31,57,31,189,31,32,31,200,31,241,31,176,31,186,31,229,31,194,31,143,31,193,31,245,31,111,31,182,31,169,31,193,31,87,31,87,30,151,31,8,31,8,30,218,31,170,31,36,31,27,31,34,31,130,31,244,31,192,31,208,31,145,31,206,31,206,30,35,31,30,31,251,31,251,30,171,31,45,31,15,31,65,31,3,31,35,31,31,31,169,31,161,31,5,31,32,31,93,31,93,30,93,29,3,31,3,30,14,31,233,31,233,30,150,31,81,31,103,31,78,31,110,31,76,31,15,31,250,31,224,31,31,31,76,31,76,30,95,31,95,30,129,31,185,31,120,31,26,31,7,31,216,31,145,31,145,30,43,31,72,31,199,31,177,31,132,31,132,30,196,31,123,31,156,31,75,31,146,31,3,31,44,31,112,31,144,31,172,31,172,30,111,31,158,31,106,31,22,31,181,31,181,30,176,31,8,31,74,31,31,31,244,31,133,31,160,31,91,31,216,31,41,31,193,31,127,31,120,31,120,30,147,31,236,31,70,31,255,31,255,30,79,31,61,31,214,31,37,31,229,31,10,31,133,31,133,30,133,29,3,31,3,30,201,31,79,31,79,30,213,31,164,31,164,30,132,31,233,31,250,31,250,30,50,31,48,31,211,31,211,30,249,31,182,31,182,30,229,31,73,31,1,31,40,31,98,31,238,31,238,30,223,31,202,31,193,31,71,31,71,30,71,29,137,31,137,30,100,31,9,31,129,31,38,31,212,31,182,31,55,31,249,31,249,30,171,31,149,31,149,30,200,31,200,30,200,29,231,31,237,31,237,30,202,31,33,31,70,31,148,31,28,31,28,30,148,31,191,31,94,31,201,31,186,31,90,31,180,31,57,31,9,31,84,31,84,30,84,29,75,31,40,31,40,30,43,31,138,31,13,31,201,31,112,31,229,31,212,31,100,31,100,30,67,31,67,30,67,29,130,31,38,31,55,31,79,31,220,31,80,31,80,30,104,31,151,31,138,31,247,31,180,31,25,31,25,30,195,31,14,31,144,31,165,31,181,31,125,31,153,31,153,30,153,29,217,31,169,31,169,30,169,29,227,31,11,31,66,31,207,31,54,31,204,31,204,30,55,31,193,31,14,31,72,31,240,31,221,31,1,31,233,31,28,31,253,31,253,30,148,31,148,30,69,31,69,31,69,30,69,29,91,31,246,31,246,30,61,31,61,30,12,31,12,30,11,31,114,31,49,31,209,31,245,31,106,31,54,31,133,31,201,31,201,30,93,31,93,30,15,31,15,30,117,31,83,31,54,31,4,31,242,31,208,31,242,31,242,30,174,31,78,31,77,31,118,31,118,30,224,31,224,30,47,31,47,30,251,31,8,31,25,31,145,31,165,31,39,31,110,31,216,31,216,30,217,31,108,31,81,31,4,31,250,31,221,31,202,31,116,31,116,30,127,31,127,30,127,29,203,31,203,30,177,31,108,31,231,31,169,31,119,31,111,31,70,31,201,31,201,30,175,31,167,31,132,31,228,31,123,31,123,30,126,31,18,31,18,30,124,31,124,30,83,31,204,31,204,30,204,29,204,28,225,31,56,31,56,30,22,31,37,31,225,31,93,31,93,30,110,31,110,30,115,31,5,31,193,31,193,30,249,31,115,31,115,30,126,31,45,31,44,31,252,31,245,31,92,31,92,30,26,31,139,31,195,31,195,30,114,31,169,31,169,30,79,31,48,31,14,31,14,30,212,31,131,31,215,31,16,31,226,31,84,31,121,31,113,31,254,31,214,31,135,31,114,31,241,31,207,31,80,31,225,31,225,30,107,31,160,31,47,31,31,31,54,31,189,31,213,31,213,30,213,29,243,31,90,31,90,30,27,31,106,31,49,31,36,31,36,30,162,31,151,31,7,31,13,31,13,30,179,31,37,31,37,30,206,31,148,31,148,30,207,31,207,30,123,31,24,31,149,31,121,31,141,31,160,31,167,31,88,31,137,31,99,31,99,30,208,31,103,31,103,30,233,31,81,31,38,31,231,31,231,30,231,29,35,31,97,31,97,30,93,31,116,31,116,30,181,31,181,30,181,29,56,31,173,31,148,31,148,30,148,29,193,31,255,31,156,31,201,31,107,31,96,31,156,31,78,31,207,31,149,31,40,31,232,31,243,31,243,30,15,31,191,31,191,30,205,31,22,31,92,31,92,30,101,31,188,31,96,31,149,31,41,31,141,31,83,31,142,31,134,31,60,31,43,31,43,30,43,29,43,28,237,31,193,31,8,31,45,31,45,30,201,31,122,31,208,31,36,31,172,31,172,30,172,29,133,31,133,30,133,29,23,31,242,31,242,30,242,29,242,28,198,31,138,31,138,30,227,31,227,30,169,31,114,31,114,30,229,31,169,31,140,31,172,31,137,31,137,30,82,31,18,31,18,30,230,31,201,31,142,31,142,31,142,30,141,31,32,31,221,31,8,31,8,30,126,31,33,31,33,30,42,31,42,30,2,31,2,30,216,31,216,30,185,31,185,30,109,31,109,30,28,31,78,31,122,31,169,31,38,31,152,31,58,31,58,30,58,29,117,31,47,31,129,31,31,31,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
