-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 317;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,253,0,249,0,127,0,75,0,64,0,186,0,44,0,56,0,119,0,233,0,89,0,50,0,68,0,190,0,0,0,172,0,162,0,6,0,0,0,78,0,231,0,0,0,187,0,0,0,0,0,138,0,88,0,202,0,118,0,124,0,0,0,93,0,137,0,244,0,211,0,51,0,0,0,241,0,201,0,7,0,44,0,157,0,217,0,178,0,78,0,115,0,44,0,242,0,0,0,44,0,0,0,0,0,181,0,27,0,124,0,26,0,0,0,69,0,195,0,0,0,0,0,0,0,0,0,47,0,51,0,98,0,214,0,78,0,133,0,167,0,183,0,62,0,194,0,121,0,225,0,96,0,120,0,62,0,7,0,4,0,17,0,140,0,108,0,234,0,117,0,112,0,0,0,71,0,212,0,97,0,62,0,136,0,181,0,0,0,240,0,209,0,0,0,92,0,0,0,8,0,235,0,242,0,0,0,0,0,205,0,73,0,208,0,108,0,126,0,115,0,56,0,244,0,222,0,153,0,0,0,141,0,125,0,77,0,108,0,0,0,148,0,76,0,0,0,233,0,67,0,0,0,76,0,140,0,140,0,251,0,162,0,160,0,222,0,57,0,169,0,191,0,75,0,0,0,203,0,245,0,123,0,0,0,100,0,140,0,179,0,168,0,6,0,229,0,100,0,104,0,0,0,225,0,33,0,52,0,42,0,100,0,147,0,110,0,163,0,216,0,0,0,149,0,7,0,21,0,0,0,212,0,54,0,170,0,158,0,86,0,20,0,47,0,48,0,0,0,0,0,72,0,39,0,154,0,17,0,212,0,0,0,224,0,126,0,202,0,242,0,10,0,94,0,0,0,149,0,67,0,29,0,227,0,65,0,206,0,0,0,147,0,198,0,68,0,105,0,0,0,200,0,59,0,148,0,0,0,200,0,59,0,155,0,13,0,111,0,0,0,16,0,252,0,0,0,236,0,202,0,56,0,113,0,0,0,0,0,229,0,0,0,63,0,156,0,135,0,145,0,0,0,58,0,230,0,0,0,139,0,0,0,136,0,165,0,127,0,115,0,245,0,190,0,74,0,208,0,195,0,1,0,0,0,0,0,119,0,1,0,69,0,123,0,99,0,92,0,196,0,0,0,0,0,10,0,240,0,76,0,0,0,246,0,0,0,170,0,211,0,161,0,218,0,22,0,23,0,51,0,130,0,156,0,248,0,123,0,221,0,221,0,62,0,166,0,0,0,0,0,255,0,210,0,54,0,166,0,0,0,197,0,59,0,206,0,131,0,106,0,0,0,87,0,0,0,115,0,233,0,196,0,62,0,140,0,40,0,155,0,39,0,210,0,252,0,187,0,28,0,81,0,43,0,59,0,2,0,180,0,104,0,0,0,43,0,245,0,23,0,175,0,195,0,151,0,10,0,49,0,22,0);
signal scenario_full  : scenario_type := (0,0,253,31,249,31,127,31,75,31,64,31,186,31,44,31,56,31,119,31,233,31,89,31,50,31,68,31,190,31,190,30,172,31,162,31,6,31,6,30,78,31,231,31,231,30,187,31,187,30,187,29,138,31,88,31,202,31,118,31,124,31,124,30,93,31,137,31,244,31,211,31,51,31,51,30,241,31,201,31,7,31,44,31,157,31,217,31,178,31,78,31,115,31,44,31,242,31,242,30,44,31,44,30,44,29,181,31,27,31,124,31,26,31,26,30,69,31,195,31,195,30,195,29,195,28,195,27,47,31,51,31,98,31,214,31,78,31,133,31,167,31,183,31,62,31,194,31,121,31,225,31,96,31,120,31,62,31,7,31,4,31,17,31,140,31,108,31,234,31,117,31,112,31,112,30,71,31,212,31,97,31,62,31,136,31,181,31,181,30,240,31,209,31,209,30,92,31,92,30,8,31,235,31,242,31,242,30,242,29,205,31,73,31,208,31,108,31,126,31,115,31,56,31,244,31,222,31,153,31,153,30,141,31,125,31,77,31,108,31,108,30,148,31,76,31,76,30,233,31,67,31,67,30,76,31,140,31,140,31,251,31,162,31,160,31,222,31,57,31,169,31,191,31,75,31,75,30,203,31,245,31,123,31,123,30,100,31,140,31,179,31,168,31,6,31,229,31,100,31,104,31,104,30,225,31,33,31,52,31,42,31,100,31,147,31,110,31,163,31,216,31,216,30,149,31,7,31,21,31,21,30,212,31,54,31,170,31,158,31,86,31,20,31,47,31,48,31,48,30,48,29,72,31,39,31,154,31,17,31,212,31,212,30,224,31,126,31,202,31,242,31,10,31,94,31,94,30,149,31,67,31,29,31,227,31,65,31,206,31,206,30,147,31,198,31,68,31,105,31,105,30,200,31,59,31,148,31,148,30,200,31,59,31,155,31,13,31,111,31,111,30,16,31,252,31,252,30,236,31,202,31,56,31,113,31,113,30,113,29,229,31,229,30,63,31,156,31,135,31,145,31,145,30,58,31,230,31,230,30,139,31,139,30,136,31,165,31,127,31,115,31,245,31,190,31,74,31,208,31,195,31,1,31,1,30,1,29,119,31,1,31,69,31,123,31,99,31,92,31,196,31,196,30,196,29,10,31,240,31,76,31,76,30,246,31,246,30,170,31,211,31,161,31,218,31,22,31,23,31,51,31,130,31,156,31,248,31,123,31,221,31,221,31,62,31,166,31,166,30,166,29,255,31,210,31,54,31,166,31,166,30,197,31,59,31,206,31,131,31,106,31,106,30,87,31,87,30,115,31,233,31,196,31,62,31,140,31,40,31,155,31,39,31,210,31,252,31,187,31,28,31,81,31,43,31,59,31,2,31,180,31,104,31,104,30,43,31,245,31,23,31,175,31,195,31,151,31,10,31,49,31,22,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
