-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 851;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (179,0,29,0,0,0,43,0,161,0,189,0,17,0,0,0,181,0,143,0,21,0,182,0,0,0,0,0,29,0,0,0,125,0,17,0,0,0,53,0,73,0,122,0,27,0,116,0,156,0,0,0,154,0,172,0,208,0,202,0,26,0,133,0,0,0,198,0,106,0,218,0,185,0,82,0,252,0,112,0,118,0,23,0,243,0,128,0,25,0,52,0,67,0,73,0,107,0,0,0,176,0,53,0,136,0,96,0,155,0,61,0,83,0,207,0,0,0,36,0,66,0,65,0,191,0,0,0,66,0,72,0,0,0,0,0,0,0,0,0,0,0,101,0,0,0,0,0,109,0,145,0,200,0,0,0,229,0,0,0,2,0,186,0,0,0,0,0,203,0,72,0,255,0,250,0,161,0,142,0,46,0,209,0,0,0,252,0,147,0,241,0,4,0,214,0,254,0,16,0,245,0,183,0,0,0,0,0,215,0,245,0,229,0,178,0,108,0,0,0,16,0,87,0,50,0,0,0,28,0,0,0,2,0,244,0,75,0,45,0,138,0,211,0,0,0,221,0,220,0,0,0,137,0,108,0,136,0,46,0,0,0,245,0,178,0,129,0,107,0,56,0,20,0,4,0,154,0,26,0,198,0,33,0,28,0,221,0,0,0,0,0,148,0,0,0,123,0,0,0,187,0,43,0,0,0,149,0,117,0,48,0,19,0,165,0,214,0,0,0,54,0,0,0,8,0,92,0,35,0,86,0,30,0,20,0,231,0,247,0,0,0,0,0,6,0,239,0,0,0,202,0,0,0,125,0,16,0,0,0,253,0,58,0,65,0,115,0,193,0,57,0,134,0,95,0,226,0,156,0,196,0,94,0,155,0,0,0,134,0,27,0,69,0,231,0,37,0,9,0,0,0,150,0,168,0,189,0,97,0,78,0,29,0,2,0,119,0,170,0,53,0,189,0,0,0,0,0,182,0,202,0,0,0,103,0,137,0,79,0,0,0,205,0,163,0,0,0,242,0,93,0,79,0,197,0,0,0,41,0,4,0,154,0,139,0,89,0,0,0,228,0,139,0,109,0,234,0,59,0,173,0,174,0,189,0,0,0,25,0,0,0,0,0,0,0,180,0,146,0,206,0,101,0,102,0,108,0,0,0,253,0,2,0,0,0,164,0,75,0,80,0,250,0,51,0,204,0,33,0,72,0,180,0,0,0,0,0,44,0,174,0,236,0,0,0,58,0,160,0,151,0,0,0,119,0,215,0,95,0,148,0,0,0,1,0,84,0,121,0,9,0,146,0,126,0,116,0,101,0,60,0,0,0,71,0,252,0,203,0,0,0,100,0,0,0,0,0,247,0,0,0,8,0,107,0,39,0,79,0,0,0,142,0,42,0,0,0,0,0,123,0,184,0,184,0,199,0,73,0,0,0,0,0,39,0,127,0,249,0,56,0,207,0,68,0,10,0,0,0,205,0,80,0,13,0,0,0,143,0,58,0,231,0,116,0,170,0,0,0,48,0,88,0,252,0,0,0,97,0,111,0,148,0,227,0,0,0,50,0,223,0,154,0,206,0,95,0,207,0,44,0,223,0,108,0,217,0,185,0,50,0,89,0,149,0,177,0,203,0,67,0,238,0,4,0,247,0,240,0,224,0,215,0,4,0,219,0,41,0,29,0,254,0,0,0,141,0,144,0,31,0,57,0,5,0,30,0,228,0,91,0,144,0,156,0,247,0,0,0,251,0,0,0,210,0,0,0,121,0,0,0,112,0,203,0,40,0,73,0,173,0,0,0,192,0,88,0,248,0,155,0,0,0,0,0,0,0,129,0,219,0,203,0,133,0,0,0,255,0,0,0,0,0,18,0,85,0,149,0,110,0,209,0,0,0,254,0,119,0,0,0,152,0,115,0,137,0,0,0,196,0,144,0,144,0,134,0,202,0,0,0,172,0,236,0,83,0,34,0,254,0,0,0,149,0,214,0,110,0,195,0,154,0,211,0,64,0,6,0,93,0,0,0,0,0,193,0,0,0,65,0,203,0,109,0,127,0,223,0,66,0,2,0,54,0,0,0,150,0,0,0,252,0,0,0,58,0,241,0,36,0,0,0,61,0,0,0,131,0,196,0,245,0,86,0,150,0,112,0,209,0,0,0,151,0,22,0,166,0,156,0,11,0,235,0,153,0,248,0,97,0,87,0,122,0,91,0,124,0,84,0,88,0,10,0,199,0,157,0,167,0,0,0,0,0,9,0,28,0,45,0,7,0,0,0,146,0,0,0,239,0,128,0,99,0,209,0,41,0,32,0,0,0,0,0,135,0,0,0,183,0,237,0,36,0,173,0,14,0,5,0,139,0,128,0,133,0,241,0,198,0,247,0,97,0,51,0,117,0,0,0,0,0,0,0,0,0,240,0,0,0,0,0,82,0,50,0,255,0,88,0,209,0,73,0,20,0,0,0,0,0,126,0,216,0,4,0,244,0,168,0,0,0,42,0,193,0,242,0,243,0,90,0,58,0,0,0,67,0,157,0,189,0,236,0,115,0,48,0,0,0,57,0,249,0,215,0,0,0,247,0,0,0,0,0,0,0,143,0,181,0,251,0,30,0,99,0,128,0,172,0,154,0,216,0,66,0,189,0,81,0,0,0,47,0,0,0,217,0,221,0,157,0,40,0,216,0,80,0,194,0,98,0,195,0,198,0,97,0,187,0,190,0,91,0,0,0,2,0,183,0,99,0,231,0,49,0,34,0,183,0,142,0,246,0,21,0,27,0,40,0,76,0,0,0,0,0,0,0,192,0,25,0,227,0,0,0,40,0,130,0,215,0,113,0,250,0,46,0,206,0,140,0,0,0,253,0,209,0,0,0,60,0,69,0,0,0,160,0,6,0,0,0,108,0,28,0,0,0,150,0,193,0,21,0,79,0,0,0,104,0,253,0,0,0,133,0,22,0,149,0,190,0,221,0,0,0,0,0,185,0,166,0,104,0,186,0,8,0,217,0,95,0,0,0,177,0,144,0,56,0,177,0,167,0,32,0,82,0,0,0,199,0,146,0,144,0,120,0,107,0,0,0,0,0,8,0,166,0,0,0,6,0,31,0,182,0,151,0,17,0,204,0,64,0,93,0,203,0,162,0,240,0,119,0,109,0,88,0,0,0,232,0,0,0,39,0,63,0,98,0,61,0,104,0,249,0,0,0,71,0,181,0,0,0,0,0,130,0,40,0,0,0,0,0,102,0,226,0,21,0,195,0,231,0,208,0,124,0,3,0,246,0,62,0,183,0,0,0,0,0,169,0,51,0,175,0,9,0,153,0,50,0,105,0,183,0,0,0,13,0,192,0,0,0,107,0,241,0,130,0,28,0,49,0,0,0,240,0,36,0,168,0,77,0,0,0,220,0,207,0,177,0,152,0,232,0,96,0,63,0,214,0,143,0,175,0,0,0,137,0,17,0,212,0,171,0,54,0,186,0,112,0,111,0,210,0,173,0,122,0,0,0,18,0,109,0,243,0,229,0,184,0,9,0,0,0,230,0,153,0,67,0,16,0,249,0,34,0,14,0,247,0,8,0,152,0,133,0,133,0,241,0,207,0,0,0,63,0,138,0,194,0,53,0,194,0,226,0,167,0,54,0,253,0,0,0,165,0,168,0,169,0,235,0,31,0,143,0,71,0,163,0,242,0,66,0,102,0,222,0,144,0,112,0,137,0,0,0,173,0,0,0,37,0,101,0,193,0,0,0,43,0,231,0,203,0,167,0,75,0,211,0,6,0,73,0,67,0,189,0,0,0,111,0,162,0,241,0,0,0,158,0,14,0,138,0,57,0,253,0);
signal scenario_full  : scenario_type := (179,31,29,31,29,30,43,31,161,31,189,31,17,31,17,30,181,31,143,31,21,31,182,31,182,30,182,29,29,31,29,30,125,31,17,31,17,30,53,31,73,31,122,31,27,31,116,31,156,31,156,30,154,31,172,31,208,31,202,31,26,31,133,31,133,30,198,31,106,31,218,31,185,31,82,31,252,31,112,31,118,31,23,31,243,31,128,31,25,31,52,31,67,31,73,31,107,31,107,30,176,31,53,31,136,31,96,31,155,31,61,31,83,31,207,31,207,30,36,31,66,31,65,31,191,31,191,30,66,31,72,31,72,30,72,29,72,28,72,27,72,26,101,31,101,30,101,29,109,31,145,31,200,31,200,30,229,31,229,30,2,31,186,31,186,30,186,29,203,31,72,31,255,31,250,31,161,31,142,31,46,31,209,31,209,30,252,31,147,31,241,31,4,31,214,31,254,31,16,31,245,31,183,31,183,30,183,29,215,31,245,31,229,31,178,31,108,31,108,30,16,31,87,31,50,31,50,30,28,31,28,30,2,31,244,31,75,31,45,31,138,31,211,31,211,30,221,31,220,31,220,30,137,31,108,31,136,31,46,31,46,30,245,31,178,31,129,31,107,31,56,31,20,31,4,31,154,31,26,31,198,31,33,31,28,31,221,31,221,30,221,29,148,31,148,30,123,31,123,30,187,31,43,31,43,30,149,31,117,31,48,31,19,31,165,31,214,31,214,30,54,31,54,30,8,31,92,31,35,31,86,31,30,31,20,31,231,31,247,31,247,30,247,29,6,31,239,31,239,30,202,31,202,30,125,31,16,31,16,30,253,31,58,31,65,31,115,31,193,31,57,31,134,31,95,31,226,31,156,31,196,31,94,31,155,31,155,30,134,31,27,31,69,31,231,31,37,31,9,31,9,30,150,31,168,31,189,31,97,31,78,31,29,31,2,31,119,31,170,31,53,31,189,31,189,30,189,29,182,31,202,31,202,30,103,31,137,31,79,31,79,30,205,31,163,31,163,30,242,31,93,31,79,31,197,31,197,30,41,31,4,31,154,31,139,31,89,31,89,30,228,31,139,31,109,31,234,31,59,31,173,31,174,31,189,31,189,30,25,31,25,30,25,29,25,28,180,31,146,31,206,31,101,31,102,31,108,31,108,30,253,31,2,31,2,30,164,31,75,31,80,31,250,31,51,31,204,31,33,31,72,31,180,31,180,30,180,29,44,31,174,31,236,31,236,30,58,31,160,31,151,31,151,30,119,31,215,31,95,31,148,31,148,30,1,31,84,31,121,31,9,31,146,31,126,31,116,31,101,31,60,31,60,30,71,31,252,31,203,31,203,30,100,31,100,30,100,29,247,31,247,30,8,31,107,31,39,31,79,31,79,30,142,31,42,31,42,30,42,29,123,31,184,31,184,31,199,31,73,31,73,30,73,29,39,31,127,31,249,31,56,31,207,31,68,31,10,31,10,30,205,31,80,31,13,31,13,30,143,31,58,31,231,31,116,31,170,31,170,30,48,31,88,31,252,31,252,30,97,31,111,31,148,31,227,31,227,30,50,31,223,31,154,31,206,31,95,31,207,31,44,31,223,31,108,31,217,31,185,31,50,31,89,31,149,31,177,31,203,31,67,31,238,31,4,31,247,31,240,31,224,31,215,31,4,31,219,31,41,31,29,31,254,31,254,30,141,31,144,31,31,31,57,31,5,31,30,31,228,31,91,31,144,31,156,31,247,31,247,30,251,31,251,30,210,31,210,30,121,31,121,30,112,31,203,31,40,31,73,31,173,31,173,30,192,31,88,31,248,31,155,31,155,30,155,29,155,28,129,31,219,31,203,31,133,31,133,30,255,31,255,30,255,29,18,31,85,31,149,31,110,31,209,31,209,30,254,31,119,31,119,30,152,31,115,31,137,31,137,30,196,31,144,31,144,31,134,31,202,31,202,30,172,31,236,31,83,31,34,31,254,31,254,30,149,31,214,31,110,31,195,31,154,31,211,31,64,31,6,31,93,31,93,30,93,29,193,31,193,30,65,31,203,31,109,31,127,31,223,31,66,31,2,31,54,31,54,30,150,31,150,30,252,31,252,30,58,31,241,31,36,31,36,30,61,31,61,30,131,31,196,31,245,31,86,31,150,31,112,31,209,31,209,30,151,31,22,31,166,31,156,31,11,31,235,31,153,31,248,31,97,31,87,31,122,31,91,31,124,31,84,31,88,31,10,31,199,31,157,31,167,31,167,30,167,29,9,31,28,31,45,31,7,31,7,30,146,31,146,30,239,31,128,31,99,31,209,31,41,31,32,31,32,30,32,29,135,31,135,30,183,31,237,31,36,31,173,31,14,31,5,31,139,31,128,31,133,31,241,31,198,31,247,31,97,31,51,31,117,31,117,30,117,29,117,28,117,27,240,31,240,30,240,29,82,31,50,31,255,31,88,31,209,31,73,31,20,31,20,30,20,29,126,31,216,31,4,31,244,31,168,31,168,30,42,31,193,31,242,31,243,31,90,31,58,31,58,30,67,31,157,31,189,31,236,31,115,31,48,31,48,30,57,31,249,31,215,31,215,30,247,31,247,30,247,29,247,28,143,31,181,31,251,31,30,31,99,31,128,31,172,31,154,31,216,31,66,31,189,31,81,31,81,30,47,31,47,30,217,31,221,31,157,31,40,31,216,31,80,31,194,31,98,31,195,31,198,31,97,31,187,31,190,31,91,31,91,30,2,31,183,31,99,31,231,31,49,31,34,31,183,31,142,31,246,31,21,31,27,31,40,31,76,31,76,30,76,29,76,28,192,31,25,31,227,31,227,30,40,31,130,31,215,31,113,31,250,31,46,31,206,31,140,31,140,30,253,31,209,31,209,30,60,31,69,31,69,30,160,31,6,31,6,30,108,31,28,31,28,30,150,31,193,31,21,31,79,31,79,30,104,31,253,31,253,30,133,31,22,31,149,31,190,31,221,31,221,30,221,29,185,31,166,31,104,31,186,31,8,31,217,31,95,31,95,30,177,31,144,31,56,31,177,31,167,31,32,31,82,31,82,30,199,31,146,31,144,31,120,31,107,31,107,30,107,29,8,31,166,31,166,30,6,31,31,31,182,31,151,31,17,31,204,31,64,31,93,31,203,31,162,31,240,31,119,31,109,31,88,31,88,30,232,31,232,30,39,31,63,31,98,31,61,31,104,31,249,31,249,30,71,31,181,31,181,30,181,29,130,31,40,31,40,30,40,29,102,31,226,31,21,31,195,31,231,31,208,31,124,31,3,31,246,31,62,31,183,31,183,30,183,29,169,31,51,31,175,31,9,31,153,31,50,31,105,31,183,31,183,30,13,31,192,31,192,30,107,31,241,31,130,31,28,31,49,31,49,30,240,31,36,31,168,31,77,31,77,30,220,31,207,31,177,31,152,31,232,31,96,31,63,31,214,31,143,31,175,31,175,30,137,31,17,31,212,31,171,31,54,31,186,31,112,31,111,31,210,31,173,31,122,31,122,30,18,31,109,31,243,31,229,31,184,31,9,31,9,30,230,31,153,31,67,31,16,31,249,31,34,31,14,31,247,31,8,31,152,31,133,31,133,31,241,31,207,31,207,30,63,31,138,31,194,31,53,31,194,31,226,31,167,31,54,31,253,31,253,30,165,31,168,31,169,31,235,31,31,31,143,31,71,31,163,31,242,31,66,31,102,31,222,31,144,31,112,31,137,31,137,30,173,31,173,30,37,31,101,31,193,31,193,30,43,31,231,31,203,31,167,31,75,31,211,31,6,31,73,31,67,31,189,31,189,30,111,31,162,31,241,31,241,30,158,31,14,31,138,31,57,31,253,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
