-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_313 is
end project_tb_313;

architecture project_tb_arch_313 of project_tb_313 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 550;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,186,0,0,0,233,0,47,0,144,0,183,0,79,0,131,0,82,0,148,0,138,0,71,0,0,0,0,0,0,0,15,0,61,0,233,0,26,0,250,0,130,0,0,0,247,0,162,0,8,0,211,0,171,0,200,0,126,0,169,0,250,0,188,0,0,0,30,0,82,0,22,0,155,0,192,0,0,0,135,0,177,0,45,0,198,0,0,0,213,0,30,0,31,0,14,0,0,0,109,0,119,0,249,0,12,0,0,0,0,0,206,0,250,0,208,0,0,0,0,0,75,0,0,0,25,0,0,0,66,0,30,0,0,0,0,0,160,0,228,0,70,0,84,0,184,0,0,0,144,0,145,0,221,0,157,0,69,0,161,0,81,0,0,0,7,0,114,0,132,0,9,0,20,0,172,0,115,0,23,0,203,0,78,0,54,0,252,0,0,0,191,0,97,0,225,0,150,0,168,0,62,0,125,0,232,0,107,0,97,0,141,0,204,0,0,0,0,0,119,0,233,0,173,0,0,0,216,0,71,0,87,0,110,0,0,0,160,0,29,0,0,0,51,0,81,0,0,0,210,0,224,0,0,0,118,0,0,0,57,0,190,0,119,0,130,0,23,0,89,0,183,0,247,0,164,0,162,0,37,0,197,0,48,0,68,0,208,0,217,0,21,0,249,0,104,0,207,0,90,0,190,0,236,0,0,0,0,0,10,0,58,0,0,0,124,0,101,0,0,0,30,0,91,0,142,0,78,0,140,0,192,0,8,0,211,0,112,0,234,0,141,0,232,0,158,0,121,0,3,0,245,0,182,0,0,0,139,0,169,0,0,0,11,0,0,0,17,0,244,0,0,0,147,0,57,0,94,0,202,0,19,0,85,0,110,0,118,0,12,0,72,0,120,0,113,0,124,0,104,0,0,0,0,0,0,0,250,0,0,0,214,0,202,0,61,0,0,0,181,0,219,0,0,0,0,0,65,0,22,0,143,0,221,0,208,0,0,0,219,0,0,0,0,0,172,0,6,0,195,0,0,0,212,0,12,0,82,0,249,0,208,0,136,0,169,0,89,0,237,0,148,0,0,0,0,0,168,0,120,0,44,0,54,0,0,0,79,0,232,0,221,0,139,0,242,0,0,0,203,0,0,0,47,0,194,0,120,0,240,0,0,0,79,0,246,0,10,0,0,0,0,0,0,0,115,0,61,0,0,0,198,0,163,0,17,0,75,0,204,0,0,0,138,0,114,0,248,0,70,0,172,0,52,0,186,0,0,0,97,0,62,0,225,0,0,0,92,0,168,0,212,0,166,0,0,0,3,0,141,0,26,0,0,0,109,0,132,0,230,0,178,0,29,0,116,0,0,0,148,0,119,0,0,0,229,0,182,0,11,0,72,0,0,0,59,0,24,0,36,0,84,0,113,0,72,0,162,0,166,0,85,0,5,0,0,0,209,0,150,0,34,0,138,0,0,0,0,0,121,0,222,0,38,0,0,0,17,0,80,0,78,0,97,0,173,0,178,0,158,0,162,0,43,0,42,0,107,0,229,0,171,0,0,0,77,0,171,0,0,0,157,0,64,0,0,0,79,0,0,0,124,0,0,0,0,0,158,0,201,0,106,0,168,0,120,0,228,0,11,0,124,0,188,0,194,0,222,0,35,0,34,0,72,0,229,0,238,0,245,0,45,0,0,0,138,0,181,0,0,0,183,0,0,0,238,0,155,0,239,0,129,0,147,0,243,0,0,0,34,0,62,0,28,0,88,0,119,0,181,0,134,0,137,0,0,0,183,0,13,0,208,0,249,0,0,0,133,0,241,0,0,0,154,0,139,0,11,0,216,0,73,0,203,0,120,0,17,0,213,0,233,0,99,0,8,0,0,0,85,0,0,0,13,0,94,0,191,0,253,0,204,0,0,0,246,0,83,0,219,0,107,0,0,0,122,0,0,0,197,0,35,0,160,0,64,0,0,0,0,0,146,0,0,0,155,0,55,0,0,0,158,0,45,0,19,0,108,0,99,0,35,0,5,0,0,0,135,0,0,0,166,0,51,0,134,0,0,0,70,0,0,0,235,0,205,0,97,0,120,0,0,0,0,0,0,0,134,0,242,0,0,0,0,0,188,0,47,0,156,0,0,0,117,0,225,0,127,0,131,0,54,0,178,0,40,0,29,0,0,0,153,0,191,0,29,0,241,0,0,0,108,0,62,0,114,0,34,0,32,0,32,0,5,0,0,0,0,0,88,0,0,0,104,0,0,0,90,0,245,0,66,0,116,0,145,0,0,0,59,0,110,0,59,0,230,0,100,0,94,0,0,0,90,0,217,0,107,0,217,0,157,0,158,0,0,0,0,0,68,0,60,0,100,0,139,0,64,0,27,0,0,0,6,0,228,0,127,0,190,0,8,0,81,0,5,0,197,0,23,0,248,0,133,0,0,0,0,0,141,0,83,0,156,0,192,0,149,0,206,0,0,0,199,0,2,0,0,0);
signal scenario_full  : scenario_type := (128,31,186,31,186,30,233,31,47,31,144,31,183,31,79,31,131,31,82,31,148,31,138,31,71,31,71,30,71,29,71,28,15,31,61,31,233,31,26,31,250,31,130,31,130,30,247,31,162,31,8,31,211,31,171,31,200,31,126,31,169,31,250,31,188,31,188,30,30,31,82,31,22,31,155,31,192,31,192,30,135,31,177,31,45,31,198,31,198,30,213,31,30,31,31,31,14,31,14,30,109,31,119,31,249,31,12,31,12,30,12,29,206,31,250,31,208,31,208,30,208,29,75,31,75,30,25,31,25,30,66,31,30,31,30,30,30,29,160,31,228,31,70,31,84,31,184,31,184,30,144,31,145,31,221,31,157,31,69,31,161,31,81,31,81,30,7,31,114,31,132,31,9,31,20,31,172,31,115,31,23,31,203,31,78,31,54,31,252,31,252,30,191,31,97,31,225,31,150,31,168,31,62,31,125,31,232,31,107,31,97,31,141,31,204,31,204,30,204,29,119,31,233,31,173,31,173,30,216,31,71,31,87,31,110,31,110,30,160,31,29,31,29,30,51,31,81,31,81,30,210,31,224,31,224,30,118,31,118,30,57,31,190,31,119,31,130,31,23,31,89,31,183,31,247,31,164,31,162,31,37,31,197,31,48,31,68,31,208,31,217,31,21,31,249,31,104,31,207,31,90,31,190,31,236,31,236,30,236,29,10,31,58,31,58,30,124,31,101,31,101,30,30,31,91,31,142,31,78,31,140,31,192,31,8,31,211,31,112,31,234,31,141,31,232,31,158,31,121,31,3,31,245,31,182,31,182,30,139,31,169,31,169,30,11,31,11,30,17,31,244,31,244,30,147,31,57,31,94,31,202,31,19,31,85,31,110,31,118,31,12,31,72,31,120,31,113,31,124,31,104,31,104,30,104,29,104,28,250,31,250,30,214,31,202,31,61,31,61,30,181,31,219,31,219,30,219,29,65,31,22,31,143,31,221,31,208,31,208,30,219,31,219,30,219,29,172,31,6,31,195,31,195,30,212,31,12,31,82,31,249,31,208,31,136,31,169,31,89,31,237,31,148,31,148,30,148,29,168,31,120,31,44,31,54,31,54,30,79,31,232,31,221,31,139,31,242,31,242,30,203,31,203,30,47,31,194,31,120,31,240,31,240,30,79,31,246,31,10,31,10,30,10,29,10,28,115,31,61,31,61,30,198,31,163,31,17,31,75,31,204,31,204,30,138,31,114,31,248,31,70,31,172,31,52,31,186,31,186,30,97,31,62,31,225,31,225,30,92,31,168,31,212,31,166,31,166,30,3,31,141,31,26,31,26,30,109,31,132,31,230,31,178,31,29,31,116,31,116,30,148,31,119,31,119,30,229,31,182,31,11,31,72,31,72,30,59,31,24,31,36,31,84,31,113,31,72,31,162,31,166,31,85,31,5,31,5,30,209,31,150,31,34,31,138,31,138,30,138,29,121,31,222,31,38,31,38,30,17,31,80,31,78,31,97,31,173,31,178,31,158,31,162,31,43,31,42,31,107,31,229,31,171,31,171,30,77,31,171,31,171,30,157,31,64,31,64,30,79,31,79,30,124,31,124,30,124,29,158,31,201,31,106,31,168,31,120,31,228,31,11,31,124,31,188,31,194,31,222,31,35,31,34,31,72,31,229,31,238,31,245,31,45,31,45,30,138,31,181,31,181,30,183,31,183,30,238,31,155,31,239,31,129,31,147,31,243,31,243,30,34,31,62,31,28,31,88,31,119,31,181,31,134,31,137,31,137,30,183,31,13,31,208,31,249,31,249,30,133,31,241,31,241,30,154,31,139,31,11,31,216,31,73,31,203,31,120,31,17,31,213,31,233,31,99,31,8,31,8,30,85,31,85,30,13,31,94,31,191,31,253,31,204,31,204,30,246,31,83,31,219,31,107,31,107,30,122,31,122,30,197,31,35,31,160,31,64,31,64,30,64,29,146,31,146,30,155,31,55,31,55,30,158,31,45,31,19,31,108,31,99,31,35,31,5,31,5,30,135,31,135,30,166,31,51,31,134,31,134,30,70,31,70,30,235,31,205,31,97,31,120,31,120,30,120,29,120,28,134,31,242,31,242,30,242,29,188,31,47,31,156,31,156,30,117,31,225,31,127,31,131,31,54,31,178,31,40,31,29,31,29,30,153,31,191,31,29,31,241,31,241,30,108,31,62,31,114,31,34,31,32,31,32,31,5,31,5,30,5,29,88,31,88,30,104,31,104,30,90,31,245,31,66,31,116,31,145,31,145,30,59,31,110,31,59,31,230,31,100,31,94,31,94,30,90,31,217,31,107,31,217,31,157,31,158,31,158,30,158,29,68,31,60,31,100,31,139,31,64,31,27,31,27,30,6,31,228,31,127,31,190,31,8,31,81,31,5,31,197,31,23,31,248,31,133,31,133,30,133,29,141,31,83,31,156,31,192,31,149,31,206,31,206,30,199,31,2,31,2,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
