-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 849;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (62,0,0,0,98,0,0,0,248,0,65,0,129,0,207,0,94,0,26,0,195,0,159,0,221,0,118,0,37,0,203,0,66,0,0,0,178,0,89,0,217,0,53,0,221,0,3,0,44,0,83,0,243,0,37,0,204,0,134,0,228,0,0,0,244,0,140,0,32,0,16,0,0,0,37,0,95,0,218,0,221,0,84,0,163,0,164,0,95,0,0,0,74,0,226,0,255,0,68,0,135,0,166,0,59,0,53,0,111,0,174,0,141,0,188,0,0,0,35,0,49,0,0,0,146,0,102,0,116,0,17,0,0,0,0,0,141,0,174,0,0,0,80,0,0,0,99,0,241,0,0,0,82,0,53,0,124,0,22,0,171,0,210,0,127,0,185,0,107,0,0,0,0,0,0,0,65,0,201,0,0,0,7,0,70,0,0,0,0,0,103,0,0,0,0,0,0,0,60,0,233,0,0,0,0,0,102,0,61,0,125,0,25,0,64,0,18,0,196,0,174,0,12,0,47,0,58,0,131,0,0,0,149,0,241,0,36,0,175,0,172,0,156,0,0,0,119,0,124,0,40,0,41,0,0,0,189,0,0,0,171,0,53,0,110,0,140,0,41,0,241,0,0,0,131,0,164,0,86,0,114,0,21,0,27,0,245,0,140,0,0,0,163,0,221,0,150,0,16,0,30,0,199,0,0,0,87,0,0,0,203,0,165,0,89,0,19,0,228,0,170,0,210,0,24,0,101,0,15,0,219,0,0,0,0,0,61,0,241,0,0,0,0,0,0,0,0,0,126,0,110,0,117,0,0,0,226,0,59,0,201,0,108,0,134,0,254,0,16,0,70,0,38,0,122,0,225,0,208,0,27,0,0,0,135,0,132,0,221,0,78,0,0,0,128,0,142,0,94,0,203,0,87,0,0,0,0,0,64,0,197,0,0,0,112,0,98,0,189,0,0,0,0,0,1,0,28,0,122,0,99,0,11,0,131,0,0,0,81,0,0,0,0,0,87,0,167,0,210,0,0,0,251,0,68,0,204,0,152,0,40,0,131,0,70,0,94,0,9,0,19,0,119,0,33,0,253,0,69,0,253,0,0,0,0,0,0,0,225,0,12,0,221,0,153,0,230,0,88,0,185,0,25,0,0,0,47,0,0,0,42,0,189,0,21,0,0,0,0,0,232,0,138,0,187,0,241,0,29,0,183,0,0,0,6,0,99,0,3,0,90,0,76,0,36,0,183,0,142,0,238,0,100,0,6,0,250,0,239,0,0,0,0,0,107,0,185,0,163,0,137,0,0,0,176,0,77,0,241,0,36,0,59,0,194,0,45,0,243,0,220,0,159,0,150,0,82,0,0,0,207,0,147,0,0,0,0,0,145,0,0,0,32,0,224,0,0,0,249,0,207,0,0,0,81,0,33,0,160,0,237,0,215,0,74,0,132,0,179,0,218,0,167,0,151,0,181,0,28,0,215,0,237,0,160,0,219,0,191,0,228,0,190,0,164,0,103,0,202,0,1,0,0,0,2,0,64,0,118,0,0,0,0,0,250,0,113,0,211,0,24,0,146,0,97,0,1,0,188,0,0,0,77,0,43,0,188,0,237,0,129,0,192,0,83,0,160,0,165,0,173,0,128,0,152,0,75,0,0,0,103,0,0,0,41,0,143,0,208,0,94,0,229,0,19,0,228,0,234,0,95,0,194,0,82,0,117,0,231,0,108,0,112,0,88,0,0,0,0,0,152,0,163,0,137,0,0,0,251,0,155,0,57,0,47,0,235,0,179,0,0,0,169,0,94,0,94,0,111,0,89,0,219,0,252,0,247,0,160,0,0,0,155,0,191,0,32,0,193,0,65,0,219,0,71,0,0,0,0,0,132,0,251,0,202,0,80,0,0,0,232,0,185,0,0,0,50,0,25,0,0,0,0,0,30,0,41,0,0,0,247,0,129,0,249,0,121,0,146,0,153,0,0,0,88,0,0,0,90,0,0,0,3,0,150,0,83,0,114,0,45,0,75,0,0,0,0,0,85,0,157,0,245,0,138,0,0,0,39,0,0,0,173,0,0,0,195,0,0,0,105,0,97,0,216,0,0,0,169,0,105,0,113,0,135,0,140,0,231,0,0,0,72,0,26,0,159,0,0,0,193,0,172,0,112,0,237,0,48,0,145,0,45,0,145,0,223,0,70,0,79,0,156,0,0,0,0,0,135,0,251,0,67,0,130,0,96,0,89,0,248,0,123,0,232,0,46,0,0,0,67,0,40,0,62,0,0,0,144,0,0,0,192,0,156,0,242,0,0,0,23,0,21,0,0,0,87,0,0,0,201,0,216,0,251,0,136,0,133,0,12,0,39,0,112,0,242,0,234,0,6,0,171,0,1,0,185,0,92,0,0,0,111,0,110,0,19,0,0,0,0,0,8,0,0,0,131,0,44,0,246,0,79,0,98,0,145,0,244,0,44,0,167,0,87,0,72,0,3,0,99,0,247,0,50,0,55,0,100,0,180,0,124,0,208,0,164,0,66,0,106,0,131,0,217,0,223,0,0,0,0,0,0,0,0,0,217,0,102,0,0,0,115,0,169,0,51,0,87,0,225,0,68,0,213,0,0,0,253,0,205,0,23,0,0,0,243,0,152,0,206,0,0,0,222,0,137,0,140,0,77,0,163,0,218,0,0,0,254,0,29,0,184,0,248,0,82,0,0,0,0,0,171,0,63,0,212,0,0,0,0,0,169,0,49,0,0,0,250,0,85,0,198,0,0,0,217,0,0,0,32,0,143,0,62,0,37,0,52,0,155,0,156,0,18,0,215,0,16,0,134,0,123,0,199,0,0,0,39,0,227,0,236,0,0,0,0,0,28,0,239,0,149,0,225,0,106,0,189,0,217,0,28,0,0,0,168,0,149,0,0,0,87,0,0,0,207,0,216,0,223,0,187,0,255,0,209,0,13,0,222,0,0,0,137,0,107,0,49,0,74,0,134,0,51,0,151,0,134,0,209,0,99,0,219,0,133,0,103,0,197,0,31,0,222,0,142,0,174,0,138,0,64,0,34,0,87,0,0,0,214,0,0,0,106,0,211,0,226,0,13,0,199,0,194,0,112,0,0,0,190,0,18,0,10,0,0,0,0,0,0,0,245,0,67,0,0,0,234,0,77,0,0,0,0,0,0,0,153,0,0,0,225,0,182,0,134,0,78,0,33,0,48,0,227,0,198,0,164,0,90,0,0,0,112,0,242,0,30,0,208,0,88,0,167,0,0,0,116,0,0,0,177,0,91,0,12,0,222,0,0,0,0,0,78,0,201,0,133,0,138,0,206,0,0,0,44,0,118,0,0,0,99,0,128,0,216,0,239,0,103,0,95,0,215,0,72,0,130,0,208,0,181,0,64,0,168,0,115,0,0,0,0,0,149,0,117,0,122,0,72,0,0,0,249,0,0,0,0,0,60,0,97,0,243,0,102,0,56,0,91,0,0,0,69,0,222,0,93,0,102,0,197,0,219,0,139,0,140,0,161,0,0,0,235,0,183,0,13,0,176,0,115,0,223,0,127,0,68,0,100,0,223,0,225,0,187,0,0,0,0,0,0,0,241,0,181,0,0,0,197,0,0,0,0,0,0,0,245,0,28,0,156,0,32,0,0,0,111,0,0,0,0,0,96,0,155,0,34,0,0,0,139,0,220,0,172,0,157,0,191,0,52,0,50,0,160,0,220,0,36,0,196,0,188,0,245,0,0,0,58,0,226,0,214,0,173,0,234,0,187,0,75,0,214,0,246,0,212,0,0,0,109,0,0,0,19,0,210,0,227,0,0,0,140,0,242,0);
signal scenario_full  : scenario_type := (62,31,62,30,98,31,98,30,248,31,65,31,129,31,207,31,94,31,26,31,195,31,159,31,221,31,118,31,37,31,203,31,66,31,66,30,178,31,89,31,217,31,53,31,221,31,3,31,44,31,83,31,243,31,37,31,204,31,134,31,228,31,228,30,244,31,140,31,32,31,16,31,16,30,37,31,95,31,218,31,221,31,84,31,163,31,164,31,95,31,95,30,74,31,226,31,255,31,68,31,135,31,166,31,59,31,53,31,111,31,174,31,141,31,188,31,188,30,35,31,49,31,49,30,146,31,102,31,116,31,17,31,17,30,17,29,141,31,174,31,174,30,80,31,80,30,99,31,241,31,241,30,82,31,53,31,124,31,22,31,171,31,210,31,127,31,185,31,107,31,107,30,107,29,107,28,65,31,201,31,201,30,7,31,70,31,70,30,70,29,103,31,103,30,103,29,103,28,60,31,233,31,233,30,233,29,102,31,61,31,125,31,25,31,64,31,18,31,196,31,174,31,12,31,47,31,58,31,131,31,131,30,149,31,241,31,36,31,175,31,172,31,156,31,156,30,119,31,124,31,40,31,41,31,41,30,189,31,189,30,171,31,53,31,110,31,140,31,41,31,241,31,241,30,131,31,164,31,86,31,114,31,21,31,27,31,245,31,140,31,140,30,163,31,221,31,150,31,16,31,30,31,199,31,199,30,87,31,87,30,203,31,165,31,89,31,19,31,228,31,170,31,210,31,24,31,101,31,15,31,219,31,219,30,219,29,61,31,241,31,241,30,241,29,241,28,241,27,126,31,110,31,117,31,117,30,226,31,59,31,201,31,108,31,134,31,254,31,16,31,70,31,38,31,122,31,225,31,208,31,27,31,27,30,135,31,132,31,221,31,78,31,78,30,128,31,142,31,94,31,203,31,87,31,87,30,87,29,64,31,197,31,197,30,112,31,98,31,189,31,189,30,189,29,1,31,28,31,122,31,99,31,11,31,131,31,131,30,81,31,81,30,81,29,87,31,167,31,210,31,210,30,251,31,68,31,204,31,152,31,40,31,131,31,70,31,94,31,9,31,19,31,119,31,33,31,253,31,69,31,253,31,253,30,253,29,253,28,225,31,12,31,221,31,153,31,230,31,88,31,185,31,25,31,25,30,47,31,47,30,42,31,189,31,21,31,21,30,21,29,232,31,138,31,187,31,241,31,29,31,183,31,183,30,6,31,99,31,3,31,90,31,76,31,36,31,183,31,142,31,238,31,100,31,6,31,250,31,239,31,239,30,239,29,107,31,185,31,163,31,137,31,137,30,176,31,77,31,241,31,36,31,59,31,194,31,45,31,243,31,220,31,159,31,150,31,82,31,82,30,207,31,147,31,147,30,147,29,145,31,145,30,32,31,224,31,224,30,249,31,207,31,207,30,81,31,33,31,160,31,237,31,215,31,74,31,132,31,179,31,218,31,167,31,151,31,181,31,28,31,215,31,237,31,160,31,219,31,191,31,228,31,190,31,164,31,103,31,202,31,1,31,1,30,2,31,64,31,118,31,118,30,118,29,250,31,113,31,211,31,24,31,146,31,97,31,1,31,188,31,188,30,77,31,43,31,188,31,237,31,129,31,192,31,83,31,160,31,165,31,173,31,128,31,152,31,75,31,75,30,103,31,103,30,41,31,143,31,208,31,94,31,229,31,19,31,228,31,234,31,95,31,194,31,82,31,117,31,231,31,108,31,112,31,88,31,88,30,88,29,152,31,163,31,137,31,137,30,251,31,155,31,57,31,47,31,235,31,179,31,179,30,169,31,94,31,94,31,111,31,89,31,219,31,252,31,247,31,160,31,160,30,155,31,191,31,32,31,193,31,65,31,219,31,71,31,71,30,71,29,132,31,251,31,202,31,80,31,80,30,232,31,185,31,185,30,50,31,25,31,25,30,25,29,30,31,41,31,41,30,247,31,129,31,249,31,121,31,146,31,153,31,153,30,88,31,88,30,90,31,90,30,3,31,150,31,83,31,114,31,45,31,75,31,75,30,75,29,85,31,157,31,245,31,138,31,138,30,39,31,39,30,173,31,173,30,195,31,195,30,105,31,97,31,216,31,216,30,169,31,105,31,113,31,135,31,140,31,231,31,231,30,72,31,26,31,159,31,159,30,193,31,172,31,112,31,237,31,48,31,145,31,45,31,145,31,223,31,70,31,79,31,156,31,156,30,156,29,135,31,251,31,67,31,130,31,96,31,89,31,248,31,123,31,232,31,46,31,46,30,67,31,40,31,62,31,62,30,144,31,144,30,192,31,156,31,242,31,242,30,23,31,21,31,21,30,87,31,87,30,201,31,216,31,251,31,136,31,133,31,12,31,39,31,112,31,242,31,234,31,6,31,171,31,1,31,185,31,92,31,92,30,111,31,110,31,19,31,19,30,19,29,8,31,8,30,131,31,44,31,246,31,79,31,98,31,145,31,244,31,44,31,167,31,87,31,72,31,3,31,99,31,247,31,50,31,55,31,100,31,180,31,124,31,208,31,164,31,66,31,106,31,131,31,217,31,223,31,223,30,223,29,223,28,223,27,217,31,102,31,102,30,115,31,169,31,51,31,87,31,225,31,68,31,213,31,213,30,253,31,205,31,23,31,23,30,243,31,152,31,206,31,206,30,222,31,137,31,140,31,77,31,163,31,218,31,218,30,254,31,29,31,184,31,248,31,82,31,82,30,82,29,171,31,63,31,212,31,212,30,212,29,169,31,49,31,49,30,250,31,85,31,198,31,198,30,217,31,217,30,32,31,143,31,62,31,37,31,52,31,155,31,156,31,18,31,215,31,16,31,134,31,123,31,199,31,199,30,39,31,227,31,236,31,236,30,236,29,28,31,239,31,149,31,225,31,106,31,189,31,217,31,28,31,28,30,168,31,149,31,149,30,87,31,87,30,207,31,216,31,223,31,187,31,255,31,209,31,13,31,222,31,222,30,137,31,107,31,49,31,74,31,134,31,51,31,151,31,134,31,209,31,99,31,219,31,133,31,103,31,197,31,31,31,222,31,142,31,174,31,138,31,64,31,34,31,87,31,87,30,214,31,214,30,106,31,211,31,226,31,13,31,199,31,194,31,112,31,112,30,190,31,18,31,10,31,10,30,10,29,10,28,245,31,67,31,67,30,234,31,77,31,77,30,77,29,77,28,153,31,153,30,225,31,182,31,134,31,78,31,33,31,48,31,227,31,198,31,164,31,90,31,90,30,112,31,242,31,30,31,208,31,88,31,167,31,167,30,116,31,116,30,177,31,91,31,12,31,222,31,222,30,222,29,78,31,201,31,133,31,138,31,206,31,206,30,44,31,118,31,118,30,99,31,128,31,216,31,239,31,103,31,95,31,215,31,72,31,130,31,208,31,181,31,64,31,168,31,115,31,115,30,115,29,149,31,117,31,122,31,72,31,72,30,249,31,249,30,249,29,60,31,97,31,243,31,102,31,56,31,91,31,91,30,69,31,222,31,93,31,102,31,197,31,219,31,139,31,140,31,161,31,161,30,235,31,183,31,13,31,176,31,115,31,223,31,127,31,68,31,100,31,223,31,225,31,187,31,187,30,187,29,187,28,241,31,181,31,181,30,197,31,197,30,197,29,197,28,245,31,28,31,156,31,32,31,32,30,111,31,111,30,111,29,96,31,155,31,34,31,34,30,139,31,220,31,172,31,157,31,191,31,52,31,50,31,160,31,220,31,36,31,196,31,188,31,245,31,245,30,58,31,226,31,214,31,173,31,234,31,187,31,75,31,214,31,246,31,212,31,212,30,109,31,109,30,19,31,210,31,227,31,227,30,140,31,242,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
