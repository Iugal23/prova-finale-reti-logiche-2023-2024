-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 713;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,51,0,0,0,253,0,163,0,0,0,17,0,0,0,86,0,56,0,122,0,124,0,92,0,0,0,245,0,72,0,0,0,0,0,0,0,0,0,166,0,231,0,125,0,0,0,54,0,45,0,144,0,0,0,77,0,209,0,119,0,77,0,36,0,229,0,176,0,177,0,3,0,52,0,33,0,0,0,169,0,0,0,0,0,2,0,0,0,129,0,12,0,82,0,0,0,36,0,124,0,225,0,202,0,80,0,128,0,0,0,103,0,234,0,108,0,48,0,0,0,22,0,109,0,46,0,115,0,139,0,128,0,160,0,0,0,119,0,110,0,0,0,217,0,207,0,140,0,3,0,106,0,103,0,43,0,108,0,76,0,181,0,0,0,196,0,0,0,215,0,0,0,90,0,156,0,64,0,134,0,0,0,0,0,21,0,122,0,75,0,220,0,23,0,0,0,0,0,248,0,117,0,41,0,227,0,68,0,135,0,199,0,211,0,0,0,66,0,191,0,55,0,198,0,65,0,58,0,93,0,0,0,239,0,10,0,0,0,13,0,230,0,198,0,113,0,0,0,144,0,242,0,43,0,35,0,232,0,0,0,32,0,0,0,57,0,165,0,139,0,145,0,67,0,19,0,94,0,0,0,70,0,146,0,39,0,237,0,92,0,48,0,123,0,241,0,7,0,26,0,0,0,132,0,0,0,187,0,128,0,127,0,183,0,0,0,109,0,4,0,212,0,91,0,205,0,114,0,233,0,0,0,34,0,13,0,243,0,221,0,93,0,50,0,110,0,0,0,0,0,168,0,229,0,233,0,0,0,127,0,177,0,246,0,79,0,217,0,131,0,23,0,26,0,11,0,0,0,107,0,33,0,101,0,214,0,181,0,0,0,84,0,90,0,142,0,0,0,100,0,127,0,0,0,156,0,187,0,0,0,229,0,126,0,7,0,0,0,164,0,99,0,91,0,0,0,67,0,220,0,76,0,158,0,202,0,155,0,75,0,224,0,98,0,221,0,108,0,146,0,22,0,0,0,231,0,105,0,51,0,222,0,209,0,183,0,0,0,0,0,0,0,21,0,0,0,71,0,100,0,216,0,238,0,87,0,26,0,59,0,32,0,178,0,0,0,0,0,148,0,0,0,167,0,176,0,91,0,212,0,0,0,0,0,29,0,31,0,92,0,243,0,176,0,197,0,127,0,132,0,71,0,180,0,0,0,43,0,179,0,186,0,56,0,114,0,0,0,44,0,76,0,33,0,0,0,236,0,171,0,45,0,67,0,227,0,0,0,181,0,27,0,80,0,26,0,205,0,176,0,0,0,137,0,0,0,106,0,133,0,92,0,104,0,103,0,113,0,0,0,113,0,0,0,234,0,0,0,179,0,9,0,0,0,120,0,44,0,125,0,0,0,44,0,203,0,22,0,222,0,0,0,0,0,43,0,184,0,63,0,0,0,27,0,0,0,121,0,11,0,70,0,218,0,47,0,0,0,213,0,97,0,137,0,172,0,92,0,165,0,62,0,30,0,106,0,0,0,119,0,111,0,7,0,150,0,143,0,205,0,124,0,137,0,96,0,113,0,31,0,16,0,0,0,128,0,0,0,0,0,123,0,0,0,0,0,0,0,1,0,184,0,4,0,175,0,51,0,253,0,196,0,13,0,0,0,100,0,39,0,82,0,50,0,203,0,186,0,0,0,90,0,188,0,242,0,66,0,135,0,158,0,163,0,64,0,186,0,187,0,3,0,98,0,17,0,0,0,235,0,44,0,94,0,245,0,51,0,44,0,0,0,212,0,144,0,185,0,104,0,214,0,173,0,89,0,89,0,49,0,29,0,234,0,0,0,79,0,240,0,168,0,137,0,0,0,51,0,140,0,0,0,150,0,67,0,30,0,14,0,17,0,18,0,83,0,82,0,85,0,188,0,172,0,49,0,0,0,169,0,50,0,208,0,155,0,130,0,0,0,77,0,50,0,0,0,191,0,0,0,0,0,53,0,0,0,0,0,0,0,17,0,157,0,0,0,168,0,233,0,87,0,144,0,92,0,185,0,195,0,210,0,198,0,0,0,0,0,64,0,153,0,149,0,0,0,68,0,69,0,0,0,196,0,122,0,80,0,62,0,74,0,0,0,0,0,0,0,14,0,111,0,91,0,0,0,230,0,191,0,0,0,54,0,186,0,34,0,181,0,4,0,154,0,61,0,141,0,0,0,210,0,90,0,0,0,182,0,3,0,192,0,3,0,151,0,0,0,121,0,0,0,5,0,40,0,143,0,33,0,0,0,87,0,175,0,67,0,40,0,52,0,0,0,38,0,128,0,119,0,92,0,55,0,49,0,58,0,196,0,239,0,215,0,50,0,19,0,153,0,206,0,194,0,182,0,5,0,0,0,174,0,15,0,117,0,195,0,20,0,134,0,0,0,177,0,84,0,189,0,0,0,180,0,222,0,178,0,104,0,124,0,26,0,0,0,19,0,212,0,0,0,239,0,0,0,34,0,124,0,121,0,153,0,0,0,135,0,0,0,189,0,117,0,5,0,145,0,0,0,73,0,0,0,182,0,213,0,50,0,157,0,0,0,0,0,84,0,196,0,87,0,0,0,238,0,64,0,222,0,0,0,0,0,0,0,188,0,172,0,190,0,233,0,160,0,113,0,119,0,173,0,0,0,164,0,21,0,148,0,0,0,22,0,175,0,0,0,0,0,153,0,56,0,69,0,0,0,204,0,179,0,161,0,10,0,43,0,84,0,0,0,0,0,77,0,253,0,3,0,77,0,0,0,0,0,250,0,124,0,85,0,127,0,173,0,18,0,182,0,178,0,75,0,165,0,0,0,254,0,206,0,33,0,0,0,0,0,129,0,140,0,160,0,251,0,175,0,67,0,82,0,15,0,44,0,58,0,117,0,137,0,254,0,224,0,226,0,91,0,209,0,161,0,178,0,192,0,234,0,150,0,151,0,166,0,236,0,0,0,53,0,0,0,4,0,134,0,248,0,169,0,136,0,247,0,0,0,42,0,34,0,147,0,107,0,240,0,134,0,185,0,187,0,139,0,0,0,248,0,11,0,170,0,87,0,80,0,188,0,50,0,88,0,116,0,0,0,0,0,130,0,0,0,0,0,120,0,1,0,34,0,52,0,48,0,142,0,132,0,104,0,0,0,209,0,0,0,114,0,97,0,193,0,31,0,227,0,163,0,120,0,0,0);
signal scenario_full  : scenario_type := (83,31,51,31,51,30,253,31,163,31,163,30,17,31,17,30,86,31,56,31,122,31,124,31,92,31,92,30,245,31,72,31,72,30,72,29,72,28,72,27,166,31,231,31,125,31,125,30,54,31,45,31,144,31,144,30,77,31,209,31,119,31,77,31,36,31,229,31,176,31,177,31,3,31,52,31,33,31,33,30,169,31,169,30,169,29,2,31,2,30,129,31,12,31,82,31,82,30,36,31,124,31,225,31,202,31,80,31,128,31,128,30,103,31,234,31,108,31,48,31,48,30,22,31,109,31,46,31,115,31,139,31,128,31,160,31,160,30,119,31,110,31,110,30,217,31,207,31,140,31,3,31,106,31,103,31,43,31,108,31,76,31,181,31,181,30,196,31,196,30,215,31,215,30,90,31,156,31,64,31,134,31,134,30,134,29,21,31,122,31,75,31,220,31,23,31,23,30,23,29,248,31,117,31,41,31,227,31,68,31,135,31,199,31,211,31,211,30,66,31,191,31,55,31,198,31,65,31,58,31,93,31,93,30,239,31,10,31,10,30,13,31,230,31,198,31,113,31,113,30,144,31,242,31,43,31,35,31,232,31,232,30,32,31,32,30,57,31,165,31,139,31,145,31,67,31,19,31,94,31,94,30,70,31,146,31,39,31,237,31,92,31,48,31,123,31,241,31,7,31,26,31,26,30,132,31,132,30,187,31,128,31,127,31,183,31,183,30,109,31,4,31,212,31,91,31,205,31,114,31,233,31,233,30,34,31,13,31,243,31,221,31,93,31,50,31,110,31,110,30,110,29,168,31,229,31,233,31,233,30,127,31,177,31,246,31,79,31,217,31,131,31,23,31,26,31,11,31,11,30,107,31,33,31,101,31,214,31,181,31,181,30,84,31,90,31,142,31,142,30,100,31,127,31,127,30,156,31,187,31,187,30,229,31,126,31,7,31,7,30,164,31,99,31,91,31,91,30,67,31,220,31,76,31,158,31,202,31,155,31,75,31,224,31,98,31,221,31,108,31,146,31,22,31,22,30,231,31,105,31,51,31,222,31,209,31,183,31,183,30,183,29,183,28,21,31,21,30,71,31,100,31,216,31,238,31,87,31,26,31,59,31,32,31,178,31,178,30,178,29,148,31,148,30,167,31,176,31,91,31,212,31,212,30,212,29,29,31,31,31,92,31,243,31,176,31,197,31,127,31,132,31,71,31,180,31,180,30,43,31,179,31,186,31,56,31,114,31,114,30,44,31,76,31,33,31,33,30,236,31,171,31,45,31,67,31,227,31,227,30,181,31,27,31,80,31,26,31,205,31,176,31,176,30,137,31,137,30,106,31,133,31,92,31,104,31,103,31,113,31,113,30,113,31,113,30,234,31,234,30,179,31,9,31,9,30,120,31,44,31,125,31,125,30,44,31,203,31,22,31,222,31,222,30,222,29,43,31,184,31,63,31,63,30,27,31,27,30,121,31,11,31,70,31,218,31,47,31,47,30,213,31,97,31,137,31,172,31,92,31,165,31,62,31,30,31,106,31,106,30,119,31,111,31,7,31,150,31,143,31,205,31,124,31,137,31,96,31,113,31,31,31,16,31,16,30,128,31,128,30,128,29,123,31,123,30,123,29,123,28,1,31,184,31,4,31,175,31,51,31,253,31,196,31,13,31,13,30,100,31,39,31,82,31,50,31,203,31,186,31,186,30,90,31,188,31,242,31,66,31,135,31,158,31,163,31,64,31,186,31,187,31,3,31,98,31,17,31,17,30,235,31,44,31,94,31,245,31,51,31,44,31,44,30,212,31,144,31,185,31,104,31,214,31,173,31,89,31,89,31,49,31,29,31,234,31,234,30,79,31,240,31,168,31,137,31,137,30,51,31,140,31,140,30,150,31,67,31,30,31,14,31,17,31,18,31,83,31,82,31,85,31,188,31,172,31,49,31,49,30,169,31,50,31,208,31,155,31,130,31,130,30,77,31,50,31,50,30,191,31,191,30,191,29,53,31,53,30,53,29,53,28,17,31,157,31,157,30,168,31,233,31,87,31,144,31,92,31,185,31,195,31,210,31,198,31,198,30,198,29,64,31,153,31,149,31,149,30,68,31,69,31,69,30,196,31,122,31,80,31,62,31,74,31,74,30,74,29,74,28,14,31,111,31,91,31,91,30,230,31,191,31,191,30,54,31,186,31,34,31,181,31,4,31,154,31,61,31,141,31,141,30,210,31,90,31,90,30,182,31,3,31,192,31,3,31,151,31,151,30,121,31,121,30,5,31,40,31,143,31,33,31,33,30,87,31,175,31,67,31,40,31,52,31,52,30,38,31,128,31,119,31,92,31,55,31,49,31,58,31,196,31,239,31,215,31,50,31,19,31,153,31,206,31,194,31,182,31,5,31,5,30,174,31,15,31,117,31,195,31,20,31,134,31,134,30,177,31,84,31,189,31,189,30,180,31,222,31,178,31,104,31,124,31,26,31,26,30,19,31,212,31,212,30,239,31,239,30,34,31,124,31,121,31,153,31,153,30,135,31,135,30,189,31,117,31,5,31,145,31,145,30,73,31,73,30,182,31,213,31,50,31,157,31,157,30,157,29,84,31,196,31,87,31,87,30,238,31,64,31,222,31,222,30,222,29,222,28,188,31,172,31,190,31,233,31,160,31,113,31,119,31,173,31,173,30,164,31,21,31,148,31,148,30,22,31,175,31,175,30,175,29,153,31,56,31,69,31,69,30,204,31,179,31,161,31,10,31,43,31,84,31,84,30,84,29,77,31,253,31,3,31,77,31,77,30,77,29,250,31,124,31,85,31,127,31,173,31,18,31,182,31,178,31,75,31,165,31,165,30,254,31,206,31,33,31,33,30,33,29,129,31,140,31,160,31,251,31,175,31,67,31,82,31,15,31,44,31,58,31,117,31,137,31,254,31,224,31,226,31,91,31,209,31,161,31,178,31,192,31,234,31,150,31,151,31,166,31,236,31,236,30,53,31,53,30,4,31,134,31,248,31,169,31,136,31,247,31,247,30,42,31,34,31,147,31,107,31,240,31,134,31,185,31,187,31,139,31,139,30,248,31,11,31,170,31,87,31,80,31,188,31,50,31,88,31,116,31,116,30,116,29,130,31,130,30,130,29,120,31,1,31,34,31,52,31,48,31,142,31,132,31,104,31,104,30,209,31,209,30,114,31,97,31,193,31,31,31,227,31,163,31,120,31,120,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
