-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 688;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,95,0,98,0,0,0,241,0,0,0,200,0,23,0,78,0,60,0,153,0,110,0,0,0,0,0,0,0,0,0,78,0,0,0,51,0,32,0,0,0,0,0,63,0,0,0,0,0,0,0,254,0,13,0,252,0,222,0,0,0,167,0,255,0,0,0,0,0,104,0,202,0,115,0,0,0,29,0,0,0,86,0,246,0,226,0,0,0,255,0,133,0,138,0,80,0,0,0,134,0,61,0,148,0,244,0,89,0,0,0,0,0,155,0,2,0,0,0,194,0,105,0,160,0,125,0,0,0,177,0,171,0,193,0,0,0,0,0,122,0,0,0,209,0,230,0,205,0,171,0,0,0,0,0,104,0,137,0,56,0,182,0,0,0,209,0,116,0,0,0,130,0,255,0,0,0,2,0,0,0,108,0,124,0,132,0,58,0,0,0,1,0,0,0,0,0,171,0,243,0,85,0,188,0,58,0,0,0,229,0,103,0,0,0,0,0,120,0,125,0,222,0,0,0,238,0,250,0,241,0,79,0,103,0,153,0,187,0,76,0,133,0,236,0,12,0,61,0,120,0,164,0,213,0,125,0,66,0,144,0,197,0,233,0,139,0,182,0,89,0,174,0,109,0,41,0,0,0,42,0,156,0,146,0,142,0,30,0,40,0,193,0,195,0,104,0,14,0,247,0,197,0,114,0,247,0,111,0,174,0,74,0,0,0,166,0,14,0,37,0,203,0,0,0,101,0,193,0,0,0,158,0,110,0,92,0,48,0,241,0,0,0,234,0,255,0,0,0,167,0,138,0,142,0,249,0,139,0,0,0,190,0,116,0,120,0,0,0,213,0,56,0,123,0,39,0,52,0,170,0,242,0,0,0,8,0,0,0,29,0,200,0,0,0,0,0,28,0,180,0,27,0,17,0,0,0,0,0,0,0,156,0,0,0,35,0,210,0,0,0,42,0,0,0,43,0,148,0,145,0,230,0,35,0,223,0,0,0,130,0,71,0,84,0,136,0,44,0,31,0,0,0,248,0,135,0,117,0,230,0,0,0,27,0,123,0,208,0,20,0,122,0,171,0,238,0,148,0,0,0,218,0,238,0,220,0,224,0,0,0,143,0,0,0,113,0,86,0,20,0,0,0,0,0,13,0,0,0,170,0,64,0,107,0,221,0,225,0,193,0,147,0,74,0,158,0,58,0,236,0,104,0,73,0,175,0,170,0,44,0,134,0,253,0,147,0,0,0,127,0,0,0,8,0,169,0,200,0,240,0,0,0,186,0,43,0,0,0,80,0,0,0,19,0,101,0,96,0,134,0,91,0,0,0,186,0,28,0,0,0,3,0,60,0,248,0,159,0,0,0,181,0,42,0,0,0,169,0,252,0,0,0,0,0,64,0,234,0,146,0,161,0,163,0,144,0,132,0,211,0,0,0,196,0,110,0,154,0,0,0,169,0,8,0,0,0,128,0,0,0,129,0,0,0,9,0,172,0,74,0,113,0,217,0,140,0,219,0,190,0,0,0,2,0,161,0,69,0,122,0,0,0,223,0,45,0,208,0,165,0,206,0,147,0,201,0,141,0,254,0,185,0,39,0,40,0,233,0,218,0,110,0,125,0,0,0,0,0,177,0,232,0,69,0,3,0,47,0,75,0,0,0,16,0,182,0,133,0,208,0,120,0,246,0,0,0,10,0,22,0,36,0,0,0,113,0,0,0,0,0,37,0,193,0,184,0,250,0,69,0,195,0,10,0,237,0,0,0,34,0,185,0,46,0,227,0,147,0,147,0,244,0,0,0,0,0,151,0,77,0,59,0,146,0,126,0,7,0,89,0,49,0,187,0,181,0,152,0,19,0,253,0,47,0,218,0,105,0,2,0,215,0,107,0,91,0,242,0,235,0,0,0,0,0,104,0,178,0,0,0,209,0,0,0,157,0,93,0,0,0,186,0,48,0,39,0,170,0,131,0,139,0,220,0,45,0,138,0,67,0,0,0,215,0,198,0,90,0,105,0,112,0,0,0,60,0,14,0,0,0,63,0,177,0,0,0,6,0,104,0,96,0,140,0,210,0,55,0,119,0,56,0,151,0,216,0,70,0,145,0,0,0,181,0,114,0,0,0,0,0,44,0,0,0,56,0,112,0,163,0,76,0,117,0,121,0,88,0,58,0,122,0,60,0,211,0,84,0,0,0,105,0,25,0,69,0,133,0,104,0,87,0,127,0,241,0,235,0,211,0,74,0,0,0,0,0,171,0,21,0,182,0,126,0,80,0,93,0,251,0,0,0,0,0,140,0,83,0,127,0,186,0,65,0,0,0,221,0,46,0,96,0,33,0,112,0,84,0,215,0,0,0,27,0,0,0,95,0,106,0,170,0,196,0,0,0,178,0,17,0,0,0,0,0,160,0,235,0,241,0,108,0,67,0,0,0,21,0,170,0,191,0,147,0,0,0,140,0,204,0,211,0,114,0,124,0,30,0,124,0,49,0,95,0,87,0,0,0,253,0,145,0,152,0,200,0,78,0,189,0,7,0,241,0,247,0,0,0,31,0,216,0,0,0,175,0,123,0,57,0,110,0,82,0,67,0,0,0,212,0,20,0,191,0,0,0,240,0,75,0,192,0,0,0,127,0,70,0,160,0,82,0,34,0,151,0,162,0,76,0,64,0,242,0,187,0,172,0,154,0,0,0,61,0,0,0,41,0,254,0,0,0,77,0,122,0,78,0,219,0,4,0,42,0,115,0,49,0,218,0,25,0,161,0,212,0,111,0,198,0,108,0,0,0,8,0,0,0,10,0,158,0,175,0,29,0,191,0,126,0,100,0,132,0,41,0,210,0,213,0,63,0,0,0,18,0,56,0,206,0,238,0,120,0,213,0,162,0,34,0,36,0,137,0,116,0,30,0,24,0,38,0,194,0,0,0,53,0,28,0,130,0,148,0,33,0,202,0,0,0,32,0,52,0,94,0,0,0,79,0,57,0,0,0,162,0,126,0,144,0,203,0,117,0,233,0,97,0,220,0,196,0,39,0,217,0,0,0,0,0,0,0,0,0,189,0,255,0,0,0,19,0,26,0,97,0,53,0,137,0,171,0,0,0);
signal scenario_full  : scenario_type := (0,0,95,31,98,31,98,30,241,31,241,30,200,31,23,31,78,31,60,31,153,31,110,31,110,30,110,29,110,28,110,27,78,31,78,30,51,31,32,31,32,30,32,29,63,31,63,30,63,29,63,28,254,31,13,31,252,31,222,31,222,30,167,31,255,31,255,30,255,29,104,31,202,31,115,31,115,30,29,31,29,30,86,31,246,31,226,31,226,30,255,31,133,31,138,31,80,31,80,30,134,31,61,31,148,31,244,31,89,31,89,30,89,29,155,31,2,31,2,30,194,31,105,31,160,31,125,31,125,30,177,31,171,31,193,31,193,30,193,29,122,31,122,30,209,31,230,31,205,31,171,31,171,30,171,29,104,31,137,31,56,31,182,31,182,30,209,31,116,31,116,30,130,31,255,31,255,30,2,31,2,30,108,31,124,31,132,31,58,31,58,30,1,31,1,30,1,29,171,31,243,31,85,31,188,31,58,31,58,30,229,31,103,31,103,30,103,29,120,31,125,31,222,31,222,30,238,31,250,31,241,31,79,31,103,31,153,31,187,31,76,31,133,31,236,31,12,31,61,31,120,31,164,31,213,31,125,31,66,31,144,31,197,31,233,31,139,31,182,31,89,31,174,31,109,31,41,31,41,30,42,31,156,31,146,31,142,31,30,31,40,31,193,31,195,31,104,31,14,31,247,31,197,31,114,31,247,31,111,31,174,31,74,31,74,30,166,31,14,31,37,31,203,31,203,30,101,31,193,31,193,30,158,31,110,31,92,31,48,31,241,31,241,30,234,31,255,31,255,30,167,31,138,31,142,31,249,31,139,31,139,30,190,31,116,31,120,31,120,30,213,31,56,31,123,31,39,31,52,31,170,31,242,31,242,30,8,31,8,30,29,31,200,31,200,30,200,29,28,31,180,31,27,31,17,31,17,30,17,29,17,28,156,31,156,30,35,31,210,31,210,30,42,31,42,30,43,31,148,31,145,31,230,31,35,31,223,31,223,30,130,31,71,31,84,31,136,31,44,31,31,31,31,30,248,31,135,31,117,31,230,31,230,30,27,31,123,31,208,31,20,31,122,31,171,31,238,31,148,31,148,30,218,31,238,31,220,31,224,31,224,30,143,31,143,30,113,31,86,31,20,31,20,30,20,29,13,31,13,30,170,31,64,31,107,31,221,31,225,31,193,31,147,31,74,31,158,31,58,31,236,31,104,31,73,31,175,31,170,31,44,31,134,31,253,31,147,31,147,30,127,31,127,30,8,31,169,31,200,31,240,31,240,30,186,31,43,31,43,30,80,31,80,30,19,31,101,31,96,31,134,31,91,31,91,30,186,31,28,31,28,30,3,31,60,31,248,31,159,31,159,30,181,31,42,31,42,30,169,31,252,31,252,30,252,29,64,31,234,31,146,31,161,31,163,31,144,31,132,31,211,31,211,30,196,31,110,31,154,31,154,30,169,31,8,31,8,30,128,31,128,30,129,31,129,30,9,31,172,31,74,31,113,31,217,31,140,31,219,31,190,31,190,30,2,31,161,31,69,31,122,31,122,30,223,31,45,31,208,31,165,31,206,31,147,31,201,31,141,31,254,31,185,31,39,31,40,31,233,31,218,31,110,31,125,31,125,30,125,29,177,31,232,31,69,31,3,31,47,31,75,31,75,30,16,31,182,31,133,31,208,31,120,31,246,31,246,30,10,31,22,31,36,31,36,30,113,31,113,30,113,29,37,31,193,31,184,31,250,31,69,31,195,31,10,31,237,31,237,30,34,31,185,31,46,31,227,31,147,31,147,31,244,31,244,30,244,29,151,31,77,31,59,31,146,31,126,31,7,31,89,31,49,31,187,31,181,31,152,31,19,31,253,31,47,31,218,31,105,31,2,31,215,31,107,31,91,31,242,31,235,31,235,30,235,29,104,31,178,31,178,30,209,31,209,30,157,31,93,31,93,30,186,31,48,31,39,31,170,31,131,31,139,31,220,31,45,31,138,31,67,31,67,30,215,31,198,31,90,31,105,31,112,31,112,30,60,31,14,31,14,30,63,31,177,31,177,30,6,31,104,31,96,31,140,31,210,31,55,31,119,31,56,31,151,31,216,31,70,31,145,31,145,30,181,31,114,31,114,30,114,29,44,31,44,30,56,31,112,31,163,31,76,31,117,31,121,31,88,31,58,31,122,31,60,31,211,31,84,31,84,30,105,31,25,31,69,31,133,31,104,31,87,31,127,31,241,31,235,31,211,31,74,31,74,30,74,29,171,31,21,31,182,31,126,31,80,31,93,31,251,31,251,30,251,29,140,31,83,31,127,31,186,31,65,31,65,30,221,31,46,31,96,31,33,31,112,31,84,31,215,31,215,30,27,31,27,30,95,31,106,31,170,31,196,31,196,30,178,31,17,31,17,30,17,29,160,31,235,31,241,31,108,31,67,31,67,30,21,31,170,31,191,31,147,31,147,30,140,31,204,31,211,31,114,31,124,31,30,31,124,31,49,31,95,31,87,31,87,30,253,31,145,31,152,31,200,31,78,31,189,31,7,31,241,31,247,31,247,30,31,31,216,31,216,30,175,31,123,31,57,31,110,31,82,31,67,31,67,30,212,31,20,31,191,31,191,30,240,31,75,31,192,31,192,30,127,31,70,31,160,31,82,31,34,31,151,31,162,31,76,31,64,31,242,31,187,31,172,31,154,31,154,30,61,31,61,30,41,31,254,31,254,30,77,31,122,31,78,31,219,31,4,31,42,31,115,31,49,31,218,31,25,31,161,31,212,31,111,31,198,31,108,31,108,30,8,31,8,30,10,31,158,31,175,31,29,31,191,31,126,31,100,31,132,31,41,31,210,31,213,31,63,31,63,30,18,31,56,31,206,31,238,31,120,31,213,31,162,31,34,31,36,31,137,31,116,31,30,31,24,31,38,31,194,31,194,30,53,31,28,31,130,31,148,31,33,31,202,31,202,30,32,31,52,31,94,31,94,30,79,31,57,31,57,30,162,31,126,31,144,31,203,31,117,31,233,31,97,31,220,31,196,31,39,31,217,31,217,30,217,29,217,28,217,27,189,31,255,31,255,30,19,31,26,31,97,31,53,31,137,31,171,31,171,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
