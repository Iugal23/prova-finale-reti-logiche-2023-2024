-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_425 is
end project_tb_425;

architecture project_tb_arch_425 of project_tb_425 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 684;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,48,0,0,0,135,0,0,0,195,0,135,0,175,0,189,0,0,0,28,0,202,0,40,0,40,0,47,0,0,0,126,0,29,0,0,0,0,0,0,0,122,0,81,0,121,0,148,0,194,0,204,0,108,0,231,0,66,0,211,0,3,0,0,0,0,0,0,0,73,0,226,0,80,0,207,0,98,0,195,0,119,0,38,0,144,0,128,0,0,0,0,0,128,0,81,0,70,0,0,0,121,0,0,0,56,0,5,0,159,0,168,0,227,0,168,0,83,0,206,0,202,0,211,0,84,0,178,0,220,0,0,0,117,0,0,0,49,0,0,0,0,0,98,0,80,0,0,0,254,0,0,0,0,0,169,0,0,0,24,0,0,0,120,0,167,0,95,0,108,0,0,0,64,0,80,0,32,0,249,0,219,0,213,0,59,0,54,0,195,0,231,0,135,0,82,0,0,0,78,0,99,0,20,0,74,0,187,0,0,0,250,0,0,0,139,0,0,0,98,0,239,0,46,0,0,0,0,0,0,0,67,0,250,0,189,0,27,0,177,0,179,0,59,0,0,0,0,0,0,0,141,0,203,0,89,0,14,0,246,0,0,0,239,0,107,0,45,0,0,0,61,0,84,0,33,0,87,0,144,0,0,0,214,0,0,0,96,0,215,0,0,0,218,0,202,0,154,0,62,0,156,0,137,0,60,0,226,0,0,0,81,0,89,0,242,0,0,0,111,0,40,0,40,0,0,0,86,0,135,0,219,0,182,0,2,0,12,0,1,0,211,0,0,0,158,0,179,0,0,0,236,0,165,0,162,0,96,0,33,0,186,0,0,0,12,0,0,0,240,0,18,0,105,0,163,0,251,0,0,0,245,0,217,0,54,0,0,0,55,0,0,0,88,0,33,0,250,0,184,0,124,0,210,0,14,0,4,0,182,0,0,0,1,0,189,0,0,0,0,0,157,0,26,0,28,0,91,0,18,0,203,0,190,0,134,0,20,0,246,0,232,0,177,0,0,0,245,0,226,0,2,0,0,0,103,0,61,0,205,0,245,0,4,0,79,0,252,0,166,0,146,0,245,0,149,0,0,0,185,0,239,0,31,0,220,0,0,0,229,0,53,0,117,0,0,0,11,0,0,0,38,0,159,0,62,0,251,0,0,0,128,0,179,0,59,0,0,0,27,0,157,0,117,0,71,0,90,0,199,0,118,0,39,0,250,0,25,0,35,0,124,0,121,0,87,0,168,0,133,0,0,0,202,0,0,0,0,0,74,0,16,0,149,0,40,0,255,0,143,0,33,0,0,0,0,0,0,0,230,0,49,0,189,0,158,0,169,0,0,0,133,0,0,0,168,0,6,0,77,0,149,0,67,0,246,0,20,0,210,0,158,0,118,0,0,0,0,0,96,0,0,0,151,0,0,0,0,0,0,0,4,0,65,0,200,0,89,0,118,0,0,0,205,0,152,0,2,0,4,0,247,0,230,0,0,0,193,0,66,0,0,0,0,0,179,0,204,0,94,0,221,0,190,0,169,0,0,0,0,0,0,0,141,0,211,0,61,0,62,0,118,0,69,0,53,0,201,0,102,0,65,0,217,0,33,0,24,0,173,0,100,0,142,0,65,0,66,0,224,0,62,0,49,0,85,0,0,0,154,0,95,0,147,0,110,0,209,0,0,0,0,0,0,0,14,0,0,0,239,0,239,0,142,0,211,0,217,0,0,0,0,0,178,0,115,0,141,0,23,0,131,0,0,0,187,0,53,0,0,0,73,0,81,0,250,0,0,0,90,0,0,0,0,0,159,0,0,0,178,0,123,0,132,0,190,0,52,0,58,0,70,0,26,0,0,0,35,0,137,0,250,0,183,0,151,0,166,0,211,0,222,0,0,0,111,0,88,0,16,0,153,0,0,0,33,0,0,0,0,0,87,0,37,0,133,0,0,0,220,0,0,0,0,0,56,0,13,0,217,0,0,0,103,0,206,0,85,0,47,0,0,0,126,0,167,0,162,0,107,0,187,0,109,0,52,0,219,0,228,0,0,0,114,0,0,0,133,0,0,0,71,0,165,0,0,0,46,0,195,0,0,0,251,0,101,0,227,0,221,0,93,0,7,0,252,0,234,0,0,0,140,0,94,0,0,0,82,0,0,0,142,0,52,0,164,0,61,0,206,0,93,0,125,0,0,0,85,0,0,0,0,0,216,0,42,0,37,0,211,0,18,0,97,0,243,0,22,0,0,0,150,0,234,0,168,0,0,0,232,0,108,0,127,0,0,0,254,0,8,0,67,0,184,0,0,0,177,0,161,0,84,0,109,0,206,0,203,0,62,0,101,0,72,0,239,0,0,0,86,0,136,0,254,0,0,0,34,0,240,0,88,0,225,0,80,0,181,0,79,0,112,0,56,0,11,0,203,0,247,0,8,0,147,0,85,0,67,0,65,0,0,0,40,0,0,0,86,0,245,0,87,0,170,0,48,0,0,0,170,0,242,0,70,0,3,0,0,0,163,0,7,0,242,0,34,0,63,0,213,0,247,0,7,0,242,0,189,0,184,0,64,0,0,0,160,0,179,0,184,0,95,0,203,0,76,0,30,0,205,0,146,0,205,0,207,0,226,0,0,0,241,0,209,0,26,0,138,0,84,0,220,0,0,0,107,0,115,0,0,0,0,0,193,0,247,0,201,0,236,0,129,0,175,0,227,0,178,0,0,0,190,0,66,0,129,0,55,0,218,0,133,0,67,0,235,0,245,0,113,0,233,0,0,0,244,0,0,0,116,0,175,0,229,0,247,0,128,0,228,0,59,0,86,0,10,0,130,0,0,0,83,0,49,0,29,0,243,0,0,0,11,0,83,0,123,0,60,0,22,0,62,0,95,0,114,0,6,0,4,0,68,0,0,0,72,0,24,0,62,0,0,0,226,0,205,0,208,0,0,0,0,0,183,0,15,0,116,0,168,0,85,0,199,0,179,0,173,0,25,0,0,0,57,0,0,0,172,0,0,0,0,0,208,0,178,0,0,0,0,0,122,0,174,0,111,0,21,0,0,0,114,0,0,0,0,0,28,0,164,0,31,0,41,0,32,0);
signal scenario_full  : scenario_type := (0,0,48,31,48,30,135,31,135,30,195,31,135,31,175,31,189,31,189,30,28,31,202,31,40,31,40,31,47,31,47,30,126,31,29,31,29,30,29,29,29,28,122,31,81,31,121,31,148,31,194,31,204,31,108,31,231,31,66,31,211,31,3,31,3,30,3,29,3,28,73,31,226,31,80,31,207,31,98,31,195,31,119,31,38,31,144,31,128,31,128,30,128,29,128,31,81,31,70,31,70,30,121,31,121,30,56,31,5,31,159,31,168,31,227,31,168,31,83,31,206,31,202,31,211,31,84,31,178,31,220,31,220,30,117,31,117,30,49,31,49,30,49,29,98,31,80,31,80,30,254,31,254,30,254,29,169,31,169,30,24,31,24,30,120,31,167,31,95,31,108,31,108,30,64,31,80,31,32,31,249,31,219,31,213,31,59,31,54,31,195,31,231,31,135,31,82,31,82,30,78,31,99,31,20,31,74,31,187,31,187,30,250,31,250,30,139,31,139,30,98,31,239,31,46,31,46,30,46,29,46,28,67,31,250,31,189,31,27,31,177,31,179,31,59,31,59,30,59,29,59,28,141,31,203,31,89,31,14,31,246,31,246,30,239,31,107,31,45,31,45,30,61,31,84,31,33,31,87,31,144,31,144,30,214,31,214,30,96,31,215,31,215,30,218,31,202,31,154,31,62,31,156,31,137,31,60,31,226,31,226,30,81,31,89,31,242,31,242,30,111,31,40,31,40,31,40,30,86,31,135,31,219,31,182,31,2,31,12,31,1,31,211,31,211,30,158,31,179,31,179,30,236,31,165,31,162,31,96,31,33,31,186,31,186,30,12,31,12,30,240,31,18,31,105,31,163,31,251,31,251,30,245,31,217,31,54,31,54,30,55,31,55,30,88,31,33,31,250,31,184,31,124,31,210,31,14,31,4,31,182,31,182,30,1,31,189,31,189,30,189,29,157,31,26,31,28,31,91,31,18,31,203,31,190,31,134,31,20,31,246,31,232,31,177,31,177,30,245,31,226,31,2,31,2,30,103,31,61,31,205,31,245,31,4,31,79,31,252,31,166,31,146,31,245,31,149,31,149,30,185,31,239,31,31,31,220,31,220,30,229,31,53,31,117,31,117,30,11,31,11,30,38,31,159,31,62,31,251,31,251,30,128,31,179,31,59,31,59,30,27,31,157,31,117,31,71,31,90,31,199,31,118,31,39,31,250,31,25,31,35,31,124,31,121,31,87,31,168,31,133,31,133,30,202,31,202,30,202,29,74,31,16,31,149,31,40,31,255,31,143,31,33,31,33,30,33,29,33,28,230,31,49,31,189,31,158,31,169,31,169,30,133,31,133,30,168,31,6,31,77,31,149,31,67,31,246,31,20,31,210,31,158,31,118,31,118,30,118,29,96,31,96,30,151,31,151,30,151,29,151,28,4,31,65,31,200,31,89,31,118,31,118,30,205,31,152,31,2,31,4,31,247,31,230,31,230,30,193,31,66,31,66,30,66,29,179,31,204,31,94,31,221,31,190,31,169,31,169,30,169,29,169,28,141,31,211,31,61,31,62,31,118,31,69,31,53,31,201,31,102,31,65,31,217,31,33,31,24,31,173,31,100,31,142,31,65,31,66,31,224,31,62,31,49,31,85,31,85,30,154,31,95,31,147,31,110,31,209,31,209,30,209,29,209,28,14,31,14,30,239,31,239,31,142,31,211,31,217,31,217,30,217,29,178,31,115,31,141,31,23,31,131,31,131,30,187,31,53,31,53,30,73,31,81,31,250,31,250,30,90,31,90,30,90,29,159,31,159,30,178,31,123,31,132,31,190,31,52,31,58,31,70,31,26,31,26,30,35,31,137,31,250,31,183,31,151,31,166,31,211,31,222,31,222,30,111,31,88,31,16,31,153,31,153,30,33,31,33,30,33,29,87,31,37,31,133,31,133,30,220,31,220,30,220,29,56,31,13,31,217,31,217,30,103,31,206,31,85,31,47,31,47,30,126,31,167,31,162,31,107,31,187,31,109,31,52,31,219,31,228,31,228,30,114,31,114,30,133,31,133,30,71,31,165,31,165,30,46,31,195,31,195,30,251,31,101,31,227,31,221,31,93,31,7,31,252,31,234,31,234,30,140,31,94,31,94,30,82,31,82,30,142,31,52,31,164,31,61,31,206,31,93,31,125,31,125,30,85,31,85,30,85,29,216,31,42,31,37,31,211,31,18,31,97,31,243,31,22,31,22,30,150,31,234,31,168,31,168,30,232,31,108,31,127,31,127,30,254,31,8,31,67,31,184,31,184,30,177,31,161,31,84,31,109,31,206,31,203,31,62,31,101,31,72,31,239,31,239,30,86,31,136,31,254,31,254,30,34,31,240,31,88,31,225,31,80,31,181,31,79,31,112,31,56,31,11,31,203,31,247,31,8,31,147,31,85,31,67,31,65,31,65,30,40,31,40,30,86,31,245,31,87,31,170,31,48,31,48,30,170,31,242,31,70,31,3,31,3,30,163,31,7,31,242,31,34,31,63,31,213,31,247,31,7,31,242,31,189,31,184,31,64,31,64,30,160,31,179,31,184,31,95,31,203,31,76,31,30,31,205,31,146,31,205,31,207,31,226,31,226,30,241,31,209,31,26,31,138,31,84,31,220,31,220,30,107,31,115,31,115,30,115,29,193,31,247,31,201,31,236,31,129,31,175,31,227,31,178,31,178,30,190,31,66,31,129,31,55,31,218,31,133,31,67,31,235,31,245,31,113,31,233,31,233,30,244,31,244,30,116,31,175,31,229,31,247,31,128,31,228,31,59,31,86,31,10,31,130,31,130,30,83,31,49,31,29,31,243,31,243,30,11,31,83,31,123,31,60,31,22,31,62,31,95,31,114,31,6,31,4,31,68,31,68,30,72,31,24,31,62,31,62,30,226,31,205,31,208,31,208,30,208,29,183,31,15,31,116,31,168,31,85,31,199,31,179,31,173,31,25,31,25,30,57,31,57,30,172,31,172,30,172,29,208,31,178,31,178,30,178,29,122,31,174,31,111,31,21,31,21,30,114,31,114,30,114,29,28,31,164,31,31,31,41,31,32,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
