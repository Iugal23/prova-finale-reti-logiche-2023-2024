-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 687;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (145,0,89,0,0,0,192,0,47,0,165,0,100,0,59,0,142,0,0,0,115,0,140,0,70,0,140,0,8,0,222,0,120,0,200,0,112,0,161,0,137,0,36,0,229,0,153,0,238,0,224,0,229,0,57,0,237,0,228,0,79,0,103,0,171,0,222,0,174,0,176,0,111,0,253,0,176,0,230,0,51,0,1,0,176,0,230,0,39,0,246,0,233,0,0,0,207,0,245,0,0,0,150,0,252,0,241,0,20,0,248,0,160,0,139,0,117,0,103,0,84,0,148,0,0,0,200,0,234,0,143,0,0,0,251,0,83,0,53,0,80,0,209,0,165,0,0,0,63,0,52,0,253,0,183,0,238,0,118,0,108,0,213,0,156,0,223,0,64,0,37,0,62,0,70,0,0,0,150,0,165,0,168,0,0,0,12,0,184,0,111,0,0,0,24,0,17,0,210,0,20,0,87,0,122,0,0,0,147,0,70,0,150,0,12,0,0,0,246,0,0,0,6,0,57,0,132,0,0,0,0,0,0,0,121,0,0,0,250,0,110,0,0,0,204,0,0,0,233,0,130,0,139,0,184,0,96,0,51,0,0,0,86,0,125,0,29,0,42,0,7,0,0,0,29,0,0,0,146,0,135,0,211,0,187,0,0,0,52,0,23,0,160,0,219,0,0,0,22,0,27,0,226,0,0,0,21,0,0,0,31,0,125,0,234,0,0,0,58,0,91,0,116,0,107,0,151,0,86,0,30,0,193,0,200,0,0,0,0,0,13,0,0,0,183,0,0,0,29,0,32,0,49,0,53,0,149,0,98,0,123,0,0,0,0,0,194,0,39,0,94,0,200,0,106,0,186,0,180,0,152,0,126,0,0,0,0,0,125,0,179,0,29,0,82,0,21,0,38,0,107,0,120,0,0,0,0,0,62,0,0,0,156,0,164,0,43,0,173,0,86,0,66,0,106,0,0,0,27,0,130,0,3,0,0,0,81,0,237,0,51,0,0,0,91,0,232,0,107,0,69,0,28,0,45,0,0,0,205,0,255,0,228,0,0,0,117,0,105,0,123,0,65,0,0,0,3,0,102,0,8,0,19,0,0,0,153,0,235,0,0,0,240,0,56,0,93,0,0,0,8,0,102,0,100,0,234,0,3,0,0,0,184,0,252,0,226,0,236,0,92,0,37,0,5,0,0,0,145,0,213,0,132,0,239,0,16,0,0,0,194,0,0,0,242,0,0,0,0,0,13,0,220,0,99,0,137,0,200,0,99,0,115,0,32,0,134,0,0,0,89,0,31,0,166,0,199,0,248,0,109,0,221,0,28,0,163,0,0,0,172,0,113,0,18,0,158,0,100,0,222,0,172,0,0,0,140,0,114,0,223,0,37,0,4,0,229,0,69,0,59,0,0,0,205,0,3,0,171,0,131,0,119,0,44,0,232,0,246,0,83,0,0,0,216,0,61,0,199,0,0,0,203,0,0,0,202,0,90,0,70,0,111,0,186,0,155,0,127,0,8,0,12,0,133,0,8,0,233,0,109,0,21,0,203,0,203,0,113,0,200,0,0,0,96,0,254,0,213,0,219,0,185,0,218,0,210,0,23,0,239,0,0,0,0,0,63,0,28,0,137,0,232,0,192,0,238,0,0,0,192,0,185,0,137,0,199,0,0,0,0,0,0,0,24,0,0,0,108,0,246,0,38,0,243,0,104,0,39,0,151,0,0,0,15,0,254,0,109,0,216,0,137,0,166,0,246,0,206,0,211,0,94,0,48,0,65,0,173,0,193,0,144,0,31,0,160,0,153,0,54,0,0,0,102,0,0,0,14,0,147,0,176,0,163,0,34,0,143,0,87,0,125,0,0,0,34,0,240,0,121,0,81,0,246,0,109,0,101,0,136,0,215,0,221,0,142,0,243,0,203,0,200,0,214,0,0,0,60,0,171,0,179,0,26,0,26,0,53,0,0,0,243,0,15,0,169,0,233,0,187,0,0,0,0,0,165,0,187,0,0,0,0,0,165,0,135,0,226,0,0,0,188,0,0,0,74,0,0,0,178,0,242,0,132,0,46,0,104,0,0,0,161,0,144,0,0,0,245,0,217,0,53,0,71,0,113,0,168,0,0,0,0,0,0,0,0,0,142,0,192,0,42,0,0,0,232,0,0,0,77,0,160,0,57,0,129,0,0,0,0,0,69,0,0,0,29,0,0,0,0,0,173,0,120,0,47,0,0,0,118,0,0,0,37,0,122,0,234,0,125,0,159,0,150,0,0,0,0,0,173,0,34,0,13,0,239,0,121,0,225,0,0,0,216,0,141,0,0,0,245,0,76,0,103,0,141,0,244,0,0,0,197,0,221,0,0,0,0,0,0,0,127,0,31,0,110,0,50,0,86,0,59,0,22,0,23,0,126,0,0,0,0,0,179,0,158,0,135,0,189,0,34,0,247,0,170,0,0,0,64,0,186,0,0,0,52,0,161,0,2,0,0,0,24,0,221,0,227,0,195,0,220,0,201,0,88,0,168,0,131,0,0,0,35,0,0,0,170,0,222,0,133,0,236,0,54,0,74,0,186,0,111,0,98,0,103,0,0,0,117,0,70,0,229,0,206,0,68,0,165,0,31,0,177,0,159,0,219,0,0,0,153,0,177,0,183,0,94,0,0,0,245,0,56,0,231,0,232,0,211,0,39,0,0,0,126,0,201,0,20,0,248,0,103,0,0,0,0,0,0,0,128,0,15,0,237,0,109,0,0,0,124,0,230,0,0,0,92,0,177,0,0,0,2,0,147,0,0,0,25,0,214,0,244,0,0,0,155,0,0,0,0,0,0,0,199,0,0,0,27,0,190,0,50,0,225,0,211,0,207,0,86,0,117,0,225,0,162,0,0,0,244,0,0,0,199,0,183,0,220,0,62,0,231,0,127,0,173,0,209,0,0,0,137,0,0,0,0,0,101,0,0,0,136,0,245,0,0,0,246,0,0,0,0,0,68,0,0,0,64,0,90,0,21,0,162,0,106,0,205,0,118,0,3,0,170,0,203,0,0,0,0,0,120,0,149,0,0,0,214,0,201,0,117,0,40,0,87,0,0,0,0,0);
signal scenario_full  : scenario_type := (145,31,89,31,89,30,192,31,47,31,165,31,100,31,59,31,142,31,142,30,115,31,140,31,70,31,140,31,8,31,222,31,120,31,200,31,112,31,161,31,137,31,36,31,229,31,153,31,238,31,224,31,229,31,57,31,237,31,228,31,79,31,103,31,171,31,222,31,174,31,176,31,111,31,253,31,176,31,230,31,51,31,1,31,176,31,230,31,39,31,246,31,233,31,233,30,207,31,245,31,245,30,150,31,252,31,241,31,20,31,248,31,160,31,139,31,117,31,103,31,84,31,148,31,148,30,200,31,234,31,143,31,143,30,251,31,83,31,53,31,80,31,209,31,165,31,165,30,63,31,52,31,253,31,183,31,238,31,118,31,108,31,213,31,156,31,223,31,64,31,37,31,62,31,70,31,70,30,150,31,165,31,168,31,168,30,12,31,184,31,111,31,111,30,24,31,17,31,210,31,20,31,87,31,122,31,122,30,147,31,70,31,150,31,12,31,12,30,246,31,246,30,6,31,57,31,132,31,132,30,132,29,132,28,121,31,121,30,250,31,110,31,110,30,204,31,204,30,233,31,130,31,139,31,184,31,96,31,51,31,51,30,86,31,125,31,29,31,42,31,7,31,7,30,29,31,29,30,146,31,135,31,211,31,187,31,187,30,52,31,23,31,160,31,219,31,219,30,22,31,27,31,226,31,226,30,21,31,21,30,31,31,125,31,234,31,234,30,58,31,91,31,116,31,107,31,151,31,86,31,30,31,193,31,200,31,200,30,200,29,13,31,13,30,183,31,183,30,29,31,32,31,49,31,53,31,149,31,98,31,123,31,123,30,123,29,194,31,39,31,94,31,200,31,106,31,186,31,180,31,152,31,126,31,126,30,126,29,125,31,179,31,29,31,82,31,21,31,38,31,107,31,120,31,120,30,120,29,62,31,62,30,156,31,164,31,43,31,173,31,86,31,66,31,106,31,106,30,27,31,130,31,3,31,3,30,81,31,237,31,51,31,51,30,91,31,232,31,107,31,69,31,28,31,45,31,45,30,205,31,255,31,228,31,228,30,117,31,105,31,123,31,65,31,65,30,3,31,102,31,8,31,19,31,19,30,153,31,235,31,235,30,240,31,56,31,93,31,93,30,8,31,102,31,100,31,234,31,3,31,3,30,184,31,252,31,226,31,236,31,92,31,37,31,5,31,5,30,145,31,213,31,132,31,239,31,16,31,16,30,194,31,194,30,242,31,242,30,242,29,13,31,220,31,99,31,137,31,200,31,99,31,115,31,32,31,134,31,134,30,89,31,31,31,166,31,199,31,248,31,109,31,221,31,28,31,163,31,163,30,172,31,113,31,18,31,158,31,100,31,222,31,172,31,172,30,140,31,114,31,223,31,37,31,4,31,229,31,69,31,59,31,59,30,205,31,3,31,171,31,131,31,119,31,44,31,232,31,246,31,83,31,83,30,216,31,61,31,199,31,199,30,203,31,203,30,202,31,90,31,70,31,111,31,186,31,155,31,127,31,8,31,12,31,133,31,8,31,233,31,109,31,21,31,203,31,203,31,113,31,200,31,200,30,96,31,254,31,213,31,219,31,185,31,218,31,210,31,23,31,239,31,239,30,239,29,63,31,28,31,137,31,232,31,192,31,238,31,238,30,192,31,185,31,137,31,199,31,199,30,199,29,199,28,24,31,24,30,108,31,246,31,38,31,243,31,104,31,39,31,151,31,151,30,15,31,254,31,109,31,216,31,137,31,166,31,246,31,206,31,211,31,94,31,48,31,65,31,173,31,193,31,144,31,31,31,160,31,153,31,54,31,54,30,102,31,102,30,14,31,147,31,176,31,163,31,34,31,143,31,87,31,125,31,125,30,34,31,240,31,121,31,81,31,246,31,109,31,101,31,136,31,215,31,221,31,142,31,243,31,203,31,200,31,214,31,214,30,60,31,171,31,179,31,26,31,26,31,53,31,53,30,243,31,15,31,169,31,233,31,187,31,187,30,187,29,165,31,187,31,187,30,187,29,165,31,135,31,226,31,226,30,188,31,188,30,74,31,74,30,178,31,242,31,132,31,46,31,104,31,104,30,161,31,144,31,144,30,245,31,217,31,53,31,71,31,113,31,168,31,168,30,168,29,168,28,168,27,142,31,192,31,42,31,42,30,232,31,232,30,77,31,160,31,57,31,129,31,129,30,129,29,69,31,69,30,29,31,29,30,29,29,173,31,120,31,47,31,47,30,118,31,118,30,37,31,122,31,234,31,125,31,159,31,150,31,150,30,150,29,173,31,34,31,13,31,239,31,121,31,225,31,225,30,216,31,141,31,141,30,245,31,76,31,103,31,141,31,244,31,244,30,197,31,221,31,221,30,221,29,221,28,127,31,31,31,110,31,50,31,86,31,59,31,22,31,23,31,126,31,126,30,126,29,179,31,158,31,135,31,189,31,34,31,247,31,170,31,170,30,64,31,186,31,186,30,52,31,161,31,2,31,2,30,24,31,221,31,227,31,195,31,220,31,201,31,88,31,168,31,131,31,131,30,35,31,35,30,170,31,222,31,133,31,236,31,54,31,74,31,186,31,111,31,98,31,103,31,103,30,117,31,70,31,229,31,206,31,68,31,165,31,31,31,177,31,159,31,219,31,219,30,153,31,177,31,183,31,94,31,94,30,245,31,56,31,231,31,232,31,211,31,39,31,39,30,126,31,201,31,20,31,248,31,103,31,103,30,103,29,103,28,128,31,15,31,237,31,109,31,109,30,124,31,230,31,230,30,92,31,177,31,177,30,2,31,147,31,147,30,25,31,214,31,244,31,244,30,155,31,155,30,155,29,155,28,199,31,199,30,27,31,190,31,50,31,225,31,211,31,207,31,86,31,117,31,225,31,162,31,162,30,244,31,244,30,199,31,183,31,220,31,62,31,231,31,127,31,173,31,209,31,209,30,137,31,137,30,137,29,101,31,101,30,136,31,245,31,245,30,246,31,246,30,246,29,68,31,68,30,64,31,90,31,21,31,162,31,106,31,205,31,118,31,3,31,170,31,203,31,203,30,203,29,120,31,149,31,149,30,214,31,201,31,117,31,40,31,87,31,87,30,87,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
