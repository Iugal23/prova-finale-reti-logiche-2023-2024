-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_941 is
end project_tb_941;

architecture project_tb_arch_941 of project_tb_941 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1018;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,145,0,1,0,112,0,0,0,186,0,182,0,155,0,184,0,176,0,0,0,7,0,240,0,0,0,154,0,169,0,41,0,87,0,34,0,135,0,173,0,0,0,139,0,97,0,0,0,0,0,83,0,19,0,0,0,245,0,147,0,83,0,68,0,38,0,172,0,74,0,251,0,0,0,42,0,222,0,0,0,20,0,227,0,63,0,136,0,234,0,0,0,248,0,0,0,195,0,7,0,178,0,248,0,16,0,0,0,0,0,74,0,210,0,6,0,6,0,90,0,170,0,241,0,0,0,60,0,212,0,210,0,0,0,255,0,44,0,253,0,67,0,105,0,181,0,92,0,121,0,239,0,71,0,186,0,0,0,59,0,178,0,217,0,244,0,77,0,49,0,198,0,192,0,185,0,0,0,148,0,47,0,117,0,119,0,0,0,165,0,188,0,0,0,0,0,174,0,42,0,15,0,0,0,0,0,224,0,0,0,4,0,33,0,30,0,208,0,0,0,0,0,117,0,0,0,253,0,66,0,211,0,200,0,0,0,177,0,127,0,134,0,26,0,120,0,26,0,0,0,95,0,250,0,135,0,247,0,248,0,0,0,137,0,135,0,9,0,250,0,202,0,108,0,224,0,178,0,0,0,236,0,242,0,44,0,177,0,184,0,195,0,121,0,161,0,170,0,164,0,0,0,0,0,78,0,160,0,171,0,155,0,251,0,98,0,230,0,89,0,139,0,48,0,67,0,169,0,141,0,0,0,212,0,0,0,39,0,10,0,109,0,169,0,109,0,19,0,221,0,3,0,0,0,202,0,114,0,0,0,0,0,57,0,30,0,217,0,115,0,33,0,135,0,151,0,180,0,0,0,130,0,1,0,219,0,157,0,250,0,29,0,120,0,126,0,218,0,207,0,25,0,142,0,0,0,0,0,162,0,0,0,154,0,237,0,197,0,0,0,5,0,135,0,26,0,0,0,214,0,32,0,167,0,0,0,249,0,0,0,0,0,171,0,146,0,145,0,143,0,144,0,220,0,194,0,100,0,214,0,163,0,0,0,0,0,233,0,175,0,127,0,0,0,88,0,179,0,217,0,0,0,193,0,208,0,180,0,73,0,15,0,0,0,49,0,21,0,241,0,7,0,75,0,156,0,18,0,111,0,34,0,30,0,210,0,177,0,145,0,223,0,12,0,209,0,251,0,185,0,46,0,122,0,126,0,122,0,73,0,56,0,100,0,122,0,7,0,0,0,186,0,63,0,187,0,4,0,69,0,0,0,237,0,43,0,110,0,87,0,60,0,30,0,168,0,10,0,0,0,56,0,0,0,116,0,247,0,53,0,5,0,72,0,0,0,143,0,0,0,0,0,0,0,67,0,76,0,0,0,58,0,203,0,23,0,0,0,0,0,0,0,197,0,77,0,222,0,42,0,31,0,128,0,59,0,211,0,93,0,255,0,171,0,167,0,104,0,154,0,242,0,135,0,51,0,133,0,232,0,87,0,248,0,224,0,0,0,14,0,50,0,137,0,65,0,200,0,72,0,244,0,112,0,177,0,206,0,0,0,153,0,227,0,222,0,123,0,201,0,201,0,0,0,109,0,29,0,30,0,231,0,181,0,72,0,249,0,67,0,247,0,0,0,200,0,1,0,211,0,74,0,243,0,148,0,172,0,208,0,54,0,94,0,122,0,200,0,0,0,0,0,101,0,72,0,131,0,0,0,0,0,0,0,184,0,36,0,171,0,26,0,200,0,53,0,0,0,47,0,0,0,0,0,153,0,94,0,60,0,234,0,115,0,205,0,217,0,0,0,184,0,103,0,221,0,207,0,5,0,96,0,245,0,101,0,189,0,4,0,237,0,0,0,16,0,149,0,98,0,199,0,184,0,191,0,245,0,0,0,181,0,29,0,14,0,127,0,3,0,43,0,32,0,0,0,12,0,163,0,65,0,171,0,103,0,171,0,167,0,196,0,97,0,62,0,16,0,254,0,231,0,192,0,160,0,0,0,46,0,205,0,0,0,55,0,17,0,34,0,61,0,30,0,187,0,30,0,249,0,14,0,18,0,85,0,140,0,117,0,235,0,251,0,236,0,0,0,75,0,104,0,183,0,228,0,49,0,143,0,123,0,110,0,55,0,117,0,21,0,35,0,136,0,202,0,26,0,187,0,0,0,222,0,60,0,0,0,1,0,0,0,122,0,124,0,191,0,0,0,103,0,218,0,54,0,32,0,0,0,40,0,0,0,125,0,57,0,72,0,87,0,233,0,181,0,0,0,108,0,101,0,70,0,205,0,0,0,81,0,212,0,123,0,0,0,32,0,0,0,0,0,77,0,0,0,200,0,203,0,186,0,255,0,191,0,59,0,68,0,26,0,105,0,208,0,103,0,168,0,70,0,119,0,67,0,22,0,0,0,158,0,162,0,152,0,141,0,181,0,81,0,192,0,0,0,0,0,107,0,219,0,203,0,13,0,200,0,169,0,201,0,143,0,225,0,90,0,111,0,239,0,119,0,128,0,122,0,134,0,0,0,0,0,178,0,0,0,129,0,0,0,209,0,0,0,90,0,176,0,30,0,0,0,200,0,122,0,0,0,120,0,99,0,63,0,248,0,161,0,4,0,35,0,193,0,99,0,44,0,118,0,31,0,8,0,55,0,0,0,112,0,106,0,204,0,0,0,126,0,0,0,47,0,166,0,183,0,237,0,0,0,233,0,8,0,227,0,119,0,83,0,90,0,62,0,161,0,112,0,0,0,0,0,231,0,111,0,192,0,0,0,0,0,179,0,0,0,84,0,150,0,154,0,133,0,6,0,10,0,0,0,0,0,101,0,219,0,187,0,142,0,192,0,0,0,182,0,53,0,42,0,234,0,129,0,142,0,0,0,232,0,0,0,249,0,198,0,170,0,63,0,117,0,227,0,0,0,0,0,221,0,55,0,205,0,99,0,26,0,185,0,0,0,96,0,0,0,50,0,47,0,0,0,0,0,63,0,43,0,55,0,184,0,17,0,74,0,0,0,220,0,45,0,0,0,173,0,2,0,96,0,0,0,250,0,203,0,0,0,92,0,164,0,0,0,183,0,248,0,0,0,42,0,2,0,12,0,38,0,0,0,19,0,219,0,80,0,187,0,0,0,41,0,54,0,87,0,46,0,133,0,0,0,202,0,123,0,51,0,207,0,18,0,36,0,51,0,0,0,85,0,0,0,0,0,115,0,102,0,198,0,12,0,0,0,100,0,0,0,235,0,168,0,49,0,0,0,0,0,231,0,231,0,104,0,102,0,121,0,0,0,190,0,187,0,124,0,230,0,89,0,222,0,153,0,203,0,114,0,128,0,0,0,27,0,0,0,40,0,183,0,158,0,11,0,0,0,66,0,240,0,77,0,68,0,195,0,140,0,62,0,141,0,250,0,0,0,81,0,165,0,12,0,0,0,57,0,101,0,189,0,33,0,0,0,206,0,166,0,0,0,0,0,0,0,228,0,87,0,122,0,0,0,104,0,98,0,142,0,155,0,80,0,237,0,162,0,128,0,120,0,154,0,0,0,149,0,0,0,98,0,33,0,164,0,183,0,204,0,219,0,145,0,0,0,135,0,86,0,66,0,80,0,6,0,78,0,157,0,0,0,0,0,233,0,4,0,192,0,116,0,226,0,214,0,184,0,162,0,80,0,74,0,250,0,103,0,148,0,40,0,55,0,0,0,39,0,250,0,13,0,126,0,229,0,207,0,191,0,0,0,73,0,73,0,191,0,23,0,66,0,14,0,128,0,79,0,49,0,192,0,243,0,0,0,54,0,254,0,0,0,148,0,121,0,159,0,106,0,244,0,114,0,0,0,81,0,39,0,13,0,0,0,54,0,89,0,22,0,0,0,0,0,220,0,0,0,253,0,9,0,149,0,246,0,211,0,0,0,0,0,147,0,0,0,46,0,140,0,113,0,146,0,5,0,0,0,237,0,212,0,97,0,0,0,152,0,8,0,68,0,43,0,85,0,175,0,67,0,51,0,0,0,148,0,118,0,85,0,145,0,0,0,164,0,28,0,160,0,67,0,226,0,0,0,0,0,16,0,2,0,254,0,29,0,162,0,16,0,84,0,25,0,182,0,148,0,173,0,174,0,230,0,24,0,224,0,121,0,106,0,200,0,145,0,91,0,122,0,85,0,151,0,130,0,221,0,53,0,158,0,239,0,0,0,174,0,240,0,0,0,7,0,149,0,24,0,55,0,20,0,62,0,0,0,0,0,37,0,213,0,125,0,213,0,0,0,52,0,80,0,0,0,174,0,0,0,76,0,53,0,136,0,251,0,205,0,154,0,221,0,212,0,138,0,108,0,0,0,0,0,185,0,0,0,10,0,0,0,180,0,167,0,77,0,27,0,37,0,0,0,213,0,138,0,135,0,0,0,236,0,0,0,184,0,46,0,39,0,167,0,0,0,233,0,76,0,0,0,242,0,147,0,211,0,175,0,105,0,0,0,240,0,170,0,75,0,202,0,251,0,61,0,0,0,208,0,3,0,9,0,97,0,52,0,88,0,189,0,19,0,0,0,119,0,180,0,138,0,17,0,63,0);
signal scenario_full  : scenario_type := (0,0,145,31,1,31,112,31,112,30,186,31,182,31,155,31,184,31,176,31,176,30,7,31,240,31,240,30,154,31,169,31,41,31,87,31,34,31,135,31,173,31,173,30,139,31,97,31,97,30,97,29,83,31,19,31,19,30,245,31,147,31,83,31,68,31,38,31,172,31,74,31,251,31,251,30,42,31,222,31,222,30,20,31,227,31,63,31,136,31,234,31,234,30,248,31,248,30,195,31,7,31,178,31,248,31,16,31,16,30,16,29,74,31,210,31,6,31,6,31,90,31,170,31,241,31,241,30,60,31,212,31,210,31,210,30,255,31,44,31,253,31,67,31,105,31,181,31,92,31,121,31,239,31,71,31,186,31,186,30,59,31,178,31,217,31,244,31,77,31,49,31,198,31,192,31,185,31,185,30,148,31,47,31,117,31,119,31,119,30,165,31,188,31,188,30,188,29,174,31,42,31,15,31,15,30,15,29,224,31,224,30,4,31,33,31,30,31,208,31,208,30,208,29,117,31,117,30,253,31,66,31,211,31,200,31,200,30,177,31,127,31,134,31,26,31,120,31,26,31,26,30,95,31,250,31,135,31,247,31,248,31,248,30,137,31,135,31,9,31,250,31,202,31,108,31,224,31,178,31,178,30,236,31,242,31,44,31,177,31,184,31,195,31,121,31,161,31,170,31,164,31,164,30,164,29,78,31,160,31,171,31,155,31,251,31,98,31,230,31,89,31,139,31,48,31,67,31,169,31,141,31,141,30,212,31,212,30,39,31,10,31,109,31,169,31,109,31,19,31,221,31,3,31,3,30,202,31,114,31,114,30,114,29,57,31,30,31,217,31,115,31,33,31,135,31,151,31,180,31,180,30,130,31,1,31,219,31,157,31,250,31,29,31,120,31,126,31,218,31,207,31,25,31,142,31,142,30,142,29,162,31,162,30,154,31,237,31,197,31,197,30,5,31,135,31,26,31,26,30,214,31,32,31,167,31,167,30,249,31,249,30,249,29,171,31,146,31,145,31,143,31,144,31,220,31,194,31,100,31,214,31,163,31,163,30,163,29,233,31,175,31,127,31,127,30,88,31,179,31,217,31,217,30,193,31,208,31,180,31,73,31,15,31,15,30,49,31,21,31,241,31,7,31,75,31,156,31,18,31,111,31,34,31,30,31,210,31,177,31,145,31,223,31,12,31,209,31,251,31,185,31,46,31,122,31,126,31,122,31,73,31,56,31,100,31,122,31,7,31,7,30,186,31,63,31,187,31,4,31,69,31,69,30,237,31,43,31,110,31,87,31,60,31,30,31,168,31,10,31,10,30,56,31,56,30,116,31,247,31,53,31,5,31,72,31,72,30,143,31,143,30,143,29,143,28,67,31,76,31,76,30,58,31,203,31,23,31,23,30,23,29,23,28,197,31,77,31,222,31,42,31,31,31,128,31,59,31,211,31,93,31,255,31,171,31,167,31,104,31,154,31,242,31,135,31,51,31,133,31,232,31,87,31,248,31,224,31,224,30,14,31,50,31,137,31,65,31,200,31,72,31,244,31,112,31,177,31,206,31,206,30,153,31,227,31,222,31,123,31,201,31,201,31,201,30,109,31,29,31,30,31,231,31,181,31,72,31,249,31,67,31,247,31,247,30,200,31,1,31,211,31,74,31,243,31,148,31,172,31,208,31,54,31,94,31,122,31,200,31,200,30,200,29,101,31,72,31,131,31,131,30,131,29,131,28,184,31,36,31,171,31,26,31,200,31,53,31,53,30,47,31,47,30,47,29,153,31,94,31,60,31,234,31,115,31,205,31,217,31,217,30,184,31,103,31,221,31,207,31,5,31,96,31,245,31,101,31,189,31,4,31,237,31,237,30,16,31,149,31,98,31,199,31,184,31,191,31,245,31,245,30,181,31,29,31,14,31,127,31,3,31,43,31,32,31,32,30,12,31,163,31,65,31,171,31,103,31,171,31,167,31,196,31,97,31,62,31,16,31,254,31,231,31,192,31,160,31,160,30,46,31,205,31,205,30,55,31,17,31,34,31,61,31,30,31,187,31,30,31,249,31,14,31,18,31,85,31,140,31,117,31,235,31,251,31,236,31,236,30,75,31,104,31,183,31,228,31,49,31,143,31,123,31,110,31,55,31,117,31,21,31,35,31,136,31,202,31,26,31,187,31,187,30,222,31,60,31,60,30,1,31,1,30,122,31,124,31,191,31,191,30,103,31,218,31,54,31,32,31,32,30,40,31,40,30,125,31,57,31,72,31,87,31,233,31,181,31,181,30,108,31,101,31,70,31,205,31,205,30,81,31,212,31,123,31,123,30,32,31,32,30,32,29,77,31,77,30,200,31,203,31,186,31,255,31,191,31,59,31,68,31,26,31,105,31,208,31,103,31,168,31,70,31,119,31,67,31,22,31,22,30,158,31,162,31,152,31,141,31,181,31,81,31,192,31,192,30,192,29,107,31,219,31,203,31,13,31,200,31,169,31,201,31,143,31,225,31,90,31,111,31,239,31,119,31,128,31,122,31,134,31,134,30,134,29,178,31,178,30,129,31,129,30,209,31,209,30,90,31,176,31,30,31,30,30,200,31,122,31,122,30,120,31,99,31,63,31,248,31,161,31,4,31,35,31,193,31,99,31,44,31,118,31,31,31,8,31,55,31,55,30,112,31,106,31,204,31,204,30,126,31,126,30,47,31,166,31,183,31,237,31,237,30,233,31,8,31,227,31,119,31,83,31,90,31,62,31,161,31,112,31,112,30,112,29,231,31,111,31,192,31,192,30,192,29,179,31,179,30,84,31,150,31,154,31,133,31,6,31,10,31,10,30,10,29,101,31,219,31,187,31,142,31,192,31,192,30,182,31,53,31,42,31,234,31,129,31,142,31,142,30,232,31,232,30,249,31,198,31,170,31,63,31,117,31,227,31,227,30,227,29,221,31,55,31,205,31,99,31,26,31,185,31,185,30,96,31,96,30,50,31,47,31,47,30,47,29,63,31,43,31,55,31,184,31,17,31,74,31,74,30,220,31,45,31,45,30,173,31,2,31,96,31,96,30,250,31,203,31,203,30,92,31,164,31,164,30,183,31,248,31,248,30,42,31,2,31,12,31,38,31,38,30,19,31,219,31,80,31,187,31,187,30,41,31,54,31,87,31,46,31,133,31,133,30,202,31,123,31,51,31,207,31,18,31,36,31,51,31,51,30,85,31,85,30,85,29,115,31,102,31,198,31,12,31,12,30,100,31,100,30,235,31,168,31,49,31,49,30,49,29,231,31,231,31,104,31,102,31,121,31,121,30,190,31,187,31,124,31,230,31,89,31,222,31,153,31,203,31,114,31,128,31,128,30,27,31,27,30,40,31,183,31,158,31,11,31,11,30,66,31,240,31,77,31,68,31,195,31,140,31,62,31,141,31,250,31,250,30,81,31,165,31,12,31,12,30,57,31,101,31,189,31,33,31,33,30,206,31,166,31,166,30,166,29,166,28,228,31,87,31,122,31,122,30,104,31,98,31,142,31,155,31,80,31,237,31,162,31,128,31,120,31,154,31,154,30,149,31,149,30,98,31,33,31,164,31,183,31,204,31,219,31,145,31,145,30,135,31,86,31,66,31,80,31,6,31,78,31,157,31,157,30,157,29,233,31,4,31,192,31,116,31,226,31,214,31,184,31,162,31,80,31,74,31,250,31,103,31,148,31,40,31,55,31,55,30,39,31,250,31,13,31,126,31,229,31,207,31,191,31,191,30,73,31,73,31,191,31,23,31,66,31,14,31,128,31,79,31,49,31,192,31,243,31,243,30,54,31,254,31,254,30,148,31,121,31,159,31,106,31,244,31,114,31,114,30,81,31,39,31,13,31,13,30,54,31,89,31,22,31,22,30,22,29,220,31,220,30,253,31,9,31,149,31,246,31,211,31,211,30,211,29,147,31,147,30,46,31,140,31,113,31,146,31,5,31,5,30,237,31,212,31,97,31,97,30,152,31,8,31,68,31,43,31,85,31,175,31,67,31,51,31,51,30,148,31,118,31,85,31,145,31,145,30,164,31,28,31,160,31,67,31,226,31,226,30,226,29,16,31,2,31,254,31,29,31,162,31,16,31,84,31,25,31,182,31,148,31,173,31,174,31,230,31,24,31,224,31,121,31,106,31,200,31,145,31,91,31,122,31,85,31,151,31,130,31,221,31,53,31,158,31,239,31,239,30,174,31,240,31,240,30,7,31,149,31,24,31,55,31,20,31,62,31,62,30,62,29,37,31,213,31,125,31,213,31,213,30,52,31,80,31,80,30,174,31,174,30,76,31,53,31,136,31,251,31,205,31,154,31,221,31,212,31,138,31,108,31,108,30,108,29,185,31,185,30,10,31,10,30,180,31,167,31,77,31,27,31,37,31,37,30,213,31,138,31,135,31,135,30,236,31,236,30,184,31,46,31,39,31,167,31,167,30,233,31,76,31,76,30,242,31,147,31,211,31,175,31,105,31,105,30,240,31,170,31,75,31,202,31,251,31,61,31,61,30,208,31,3,31,9,31,97,31,52,31,88,31,189,31,19,31,19,30,119,31,180,31,138,31,17,31,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
