-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 405;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (66,0,228,0,126,0,217,0,1,0,0,0,0,0,94,0,163,0,4,0,0,0,9,0,227,0,148,0,0,0,169,0,161,0,191,0,11,0,123,0,180,0,160,0,144,0,146,0,249,0,36,0,207,0,112,0,206,0,223,0,237,0,60,0,0,0,0,0,183,0,68,0,88,0,198,0,214,0,116,0,20,0,98,0,62,0,18,0,150,0,234,0,238,0,119,0,40,0,21,0,77,0,0,0,0,0,86,0,96,0,252,0,0,0,88,0,50,0,42,0,89,0,0,0,255,0,171,0,54,0,33,0,49,0,235,0,120,0,13,0,7,0,0,0,21,0,65,0,206,0,0,0,0,0,48,0,27,0,0,0,0,0,228,0,64,0,0,0,0,0,0,0,65,0,26,0,147,0,0,0,0,0,179,0,94,0,118,0,0,0,26,0,27,0,91,0,255,0,205,0,232,0,44,0,235,0,179,0,54,0,39,0,32,0,0,0,0,0,193,0,100,0,213,0,0,0,95,0,0,0,228,0,99,0,179,0,30,0,54,0,224,0,179,0,236,0,6,0,0,0,99,0,108,0,0,0,221,0,43,0,0,0,163,0,73,0,96,0,0,0,0,0,0,0,0,0,205,0,0,0,61,0,145,0,0,0,249,0,0,0,237,0,0,0,143,0,175,0,59,0,211,0,74,0,160,0,207,0,254,0,135,0,0,0,1,0,84,0,159,0,47,0,60,0,244,0,145,0,75,0,241,0,0,0,118,0,0,0,0,0,113,0,12,0,0,0,0,0,136,0,108,0,0,0,101,0,27,0,54,0,45,0,0,0,0,0,166,0,202,0,167,0,0,0,99,0,18,0,166,0,67,0,161,0,229,0,200,0,87,0,196,0,200,0,87,0,0,0,71,0,131,0,106,0,26,0,254,0,0,0,226,0,121,0,72,0,0,0,183,0,246,0,153,0,52,0,140,0,72,0,27,0,119,0,128,0,123,0,152,0,158,0,149,0,159,0,19,0,183,0,130,0,166,0,253,0,129,0,164,0,147,0,0,0,84,0,173,0,4,0,20,0,89,0,122,0,0,0,142,0,127,0,0,0,123,0,70,0,11,0,200,0,163,0,0,0,45,0,205,0,203,0,54,0,0,0,49,0,205,0,223,0,181,0,230,0,221,0,139,0,97,0,0,0,114,0,109,0,158,0,222,0,202,0,23,0,231,0,137,0,76,0,171,0,233,0,50,0,114,0,195,0,0,0,184,0,246,0,56,0,0,0,86,0,88,0,231,0,0,0,77,0,225,0,134,0,131,0,238,0,55,0,48,0,0,0,89,0,117,0,60,0,163,0,192,0,251,0,48,0,67,0,144,0,30,0,0,0,29,0,190,0,103,0,147,0,125,0,207,0,0,0,173,0,0,0,205,0,49,0,0,0,255,0,230,0,0,0,0,0,195,0,133,0,128,0,0,0,28,0,144,0,72,0,80,0,184,0,194,0,60,0,34,0,138,0,78,0,0,0,150,0,31,0,183,0,121,0,45,0,0,0,182,0,55,0,185,0,251,0,0,0,105,0,94,0,0,0,0,0,0,0,58,0,85,0,28,0,26,0,178,0,177,0,99,0,31,0,49,0,0,0,106,0,134,0,193,0,0,0,98,0,0,0,0,0,114,0,137,0,42,0,180,0,39,0,193,0,158,0,0,0,185,0,50,0,168,0,39,0,0,0,174,0,202,0,190,0,0,0,240,0,40,0,180,0,168,0,254,0,206,0,221,0,83,0,100,0,149,0,142,0,0,0,21,0,16,0,50,0,138,0,167,0,109,0,208,0,29,0);
signal scenario_full  : scenario_type := (66,31,228,31,126,31,217,31,1,31,1,30,1,29,94,31,163,31,4,31,4,30,9,31,227,31,148,31,148,30,169,31,161,31,191,31,11,31,123,31,180,31,160,31,144,31,146,31,249,31,36,31,207,31,112,31,206,31,223,31,237,31,60,31,60,30,60,29,183,31,68,31,88,31,198,31,214,31,116,31,20,31,98,31,62,31,18,31,150,31,234,31,238,31,119,31,40,31,21,31,77,31,77,30,77,29,86,31,96,31,252,31,252,30,88,31,50,31,42,31,89,31,89,30,255,31,171,31,54,31,33,31,49,31,235,31,120,31,13,31,7,31,7,30,21,31,65,31,206,31,206,30,206,29,48,31,27,31,27,30,27,29,228,31,64,31,64,30,64,29,64,28,65,31,26,31,147,31,147,30,147,29,179,31,94,31,118,31,118,30,26,31,27,31,91,31,255,31,205,31,232,31,44,31,235,31,179,31,54,31,39,31,32,31,32,30,32,29,193,31,100,31,213,31,213,30,95,31,95,30,228,31,99,31,179,31,30,31,54,31,224,31,179,31,236,31,6,31,6,30,99,31,108,31,108,30,221,31,43,31,43,30,163,31,73,31,96,31,96,30,96,29,96,28,96,27,205,31,205,30,61,31,145,31,145,30,249,31,249,30,237,31,237,30,143,31,175,31,59,31,211,31,74,31,160,31,207,31,254,31,135,31,135,30,1,31,84,31,159,31,47,31,60,31,244,31,145,31,75,31,241,31,241,30,118,31,118,30,118,29,113,31,12,31,12,30,12,29,136,31,108,31,108,30,101,31,27,31,54,31,45,31,45,30,45,29,166,31,202,31,167,31,167,30,99,31,18,31,166,31,67,31,161,31,229,31,200,31,87,31,196,31,200,31,87,31,87,30,71,31,131,31,106,31,26,31,254,31,254,30,226,31,121,31,72,31,72,30,183,31,246,31,153,31,52,31,140,31,72,31,27,31,119,31,128,31,123,31,152,31,158,31,149,31,159,31,19,31,183,31,130,31,166,31,253,31,129,31,164,31,147,31,147,30,84,31,173,31,4,31,20,31,89,31,122,31,122,30,142,31,127,31,127,30,123,31,70,31,11,31,200,31,163,31,163,30,45,31,205,31,203,31,54,31,54,30,49,31,205,31,223,31,181,31,230,31,221,31,139,31,97,31,97,30,114,31,109,31,158,31,222,31,202,31,23,31,231,31,137,31,76,31,171,31,233,31,50,31,114,31,195,31,195,30,184,31,246,31,56,31,56,30,86,31,88,31,231,31,231,30,77,31,225,31,134,31,131,31,238,31,55,31,48,31,48,30,89,31,117,31,60,31,163,31,192,31,251,31,48,31,67,31,144,31,30,31,30,30,29,31,190,31,103,31,147,31,125,31,207,31,207,30,173,31,173,30,205,31,49,31,49,30,255,31,230,31,230,30,230,29,195,31,133,31,128,31,128,30,28,31,144,31,72,31,80,31,184,31,194,31,60,31,34,31,138,31,78,31,78,30,150,31,31,31,183,31,121,31,45,31,45,30,182,31,55,31,185,31,251,31,251,30,105,31,94,31,94,30,94,29,94,28,58,31,85,31,28,31,26,31,178,31,177,31,99,31,31,31,49,31,49,30,106,31,134,31,193,31,193,30,98,31,98,30,98,29,114,31,137,31,42,31,180,31,39,31,193,31,158,31,158,30,185,31,50,31,168,31,39,31,39,30,174,31,202,31,190,31,190,30,240,31,40,31,180,31,168,31,254,31,206,31,221,31,83,31,100,31,149,31,142,31,142,30,21,31,16,31,50,31,138,31,167,31,109,31,208,31,29,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
