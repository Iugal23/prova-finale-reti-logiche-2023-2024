-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_110 is
end project_tb_110;

architecture project_tb_arch_110 of project_tb_110 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 278;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,66,0,180,0,32,0,23,0,83,0,182,0,213,0,48,0,194,0,81,0,4,0,143,0,243,0,127,0,0,0,198,0,136,0,230,0,69,0,159,0,148,0,167,0,186,0,240,0,54,0,111,0,182,0,1,0,0,0,102,0,0,0,118,0,65,0,210,0,0,0,79,0,223,0,74,0,0,0,160,0,0,0,16,0,140,0,50,0,0,0,64,0,59,0,26,0,77,0,173,0,0,0,6,0,17,0,0,0,166,0,0,0,0,0,32,0,203,0,0,0,105,0,99,0,219,0,0,0,179,0,177,0,87,0,16,0,0,0,0,0,35,0,0,0,0,0,98,0,8,0,205,0,0,0,241,0,230,0,0,0,21,0,67,0,164,0,147,0,101,0,92,0,4,0,0,0,199,0,246,0,0,0,229,0,195,0,0,0,85,0,232,0,90,0,2,0,128,0,16,0,0,0,86,0,71,0,219,0,242,0,176,0,18,0,238,0,200,0,227,0,0,0,46,0,107,0,144,0,82,0,251,0,124,0,20,0,0,0,124,0,5,0,15,0,50,0,234,0,70,0,129,0,96,0,0,0,125,0,105,0,57,0,135,0,160,0,16,0,112,0,130,0,59,0,172,0,237,0,0,0,13,0,0,0,212,0,188,0,35,0,209,0,114,0,54,0,51,0,179,0,180,0,231,0,12,0,30,0,233,0,130,0,0,0,0,0,241,0,47,0,0,0,243,0,130,0,207,0,0,0,252,0,62,0,93,0,68,0,0,0,229,0,165,0,154,0,212,0,114,0,63,0,4,0,98,0,120,0,0,0,0,0,213,0,0,0,0,0,199,0,129,0,55,0,45,0,12,0,17,0,90,0,195,0,41,0,22,0,141,0,228,0,201,0,47,0,55,0,239,0,0,0,20,0,249,0,93,0,75,0,76,0,0,0,133,0,78,0,211,0,218,0,179,0,103,0,221,0,41,0,195,0,71,0,158,0,100,0,234,0,207,0,220,0,45,0,77,0,0,0,189,0,0,0,141,0,27,0,0,0,0,0,123,0,152,0,115,0,156,0,95,0,157,0,56,0,16,0,68,0,207,0,15,0,0,0,179,0,2,0,132,0,0,0,0,0,187,0,67,0,21,0,73,0,28,0,175,0,211,0,241,0,189,0,96,0,126,0,170,0,0,0,56,0,188,0,44,0,9,0,1,0,0,0,149,0,0,0,204,0,89,0,0,0,113,0,0,0,119,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,66,31,180,31,32,31,23,31,83,31,182,31,213,31,48,31,194,31,81,31,4,31,143,31,243,31,127,31,127,30,198,31,136,31,230,31,69,31,159,31,148,31,167,31,186,31,240,31,54,31,111,31,182,31,1,31,1,30,102,31,102,30,118,31,65,31,210,31,210,30,79,31,223,31,74,31,74,30,160,31,160,30,16,31,140,31,50,31,50,30,64,31,59,31,26,31,77,31,173,31,173,30,6,31,17,31,17,30,166,31,166,30,166,29,32,31,203,31,203,30,105,31,99,31,219,31,219,30,179,31,177,31,87,31,16,31,16,30,16,29,35,31,35,30,35,29,98,31,8,31,205,31,205,30,241,31,230,31,230,30,21,31,67,31,164,31,147,31,101,31,92,31,4,31,4,30,199,31,246,31,246,30,229,31,195,31,195,30,85,31,232,31,90,31,2,31,128,31,16,31,16,30,86,31,71,31,219,31,242,31,176,31,18,31,238,31,200,31,227,31,227,30,46,31,107,31,144,31,82,31,251,31,124,31,20,31,20,30,124,31,5,31,15,31,50,31,234,31,70,31,129,31,96,31,96,30,125,31,105,31,57,31,135,31,160,31,16,31,112,31,130,31,59,31,172,31,237,31,237,30,13,31,13,30,212,31,188,31,35,31,209,31,114,31,54,31,51,31,179,31,180,31,231,31,12,31,30,31,233,31,130,31,130,30,130,29,241,31,47,31,47,30,243,31,130,31,207,31,207,30,252,31,62,31,93,31,68,31,68,30,229,31,165,31,154,31,212,31,114,31,63,31,4,31,98,31,120,31,120,30,120,29,213,31,213,30,213,29,199,31,129,31,55,31,45,31,12,31,17,31,90,31,195,31,41,31,22,31,141,31,228,31,201,31,47,31,55,31,239,31,239,30,20,31,249,31,93,31,75,31,76,31,76,30,133,31,78,31,211,31,218,31,179,31,103,31,221,31,41,31,195,31,71,31,158,31,100,31,234,31,207,31,220,31,45,31,77,31,77,30,189,31,189,30,141,31,27,31,27,30,27,29,123,31,152,31,115,31,156,31,95,31,157,31,56,31,16,31,68,31,207,31,15,31,15,30,179,31,2,31,132,31,132,30,132,29,187,31,67,31,21,31,73,31,28,31,175,31,211,31,241,31,189,31,96,31,126,31,170,31,170,30,56,31,188,31,44,31,9,31,1,31,1,30,149,31,149,30,204,31,89,31,89,30,113,31,113,30,119,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
