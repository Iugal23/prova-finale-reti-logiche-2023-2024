-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_894 is
end project_tb_894;

architecture project_tb_arch_894 of project_tb_894 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 486;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (176,0,0,0,126,0,67,0,139,0,231,0,93,0,24,0,29,0,73,0,0,0,58,0,0,0,239,0,132,0,113,0,146,0,219,0,0,0,225,0,53,0,52,0,202,0,148,0,188,0,93,0,160,0,178,0,0,0,0,0,7,0,35,0,0,0,145,0,127,0,66,0,140,0,0,0,110,0,0,0,5,0,230,0,78,0,0,0,87,0,79,0,77,0,0,0,202,0,74,0,0,0,98,0,131,0,173,0,217,0,218,0,100,0,0,0,152,0,154,0,184,0,80,0,99,0,22,0,0,0,0,0,53,0,71,0,12,0,153,0,95,0,157,0,127,0,108,0,86,0,37,0,47,0,200,0,235,0,34,0,115,0,181,0,0,0,87,0,152,0,75,0,0,0,12,0,208,0,237,0,39,0,0,0,143,0,247,0,146,0,0,0,183,0,5,0,0,0,228,0,0,0,11,0,249,0,39,0,53,0,0,0,231,0,181,0,154,0,137,0,0,0,43,0,103,0,57,0,196,0,97,0,0,0,56,0,96,0,101,0,171,0,166,0,0,0,14,0,42,0,158,0,0,0,49,0,0,0,194,0,243,0,84,0,0,0,117,0,93,0,0,0,16,0,0,0,142,0,228,0,141,0,51,0,61,0,59,0,160,0,0,0,75,0,14,0,0,0,214,0,181,0,199,0,0,0,221,0,157,0,0,0,126,0,125,0,11,0,50,0,46,0,19,0,215,0,122,0,71,0,159,0,238,0,0,0,0,0,149,0,93,0,195,0,66,0,90,0,0,0,0,0,0,0,0,0,39,0,176,0,129,0,0,0,100,0,207,0,0,0,171,0,0,0,45,0,132,0,6,0,0,0,47,0,0,0,36,0,98,0,240,0,114,0,21,0,0,0,161,0,0,0,0,0,244,0,62,0,146,0,0,0,147,0,0,0,0,0,0,0,138,0,173,0,0,0,98,0,0,0,0,0,48,0,26,0,49,0,119,0,0,0,163,0,0,0,223,0,95,0,0,0,155,0,51,0,7,0,114,0,190,0,52,0,0,0,196,0,8,0,4,0,209,0,0,0,88,0,143,0,72,0,106,0,52,0,79,0,0,0,110,0,92,0,165,0,0,0,136,0,0,0,47,0,138,0,3,0,129,0,0,0,143,0,77,0,24,0,230,0,30,0,33,0,195,0,26,0,159,0,0,0,144,0,0,0,202,0,57,0,243,0,55,0,0,0,53,0,243,0,195,0,242,0,0,0,0,0,244,0,32,0,194,0,198,0,0,0,75,0,0,0,0,0,151,0,165,0,103,0,83,0,161,0,30,0,63,0,144,0,212,0,54,0,56,0,92,0,0,0,16,0,57,0,126,0,182,0,174,0,0,0,158,0,194,0,22,0,171,0,80,0,121,0,82,0,224,0,85,0,132,0,37,0,64,0,147,0,121,0,161,0,151,0,90,0,154,0,195,0,229,0,175,0,64,0,26,0,0,0,85,0,0,0,44,0,0,0,253,0,248,0,0,0,68,0,85,0,242,0,249,0,119,0,195,0,0,0,193,0,123,0,0,0,0,0,0,0,118,0,87,0,0,0,91,0,233,0,134,0,215,0,0,0,0,0,209,0,140,0,70,0,183,0,137,0,79,0,3,0,241,0,0,0,200,0,32,0,165,0,202,0,103,0,236,0,86,0,27,0,229,0,237,0,0,0,34,0,2,0,158,0,205,0,105,0,124,0,0,0,94,0,119,0,88,0,57,0,191,0,0,0,134,0,121,0,0,0,184,0,0,0,0,0,22,0,73,0,172,0,0,0,128,0,24,0,71,0,123,0,204,0,104,0,132,0,40,0,38,0,194,0,224,0,6,0,49,0,146,0,169,0,110,0,60,0,150,0,233,0,233,0,15,0,238,0,69,0,142,0,0,0,82,0,0,0,172,0,217,0,46,0,147,0,193,0,113,0,0,0,0,0,0,0,63,0,115,0,0,0,180,0,0,0,202,0,0,0,103,0,163,0,126,0,150,0,240,0,0,0,0,0,0,0,153,0,97,0,32,0,214,0,16,0,120,0,209,0,101,0,182,0,65,0,162,0,24,0,0,0,197,0,34,0,0,0,227,0,11,0,235,0,139,0,72,0,55,0,29,0,252,0,0,0,0,0,127,0,134,0,249,0,35,0,42,0,0,0,197,0,168,0);
signal scenario_full  : scenario_type := (176,31,176,30,126,31,67,31,139,31,231,31,93,31,24,31,29,31,73,31,73,30,58,31,58,30,239,31,132,31,113,31,146,31,219,31,219,30,225,31,53,31,52,31,202,31,148,31,188,31,93,31,160,31,178,31,178,30,178,29,7,31,35,31,35,30,145,31,127,31,66,31,140,31,140,30,110,31,110,30,5,31,230,31,78,31,78,30,87,31,79,31,77,31,77,30,202,31,74,31,74,30,98,31,131,31,173,31,217,31,218,31,100,31,100,30,152,31,154,31,184,31,80,31,99,31,22,31,22,30,22,29,53,31,71,31,12,31,153,31,95,31,157,31,127,31,108,31,86,31,37,31,47,31,200,31,235,31,34,31,115,31,181,31,181,30,87,31,152,31,75,31,75,30,12,31,208,31,237,31,39,31,39,30,143,31,247,31,146,31,146,30,183,31,5,31,5,30,228,31,228,30,11,31,249,31,39,31,53,31,53,30,231,31,181,31,154,31,137,31,137,30,43,31,103,31,57,31,196,31,97,31,97,30,56,31,96,31,101,31,171,31,166,31,166,30,14,31,42,31,158,31,158,30,49,31,49,30,194,31,243,31,84,31,84,30,117,31,93,31,93,30,16,31,16,30,142,31,228,31,141,31,51,31,61,31,59,31,160,31,160,30,75,31,14,31,14,30,214,31,181,31,199,31,199,30,221,31,157,31,157,30,126,31,125,31,11,31,50,31,46,31,19,31,215,31,122,31,71,31,159,31,238,31,238,30,238,29,149,31,93,31,195,31,66,31,90,31,90,30,90,29,90,28,90,27,39,31,176,31,129,31,129,30,100,31,207,31,207,30,171,31,171,30,45,31,132,31,6,31,6,30,47,31,47,30,36,31,98,31,240,31,114,31,21,31,21,30,161,31,161,30,161,29,244,31,62,31,146,31,146,30,147,31,147,30,147,29,147,28,138,31,173,31,173,30,98,31,98,30,98,29,48,31,26,31,49,31,119,31,119,30,163,31,163,30,223,31,95,31,95,30,155,31,51,31,7,31,114,31,190,31,52,31,52,30,196,31,8,31,4,31,209,31,209,30,88,31,143,31,72,31,106,31,52,31,79,31,79,30,110,31,92,31,165,31,165,30,136,31,136,30,47,31,138,31,3,31,129,31,129,30,143,31,77,31,24,31,230,31,30,31,33,31,195,31,26,31,159,31,159,30,144,31,144,30,202,31,57,31,243,31,55,31,55,30,53,31,243,31,195,31,242,31,242,30,242,29,244,31,32,31,194,31,198,31,198,30,75,31,75,30,75,29,151,31,165,31,103,31,83,31,161,31,30,31,63,31,144,31,212,31,54,31,56,31,92,31,92,30,16,31,57,31,126,31,182,31,174,31,174,30,158,31,194,31,22,31,171,31,80,31,121,31,82,31,224,31,85,31,132,31,37,31,64,31,147,31,121,31,161,31,151,31,90,31,154,31,195,31,229,31,175,31,64,31,26,31,26,30,85,31,85,30,44,31,44,30,253,31,248,31,248,30,68,31,85,31,242,31,249,31,119,31,195,31,195,30,193,31,123,31,123,30,123,29,123,28,118,31,87,31,87,30,91,31,233,31,134,31,215,31,215,30,215,29,209,31,140,31,70,31,183,31,137,31,79,31,3,31,241,31,241,30,200,31,32,31,165,31,202,31,103,31,236,31,86,31,27,31,229,31,237,31,237,30,34,31,2,31,158,31,205,31,105,31,124,31,124,30,94,31,119,31,88,31,57,31,191,31,191,30,134,31,121,31,121,30,184,31,184,30,184,29,22,31,73,31,172,31,172,30,128,31,24,31,71,31,123,31,204,31,104,31,132,31,40,31,38,31,194,31,224,31,6,31,49,31,146,31,169,31,110,31,60,31,150,31,233,31,233,31,15,31,238,31,69,31,142,31,142,30,82,31,82,30,172,31,217,31,46,31,147,31,193,31,113,31,113,30,113,29,113,28,63,31,115,31,115,30,180,31,180,30,202,31,202,30,103,31,163,31,126,31,150,31,240,31,240,30,240,29,240,28,153,31,97,31,32,31,214,31,16,31,120,31,209,31,101,31,182,31,65,31,162,31,24,31,24,30,197,31,34,31,34,30,227,31,11,31,235,31,139,31,72,31,55,31,29,31,252,31,252,30,252,29,127,31,134,31,249,31,35,31,42,31,42,30,197,31,168,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
