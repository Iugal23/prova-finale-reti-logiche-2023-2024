-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 866;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (170,0,212,0,88,0,242,0,0,0,0,0,0,0,64,0,90,0,231,0,117,0,17,0,47,0,235,0,93,0,191,0,137,0,245,0,131,0,0,0,156,0,226,0,185,0,255,0,120,0,14,0,89,0,24,0,0,0,0,0,171,0,28,0,96,0,231,0,97,0,209,0,111,0,110,0,103,0,158,0,70,0,74,0,146,0,73,0,100,0,0,0,31,0,27,0,26,0,215,0,49,0,78,0,62,0,87,0,243,0,0,0,224,0,8,0,30,0,110,0,161,0,239,0,94,0,158,0,91,0,186,0,210,0,101,0,66,0,115,0,41,0,0,0,46,0,202,0,149,0,0,0,248,0,0,0,18,0,145,0,93,0,50,0,193,0,237,0,117,0,0,0,0,0,0,0,117,0,186,0,72,0,83,0,0,0,186,0,133,0,219,0,0,0,194,0,47,0,251,0,99,0,167,0,7,0,152,0,0,0,26,0,191,0,223,0,0,0,172,0,0,0,226,0,156,0,239,0,107,0,199,0,185,0,126,0,145,0,68,0,30,0,172,0,224,0,236,0,56,0,228,0,188,0,137,0,228,0,0,0,58,0,255,0,0,0,28,0,27,0,223,0,167,0,0,0,0,0,172,0,236,0,129,0,0,0,148,0,180,0,0,0,203,0,0,0,18,0,224,0,237,0,99,0,239,0,138,0,0,0,90,0,129,0,0,0,228,0,0,0,0,0,209,0,170,0,145,0,0,0,5,0,0,0,17,0,121,0,199,0,86,0,12,0,219,0,215,0,99,0,142,0,13,0,73,0,118,0,75,0,195,0,222,0,62,0,143,0,181,0,0,0,255,0,23,0,184,0,0,0,168,0,149,0,134,0,109,0,250,0,0,0,192,0,0,0,222,0,108,0,103,0,176,0,240,0,0,0,229,0,0,0,254,0,133,0,30,0,0,0,243,0,111,0,197,0,167,0,135,0,0,0,114,0,181,0,61,0,208,0,216,0,27,0,0,0,0,0,86,0,237,0,152,0,18,0,20,0,243,0,96,0,0,0,165,0,190,0,13,0,123,0,239,0,189,0,124,0,217,0,226,0,120,0,182,0,0,0,45,0,201,0,37,0,0,0,199,0,89,0,169,0,0,0,187,0,121,0,37,0,92,0,229,0,0,0,87,0,168,0,0,0,82,0,199,0,236,0,105,0,72,0,145,0,0,0,80,0,0,0,0,0,0,0,71,0,167,0,97,0,0,0,102,0,26,0,140,0,0,0,113,0,60,0,0,0,0,0,115,0,19,0,0,0,0,0,228,0,249,0,0,0,249,0,103,0,0,0,77,0,42,0,205,0,150,0,122,0,0,0,137,0,0,0,100,0,67,0,79,0,208,0,210,0,34,0,35,0,0,0,0,0,0,0,0,0,0,0,103,0,178,0,162,0,0,0,32,0,0,0,2,0,68,0,165,0,5,0,63,0,160,0,0,0,56,0,80,0,0,0,250,0,76,0,232,0,0,0,100,0,13,0,104,0,197,0,24,0,253,0,42,0,230,0,17,0,97,0,0,0,0,0,3,0,235,0,95,0,159,0,37,0,2,0,0,0,201,0,176,0,0,0,53,0,84,0,31,0,190,0,89,0,30,0,144,0,0,0,39,0,114,0,56,0,0,0,123,0,249,0,232,0,0,0,35,0,166,0,0,0,212,0,182,0,55,0,153,0,16,0,128,0,255,0,69,0,0,0,0,0,157,0,168,0,0,0,228,0,152,0,241,0,0,0,229,0,211,0,233,0,0,0,0,0,182,0,0,0,0,0,0,0,0,0,134,0,231,0,49,0,64,0,232,0,92,0,93,0,94,0,40,0,0,0,139,0,69,0,190,0,72,0,19,0,24,0,74,0,80,0,76,0,230,0,46,0,130,0,109,0,0,0,189,0,0,0,0,0,22,0,35,0,36,0,144,0,139,0,26,0,89,0,5,0,203,0,0,0,0,0,179,0,62,0,0,0,230,0,0,0,254,0,0,0,0,0,0,0,12,0,238,0,83,0,246,0,151,0,233,0,42,0,248,0,129,0,0,0,0,0,0,0,0,0,124,0,93,0,144,0,8,0,164,0,92,0,251,0,188,0,199,0,254,0,0,0,207,0,173,0,88,0,72,0,104,0,34,0,207,0,23,0,151,0,99,0,140,0,86,0,6,0,0,0,90,0,245,0,77,0,0,0,0,0,229,0,78,0,0,0,239,0,241,0,142,0,99,0,136,0,28,0,141,0,70,0,82,0,116,0,99,0,148,0,8,0,215,0,215,0,204,0,152,0,197,0,39,0,146,0,129,0,0,0,150,0,155,0,181,0,64,0,78,0,0,0,168,0,190,0,255,0,8,0,248,0,185,0,250,0,187,0,51,0,148,0,80,0,130,0,73,0,246,0,143,0,0,0,144,0,143,0,196,0,0,0,241,0,153,0,149,0,0,0,72,0,166,0,85,0,176,0,178,0,54,0,98,0,228,0,149,0,95,0,250,0,0,0,176,0,37,0,130,0,198,0,223,0,0,0,0,0,15,0,93,0,112,0,107,0,0,0,156,0,235,0,4,0,66,0,50,0,103,0,209,0,0,0,0,0,7,0,221,0,61,0,107,0,0,0,69,0,61,0,0,0,150,0,128,0,0,0,175,0,77,0,3,0,211,0,60,0,153,0,133,0,141,0,159,0,0,0,50,0,198,0,0,0,0,0,34,0,182,0,68,0,77,0,223,0,197,0,157,0,110,0,193,0,190,0,0,0,0,0,222,0,238,0,204,0,224,0,12,0,223,0,60,0,236,0,215,0,229,0,159,0,194,0,188,0,6,0,98,0,0,0,108,0,162,0,121,0,17,0,157,0,204,0,0,0,243,0,77,0,95,0,173,0,111,0,77,0,167,0,25,0,249,0,2,0,188,0,0,0,45,0,69,0,200,0,0,0,206,0,139,0,0,0,200,0,156,0,173,0,153,0,22,0,42,0,120,0,18,0,223,0,92,0,104,0,214,0,0,0,31,0,61,0,128,0,183,0,22,0,0,0,58,0,0,0,243,0,243,0,35,0,120,0,218,0,17,0,156,0,27,0,78,0,0,0,55,0,147,0,100,0,0,0,149,0,93,0,141,0,0,0,189,0,120,0,11,0,0,0,248,0,0,0,23,0,15,0,154,0,0,0,33,0,144,0,79,0,180,0,36,0,77,0,28,0,102,0,0,0,213,0,111,0,234,0,132,0,240,0,69,0,251,0,192,0,0,0,220,0,49,0,41,0,93,0,61,0,219,0,133,0,246,0,191,0,0,0,10,0,0,0,168,0,86,0,69,0,206,0,55,0,117,0,80,0,0,0,158,0,55,0,76,0,216,0,128,0,131,0,223,0,0,0,0,0,0,0,127,0,140,0,169,0,190,0,0,0,0,0,80,0,67,0,119,0,221,0,42,0,0,0,39,0,217,0,6,0,107,0,135,0,44,0,67,0,0,0,166,0,84,0,141,0,165,0,0,0,83,0,183,0,35,0,76,0,97,0,0,0,42,0,71,0,127,0,107,0,49,0,138,0,0,0,195,0,189,0,0,0,135,0,120,0,97,0,116,0,200,0,9,0,206,0,207,0,207,0,0,0,62,0,111,0,205,0,219,0,205,0,99,0,217,0,0,0,85,0,196,0,106,0,0,0,168,0,145,0,0,0,212,0,0,0,0,0,69,0,61,0,159,0,54,0,119,0,114,0,228,0,6,0,0,0,97,0,0,0,84,0,51,0,57,0,100,0,81,0,186,0,11,0,0,0,0,0,199,0,50,0,164,0,221,0,65,0,50,0,87,0,181,0,160,0,0,0,0,0,113,0,100,0,78,0,239,0,222,0,137,0,216,0,127,0,65,0,0,0);
signal scenario_full  : scenario_type := (170,31,212,31,88,31,242,31,242,30,242,29,242,28,64,31,90,31,231,31,117,31,17,31,47,31,235,31,93,31,191,31,137,31,245,31,131,31,131,30,156,31,226,31,185,31,255,31,120,31,14,31,89,31,24,31,24,30,24,29,171,31,28,31,96,31,231,31,97,31,209,31,111,31,110,31,103,31,158,31,70,31,74,31,146,31,73,31,100,31,100,30,31,31,27,31,26,31,215,31,49,31,78,31,62,31,87,31,243,31,243,30,224,31,8,31,30,31,110,31,161,31,239,31,94,31,158,31,91,31,186,31,210,31,101,31,66,31,115,31,41,31,41,30,46,31,202,31,149,31,149,30,248,31,248,30,18,31,145,31,93,31,50,31,193,31,237,31,117,31,117,30,117,29,117,28,117,31,186,31,72,31,83,31,83,30,186,31,133,31,219,31,219,30,194,31,47,31,251,31,99,31,167,31,7,31,152,31,152,30,26,31,191,31,223,31,223,30,172,31,172,30,226,31,156,31,239,31,107,31,199,31,185,31,126,31,145,31,68,31,30,31,172,31,224,31,236,31,56,31,228,31,188,31,137,31,228,31,228,30,58,31,255,31,255,30,28,31,27,31,223,31,167,31,167,30,167,29,172,31,236,31,129,31,129,30,148,31,180,31,180,30,203,31,203,30,18,31,224,31,237,31,99,31,239,31,138,31,138,30,90,31,129,31,129,30,228,31,228,30,228,29,209,31,170,31,145,31,145,30,5,31,5,30,17,31,121,31,199,31,86,31,12,31,219,31,215,31,99,31,142,31,13,31,73,31,118,31,75,31,195,31,222,31,62,31,143,31,181,31,181,30,255,31,23,31,184,31,184,30,168,31,149,31,134,31,109,31,250,31,250,30,192,31,192,30,222,31,108,31,103,31,176,31,240,31,240,30,229,31,229,30,254,31,133,31,30,31,30,30,243,31,111,31,197,31,167,31,135,31,135,30,114,31,181,31,61,31,208,31,216,31,27,31,27,30,27,29,86,31,237,31,152,31,18,31,20,31,243,31,96,31,96,30,165,31,190,31,13,31,123,31,239,31,189,31,124,31,217,31,226,31,120,31,182,31,182,30,45,31,201,31,37,31,37,30,199,31,89,31,169,31,169,30,187,31,121,31,37,31,92,31,229,31,229,30,87,31,168,31,168,30,82,31,199,31,236,31,105,31,72,31,145,31,145,30,80,31,80,30,80,29,80,28,71,31,167,31,97,31,97,30,102,31,26,31,140,31,140,30,113,31,60,31,60,30,60,29,115,31,19,31,19,30,19,29,228,31,249,31,249,30,249,31,103,31,103,30,77,31,42,31,205,31,150,31,122,31,122,30,137,31,137,30,100,31,67,31,79,31,208,31,210,31,34,31,35,31,35,30,35,29,35,28,35,27,35,26,103,31,178,31,162,31,162,30,32,31,32,30,2,31,68,31,165,31,5,31,63,31,160,31,160,30,56,31,80,31,80,30,250,31,76,31,232,31,232,30,100,31,13,31,104,31,197,31,24,31,253,31,42,31,230,31,17,31,97,31,97,30,97,29,3,31,235,31,95,31,159,31,37,31,2,31,2,30,201,31,176,31,176,30,53,31,84,31,31,31,190,31,89,31,30,31,144,31,144,30,39,31,114,31,56,31,56,30,123,31,249,31,232,31,232,30,35,31,166,31,166,30,212,31,182,31,55,31,153,31,16,31,128,31,255,31,69,31,69,30,69,29,157,31,168,31,168,30,228,31,152,31,241,31,241,30,229,31,211,31,233,31,233,30,233,29,182,31,182,30,182,29,182,28,182,27,134,31,231,31,49,31,64,31,232,31,92,31,93,31,94,31,40,31,40,30,139,31,69,31,190,31,72,31,19,31,24,31,74,31,80,31,76,31,230,31,46,31,130,31,109,31,109,30,189,31,189,30,189,29,22,31,35,31,36,31,144,31,139,31,26,31,89,31,5,31,203,31,203,30,203,29,179,31,62,31,62,30,230,31,230,30,254,31,254,30,254,29,254,28,12,31,238,31,83,31,246,31,151,31,233,31,42,31,248,31,129,31,129,30,129,29,129,28,129,27,124,31,93,31,144,31,8,31,164,31,92,31,251,31,188,31,199,31,254,31,254,30,207,31,173,31,88,31,72,31,104,31,34,31,207,31,23,31,151,31,99,31,140,31,86,31,6,31,6,30,90,31,245,31,77,31,77,30,77,29,229,31,78,31,78,30,239,31,241,31,142,31,99,31,136,31,28,31,141,31,70,31,82,31,116,31,99,31,148,31,8,31,215,31,215,31,204,31,152,31,197,31,39,31,146,31,129,31,129,30,150,31,155,31,181,31,64,31,78,31,78,30,168,31,190,31,255,31,8,31,248,31,185,31,250,31,187,31,51,31,148,31,80,31,130,31,73,31,246,31,143,31,143,30,144,31,143,31,196,31,196,30,241,31,153,31,149,31,149,30,72,31,166,31,85,31,176,31,178,31,54,31,98,31,228,31,149,31,95,31,250,31,250,30,176,31,37,31,130,31,198,31,223,31,223,30,223,29,15,31,93,31,112,31,107,31,107,30,156,31,235,31,4,31,66,31,50,31,103,31,209,31,209,30,209,29,7,31,221,31,61,31,107,31,107,30,69,31,61,31,61,30,150,31,128,31,128,30,175,31,77,31,3,31,211,31,60,31,153,31,133,31,141,31,159,31,159,30,50,31,198,31,198,30,198,29,34,31,182,31,68,31,77,31,223,31,197,31,157,31,110,31,193,31,190,31,190,30,190,29,222,31,238,31,204,31,224,31,12,31,223,31,60,31,236,31,215,31,229,31,159,31,194,31,188,31,6,31,98,31,98,30,108,31,162,31,121,31,17,31,157,31,204,31,204,30,243,31,77,31,95,31,173,31,111,31,77,31,167,31,25,31,249,31,2,31,188,31,188,30,45,31,69,31,200,31,200,30,206,31,139,31,139,30,200,31,156,31,173,31,153,31,22,31,42,31,120,31,18,31,223,31,92,31,104,31,214,31,214,30,31,31,61,31,128,31,183,31,22,31,22,30,58,31,58,30,243,31,243,31,35,31,120,31,218,31,17,31,156,31,27,31,78,31,78,30,55,31,147,31,100,31,100,30,149,31,93,31,141,31,141,30,189,31,120,31,11,31,11,30,248,31,248,30,23,31,15,31,154,31,154,30,33,31,144,31,79,31,180,31,36,31,77,31,28,31,102,31,102,30,213,31,111,31,234,31,132,31,240,31,69,31,251,31,192,31,192,30,220,31,49,31,41,31,93,31,61,31,219,31,133,31,246,31,191,31,191,30,10,31,10,30,168,31,86,31,69,31,206,31,55,31,117,31,80,31,80,30,158,31,55,31,76,31,216,31,128,31,131,31,223,31,223,30,223,29,223,28,127,31,140,31,169,31,190,31,190,30,190,29,80,31,67,31,119,31,221,31,42,31,42,30,39,31,217,31,6,31,107,31,135,31,44,31,67,31,67,30,166,31,84,31,141,31,165,31,165,30,83,31,183,31,35,31,76,31,97,31,97,30,42,31,71,31,127,31,107,31,49,31,138,31,138,30,195,31,189,31,189,30,135,31,120,31,97,31,116,31,200,31,9,31,206,31,207,31,207,31,207,30,62,31,111,31,205,31,219,31,205,31,99,31,217,31,217,30,85,31,196,31,106,31,106,30,168,31,145,31,145,30,212,31,212,30,212,29,69,31,61,31,159,31,54,31,119,31,114,31,228,31,6,31,6,30,97,31,97,30,84,31,51,31,57,31,100,31,81,31,186,31,11,31,11,30,11,29,199,31,50,31,164,31,221,31,65,31,50,31,87,31,181,31,160,31,160,30,160,29,113,31,100,31,78,31,239,31,222,31,137,31,216,31,127,31,65,31,65,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
