-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 910;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,116,0,125,0,194,0,134,0,17,0,23,0,0,0,13,0,0,0,101,0,39,0,26,0,68,0,130,0,205,0,56,0,197,0,182,0,174,0,35,0,35,0,0,0,0,0,30,0,12,0,161,0,62,0,164,0,0,0,34,0,173,0,200,0,220,0,40,0,0,0,102,0,0,0,0,0,211,0,0,0,179,0,125,0,18,0,104,0,136,0,206,0,35,0,241,0,226,0,0,0,33,0,127,0,62,0,229,0,253,0,48,0,137,0,58,0,62,0,255,0,223,0,122,0,55,0,29,0,190,0,128,0,217,0,105,0,234,0,55,0,20,0,29,0,1,0,0,0,97,0,222,0,34,0,0,0,122,0,150,0,87,0,202,0,249,0,0,0,132,0,26,0,56,0,142,0,183,0,63,0,168,0,255,0,233,0,82,0,177,0,0,0,0,0,185,0,201,0,66,0,246,0,210,0,119,0,17,0,170,0,0,0,24,0,136,0,73,0,242,0,28,0,0,0,49,0,193,0,147,0,218,0,8,0,206,0,0,0,95,0,0,0,0,0,0,0,11,0,73,0,116,0,156,0,226,0,0,0,186,0,91,0,247,0,123,0,207,0,119,0,226,0,57,0,180,0,35,0,108,0,0,0,100,0,0,0,5,0,0,0,0,0,16,0,27,0,0,0,93,0,249,0,208,0,230,0,23,0,254,0,0,0,230,0,228,0,0,0,110,0,141,0,238,0,0,0,93,0,166,0,0,0,220,0,57,0,2,0,37,0,0,0,146,0,0,0,223,0,233,0,14,0,50,0,150,0,242,0,142,0,0,0,226,0,247,0,46,0,18,0,26,0,121,0,185,0,6,0,0,0,9,0,45,0,11,0,154,0,34,0,219,0,86,0,215,0,244,0,0,0,238,0,0,0,0,0,248,0,0,0,236,0,192,0,144,0,156,0,60,0,3,0,44,0,117,0,0,0,219,0,208,0,39,0,95,0,61,0,218,0,0,0,4,0,50,0,13,0,161,0,47,0,212,0,123,0,0,0,133,0,0,0,0,0,163,0,196,0,0,0,185,0,0,0,163,0,224,0,108,0,214,0,204,0,0,0,191,0,252,0,206,0,141,0,75,0,26,0,0,0,67,0,0,0,250,0,51,0,228,0,230,0,153,0,199,0,181,0,68,0,221,0,0,0,206,0,23,0,248,0,83,0,211,0,0,0,0,0,206,0,34,0,40,0,0,0,133,0,2,0,0,0,130,0,0,0,1,0,112,0,0,0,0,0,79,0,89,0,0,0,0,0,212,0,27,0,0,0,233,0,209,0,0,0,0,0,252,0,232,0,114,0,98,0,129,0,204,0,73,0,0,0,27,0,111,0,69,0,137,0,231,0,198,0,175,0,0,0,102,0,108,0,233,0,131,0,65,0,218,0,72,0,208,0,61,0,24,0,102,0,0,0,81,0,229,0,0,0,0,0,252,0,61,0,214,0,234,0,45,0,75,0,130,0,0,0,34,0,2,0,0,0,243,0,255,0,188,0,0,0,250,0,162,0,177,0,236,0,44,0,82,0,82,0,139,0,133,0,212,0,171,0,24,0,52,0,106,0,118,0,30,0,194,0,191,0,217,0,156,0,0,0,100,0,60,0,0,0,193,0,174,0,86,0,40,0,161,0,92,0,0,0,102,0,190,0,0,0,94,0,62,0,188,0,190,0,77,0,95,0,83,0,221,0,232,0,0,0,201,0,87,0,136,0,58,0,106,0,191,0,0,0,61,0,211,0,0,0,117,0,52,0,156,0,168,0,210,0,0,0,155,0,0,0,31,0,88,0,0,0,176,0,13,0,252,0,0,0,58,0,177,0,198,0,0,0,0,0,219,0,0,0,30,0,0,0,105,0,110,0,108,0,131,0,103,0,162,0,142,0,25,0,0,0,0,0,239,0,196,0,120,0,196,0,10,0,230,0,0,0,6,0,175,0,0,0,134,0,121,0,89,0,211,0,118,0,0,0,51,0,61,0,0,0,159,0,30,0,250,0,211,0,0,0,22,0,206,0,17,0,157,0,108,0,194,0,29,0,21,0,96,0,159,0,175,0,72,0,80,0,0,0,20,0,208,0,6,0,0,0,31,0,186,0,216,0,187,0,94,0,144,0,228,0,170,0,117,0,15,0,62,0,0,0,3,0,0,0,90,0,193,0,234,0,0,0,71,0,127,0,77,0,149,0,61,0,0,0,233,0,0,0,47,0,0,0,0,0,160,0,42,0,128,0,0,0,203,0,64,0,0,0,5,0,233,0,140,0,34,0,140,0,99,0,186,0,44,0,188,0,160,0,226,0,96,0,62,0,162,0,161,0,229,0,161,0,0,0,105,0,21,0,14,0,159,0,0,0,53,0,252,0,0,0,12,0,74,0,70,0,222,0,41,0,0,0,63,0,98,0,78,0,23,0,38,0,62,0,33,0,201,0,0,0,135,0,136,0,23,0,22,0,70,0,117,0,22,0,144,0,0,0,139,0,153,0,137,0,0,0,158,0,136,0,74,0,88,0,8,0,140,0,44,0,247,0,0,0,204,0,165,0,13,0,0,0,223,0,241,0,167,0,232,0,60,0,80,0,181,0,0,0,0,0,132,0,49,0,41,0,123,0,0,0,199,0,61,0,239,0,227,0,100,0,92,0,54,0,190,0,24,0,10,0,215,0,157,0,161,0,176,0,0,0,86,0,73,0,66,0,102,0,230,0,125,0,0,0,36,0,234,0,123,0,0,0,0,0,255,0,0,0,26,0,89,0,41,0,254,0,96,0,81,0,158,0,195,0,245,0,131,0,101,0,10,0,134,0,50,0,213,0,224,0,62,0,0,0,0,0,0,0,218,0,238,0,0,0,168,0,0,0,16,0,0,0,143,0,201,0,66,0,26,0,158,0,138,0,149,0,176,0,234,0,11,0,64,0,219,0,24,0,3,0,247,0,114,0,0,0,129,0,109,0,147,0,193,0,4,0,74,0,133,0,0,0,12,0,146,0,145,0,225,0,4,0,74,0,0,0,90,0,219,0,0,0,111,0,233,0,156,0,0,0,0,0,187,0,150,0,0,0,0,0,87,0,232,0,165,0,78,0,0,0,144,0,150,0,25,0,201,0,74,0,68,0,67,0,4,0,0,0,101,0,220,0,163,0,0,0,13,0,0,0,141,0,253,0,163,0,0,0,4,0,9,0,33,0,0,0,217,0,154,0,72,0,0,0,94,0,127,0,82,0,252,0,233,0,0,0,32,0,21,0,0,0,123,0,7,0,55,0,0,0,214,0,0,0,28,0,36,0,0,0,110,0,195,0,58,0,45,0,0,0,82,0,86,0,159,0,72,0,0,0,0,0,54,0,167,0,0,0,79,0,93,0,4,0,24,0,200,0,21,0,254,0,167,0,98,0,94,0,90,0,63,0,51,0,199,0,85,0,62,0,114,0,0,0,152,0,77,0,231,0,0,0,41,0,0,0,234,0,29,0,104,0,0,0,230,0,129,0,201,0,3,0,186,0,140,0,246,0,50,0,203,0,149,0,136,0,180,0,212,0,122,0,193,0,104,0,87,0,104,0,63,0,153,0,164,0,193,0,72,0,119,0,166,0,0,0,236,0,239,0,114,0,0,0,0,0,209,0,81,0,46,0,237,0,0,0,0,0,53,0,249,0,209,0,197,0,219,0,230,0,0,0,210,0,221,0,109,0,0,0,0,0,55,0,207,0,250,0,141,0,252,0,64,0,106,0,161,0,235,0,0,0,190,0,63,0,112,0,3,0,241,0,16,0,118,0,71,0,102,0,99,0,62,0,195,0,178,0,0,0,174,0,207,0,236,0,131,0,144,0,142,0,247,0,15,0,146,0,255,0,108,0,0,0,92,0,90,0,91,0,229,0,173,0,37,0,0,0,113,0,0,0,127,0,34,0,0,0,76,0,18,0,0,0,0,0,255,0,129,0,238,0,0,0,200,0,190,0,184,0,217,0,107,0,95,0,70,0,41,0,8,0,0,0,68,0,107,0,0,0,218,0,8,0,68,0,0,0,118,0,253,0,88,0,161,0,134,0,142,0,192,0,88,0);
signal scenario_full  : scenario_type := (245,31,116,31,125,31,194,31,134,31,17,31,23,31,23,30,13,31,13,30,101,31,39,31,26,31,68,31,130,31,205,31,56,31,197,31,182,31,174,31,35,31,35,31,35,30,35,29,30,31,12,31,161,31,62,31,164,31,164,30,34,31,173,31,200,31,220,31,40,31,40,30,102,31,102,30,102,29,211,31,211,30,179,31,125,31,18,31,104,31,136,31,206,31,35,31,241,31,226,31,226,30,33,31,127,31,62,31,229,31,253,31,48,31,137,31,58,31,62,31,255,31,223,31,122,31,55,31,29,31,190,31,128,31,217,31,105,31,234,31,55,31,20,31,29,31,1,31,1,30,97,31,222,31,34,31,34,30,122,31,150,31,87,31,202,31,249,31,249,30,132,31,26,31,56,31,142,31,183,31,63,31,168,31,255,31,233,31,82,31,177,31,177,30,177,29,185,31,201,31,66,31,246,31,210,31,119,31,17,31,170,31,170,30,24,31,136,31,73,31,242,31,28,31,28,30,49,31,193,31,147,31,218,31,8,31,206,31,206,30,95,31,95,30,95,29,95,28,11,31,73,31,116,31,156,31,226,31,226,30,186,31,91,31,247,31,123,31,207,31,119,31,226,31,57,31,180,31,35,31,108,31,108,30,100,31,100,30,5,31,5,30,5,29,16,31,27,31,27,30,93,31,249,31,208,31,230,31,23,31,254,31,254,30,230,31,228,31,228,30,110,31,141,31,238,31,238,30,93,31,166,31,166,30,220,31,57,31,2,31,37,31,37,30,146,31,146,30,223,31,233,31,14,31,50,31,150,31,242,31,142,31,142,30,226,31,247,31,46,31,18,31,26,31,121,31,185,31,6,31,6,30,9,31,45,31,11,31,154,31,34,31,219,31,86,31,215,31,244,31,244,30,238,31,238,30,238,29,248,31,248,30,236,31,192,31,144,31,156,31,60,31,3,31,44,31,117,31,117,30,219,31,208,31,39,31,95,31,61,31,218,31,218,30,4,31,50,31,13,31,161,31,47,31,212,31,123,31,123,30,133,31,133,30,133,29,163,31,196,31,196,30,185,31,185,30,163,31,224,31,108,31,214,31,204,31,204,30,191,31,252,31,206,31,141,31,75,31,26,31,26,30,67,31,67,30,250,31,51,31,228,31,230,31,153,31,199,31,181,31,68,31,221,31,221,30,206,31,23,31,248,31,83,31,211,31,211,30,211,29,206,31,34,31,40,31,40,30,133,31,2,31,2,30,130,31,130,30,1,31,112,31,112,30,112,29,79,31,89,31,89,30,89,29,212,31,27,31,27,30,233,31,209,31,209,30,209,29,252,31,232,31,114,31,98,31,129,31,204,31,73,31,73,30,27,31,111,31,69,31,137,31,231,31,198,31,175,31,175,30,102,31,108,31,233,31,131,31,65,31,218,31,72,31,208,31,61,31,24,31,102,31,102,30,81,31,229,31,229,30,229,29,252,31,61,31,214,31,234,31,45,31,75,31,130,31,130,30,34,31,2,31,2,30,243,31,255,31,188,31,188,30,250,31,162,31,177,31,236,31,44,31,82,31,82,31,139,31,133,31,212,31,171,31,24,31,52,31,106,31,118,31,30,31,194,31,191,31,217,31,156,31,156,30,100,31,60,31,60,30,193,31,174,31,86,31,40,31,161,31,92,31,92,30,102,31,190,31,190,30,94,31,62,31,188,31,190,31,77,31,95,31,83,31,221,31,232,31,232,30,201,31,87,31,136,31,58,31,106,31,191,31,191,30,61,31,211,31,211,30,117,31,52,31,156,31,168,31,210,31,210,30,155,31,155,30,31,31,88,31,88,30,176,31,13,31,252,31,252,30,58,31,177,31,198,31,198,30,198,29,219,31,219,30,30,31,30,30,105,31,110,31,108,31,131,31,103,31,162,31,142,31,25,31,25,30,25,29,239,31,196,31,120,31,196,31,10,31,230,31,230,30,6,31,175,31,175,30,134,31,121,31,89,31,211,31,118,31,118,30,51,31,61,31,61,30,159,31,30,31,250,31,211,31,211,30,22,31,206,31,17,31,157,31,108,31,194,31,29,31,21,31,96,31,159,31,175,31,72,31,80,31,80,30,20,31,208,31,6,31,6,30,31,31,186,31,216,31,187,31,94,31,144,31,228,31,170,31,117,31,15,31,62,31,62,30,3,31,3,30,90,31,193,31,234,31,234,30,71,31,127,31,77,31,149,31,61,31,61,30,233,31,233,30,47,31,47,30,47,29,160,31,42,31,128,31,128,30,203,31,64,31,64,30,5,31,233,31,140,31,34,31,140,31,99,31,186,31,44,31,188,31,160,31,226,31,96,31,62,31,162,31,161,31,229,31,161,31,161,30,105,31,21,31,14,31,159,31,159,30,53,31,252,31,252,30,12,31,74,31,70,31,222,31,41,31,41,30,63,31,98,31,78,31,23,31,38,31,62,31,33,31,201,31,201,30,135,31,136,31,23,31,22,31,70,31,117,31,22,31,144,31,144,30,139,31,153,31,137,31,137,30,158,31,136,31,74,31,88,31,8,31,140,31,44,31,247,31,247,30,204,31,165,31,13,31,13,30,223,31,241,31,167,31,232,31,60,31,80,31,181,31,181,30,181,29,132,31,49,31,41,31,123,31,123,30,199,31,61,31,239,31,227,31,100,31,92,31,54,31,190,31,24,31,10,31,215,31,157,31,161,31,176,31,176,30,86,31,73,31,66,31,102,31,230,31,125,31,125,30,36,31,234,31,123,31,123,30,123,29,255,31,255,30,26,31,89,31,41,31,254,31,96,31,81,31,158,31,195,31,245,31,131,31,101,31,10,31,134,31,50,31,213,31,224,31,62,31,62,30,62,29,62,28,218,31,238,31,238,30,168,31,168,30,16,31,16,30,143,31,201,31,66,31,26,31,158,31,138,31,149,31,176,31,234,31,11,31,64,31,219,31,24,31,3,31,247,31,114,31,114,30,129,31,109,31,147,31,193,31,4,31,74,31,133,31,133,30,12,31,146,31,145,31,225,31,4,31,74,31,74,30,90,31,219,31,219,30,111,31,233,31,156,31,156,30,156,29,187,31,150,31,150,30,150,29,87,31,232,31,165,31,78,31,78,30,144,31,150,31,25,31,201,31,74,31,68,31,67,31,4,31,4,30,101,31,220,31,163,31,163,30,13,31,13,30,141,31,253,31,163,31,163,30,4,31,9,31,33,31,33,30,217,31,154,31,72,31,72,30,94,31,127,31,82,31,252,31,233,31,233,30,32,31,21,31,21,30,123,31,7,31,55,31,55,30,214,31,214,30,28,31,36,31,36,30,110,31,195,31,58,31,45,31,45,30,82,31,86,31,159,31,72,31,72,30,72,29,54,31,167,31,167,30,79,31,93,31,4,31,24,31,200,31,21,31,254,31,167,31,98,31,94,31,90,31,63,31,51,31,199,31,85,31,62,31,114,31,114,30,152,31,77,31,231,31,231,30,41,31,41,30,234,31,29,31,104,31,104,30,230,31,129,31,201,31,3,31,186,31,140,31,246,31,50,31,203,31,149,31,136,31,180,31,212,31,122,31,193,31,104,31,87,31,104,31,63,31,153,31,164,31,193,31,72,31,119,31,166,31,166,30,236,31,239,31,114,31,114,30,114,29,209,31,81,31,46,31,237,31,237,30,237,29,53,31,249,31,209,31,197,31,219,31,230,31,230,30,210,31,221,31,109,31,109,30,109,29,55,31,207,31,250,31,141,31,252,31,64,31,106,31,161,31,235,31,235,30,190,31,63,31,112,31,3,31,241,31,16,31,118,31,71,31,102,31,99,31,62,31,195,31,178,31,178,30,174,31,207,31,236,31,131,31,144,31,142,31,247,31,15,31,146,31,255,31,108,31,108,30,92,31,90,31,91,31,229,31,173,31,37,31,37,30,113,31,113,30,127,31,34,31,34,30,76,31,18,31,18,30,18,29,255,31,129,31,238,31,238,30,200,31,190,31,184,31,217,31,107,31,95,31,70,31,41,31,8,31,8,30,68,31,107,31,107,30,218,31,8,31,68,31,68,30,118,31,253,31,88,31,161,31,134,31,142,31,192,31,88,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
