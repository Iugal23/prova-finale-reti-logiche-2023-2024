-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 365;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,195,0,97,0,34,0,111,0,156,0,222,0,106,0,0,0,56,0,204,0,86,0,132,0,56,0,158,0,54,0,157,0,254,0,54,0,0,0,229,0,208,0,121,0,254,0,13,0,62,0,66,0,252,0,0,0,174,0,0,0,212,0,176,0,142,0,180,0,162,0,118,0,249,0,0,0,162,0,0,0,0,0,0,0,223,0,246,0,110,0,0,0,139,0,157,0,238,0,0,0,79,0,229,0,0,0,165,0,74,0,108,0,241,0,138,0,101,0,3,0,183,0,20,0,156,0,234,0,197,0,67,0,0,0,6,0,147,0,209,0,223,0,192,0,154,0,34,0,140,0,20,0,47,0,135,0,91,0,69,0,76,0,45,0,255,0,0,0,101,0,85,0,175,0,60,0,247,0,0,0,0,0,250,0,232,0,0,0,63,0,142,0,172,0,54,0,50,0,242,0,125,0,179,0,77,0,0,0,45,0,153,0,59,0,39,0,159,0,50,0,176,0,6,0,152,0,24,0,46,0,112,0,130,0,102,0,193,0,200,0,101,0,21,0,10,0,239,0,130,0,0,0,55,0,201,0,227,0,120,0,0,0,254,0,0,0,219,0,177,0,204,0,199,0,4,0,211,0,92,0,253,0,0,0,0,0,0,0,228,0,236,0,0,0,0,0,181,0,159,0,210,0,33,0,0,0,56,0,120,0,58,0,2,0,130,0,0,0,241,0,119,0,71,0,183,0,46,0,244,0,188,0,0,0,47,0,179,0,31,0,65,0,0,0,0,0,99,0,249,0,212,0,95,0,0,0,0,0,170,0,0,0,0,0,93,0,57,0,0,0,70,0,189,0,233,0,182,0,227,0,0,0,205,0,69,0,0,0,147,0,161,0,0,0,187,0,214,0,187,0,78,0,194,0,13,0,0,0,194,0,68,0,4,0,27,0,0,0,99,0,0,0,249,0,30,0,93,0,91,0,141,0,0,0,77,0,160,0,10,0,49,0,86,0,48,0,95,0,91,0,0,0,227,0,74,0,0,0,0,0,0,0,233,0,181,0,0,0,201,0,182,0,23,0,228,0,216,0,238,0,76,0,60,0,150,0,127,0,0,0,142,0,0,0,186,0,234,0,251,0,76,0,96,0,71,0,0,0,0,0,152,0,0,0,204,0,40,0,0,0,32,0,2,0,45,0,0,0,202,0,17,0,0,0,161,0,225,0,15,0,0,0,134,0,0,0,121,0,196,0,0,0,0,0,17,0,94,0,182,0,127,0,37,0,94,0,222,0,50,0,0,0,2,0,146,0,165,0,92,0,206,0,17,0,191,0,57,0,124,0,35,0,100,0,199,0,0,0,0,0,0,0,0,0,176,0,41,0,43,0,205,0,70,0,122,0,0,0,171,0,63,0,75,0,150,0,9,0,0,0,77,0,89,0,0,0,128,0,0,0,15,0,119,0,72,0,0,0,0,0,135,0,219,0,200,0,166,0,174,0,207,0,0,0,76,0,138,0,107,0,159,0,102,0,206,0,175,0,0,0,157,0,66,0,161,0,213,0,0,0,0,0,238,0,163,0,203,0,208,0,142,0,163,0,0,0,175,0,113,0,254,0,0,0,206,0,47,0,37,0,84,0,249,0,83,0,76,0);
signal scenario_full  : scenario_type := (0,0,195,31,97,31,34,31,111,31,156,31,222,31,106,31,106,30,56,31,204,31,86,31,132,31,56,31,158,31,54,31,157,31,254,31,54,31,54,30,229,31,208,31,121,31,254,31,13,31,62,31,66,31,252,31,252,30,174,31,174,30,212,31,176,31,142,31,180,31,162,31,118,31,249,31,249,30,162,31,162,30,162,29,162,28,223,31,246,31,110,31,110,30,139,31,157,31,238,31,238,30,79,31,229,31,229,30,165,31,74,31,108,31,241,31,138,31,101,31,3,31,183,31,20,31,156,31,234,31,197,31,67,31,67,30,6,31,147,31,209,31,223,31,192,31,154,31,34,31,140,31,20,31,47,31,135,31,91,31,69,31,76,31,45,31,255,31,255,30,101,31,85,31,175,31,60,31,247,31,247,30,247,29,250,31,232,31,232,30,63,31,142,31,172,31,54,31,50,31,242,31,125,31,179,31,77,31,77,30,45,31,153,31,59,31,39,31,159,31,50,31,176,31,6,31,152,31,24,31,46,31,112,31,130,31,102,31,193,31,200,31,101,31,21,31,10,31,239,31,130,31,130,30,55,31,201,31,227,31,120,31,120,30,254,31,254,30,219,31,177,31,204,31,199,31,4,31,211,31,92,31,253,31,253,30,253,29,253,28,228,31,236,31,236,30,236,29,181,31,159,31,210,31,33,31,33,30,56,31,120,31,58,31,2,31,130,31,130,30,241,31,119,31,71,31,183,31,46,31,244,31,188,31,188,30,47,31,179,31,31,31,65,31,65,30,65,29,99,31,249,31,212,31,95,31,95,30,95,29,170,31,170,30,170,29,93,31,57,31,57,30,70,31,189,31,233,31,182,31,227,31,227,30,205,31,69,31,69,30,147,31,161,31,161,30,187,31,214,31,187,31,78,31,194,31,13,31,13,30,194,31,68,31,4,31,27,31,27,30,99,31,99,30,249,31,30,31,93,31,91,31,141,31,141,30,77,31,160,31,10,31,49,31,86,31,48,31,95,31,91,31,91,30,227,31,74,31,74,30,74,29,74,28,233,31,181,31,181,30,201,31,182,31,23,31,228,31,216,31,238,31,76,31,60,31,150,31,127,31,127,30,142,31,142,30,186,31,234,31,251,31,76,31,96,31,71,31,71,30,71,29,152,31,152,30,204,31,40,31,40,30,32,31,2,31,45,31,45,30,202,31,17,31,17,30,161,31,225,31,15,31,15,30,134,31,134,30,121,31,196,31,196,30,196,29,17,31,94,31,182,31,127,31,37,31,94,31,222,31,50,31,50,30,2,31,146,31,165,31,92,31,206,31,17,31,191,31,57,31,124,31,35,31,100,31,199,31,199,30,199,29,199,28,199,27,176,31,41,31,43,31,205,31,70,31,122,31,122,30,171,31,63,31,75,31,150,31,9,31,9,30,77,31,89,31,89,30,128,31,128,30,15,31,119,31,72,31,72,30,72,29,135,31,219,31,200,31,166,31,174,31,207,31,207,30,76,31,138,31,107,31,159,31,102,31,206,31,175,31,175,30,157,31,66,31,161,31,213,31,213,30,213,29,238,31,163,31,203,31,208,31,142,31,163,31,163,30,175,31,113,31,254,31,254,30,206,31,47,31,37,31,84,31,249,31,83,31,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
