-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 637;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,72,0,178,0,217,0,217,0,188,0,0,0,0,0,0,0,55,0,188,0,0,0,210,0,98,0,16,0,112,0,18,0,233,0,190,0,198,0,206,0,31,0,0,0,106,0,37,0,169,0,58,0,212,0,90,0,135,0,131,0,211,0,157,0,57,0,146,0,92,0,9,0,71,0,218,0,0,0,182,0,185,0,206,0,0,0,123,0,202,0,132,0,0,0,0,0,172,0,244,0,26,0,90,0,119,0,136,0,0,0,254,0,113,0,82,0,108,0,0,0,236,0,246,0,88,0,9,0,88,0,196,0,225,0,242,0,108,0,234,0,106,0,178,0,0,0,156,0,237,0,3,0,48,0,0,0,17,0,25,0,106,0,0,0,224,0,8,0,0,0,100,0,56,0,216,0,16,0,0,0,222,0,0,0,9,0,0,0,0,0,0,0,194,0,0,0,18,0,163,0,244,0,0,0,0,0,150,0,35,0,45,0,204,0,245,0,157,0,125,0,0,0,0,0,138,0,154,0,132,0,190,0,122,0,0,0,168,0,231,0,0,0,0,0,242,0,195,0,27,0,0,0,140,0,0,0,201,0,146,0,110,0,205,0,152,0,59,0,94,0,123,0,0,0,176,0,40,0,130,0,52,0,223,0,189,0,7,0,96,0,123,0,62,0,80,0,0,0,199,0,179,0,181,0,88,0,203,0,202,0,25,0,173,0,146,0,46,0,66,0,69,0,42,0,203,0,209,0,187,0,0,0,0,0,123,0,0,0,104,0,72,0,0,0,196,0,144,0,222,0,206,0,139,0,66,0,146,0,0,0,5,0,74,0,157,0,0,0,237,0,117,0,87,0,137,0,0,0,52,0,61,0,86,0,250,0,213,0,0,0,0,0,70,0,0,0,0,0,33,0,7,0,246,0,112,0,46,0,151,0,42,0,35,0,158,0,94,0,10,0,0,0,128,0,0,0,81,0,79,0,205,0,248,0,0,0,22,0,6,0,0,0,0,0,0,0,253,0,143,0,206,0,0,0,237,0,24,0,101,0,0,0,0,0,138,0,105,0,0,0,0,0,176,0,74,0,170,0,120,0,79,0,156,0,0,0,0,0,0,0,117,0,40,0,11,0,134,0,132,0,40,0,0,0,105,0,14,0,217,0,129,0,174,0,43,0,0,0,48,0,85,0,215,0,3,0,175,0,215,0,176,0,0,0,41,0,5,0,251,0,76,0,161,0,83,0,22,0,173,0,214,0,173,0,133,0,42,0,169,0,253,0,224,0,190,0,133,0,220,0,199,0,0,0,0,0,160,0,177,0,98,0,201,0,113,0,157,0,68,0,173,0,32,0,0,0,101,0,209,0,96,0,236,0,123,0,0,0,7,0,172,0,20,0,102,0,78,0,225,0,107,0,3,0,83,0,194,0,20,0,9,0,216,0,232,0,40,0,48,0,194,0,86,0,13,0,243,0,0,0,182,0,0,0,134,0,0,0,0,0,245,0,178,0,0,0,48,0,179,0,222,0,232,0,194,0,16,0,0,0,98,0,115,0,57,0,50,0,178,0,39,0,131,0,233,0,21,0,188,0,190,0,194,0,54,0,224,0,71,0,82,0,173,0,0,0,238,0,175,0,59,0,238,0,63,0,87,0,181,0,37,0,0,0,125,0,23,0,201,0,220,0,0,0,108,0,217,0,154,0,0,0,0,0,0,0,0,0,6,0,102,0,0,0,48,0,16,0,197,0,0,0,39,0,226,0,99,0,163,0,253,0,29,0,246,0,0,0,33,0,128,0,191,0,145,0,160,0,0,0,153,0,0,0,95,0,0,0,0,0,48,0,249,0,169,0,119,0,240,0,135,0,0,0,244,0,0,0,96,0,0,0,18,0,86,0,161,0,133,0,74,0,97,0,119,0,51,0,179,0,229,0,83,0,217,0,206,0,0,0,64,0,0,0,17,0,0,0,190,0,134,0,234,0,0,0,74,0,98,0,211,0,5,0,61,0,53,0,0,0,147,0,45,0,121,0,89,0,206,0,228,0,188,0,6,0,200,0,0,0,37,0,227,0,176,0,50,0,225,0,196,0,16,0,171,0,1,0,175,0,0,0,36,0,203,0,72,0,0,0,136,0,44,0,169,0,54,0,33,0,208,0,239,0,184,0,124,0,9,0,36,0,0,0,219,0,137,0,208,0,154,0,0,0,106,0,0,0,85,0,147,0,59,0,0,0,0,0,234,0,175,0,106,0,215,0,57,0,238,0,166,0,100,0,240,0,234,0,27,0,115,0,165,0,176,0,237,0,0,0,0,0,0,0,0,0,115,0,0,0,165,0,99,0,114,0,224,0,91,0,201,0,42,0,0,0,0,0,140,0,7,0,201,0,96,0,180,0,224,0,9,0,215,0,128,0,0,0,151,0,30,0,192,0,210,0,117,0,0,0,232,0,0,0,131,0,76,0,97,0,56,0,137,0,0,0,171,0,73,0,188,0,124,0,252,0,105,0,201,0,43,0,154,0,2,0,203,0,206,0,0,0,67,0,159,0,0,0,0,0,0,0,0,0,22,0,73,0,219,0,94,0,0,0,0,0,0,0,205,0,0,0,210,0,24,0,95,0,34,0,22,0,38,0,211,0,143,0,170,0,0,0,21,0,54,0,176,0,45,0,233,0,55,0,0,0,224,0,57,0,130,0,100,0,214,0,207,0,64,0,79,0,222,0,206,0,0,0,141,0,5,0,223,0,0,0,46,0,248,0,212,0,81,0,0,0,37,0,0,0,158,0,130,0,26,0,54,0,36,0,250,0,166,0,146,0,25,0,45,0,75,0,54,0,182,0,0,0,252,0,29,0,53,0,157,0,178,0,0,0,38,0);
signal scenario_full  : scenario_type := (0,0,72,31,178,31,217,31,217,31,188,31,188,30,188,29,188,28,55,31,188,31,188,30,210,31,98,31,16,31,112,31,18,31,233,31,190,31,198,31,206,31,31,31,31,30,106,31,37,31,169,31,58,31,212,31,90,31,135,31,131,31,211,31,157,31,57,31,146,31,92,31,9,31,71,31,218,31,218,30,182,31,185,31,206,31,206,30,123,31,202,31,132,31,132,30,132,29,172,31,244,31,26,31,90,31,119,31,136,31,136,30,254,31,113,31,82,31,108,31,108,30,236,31,246,31,88,31,9,31,88,31,196,31,225,31,242,31,108,31,234,31,106,31,178,31,178,30,156,31,237,31,3,31,48,31,48,30,17,31,25,31,106,31,106,30,224,31,8,31,8,30,100,31,56,31,216,31,16,31,16,30,222,31,222,30,9,31,9,30,9,29,9,28,194,31,194,30,18,31,163,31,244,31,244,30,244,29,150,31,35,31,45,31,204,31,245,31,157,31,125,31,125,30,125,29,138,31,154,31,132,31,190,31,122,31,122,30,168,31,231,31,231,30,231,29,242,31,195,31,27,31,27,30,140,31,140,30,201,31,146,31,110,31,205,31,152,31,59,31,94,31,123,31,123,30,176,31,40,31,130,31,52,31,223,31,189,31,7,31,96,31,123,31,62,31,80,31,80,30,199,31,179,31,181,31,88,31,203,31,202,31,25,31,173,31,146,31,46,31,66,31,69,31,42,31,203,31,209,31,187,31,187,30,187,29,123,31,123,30,104,31,72,31,72,30,196,31,144,31,222,31,206,31,139,31,66,31,146,31,146,30,5,31,74,31,157,31,157,30,237,31,117,31,87,31,137,31,137,30,52,31,61,31,86,31,250,31,213,31,213,30,213,29,70,31,70,30,70,29,33,31,7,31,246,31,112,31,46,31,151,31,42,31,35,31,158,31,94,31,10,31,10,30,128,31,128,30,81,31,79,31,205,31,248,31,248,30,22,31,6,31,6,30,6,29,6,28,253,31,143,31,206,31,206,30,237,31,24,31,101,31,101,30,101,29,138,31,105,31,105,30,105,29,176,31,74,31,170,31,120,31,79,31,156,31,156,30,156,29,156,28,117,31,40,31,11,31,134,31,132,31,40,31,40,30,105,31,14,31,217,31,129,31,174,31,43,31,43,30,48,31,85,31,215,31,3,31,175,31,215,31,176,31,176,30,41,31,5,31,251,31,76,31,161,31,83,31,22,31,173,31,214,31,173,31,133,31,42,31,169,31,253,31,224,31,190,31,133,31,220,31,199,31,199,30,199,29,160,31,177,31,98,31,201,31,113,31,157,31,68,31,173,31,32,31,32,30,101,31,209,31,96,31,236,31,123,31,123,30,7,31,172,31,20,31,102,31,78,31,225,31,107,31,3,31,83,31,194,31,20,31,9,31,216,31,232,31,40,31,48,31,194,31,86,31,13,31,243,31,243,30,182,31,182,30,134,31,134,30,134,29,245,31,178,31,178,30,48,31,179,31,222,31,232,31,194,31,16,31,16,30,98,31,115,31,57,31,50,31,178,31,39,31,131,31,233,31,21,31,188,31,190,31,194,31,54,31,224,31,71,31,82,31,173,31,173,30,238,31,175,31,59,31,238,31,63,31,87,31,181,31,37,31,37,30,125,31,23,31,201,31,220,31,220,30,108,31,217,31,154,31,154,30,154,29,154,28,154,27,6,31,102,31,102,30,48,31,16,31,197,31,197,30,39,31,226,31,99,31,163,31,253,31,29,31,246,31,246,30,33,31,128,31,191,31,145,31,160,31,160,30,153,31,153,30,95,31,95,30,95,29,48,31,249,31,169,31,119,31,240,31,135,31,135,30,244,31,244,30,96,31,96,30,18,31,86,31,161,31,133,31,74,31,97,31,119,31,51,31,179,31,229,31,83,31,217,31,206,31,206,30,64,31,64,30,17,31,17,30,190,31,134,31,234,31,234,30,74,31,98,31,211,31,5,31,61,31,53,31,53,30,147,31,45,31,121,31,89,31,206,31,228,31,188,31,6,31,200,31,200,30,37,31,227,31,176,31,50,31,225,31,196,31,16,31,171,31,1,31,175,31,175,30,36,31,203,31,72,31,72,30,136,31,44,31,169,31,54,31,33,31,208,31,239,31,184,31,124,31,9,31,36,31,36,30,219,31,137,31,208,31,154,31,154,30,106,31,106,30,85,31,147,31,59,31,59,30,59,29,234,31,175,31,106,31,215,31,57,31,238,31,166,31,100,31,240,31,234,31,27,31,115,31,165,31,176,31,237,31,237,30,237,29,237,28,237,27,115,31,115,30,165,31,99,31,114,31,224,31,91,31,201,31,42,31,42,30,42,29,140,31,7,31,201,31,96,31,180,31,224,31,9,31,215,31,128,31,128,30,151,31,30,31,192,31,210,31,117,31,117,30,232,31,232,30,131,31,76,31,97,31,56,31,137,31,137,30,171,31,73,31,188,31,124,31,252,31,105,31,201,31,43,31,154,31,2,31,203,31,206,31,206,30,67,31,159,31,159,30,159,29,159,28,159,27,22,31,73,31,219,31,94,31,94,30,94,29,94,28,205,31,205,30,210,31,24,31,95,31,34,31,22,31,38,31,211,31,143,31,170,31,170,30,21,31,54,31,176,31,45,31,233,31,55,31,55,30,224,31,57,31,130,31,100,31,214,31,207,31,64,31,79,31,222,31,206,31,206,30,141,31,5,31,223,31,223,30,46,31,248,31,212,31,81,31,81,30,37,31,37,30,158,31,130,31,26,31,54,31,36,31,250,31,166,31,146,31,25,31,45,31,75,31,54,31,182,31,182,30,252,31,29,31,53,31,157,31,178,31,178,30,38,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
