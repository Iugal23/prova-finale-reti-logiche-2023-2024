-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 960;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,61,0,0,0,118,0,162,0,165,0,165,0,178,0,247,0,156,0,97,0,234,0,173,0,244,0,94,0,19,0,46,0,193,0,2,0,69,0,66,0,159,0,185,0,121,0,58,0,0,0,128,0,185,0,7,0,123,0,188,0,27,0,228,0,0,0,0,0,180,0,142,0,0,0,166,0,183,0,206,0,107,0,80,0,117,0,22,0,0,0,51,0,32,0,59,0,152,0,46,0,236,0,136,0,88,0,248,0,98,0,112,0,121,0,128,0,113,0,58,0,35,0,27,0,184,0,49,0,204,0,208,0,77,0,97,0,86,0,0,0,133,0,162,0,0,0,163,0,0,0,173,0,163,0,223,0,17,0,0,0,0,0,187,0,41,0,94,0,0,0,139,0,209,0,133,0,244,0,107,0,184,0,61,0,170,0,141,0,133,0,56,0,100,0,120,0,180,0,42,0,176,0,86,0,192,0,29,0,0,0,0,0,91,0,228,0,0,0,197,0,0,0,156,0,135,0,97,0,112,0,232,0,206,0,150,0,250,0,246,0,0,0,0,0,197,0,169,0,0,0,154,0,157,0,125,0,102,0,172,0,99,0,97,0,83,0,54,0,0,0,75,0,83,0,71,0,153,0,207,0,71,0,25,0,230,0,0,0,120,0,233,0,24,0,110,0,204,0,198,0,12,0,100,0,36,0,106,0,232,0,253,0,147,0,0,0,0,0,0,0,0,0,44,0,154,0,238,0,111,0,70,0,40,0,169,0,141,0,106,0,0,0,36,0,193,0,0,0,146,0,31,0,96,0,221,0,161,0,0,0,217,0,71,0,13,0,145,0,17,0,246,0,102,0,23,0,174,0,206,0,0,0,20,0,240,0,36,0,49,0,145,0,0,0,10,0,82,0,236,0,14,0,0,0,31,0,90,0,0,0,184,0,157,0,210,0,73,0,0,0,127,0,98,0,58,0,188,0,20,0,127,0,125,0,0,0,154,0,0,0,9,0,176,0,173,0,200,0,112,0,0,0,0,0,140,0,49,0,107,0,110,0,232,0,93,0,184,0,0,0,0,0,153,0,14,0,201,0,0,0,121,0,19,0,90,0,171,0,177,0,95,0,243,0,72,0,134,0,202,0,247,0,26,0,212,0,229,0,179,0,58,0,15,0,88,0,33,0,100,0,218,0,0,0,207,0,0,0,83,0,217,0,113,0,87,0,0,0,240,0,26,0,234,0,243,0,121,0,0,0,250,0,222,0,152,0,0,0,16,0,0,0,241,0,0,0,0,0,187,0,1,0,0,0,95,0,0,0,218,0,87,0,108,0,67,0,0,0,45,0,107,0,243,0,225,0,178,0,6,0,68,0,51,0,100,0,54,0,0,0,0,0,165,0,113,0,236,0,0,0,175,0,153,0,108,0,0,0,0,0,225,0,219,0,240,0,126,0,242,0,68,0,34,0,0,0,0,0,187,0,202,0,47,0,18,0,179,0,0,0,229,0,0,0,126,0,0,0,0,0,24,0,23,0,53,0,0,0,56,0,177,0,131,0,0,0,0,0,0,0,119,0,241,0,150,0,0,0,59,0,2,0,0,0,232,0,90,0,188,0,121,0,90,0,15,0,0,0,0,0,146,0,193,0,75,0,176,0,204,0,250,0,36,0,73,0,224,0,0,0,237,0,186,0,199,0,164,0,0,0,0,0,182,0,14,0,36,0,78,0,0,0,212,0,18,0,113,0,73,0,13,0,0,0,109,0,146,0,215,0,149,0,0,0,90,0,0,0,203,0,10,0,100,0,237,0,0,0,95,0,246,0,232,0,66,0,181,0,164,0,251,0,0,0,108,0,154,0,58,0,0,0,0,0,223,0,0,0,116,0,192,0,146,0,39,0,140,0,123,0,0,0,49,0,233,0,34,0,135,0,0,0,60,0,161,0,230,0,172,0,216,0,26,0,0,0,199,0,253,0,128,0,192,0,66,0,109,0,118,0,38,0,17,0,99,0,0,0,65,0,128,0,57,0,0,0,61,0,0,0,203,0,188,0,0,0,163,0,250,0,71,0,136,0,137,0,152,0,185,0,62,0,64,0,79,0,0,0,133,0,115,0,0,0,254,0,196,0,0,0,148,0,0,0,112,0,147,0,41,0,164,0,77,0,48,0,144,0,0,0,0,0,246,0,121,0,0,0,140,0,25,0,0,0,59,0,146,0,237,0,183,0,0,0,9,0,161,0,0,0,203,0,0,0,243,0,118,0,0,0,11,0,75,0,0,0,0,0,0,0,170,0,0,0,138,0,0,0,131,0,178,0,0,0,13,0,248,0,119,0,0,0,203,0,120,0,0,0,0,0,213,0,147,0,0,0,43,0,142,0,211,0,53,0,0,0,190,0,119,0,159,0,85,0,111,0,254,0,103,0,0,0,38,0,3,0,149,0,0,0,18,0,0,0,143,0,65,0,222,0,0,0,72,0,0,0,159,0,88,0,203,0,180,0,120,0,128,0,0,0,122,0,216,0,78,0,0,0,86,0,0,0,183,0,237,0,159,0,96,0,94,0,111,0,129,0,114,0,8,0,0,0,214,0,28,0,152,0,0,0,128,0,161,0,182,0,211,0,205,0,44,0,49,0,66,0,116,0,226,0,64,0,57,0,144,0,0,0,0,0,210,0,31,0,152,0,0,0,0,0,160,0,0,0,58,0,0,0,201,0,40,0,188,0,72,0,167,0,195,0,222,0,90,0,109,0,10,0,226,0,0,0,203,0,17,0,56,0,187,0,0,0,228,0,108,0,227,0,3,0,226,0,2,0,207,0,8,0,98,0,57,0,7,0,253,0,0,0,131,0,236,0,235,0,96,0,0,0,85,0,13,0,0,0,131,0,1,0,254,0,159,0,235,0,241,0,71,0,247,0,0,0,140,0,241,0,0,0,0,0,216,0,70,0,0,0,89,0,73,0,209,0,253,0,23,0,70,0,23,0,110,0,215,0,44,0,17,0,226,0,87,0,237,0,158,0,0,0,225,0,0,0,244,0,157,0,188,0,47,0,185,0,91,0,29,0,115,0,200,0,218,0,73,0,145,0,170,0,235,0,0,0,223,0,124,0,0,0,0,0,141,0,127,0,99,0,166,0,162,0,66,0,141,0,154,0,84,0,0,0,141,0,45,0,0,0,41,0,225,0,6,0,0,0,218,0,6,0,11,0,0,0,11,0,65,0,0,0,106,0,55,0,22,0,87,0,122,0,243,0,75,0,127,0,3,0,213,0,17,0,84,0,58,0,11,0,83,0,182,0,224,0,22,0,255,0,241,0,135,0,205,0,26,0,0,0,57,0,0,0,117,0,36,0,150,0,179,0,84,0,244,0,98,0,242,0,0,0,18,0,103,0,76,0,0,0,94,0,0,0,0,0,0,0,35,0,66,0,159,0,0,0,52,0,234,0,0,0,242,0,198,0,185,0,0,0,133,0,0,0,105,0,36,0,0,0,0,0,71,0,24,0,142,0,138,0,0,0,209,0,184,0,222,0,238,0,200,0,121,0,0,0,0,0,39,0,227,0,59,0,113,0,0,0,0,0,68,0,151,0,224,0,147,0,58,0,0,0,146,0,245,0,16,0,207,0,23,0,58,0,0,0,171,0,112,0,7,0,229,0,246,0,87,0,3,0,0,0,0,0,68,0,24,0,36,0,254,0,234,0,0,0,101,0,0,0,77,0,77,0,228,0,170,0,235,0,0,0,54,0,168,0,0,0,0,0,203,0,248,0,172,0,22,0,228,0,211,0,32,0,215,0,212,0,107,0,0,0,225,0,21,0,25,0,7,0,206,0,162,0,187,0,11,0,20,0,159,0,39,0,149,0,123,0,96,0,0,0,4,0,224,0,144,0,102,0,102,0,0,0,159,0,217,0,77,0,119,0,17,0,161,0,0,0,230,0,223,0,58,0,102,0,166,0,0,0,119,0,152,0,234,0,5,0,61,0,183,0,0,0,186,0,182,0,38,0,67,0,0,0,95,0,144,0,0,0,10,0,21,0,134,0,0,0,155,0,251,0,85,0,237,0,0,0,0,0,223,0,0,0,155,0,0,0,137,0,107,0,66,0,227,0,46,0,0,0,192,0,0,0,0,0,14,0,43,0,72,0,0,0,180,0,232,0,19,0,138,0,104,0,79,0,13,0,0,0,0,0,0,0,21,0,123,0,170,0,167,0,113,0,59,0,250,0,0,0,0,0,253,0,254,0,0,0,126,0,65,0,15,0,106,0,247,0,78,0,0,0,147,0,43,0,241,0,131,0,166,0,0,0,0,0,166,0,0,0,103,0);
signal scenario_full  : scenario_type := (0,0,61,31,61,30,118,31,162,31,165,31,165,31,178,31,247,31,156,31,97,31,234,31,173,31,244,31,94,31,19,31,46,31,193,31,2,31,69,31,66,31,159,31,185,31,121,31,58,31,58,30,128,31,185,31,7,31,123,31,188,31,27,31,228,31,228,30,228,29,180,31,142,31,142,30,166,31,183,31,206,31,107,31,80,31,117,31,22,31,22,30,51,31,32,31,59,31,152,31,46,31,236,31,136,31,88,31,248,31,98,31,112,31,121,31,128,31,113,31,58,31,35,31,27,31,184,31,49,31,204,31,208,31,77,31,97,31,86,31,86,30,133,31,162,31,162,30,163,31,163,30,173,31,163,31,223,31,17,31,17,30,17,29,187,31,41,31,94,31,94,30,139,31,209,31,133,31,244,31,107,31,184,31,61,31,170,31,141,31,133,31,56,31,100,31,120,31,180,31,42,31,176,31,86,31,192,31,29,31,29,30,29,29,91,31,228,31,228,30,197,31,197,30,156,31,135,31,97,31,112,31,232,31,206,31,150,31,250,31,246,31,246,30,246,29,197,31,169,31,169,30,154,31,157,31,125,31,102,31,172,31,99,31,97,31,83,31,54,31,54,30,75,31,83,31,71,31,153,31,207,31,71,31,25,31,230,31,230,30,120,31,233,31,24,31,110,31,204,31,198,31,12,31,100,31,36,31,106,31,232,31,253,31,147,31,147,30,147,29,147,28,147,27,44,31,154,31,238,31,111,31,70,31,40,31,169,31,141,31,106,31,106,30,36,31,193,31,193,30,146,31,31,31,96,31,221,31,161,31,161,30,217,31,71,31,13,31,145,31,17,31,246,31,102,31,23,31,174,31,206,31,206,30,20,31,240,31,36,31,49,31,145,31,145,30,10,31,82,31,236,31,14,31,14,30,31,31,90,31,90,30,184,31,157,31,210,31,73,31,73,30,127,31,98,31,58,31,188,31,20,31,127,31,125,31,125,30,154,31,154,30,9,31,176,31,173,31,200,31,112,31,112,30,112,29,140,31,49,31,107,31,110,31,232,31,93,31,184,31,184,30,184,29,153,31,14,31,201,31,201,30,121,31,19,31,90,31,171,31,177,31,95,31,243,31,72,31,134,31,202,31,247,31,26,31,212,31,229,31,179,31,58,31,15,31,88,31,33,31,100,31,218,31,218,30,207,31,207,30,83,31,217,31,113,31,87,31,87,30,240,31,26,31,234,31,243,31,121,31,121,30,250,31,222,31,152,31,152,30,16,31,16,30,241,31,241,30,241,29,187,31,1,31,1,30,95,31,95,30,218,31,87,31,108,31,67,31,67,30,45,31,107,31,243,31,225,31,178,31,6,31,68,31,51,31,100,31,54,31,54,30,54,29,165,31,113,31,236,31,236,30,175,31,153,31,108,31,108,30,108,29,225,31,219,31,240,31,126,31,242,31,68,31,34,31,34,30,34,29,187,31,202,31,47,31,18,31,179,31,179,30,229,31,229,30,126,31,126,30,126,29,24,31,23,31,53,31,53,30,56,31,177,31,131,31,131,30,131,29,131,28,119,31,241,31,150,31,150,30,59,31,2,31,2,30,232,31,90,31,188,31,121,31,90,31,15,31,15,30,15,29,146,31,193,31,75,31,176,31,204,31,250,31,36,31,73,31,224,31,224,30,237,31,186,31,199,31,164,31,164,30,164,29,182,31,14,31,36,31,78,31,78,30,212,31,18,31,113,31,73,31,13,31,13,30,109,31,146,31,215,31,149,31,149,30,90,31,90,30,203,31,10,31,100,31,237,31,237,30,95,31,246,31,232,31,66,31,181,31,164,31,251,31,251,30,108,31,154,31,58,31,58,30,58,29,223,31,223,30,116,31,192,31,146,31,39,31,140,31,123,31,123,30,49,31,233,31,34,31,135,31,135,30,60,31,161,31,230,31,172,31,216,31,26,31,26,30,199,31,253,31,128,31,192,31,66,31,109,31,118,31,38,31,17,31,99,31,99,30,65,31,128,31,57,31,57,30,61,31,61,30,203,31,188,31,188,30,163,31,250,31,71,31,136,31,137,31,152,31,185,31,62,31,64,31,79,31,79,30,133,31,115,31,115,30,254,31,196,31,196,30,148,31,148,30,112,31,147,31,41,31,164,31,77,31,48,31,144,31,144,30,144,29,246,31,121,31,121,30,140,31,25,31,25,30,59,31,146,31,237,31,183,31,183,30,9,31,161,31,161,30,203,31,203,30,243,31,118,31,118,30,11,31,75,31,75,30,75,29,75,28,170,31,170,30,138,31,138,30,131,31,178,31,178,30,13,31,248,31,119,31,119,30,203,31,120,31,120,30,120,29,213,31,147,31,147,30,43,31,142,31,211,31,53,31,53,30,190,31,119,31,159,31,85,31,111,31,254,31,103,31,103,30,38,31,3,31,149,31,149,30,18,31,18,30,143,31,65,31,222,31,222,30,72,31,72,30,159,31,88,31,203,31,180,31,120,31,128,31,128,30,122,31,216,31,78,31,78,30,86,31,86,30,183,31,237,31,159,31,96,31,94,31,111,31,129,31,114,31,8,31,8,30,214,31,28,31,152,31,152,30,128,31,161,31,182,31,211,31,205,31,44,31,49,31,66,31,116,31,226,31,64,31,57,31,144,31,144,30,144,29,210,31,31,31,152,31,152,30,152,29,160,31,160,30,58,31,58,30,201,31,40,31,188,31,72,31,167,31,195,31,222,31,90,31,109,31,10,31,226,31,226,30,203,31,17,31,56,31,187,31,187,30,228,31,108,31,227,31,3,31,226,31,2,31,207,31,8,31,98,31,57,31,7,31,253,31,253,30,131,31,236,31,235,31,96,31,96,30,85,31,13,31,13,30,131,31,1,31,254,31,159,31,235,31,241,31,71,31,247,31,247,30,140,31,241,31,241,30,241,29,216,31,70,31,70,30,89,31,73,31,209,31,253,31,23,31,70,31,23,31,110,31,215,31,44,31,17,31,226,31,87,31,237,31,158,31,158,30,225,31,225,30,244,31,157,31,188,31,47,31,185,31,91,31,29,31,115,31,200,31,218,31,73,31,145,31,170,31,235,31,235,30,223,31,124,31,124,30,124,29,141,31,127,31,99,31,166,31,162,31,66,31,141,31,154,31,84,31,84,30,141,31,45,31,45,30,41,31,225,31,6,31,6,30,218,31,6,31,11,31,11,30,11,31,65,31,65,30,106,31,55,31,22,31,87,31,122,31,243,31,75,31,127,31,3,31,213,31,17,31,84,31,58,31,11,31,83,31,182,31,224,31,22,31,255,31,241,31,135,31,205,31,26,31,26,30,57,31,57,30,117,31,36,31,150,31,179,31,84,31,244,31,98,31,242,31,242,30,18,31,103,31,76,31,76,30,94,31,94,30,94,29,94,28,35,31,66,31,159,31,159,30,52,31,234,31,234,30,242,31,198,31,185,31,185,30,133,31,133,30,105,31,36,31,36,30,36,29,71,31,24,31,142,31,138,31,138,30,209,31,184,31,222,31,238,31,200,31,121,31,121,30,121,29,39,31,227,31,59,31,113,31,113,30,113,29,68,31,151,31,224,31,147,31,58,31,58,30,146,31,245,31,16,31,207,31,23,31,58,31,58,30,171,31,112,31,7,31,229,31,246,31,87,31,3,31,3,30,3,29,68,31,24,31,36,31,254,31,234,31,234,30,101,31,101,30,77,31,77,31,228,31,170,31,235,31,235,30,54,31,168,31,168,30,168,29,203,31,248,31,172,31,22,31,228,31,211,31,32,31,215,31,212,31,107,31,107,30,225,31,21,31,25,31,7,31,206,31,162,31,187,31,11,31,20,31,159,31,39,31,149,31,123,31,96,31,96,30,4,31,224,31,144,31,102,31,102,31,102,30,159,31,217,31,77,31,119,31,17,31,161,31,161,30,230,31,223,31,58,31,102,31,166,31,166,30,119,31,152,31,234,31,5,31,61,31,183,31,183,30,186,31,182,31,38,31,67,31,67,30,95,31,144,31,144,30,10,31,21,31,134,31,134,30,155,31,251,31,85,31,237,31,237,30,237,29,223,31,223,30,155,31,155,30,137,31,107,31,66,31,227,31,46,31,46,30,192,31,192,30,192,29,14,31,43,31,72,31,72,30,180,31,232,31,19,31,138,31,104,31,79,31,13,31,13,30,13,29,13,28,21,31,123,31,170,31,167,31,113,31,59,31,250,31,250,30,250,29,253,31,254,31,254,30,126,31,65,31,15,31,106,31,247,31,78,31,78,30,147,31,43,31,241,31,131,31,166,31,166,30,166,29,166,31,166,30,103,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
