-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_480 is
end project_tb_480;

architecture project_tb_arch_480 of project_tb_480 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 485;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (210,0,218,0,37,0,240,0,0,0,65,0,196,0,53,0,0,0,0,0,240,0,222,0,112,0,18,0,132,0,214,0,25,0,218,0,128,0,158,0,0,0,235,0,107,0,0,0,30,0,7,0,95,0,0,0,203,0,186,0,0,0,23,0,18,0,42,0,0,0,163,0,67,0,136,0,211,0,246,0,194,0,24,0,208,0,190,0,0,0,240,0,193,0,80,0,111,0,10,0,25,0,169,0,0,0,68,0,206,0,166,0,82,0,201,0,74,0,43,0,107,0,197,0,23,0,0,0,185,0,31,0,93,0,182,0,150,0,0,0,1,0,234,0,25,0,99,0,214,0,160,0,252,0,0,0,0,0,204,0,82,0,221,0,18,0,69,0,121,0,122,0,45,0,0,0,200,0,114,0,219,0,0,0,134,0,233,0,191,0,52,0,151,0,9,0,151,0,102,0,0,0,156,0,15,0,80,0,0,0,22,0,144,0,214,0,192,0,84,0,0,0,197,0,0,0,113,0,246,0,36,0,27,0,185,0,235,0,47,0,0,0,220,0,187,0,249,0,234,0,191,0,195,0,0,0,81,0,0,0,62,0,0,0,0,0,208,0,47,0,0,0,0,0,7,0,0,0,147,0,97,0,255,0,0,0,70,0,241,0,32,0,209,0,0,0,0,0,223,0,56,0,16,0,244,0,203,0,161,0,85,0,0,0,25,0,2,0,57,0,255,0,35,0,10,0,19,0,244,0,125,0,248,0,10,0,36,0,241,0,47,0,0,0,69,0,249,0,125,0,49,0,0,0,191,0,0,0,206,0,0,0,63,0,96,0,0,0,128,0,0,0,0,0,91,0,0,0,247,0,101,0,3,0,252,0,252,0,78,0,41,0,117,0,122,0,86,0,145,0,148,0,0,0,153,0,19,0,203,0,238,0,110,0,155,0,53,0,28,0,0,0,0,0,127,0,62,0,131,0,248,0,97,0,178,0,212,0,0,0,135,0,250,0,127,0,158,0,103,0,13,0,25,0,73,0,108,0,120,0,24,0,29,0,112,0,184,0,144,0,0,0,77,0,0,0,165,0,87,0,99,0,50,0,1,0,85,0,130,0,31,0,13,0,21,0,0,0,253,0,214,0,79,0,0,0,210,0,78,0,212,0,243,0,0,0,195,0,0,0,239,0,0,0,0,0,251,0,170,0,162,0,230,0,67,0,157,0,33,0,244,0,23,0,190,0,209,0,116,0,153,0,106,0,100,0,96,0,131,0,0,0,0,0,128,0,42,0,44,0,145,0,0,0,151,0,42,0,253,0,0,0,5,0,131,0,0,0,154,0,185,0,165,0,40,0,0,0,0,0,141,0,166,0,63,0,68,0,94,0,0,0,83,0,226,0,0,0,250,0,228,0,214,0,212,0,199,0,168,0,1,0,7,0,161,0,0,0,0,0,0,0,176,0,0,0,45,0,238,0,0,0,254,0,130,0,0,0,147,0,20,0,37,0,159,0,95,0,149,0,0,0,60,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,123,0,170,0,0,0,67,0,22,0,166,0,210,0,150,0,176,0,44,0,219,0,141,0,250,0,97,0,159,0,107,0,27,0,45,0,244,0,43,0,221,0,89,0,41,0,51,0,184,0,0,0,123,0,77,0,163,0,242,0,64,0,13,0,0,0,0,0,125,0,81,0,0,0,201,0,68,0,43,0,2,0,183,0,117,0,0,0,170,0,101,0,107,0,242,0,0,0,237,0,0,0,78,0,250,0,135,0,157,0,83,0,40,0,93,0,0,0,190,0,62,0,142,0,90,0,214,0,189,0,84,0,207,0,215,0,254,0,34,0,215,0,88,0,204,0,0,0,95,0,0,0,26,0,0,0,184,0,109,0,200,0,18,0,112,0,213,0,219,0,158,0,224,0,112,0,0,0,0,0,81,0,88,0,98,0,0,0,0,0,172,0,35,0,0,0,104,0,176,0,0,0,0,0,165,0,0,0,0,0,66,0,14,0,104,0,196,0,181,0,86,0,0,0,99,0,3,0,100,0,178,0,0,0,185,0,0,0,129,0,224,0,28,0,217,0,207,0,187,0,172,0,196,0,0,0,157,0,137,0,80,0,0,0,18,0,0,0,152,0,49,0,209,0,224,0,18,0,0,0,224,0);
signal scenario_full  : scenario_type := (210,31,218,31,37,31,240,31,240,30,65,31,196,31,53,31,53,30,53,29,240,31,222,31,112,31,18,31,132,31,214,31,25,31,218,31,128,31,158,31,158,30,235,31,107,31,107,30,30,31,7,31,95,31,95,30,203,31,186,31,186,30,23,31,18,31,42,31,42,30,163,31,67,31,136,31,211,31,246,31,194,31,24,31,208,31,190,31,190,30,240,31,193,31,80,31,111,31,10,31,25,31,169,31,169,30,68,31,206,31,166,31,82,31,201,31,74,31,43,31,107,31,197,31,23,31,23,30,185,31,31,31,93,31,182,31,150,31,150,30,1,31,234,31,25,31,99,31,214,31,160,31,252,31,252,30,252,29,204,31,82,31,221,31,18,31,69,31,121,31,122,31,45,31,45,30,200,31,114,31,219,31,219,30,134,31,233,31,191,31,52,31,151,31,9,31,151,31,102,31,102,30,156,31,15,31,80,31,80,30,22,31,144,31,214,31,192,31,84,31,84,30,197,31,197,30,113,31,246,31,36,31,27,31,185,31,235,31,47,31,47,30,220,31,187,31,249,31,234,31,191,31,195,31,195,30,81,31,81,30,62,31,62,30,62,29,208,31,47,31,47,30,47,29,7,31,7,30,147,31,97,31,255,31,255,30,70,31,241,31,32,31,209,31,209,30,209,29,223,31,56,31,16,31,244,31,203,31,161,31,85,31,85,30,25,31,2,31,57,31,255,31,35,31,10,31,19,31,244,31,125,31,248,31,10,31,36,31,241,31,47,31,47,30,69,31,249,31,125,31,49,31,49,30,191,31,191,30,206,31,206,30,63,31,96,31,96,30,128,31,128,30,128,29,91,31,91,30,247,31,101,31,3,31,252,31,252,31,78,31,41,31,117,31,122,31,86,31,145,31,148,31,148,30,153,31,19,31,203,31,238,31,110,31,155,31,53,31,28,31,28,30,28,29,127,31,62,31,131,31,248,31,97,31,178,31,212,31,212,30,135,31,250,31,127,31,158,31,103,31,13,31,25,31,73,31,108,31,120,31,24,31,29,31,112,31,184,31,144,31,144,30,77,31,77,30,165,31,87,31,99,31,50,31,1,31,85,31,130,31,31,31,13,31,21,31,21,30,253,31,214,31,79,31,79,30,210,31,78,31,212,31,243,31,243,30,195,31,195,30,239,31,239,30,239,29,251,31,170,31,162,31,230,31,67,31,157,31,33,31,244,31,23,31,190,31,209,31,116,31,153,31,106,31,100,31,96,31,131,31,131,30,131,29,128,31,42,31,44,31,145,31,145,30,151,31,42,31,253,31,253,30,5,31,131,31,131,30,154,31,185,31,165,31,40,31,40,30,40,29,141,31,166,31,63,31,68,31,94,31,94,30,83,31,226,31,226,30,250,31,228,31,214,31,212,31,199,31,168,31,1,31,7,31,161,31,161,30,161,29,161,28,176,31,176,30,45,31,238,31,238,30,254,31,130,31,130,30,147,31,20,31,37,31,159,31,95,31,149,31,149,30,60,31,60,30,60,29,60,31,60,30,60,29,60,28,60,27,123,31,170,31,170,30,67,31,22,31,166,31,210,31,150,31,176,31,44,31,219,31,141,31,250,31,97,31,159,31,107,31,27,31,45,31,244,31,43,31,221,31,89,31,41,31,51,31,184,31,184,30,123,31,77,31,163,31,242,31,64,31,13,31,13,30,13,29,125,31,81,31,81,30,201,31,68,31,43,31,2,31,183,31,117,31,117,30,170,31,101,31,107,31,242,31,242,30,237,31,237,30,78,31,250,31,135,31,157,31,83,31,40,31,93,31,93,30,190,31,62,31,142,31,90,31,214,31,189,31,84,31,207,31,215,31,254,31,34,31,215,31,88,31,204,31,204,30,95,31,95,30,26,31,26,30,184,31,109,31,200,31,18,31,112,31,213,31,219,31,158,31,224,31,112,31,112,30,112,29,81,31,88,31,98,31,98,30,98,29,172,31,35,31,35,30,104,31,176,31,176,30,176,29,165,31,165,30,165,29,66,31,14,31,104,31,196,31,181,31,86,31,86,30,99,31,3,31,100,31,178,31,178,30,185,31,185,30,129,31,224,31,28,31,217,31,207,31,187,31,172,31,196,31,196,30,157,31,137,31,80,31,80,30,18,31,18,30,152,31,49,31,209,31,224,31,18,31,18,30,224,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
