-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 812;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,235,0,31,0,218,0,162,0,209,0,48,0,39,0,248,0,127,0,226,0,85,0,77,0,77,0,248,0,0,0,75,0,0,0,133,0,79,0,106,0,128,0,191,0,0,0,57,0,27,0,203,0,63,0,0,0,123,0,148,0,0,0,148,0,107,0,175,0,0,0,83,0,119,0,172,0,226,0,41,0,46,0,124,0,148,0,0,0,42,0,0,0,100,0,129,0,0,0,0,0,49,0,105,0,27,0,30,0,137,0,5,0,163,0,142,0,198,0,170,0,242,0,249,0,122,0,88,0,118,0,143,0,105,0,52,0,226,0,14,0,1,0,51,0,70,0,237,0,212,0,71,0,248,0,105,0,137,0,252,0,242,0,255,0,5,0,190,0,200,0,217,0,210,0,0,0,157,0,75,0,73,0,170,0,69,0,134,0,54,0,85,0,0,0,0,0,64,0,59,0,101,0,82,0,0,0,108,0,44,0,0,0,166,0,0,0,1,0,26,0,2,0,150,0,2,0,198,0,0,0,255,0,94,0,0,0,249,0,153,0,70,0,8,0,0,0,0,0,0,0,49,0,10,0,157,0,95,0,22,0,42,0,206,0,17,0,12,0,0,0,211,0,53,0,75,0,0,0,144,0,174,0,0,0,26,0,222,0,82,0,0,0,0,0,193,0,224,0,27,0,67,0,189,0,106,0,0,0,0,0,47,0,40,0,3,0,251,0,61,0,135,0,124,0,0,0,0,0,53,0,124,0,154,0,66,0,10,0,222,0,144,0,0,0,243,0,253,0,79,0,243,0,71,0,197,0,189,0,11,0,84,0,146,0,171,0,104,0,0,0,137,0,0,0,110,0,204,0,0,0,211,0,51,0,177,0,157,0,0,0,61,0,0,0,189,0,45,0,83,0,74,0,0,0,20,0,0,0,242,0,183,0,2,0,55,0,214,0,0,0,196,0,91,0,136,0,70,0,14,0,85,0,70,0,10,0,146,0,58,0,106,0,114,0,187,0,0,0,160,0,134,0,71,0,237,0,83,0,235,0,237,0,105,0,4,0,85,0,170,0,140,0,154,0,0,0,203,0,129,0,0,0,5,0,245,0,138,0,150,0,175,0,107,0,248,0,32,0,173,0,243,0,195,0,114,0,82,0,0,0,155,0,114,0,216,0,35,0,160,0,0,0,0,0,156,0,207,0,0,0,204,0,185,0,12,0,176,0,13,0,132,0,253,0,0,0,210,0,0,0,0,0,0,0,0,0,59,0,102,0,166,0,76,0,139,0,136,0,0,0,0,0,163,0,0,0,0,0,30,0,24,0,204,0,0,0,19,0,85,0,242,0,101,0,83,0,117,0,163,0,126,0,40,0,200,0,210,0,233,0,165,0,173,0,111,0,46,0,102,0,0,0,221,0,254,0,0,0,218,0,1,0,89,0,122,0,130,0,39,0,66,0,154,0,120,0,0,0,0,0,0,0,195,0,72,0,255,0,0,0,45,0,203,0,206,0,197,0,93,0,240,0,0,0,5,0,0,0,103,0,97,0,0,0,177,0,228,0,0,0,108,0,189,0,152,0,239,0,199,0,40,0,219,0,107,0,95,0,226,0,46,0,236,0,68,0,73,0,119,0,195,0,173,0,114,0,43,0,1,0,241,0,23,0,43,0,142,0,157,0,54,0,0,0,124,0,212,0,0,0,2,0,0,0,213,0,110,0,209,0,0,0,53,0,0,0,151,0,172,0,0,0,163,0,193,0,150,0,149,0,251,0,161,0,95,0,0,0,130,0,212,0,40,0,0,0,198,0,0,0,72,0,197,0,25,0,213,0,0,0,0,0,0,0,55,0,0,0,36,0,238,0,0,0,212,0,0,0,0,0,167,0,218,0,226,0,30,0,18,0,239,0,12,0,211,0,162,0,83,0,87,0,49,0,217,0,184,0,234,0,70,0,0,0,68,0,177,0,193,0,23,0,115,0,69,0,4,0,104,0,57,0,210,0,54,0,0,0,161,0,147,0,0,0,215,0,131,0,197,0,172,0,106,0,35,0,52,0,235,0,140,0,23,0,28,0,0,0,172,0,96,0,198,0,105,0,65,0,62,0,0,0,250,0,0,0,144,0,27,0,90,0,235,0,44,0,0,0,43,0,251,0,187,0,225,0,0,0,53,0,18,0,179,0,169,0,0,0,33,0,39,0,19,0,31,0,108,0,198,0,239,0,21,0,3,0,52,0,142,0,80,0,255,0,107,0,18,0,61,0,55,0,32,0,125,0,0,0,0,0,95,0,0,0,0,0,174,0,0,0,50,0,229,0,219,0,186,0,8,0,128,0,138,0,10,0,170,0,45,0,132,0,110,0,111,0,154,0,137,0,102,0,236,0,152,0,19,0,58,0,94,0,80,0,91,0,110,0,184,0,103,0,224,0,136,0,250,0,203,0,1,0,25,0,156,0,0,0,127,0,65,0,0,0,90,0,73,0,166,0,0,0,227,0,123,0,0,0,189,0,162,0,0,0,249,0,47,0,16,0,36,0,75,0,163,0,118,0,34,0,97,0,18,0,126,0,89,0,10,0,138,0,0,0,56,0,0,0,178,0,31,0,198,0,201,0,224,0,181,0,81,0,0,0,246,0,248,0,0,0,179,0,149,0,243,0,208,0,78,0,0,0,64,0,179,0,101,0,159,0,35,0,157,0,153,0,113,0,27,0,21,0,156,0,30,0,111,0,0,0,0,0,0,0,53,0,0,0,76,0,169,0,163,0,40,0,67,0,0,0,194,0,111,0,0,0,221,0,228,0,0,0,128,0,180,0,185,0,95,0,217,0,6,0,91,0,0,0,40,0,3,0,228,0,194,0,209,0,250,0,102,0,45,0,209,0,99,0,168,0,0,0,147,0,117,0,227,0,0,0,0,0,41,0,0,0,94,0,196,0,0,0,0,0,71,0,225,0,77,0,169,0,193,0,79,0,196,0,13,0,7,0,42,0,129,0,191,0,11,0,49,0,13,0,184,0,174,0,239,0,238,0,144,0,0,0,207,0,2,0,175,0,101,0,0,0,149,0,147,0,134,0,42,0,41,0,223,0,186,0,82,0,141,0,92,0,72,0,84,0,79,0,0,0,224,0,225,0,39,0,0,0,170,0,201,0,161,0,116,0,179,0,0,0,0,0,26,0,40,0,0,0,41,0,22,0,163,0,161,0,140,0,0,0,171,0,126,0,24,0,127,0,206,0,92,0,0,0,87,0,0,0,253,0,141,0,238,0,248,0,141,0,244,0,1,0,8,0,43,0,0,0,0,0,57,0,49,0,219,0,13,0,55,0,145,0,13,0,0,0,248,0,239,0,219,0,8,0,0,0,109,0,203,0,0,0,247,0,242,0,213,0,182,0,167,0,161,0,53,0,0,0,164,0,76,0,52,0,166,0,253,0,215,0,112,0,3,0,76,0,87,0,208,0,168,0,42,0,59,0,0,0,0,0,147,0,0,0,148,0,106,0,214,0,0,0,94,0,63,0,18,0,96,0,188,0,225,0,0,0,0,0,35,0,51,0,31,0,241,0,100,0,140,0,139,0,18,0,0,0,31,0,0,0,254,0,136,0,5,0,56,0,6,0,0,0,16,0,191,0,36,0,15,0,202,0,209,0,132,0,41,0);
signal scenario_full  : scenario_type := (0,0,235,31,31,31,218,31,162,31,209,31,48,31,39,31,248,31,127,31,226,31,85,31,77,31,77,31,248,31,248,30,75,31,75,30,133,31,79,31,106,31,128,31,191,31,191,30,57,31,27,31,203,31,63,31,63,30,123,31,148,31,148,30,148,31,107,31,175,31,175,30,83,31,119,31,172,31,226,31,41,31,46,31,124,31,148,31,148,30,42,31,42,30,100,31,129,31,129,30,129,29,49,31,105,31,27,31,30,31,137,31,5,31,163,31,142,31,198,31,170,31,242,31,249,31,122,31,88,31,118,31,143,31,105,31,52,31,226,31,14,31,1,31,51,31,70,31,237,31,212,31,71,31,248,31,105,31,137,31,252,31,242,31,255,31,5,31,190,31,200,31,217,31,210,31,210,30,157,31,75,31,73,31,170,31,69,31,134,31,54,31,85,31,85,30,85,29,64,31,59,31,101,31,82,31,82,30,108,31,44,31,44,30,166,31,166,30,1,31,26,31,2,31,150,31,2,31,198,31,198,30,255,31,94,31,94,30,249,31,153,31,70,31,8,31,8,30,8,29,8,28,49,31,10,31,157,31,95,31,22,31,42,31,206,31,17,31,12,31,12,30,211,31,53,31,75,31,75,30,144,31,174,31,174,30,26,31,222,31,82,31,82,30,82,29,193,31,224,31,27,31,67,31,189,31,106,31,106,30,106,29,47,31,40,31,3,31,251,31,61,31,135,31,124,31,124,30,124,29,53,31,124,31,154,31,66,31,10,31,222,31,144,31,144,30,243,31,253,31,79,31,243,31,71,31,197,31,189,31,11,31,84,31,146,31,171,31,104,31,104,30,137,31,137,30,110,31,204,31,204,30,211,31,51,31,177,31,157,31,157,30,61,31,61,30,189,31,45,31,83,31,74,31,74,30,20,31,20,30,242,31,183,31,2,31,55,31,214,31,214,30,196,31,91,31,136,31,70,31,14,31,85,31,70,31,10,31,146,31,58,31,106,31,114,31,187,31,187,30,160,31,134,31,71,31,237,31,83,31,235,31,237,31,105,31,4,31,85,31,170,31,140,31,154,31,154,30,203,31,129,31,129,30,5,31,245,31,138,31,150,31,175,31,107,31,248,31,32,31,173,31,243,31,195,31,114,31,82,31,82,30,155,31,114,31,216,31,35,31,160,31,160,30,160,29,156,31,207,31,207,30,204,31,185,31,12,31,176,31,13,31,132,31,253,31,253,30,210,31,210,30,210,29,210,28,210,27,59,31,102,31,166,31,76,31,139,31,136,31,136,30,136,29,163,31,163,30,163,29,30,31,24,31,204,31,204,30,19,31,85,31,242,31,101,31,83,31,117,31,163,31,126,31,40,31,200,31,210,31,233,31,165,31,173,31,111,31,46,31,102,31,102,30,221,31,254,31,254,30,218,31,1,31,89,31,122,31,130,31,39,31,66,31,154,31,120,31,120,30,120,29,120,28,195,31,72,31,255,31,255,30,45,31,203,31,206,31,197,31,93,31,240,31,240,30,5,31,5,30,103,31,97,31,97,30,177,31,228,31,228,30,108,31,189,31,152,31,239,31,199,31,40,31,219,31,107,31,95,31,226,31,46,31,236,31,68,31,73,31,119,31,195,31,173,31,114,31,43,31,1,31,241,31,23,31,43,31,142,31,157,31,54,31,54,30,124,31,212,31,212,30,2,31,2,30,213,31,110,31,209,31,209,30,53,31,53,30,151,31,172,31,172,30,163,31,193,31,150,31,149,31,251,31,161,31,95,31,95,30,130,31,212,31,40,31,40,30,198,31,198,30,72,31,197,31,25,31,213,31,213,30,213,29,213,28,55,31,55,30,36,31,238,31,238,30,212,31,212,30,212,29,167,31,218,31,226,31,30,31,18,31,239,31,12,31,211,31,162,31,83,31,87,31,49,31,217,31,184,31,234,31,70,31,70,30,68,31,177,31,193,31,23,31,115,31,69,31,4,31,104,31,57,31,210,31,54,31,54,30,161,31,147,31,147,30,215,31,131,31,197,31,172,31,106,31,35,31,52,31,235,31,140,31,23,31,28,31,28,30,172,31,96,31,198,31,105,31,65,31,62,31,62,30,250,31,250,30,144,31,27,31,90,31,235,31,44,31,44,30,43,31,251,31,187,31,225,31,225,30,53,31,18,31,179,31,169,31,169,30,33,31,39,31,19,31,31,31,108,31,198,31,239,31,21,31,3,31,52,31,142,31,80,31,255,31,107,31,18,31,61,31,55,31,32,31,125,31,125,30,125,29,95,31,95,30,95,29,174,31,174,30,50,31,229,31,219,31,186,31,8,31,128,31,138,31,10,31,170,31,45,31,132,31,110,31,111,31,154,31,137,31,102,31,236,31,152,31,19,31,58,31,94,31,80,31,91,31,110,31,184,31,103,31,224,31,136,31,250,31,203,31,1,31,25,31,156,31,156,30,127,31,65,31,65,30,90,31,73,31,166,31,166,30,227,31,123,31,123,30,189,31,162,31,162,30,249,31,47,31,16,31,36,31,75,31,163,31,118,31,34,31,97,31,18,31,126,31,89,31,10,31,138,31,138,30,56,31,56,30,178,31,31,31,198,31,201,31,224,31,181,31,81,31,81,30,246,31,248,31,248,30,179,31,149,31,243,31,208,31,78,31,78,30,64,31,179,31,101,31,159,31,35,31,157,31,153,31,113,31,27,31,21,31,156,31,30,31,111,31,111,30,111,29,111,28,53,31,53,30,76,31,169,31,163,31,40,31,67,31,67,30,194,31,111,31,111,30,221,31,228,31,228,30,128,31,180,31,185,31,95,31,217,31,6,31,91,31,91,30,40,31,3,31,228,31,194,31,209,31,250,31,102,31,45,31,209,31,99,31,168,31,168,30,147,31,117,31,227,31,227,30,227,29,41,31,41,30,94,31,196,31,196,30,196,29,71,31,225,31,77,31,169,31,193,31,79,31,196,31,13,31,7,31,42,31,129,31,191,31,11,31,49,31,13,31,184,31,174,31,239,31,238,31,144,31,144,30,207,31,2,31,175,31,101,31,101,30,149,31,147,31,134,31,42,31,41,31,223,31,186,31,82,31,141,31,92,31,72,31,84,31,79,31,79,30,224,31,225,31,39,31,39,30,170,31,201,31,161,31,116,31,179,31,179,30,179,29,26,31,40,31,40,30,41,31,22,31,163,31,161,31,140,31,140,30,171,31,126,31,24,31,127,31,206,31,92,31,92,30,87,31,87,30,253,31,141,31,238,31,248,31,141,31,244,31,1,31,8,31,43,31,43,30,43,29,57,31,49,31,219,31,13,31,55,31,145,31,13,31,13,30,248,31,239,31,219,31,8,31,8,30,109,31,203,31,203,30,247,31,242,31,213,31,182,31,167,31,161,31,53,31,53,30,164,31,76,31,52,31,166,31,253,31,215,31,112,31,3,31,76,31,87,31,208,31,168,31,42,31,59,31,59,30,59,29,147,31,147,30,148,31,106,31,214,31,214,30,94,31,63,31,18,31,96,31,188,31,225,31,225,30,225,29,35,31,51,31,31,31,241,31,100,31,140,31,139,31,18,31,18,30,31,31,31,30,254,31,136,31,5,31,56,31,6,31,6,30,16,31,191,31,36,31,15,31,202,31,209,31,132,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
