-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 489;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,10,0,0,0,70,0,115,0,89,0,150,0,81,0,207,0,104,0,248,0,63,0,0,0,232,0,0,0,121,0,0,0,235,0,49,0,108,0,144,0,219,0,205,0,0,0,26,0,18,0,202,0,0,0,25,0,17,0,111,0,43,0,243,0,190,0,76,0,58,0,181,0,117,0,146,0,191,0,81,0,63,0,32,0,188,0,246,0,170,0,88,0,0,0,252,0,111,0,0,0,186,0,0,0,88,0,147,0,108,0,108,0,121,0,210,0,182,0,0,0,115,0,23,0,224,0,218,0,37,0,210,0,193,0,38,0,112,0,227,0,55,0,0,0,118,0,0,0,249,0,0,0,79,0,0,0,64,0,112,0,50,0,91,0,8,0,0,0,47,0,0,0,0,0,165,0,72,0,0,0,94,0,55,0,34,0,0,0,1,0,195,0,132,0,12,0,56,0,92,0,240,0,167,0,0,0,46,0,162,0,0,0,143,0,0,0,0,0,78,0,0,0,117,0,198,0,48,0,14,0,224,0,156,0,0,0,73,0,129,0,87,0,89,0,187,0,29,0,237,0,4,0,122,0,17,0,182,0,153,0,254,0,26,0,0,0,162,0,194,0,100,0,174,0,49,0,31,0,8,0,162,0,116,0,150,0,0,0,81,0,56,0,0,0,188,0,120,0,187,0,175,0,80,0,26,0,0,0,105,0,15,0,24,0,169,0,165,0,114,0,77,0,0,0,185,0,211,0,152,0,221,0,0,0,222,0,49,0,0,0,213,0,0,0,131,0,185,0,0,0,51,0,174,0,191,0,0,0,84,0,81,0,60,0,220,0,207,0,60,0,221,0,7,0,94,0,41,0,0,0,33,0,74,0,145,0,186,0,79,0,80,0,112,0,212,0,0,0,230,0,70,0,231,0,13,0,121,0,0,0,0,0,111,0,0,0,140,0,0,0,148,0,108,0,206,0,219,0,11,0,86,0,26,0,181,0,94,0,242,0,105,0,163,0,37,0,74,0,57,0,0,0,249,0,148,0,177,0,246,0,0,0,50,0,194,0,8,0,0,0,0,0,104,0,0,0,193,0,31,0,0,0,227,0,0,0,0,0,51,0,165,0,137,0,229,0,172,0,125,0,9,0,143,0,21,0,93,0,185,0,122,0,130,0,214,0,201,0,130,0,62,0,180,0,191,0,9,0,209,0,0,0,23,0,198,0,83,0,0,0,4,0,51,0,15,0,232,0,0,0,11,0,245,0,18,0,202,0,0,0,14,0,208,0,245,0,21,0,255,0,148,0,139,0,183,0,235,0,160,0,102,0,65,0,236,0,68,0,74,0,137,0,0,0,84,0,224,0,35,0,59,0,88,0,60,0,47,0,0,0,186,0,253,0,97,0,0,0,96,0,89,0,5,0,161,0,107,0,54,0,219,0,47,0,0,0,36,0,0,0,162,0,0,0,13,0,0,0,0,0,237,0,237,0,83,0,0,0,222,0,0,0,117,0,47,0,191,0,158,0,18,0,207,0,127,0,128,0,88,0,152,0,64,0,134,0,161,0,211,0,138,0,0,0,247,0,0,0,207,0,84,0,25,0,67,0,0,0,241,0,0,0,125,0,160,0,27,0,32,0,0,0,232,0,40,0,0,0,255,0,228,0,205,0,204,0,22,0,170,0,0,0,0,0,186,0,0,0,0,0,100,0,218,0,180,0,189,0,37,0,92,0,100,0,243,0,96,0,141,0,22,0,153,0,212,0,33,0,178,0,221,0,112,0,0,0,163,0,76,0,67,0,137,0,51,0,132,0,183,0,12,0,101,0,133,0,26,0,128,0,70,0,250,0,123,0,120,0,107,0,15,0,35,0,211,0,39,0,20,0,0,0,152,0,0,0,217,0,46,0,107,0,114,0,221,0,212,0,46,0,163,0,197,0,0,0,49,0,0,0,0,0,40,0,4,0,185,0,0,0,232,0,67,0,0,0,156,0,180,0,0,0,51,0,67,0,39,0,137,0,152,0,22,0,210,0,172,0,37,0,85,0,0,0,176,0,201,0,247,0,54,0,0,0,0,0,111,0,99,0,23,0,176,0,148,0,101,0,153,0,98,0,0,0,104,0,178,0,0,0,133,0,175,0,191,0,51,0,201,0,223,0,163,0,83,0,115,0,111,0,206,0,212,0,249,0,0,0,14,0,63,0,94,0,187,0);
signal scenario_full  : scenario_type := (102,31,10,31,10,30,70,31,115,31,89,31,150,31,81,31,207,31,104,31,248,31,63,31,63,30,232,31,232,30,121,31,121,30,235,31,49,31,108,31,144,31,219,31,205,31,205,30,26,31,18,31,202,31,202,30,25,31,17,31,111,31,43,31,243,31,190,31,76,31,58,31,181,31,117,31,146,31,191,31,81,31,63,31,32,31,188,31,246,31,170,31,88,31,88,30,252,31,111,31,111,30,186,31,186,30,88,31,147,31,108,31,108,31,121,31,210,31,182,31,182,30,115,31,23,31,224,31,218,31,37,31,210,31,193,31,38,31,112,31,227,31,55,31,55,30,118,31,118,30,249,31,249,30,79,31,79,30,64,31,112,31,50,31,91,31,8,31,8,30,47,31,47,30,47,29,165,31,72,31,72,30,94,31,55,31,34,31,34,30,1,31,195,31,132,31,12,31,56,31,92,31,240,31,167,31,167,30,46,31,162,31,162,30,143,31,143,30,143,29,78,31,78,30,117,31,198,31,48,31,14,31,224,31,156,31,156,30,73,31,129,31,87,31,89,31,187,31,29,31,237,31,4,31,122,31,17,31,182,31,153,31,254,31,26,31,26,30,162,31,194,31,100,31,174,31,49,31,31,31,8,31,162,31,116,31,150,31,150,30,81,31,56,31,56,30,188,31,120,31,187,31,175,31,80,31,26,31,26,30,105,31,15,31,24,31,169,31,165,31,114,31,77,31,77,30,185,31,211,31,152,31,221,31,221,30,222,31,49,31,49,30,213,31,213,30,131,31,185,31,185,30,51,31,174,31,191,31,191,30,84,31,81,31,60,31,220,31,207,31,60,31,221,31,7,31,94,31,41,31,41,30,33,31,74,31,145,31,186,31,79,31,80,31,112,31,212,31,212,30,230,31,70,31,231,31,13,31,121,31,121,30,121,29,111,31,111,30,140,31,140,30,148,31,108,31,206,31,219,31,11,31,86,31,26,31,181,31,94,31,242,31,105,31,163,31,37,31,74,31,57,31,57,30,249,31,148,31,177,31,246,31,246,30,50,31,194,31,8,31,8,30,8,29,104,31,104,30,193,31,31,31,31,30,227,31,227,30,227,29,51,31,165,31,137,31,229,31,172,31,125,31,9,31,143,31,21,31,93,31,185,31,122,31,130,31,214,31,201,31,130,31,62,31,180,31,191,31,9,31,209,31,209,30,23,31,198,31,83,31,83,30,4,31,51,31,15,31,232,31,232,30,11,31,245,31,18,31,202,31,202,30,14,31,208,31,245,31,21,31,255,31,148,31,139,31,183,31,235,31,160,31,102,31,65,31,236,31,68,31,74,31,137,31,137,30,84,31,224,31,35,31,59,31,88,31,60,31,47,31,47,30,186,31,253,31,97,31,97,30,96,31,89,31,5,31,161,31,107,31,54,31,219,31,47,31,47,30,36,31,36,30,162,31,162,30,13,31,13,30,13,29,237,31,237,31,83,31,83,30,222,31,222,30,117,31,47,31,191,31,158,31,18,31,207,31,127,31,128,31,88,31,152,31,64,31,134,31,161,31,211,31,138,31,138,30,247,31,247,30,207,31,84,31,25,31,67,31,67,30,241,31,241,30,125,31,160,31,27,31,32,31,32,30,232,31,40,31,40,30,255,31,228,31,205,31,204,31,22,31,170,31,170,30,170,29,186,31,186,30,186,29,100,31,218,31,180,31,189,31,37,31,92,31,100,31,243,31,96,31,141,31,22,31,153,31,212,31,33,31,178,31,221,31,112,31,112,30,163,31,76,31,67,31,137,31,51,31,132,31,183,31,12,31,101,31,133,31,26,31,128,31,70,31,250,31,123,31,120,31,107,31,15,31,35,31,211,31,39,31,20,31,20,30,152,31,152,30,217,31,46,31,107,31,114,31,221,31,212,31,46,31,163,31,197,31,197,30,49,31,49,30,49,29,40,31,4,31,185,31,185,30,232,31,67,31,67,30,156,31,180,31,180,30,51,31,67,31,39,31,137,31,152,31,22,31,210,31,172,31,37,31,85,31,85,30,176,31,201,31,247,31,54,31,54,30,54,29,111,31,99,31,23,31,176,31,148,31,101,31,153,31,98,31,98,30,104,31,178,31,178,30,133,31,175,31,191,31,51,31,201,31,223,31,163,31,83,31,115,31,111,31,206,31,212,31,249,31,249,30,14,31,63,31,94,31,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
