-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_814 is
end project_tb_814;

architecture project_tb_arch_814 of project_tb_814 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1014;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (210,0,45,0,207,0,0,0,230,0,0,0,3,0,0,0,0,0,197,0,0,0,43,0,171,0,124,0,0,0,166,0,134,0,184,0,185,0,47,0,0,0,166,0,0,0,236,0,0,0,0,0,19,0,0,0,57,0,86,0,89,0,252,0,233,0,0,0,141,0,0,0,235,0,154,0,0,0,90,0,208,0,14,0,81,0,73,0,54,0,111,0,167,0,39,0,140,0,146,0,0,0,0,0,238,0,89,0,0,0,0,0,124,0,0,0,179,0,46,0,21,0,180,0,39,0,85,0,6,0,4,0,0,0,223,0,60,0,185,0,157,0,234,0,0,0,0,0,145,0,127,0,107,0,225,0,144,0,97,0,188,0,66,0,118,0,113,0,63,0,147,0,163,0,142,0,174,0,135,0,0,0,93,0,245,0,175,0,0,0,169,0,0,0,123,0,42,0,27,0,81,0,73,0,144,0,201,0,218,0,154,0,28,0,14,0,186,0,114,0,239,0,0,0,192,0,53,0,246,0,218,0,157,0,0,0,158,0,176,0,106,0,148,0,175,0,0,0,43,0,199,0,0,0,190,0,185,0,0,0,189,0,59,0,222,0,62,0,255,0,152,0,6,0,29,0,142,0,229,0,241,0,58,0,42,0,4,0,96,0,223,0,48,0,171,0,185,0,93,0,155,0,17,0,77,0,168,0,57,0,182,0,0,0,248,0,0,0,0,0,232,0,0,0,49,0,229,0,110,0,0,0,147,0,0,0,121,0,252,0,200,0,117,0,96,0,140,0,204,0,121,0,178,0,13,0,0,0,89,0,142,0,0,0,73,0,0,0,46,0,0,0,71,0,253,0,17,0,19,0,0,0,175,0,7,0,0,0,187,0,195,0,0,0,8,0,234,0,59,0,237,0,249,0,223,0,202,0,115,0,0,0,189,0,0,0,2,0,0,0,105,0,0,0,2,0,210,0,214,0,102,0,119,0,250,0,5,0,115,0,34,0,246,0,245,0,244,0,219,0,10,0,0,0,225,0,145,0,137,0,123,0,248,0,224,0,2,0,167,0,0,0,203,0,255,0,0,0,163,0,177,0,2,0,0,0,79,0,82,0,238,0,127,0,176,0,237,0,108,0,25,0,76,0,152,0,66,0,182,0,0,0,0,0,18,0,235,0,48,0,77,0,25,0,89,0,200,0,0,0,222,0,18,0,127,0,81,0,168,0,0,0,166,0,0,0,218,0,122,0,165,0,53,0,173,0,90,0,173,0,195,0,113,0,0,0,0,0,108,0,170,0,165,0,0,0,50,0,170,0,0,0,52,0,25,0,172,0,109,0,185,0,157,0,223,0,13,0,66,0,243,0,211,0,109,0,0,0,185,0,204,0,27,0,98,0,248,0,0,0,246,0,0,0,179,0,154,0,0,0,209,0,96,0,0,0,51,0,0,0,166,0,0,0,130,0,49,0,136,0,45,0,129,0,58,0,244,0,25,0,56,0,0,0,99,0,232,0,159,0,195,0,148,0,0,0,35,0,0,0,233,0,20,0,35,0,167,0,214,0,94,0,198,0,35,0,96,0,4,0,90,0,0,0,0,0,44,0,19,0,191,0,218,0,241,0,178,0,0,0,0,0,99,0,181,0,109,0,0,0,217,0,18,0,143,0,38,0,0,0,179,0,122,0,208,0,136,0,0,0,28,0,8,0,52,0,185,0,0,0,211,0,76,0,162,0,160,0,241,0,72,0,164,0,152,0,224,0,82,0,192,0,0,0,170,0,200,0,158,0,129,0,76,0,145,0,138,0,0,0,186,0,0,0,100,0,154,0,0,0,44,0,65,0,93,0,0,0,0,0,0,0,52,0,254,0,0,0,232,0,80,0,157,0,186,0,162,0,192,0,138,0,73,0,0,0,234,0,14,0,89,0,0,0,92,0,161,0,220,0,253,0,0,0,107,0,166,0,180,0,0,0,99,0,119,0,106,0,0,0,211,0,198,0,8,0,196,0,65,0,39,0,62,0,142,0,42,0,90,0,109,0,0,0,0,0,222,0,126,0,15,0,179,0,190,0,239,0,254,0,208,0,0,0,0,0,218,0,255,0,224,0,96,0,58,0,127,0,124,0,87,0,0,0,53,0,13,0,237,0,39,0,20,0,123,0,187,0,54,0,146,0,146,0,128,0,141,0,0,0,122,0,0,0,24,0,0,0,97,0,6,0,190,0,26,0,34,0,0,0,228,0,129,0,159,0,64,0,16,0,16,0,142,0,221,0,102,0,28,0,0,0,244,0,6,0,169,0,11,0,0,0,252,0,84,0,3,0,40,0,170,0,0,0,102,0,46,0,118,0,252,0,54,0,108,0,172,0,119,0,0,0,80,0,163,0,196,0,42,0,151,0,115,0,164,0,155,0,184,0,138,0,197,0,138,0,73,0,69,0,0,0,55,0,13,0,98,0,0,0,0,0,0,0,26,0,152,0,179,0,25,0,0,0,0,0,0,0,0,0,110,0,0,0,0,0,78,0,0,0,39,0,97,0,73,0,223,0,176,0,7,0,118,0,240,0,0,0,141,0,0,0,0,0,12,0,0,0,0,0,115,0,206,0,222,0,0,0,91,0,166,0,53,0,220,0,112,0,112,0,0,0,160,0,0,0,132,0,6,0,0,0,24,0,0,0,155,0,96,0,252,0,0,0,13,0,109,0,80,0,0,0,22,0,37,0,255,0,216,0,38,0,85,0,61,0,165,0,0,0,0,0,0,0,220,0,101,0,124,0,170,0,135,0,240,0,234,0,0,0,0,0,144,0,134,0,64,0,0,0,184,0,243,0,188,0,132,0,191,0,0,0,125,0,1,0,112,0,239,0,72,0,208,0,114,0,249,0,67,0,0,0,44,0,193,0,185,0,140,0,159,0,0,0,6,0,24,0,6,0,111,0,29,0,202,0,0,0,38,0,169,0,0,0,203,0,247,0,0,0,20,0,89,0,69,0,53,0,83,0,0,0,36,0,90,0,0,0,55,0,94,0,193,0,189,0,0,0,239,0,45,0,27,0,144,0,51,0,132,0,20,0,206,0,206,0,0,0,83,0,14,0,157,0,162,0,102,0,203,0,103,0,0,0,0,0,103,0,122,0,176,0,248,0,220,0,0,0,37,0,200,0,0,0,78,0,18,0,109,0,210,0,0,0,72,0,237,0,223,0,151,0,29,0,197,0,172,0,0,0,57,0,222,0,14,0,123,0,101,0,237,0,19,0,0,0,0,0,33,0,0,0,230,0,194,0,47,0,134,0,46,0,0,0,77,0,37,0,24,0,33,0,20,0,213,0,175,0,0,0,166,0,0,0,51,0,0,0,68,0,0,0,158,0,224,0,133,0,0,0,21,0,121,0,0,0,104,0,0,0,0,0,162,0,223,0,252,0,174,0,6,0,180,0,0,0,178,0,0,0,149,0,43,0,148,0,0,0,60,0,114,0,168,0,0,0,59,0,0,0,84,0,241,0,167,0,147,0,109,0,252,0,59,0,72,0,220,0,0,0,173,0,222,0,97,0,240,0,150,0,73,0,49,0,183,0,229,0,0,0,0,0,179,0,220,0,204,0,240,0,35,0,35,0,82,0,200,0,236,0,93,0,25,0,173,0,0,0,255,0,0,0,0,0,172,0,110,0,204,0,0,0,22,0,89,0,209,0,54,0,235,0,161,0,90,0,62,0,95,0,36,0,4,0,28,0,209,0,27,0,116,0,129,0,146,0,46,0,223,0,0,0,0,0,0,0,252,0,30,0,108,0,0,0,57,0,253,0,160,0,248,0,0,0,49,0,125,0,41,0,175,0,0,0,134,0,231,0,62,0,38,0,69,0,157,0,196,0,6,0,58,0,104,0,73,0,0,0,16,0,80,0,13,0,222,0,241,0,56,0,200,0,119,0,161,0,182,0,132,0,193,0,210,0,0,0,129,0,0,0,244,0,219,0,226,0,229,0,40,0,0,0,14,0,0,0,0,0,164,0,0,0,92,0,170,0,138,0,0,0,96,0,23,0,0,0,100,0,0,0,98,0,106,0,165,0,116,0,228,0,215,0,98,0,24,0,0,0,0,0,90,0,237,0,103,0,252,0,179,0,246,0,98,0,148,0,186,0,0,0,10,0,21,0,77,0,53,0,148,0,25,0,185,0,0,0,0,0,114,0,219,0,165,0,65,0,0,0,29,0,12,0,195,0,172,0,14,0,90,0,204,0,68,0,118,0,0,0,150,0,0,0,22,0,131,0,178,0,28,0,0,0,0,0,81,0,0,0,141,0,74,0,173,0,0,0,65,0,100,0,18,0,141,0,56,0,161,0,11,0,240,0,205,0,47,0,63,0,161,0,59,0,172,0,249,0,253,0,181,0,173,0,56,0,224,0,246,0,203,0,0,0,60,0,64,0,70,0,68,0,143,0,251,0,248,0,90,0,152,0,115,0,0,0,251,0,0,0,68,0,0,0,97,0,169,0,0,0,114,0,78,0,26,0,0,0,205,0,158,0,127,0,19,0,209,0,70,0,255,0,47,0,103,0,176,0,255,0);
signal scenario_full  : scenario_type := (210,31,45,31,207,31,207,30,230,31,230,30,3,31,3,30,3,29,197,31,197,30,43,31,171,31,124,31,124,30,166,31,134,31,184,31,185,31,47,31,47,30,166,31,166,30,236,31,236,30,236,29,19,31,19,30,57,31,86,31,89,31,252,31,233,31,233,30,141,31,141,30,235,31,154,31,154,30,90,31,208,31,14,31,81,31,73,31,54,31,111,31,167,31,39,31,140,31,146,31,146,30,146,29,238,31,89,31,89,30,89,29,124,31,124,30,179,31,46,31,21,31,180,31,39,31,85,31,6,31,4,31,4,30,223,31,60,31,185,31,157,31,234,31,234,30,234,29,145,31,127,31,107,31,225,31,144,31,97,31,188,31,66,31,118,31,113,31,63,31,147,31,163,31,142,31,174,31,135,31,135,30,93,31,245,31,175,31,175,30,169,31,169,30,123,31,42,31,27,31,81,31,73,31,144,31,201,31,218,31,154,31,28,31,14,31,186,31,114,31,239,31,239,30,192,31,53,31,246,31,218,31,157,31,157,30,158,31,176,31,106,31,148,31,175,31,175,30,43,31,199,31,199,30,190,31,185,31,185,30,189,31,59,31,222,31,62,31,255,31,152,31,6,31,29,31,142,31,229,31,241,31,58,31,42,31,4,31,96,31,223,31,48,31,171,31,185,31,93,31,155,31,17,31,77,31,168,31,57,31,182,31,182,30,248,31,248,30,248,29,232,31,232,30,49,31,229,31,110,31,110,30,147,31,147,30,121,31,252,31,200,31,117,31,96,31,140,31,204,31,121,31,178,31,13,31,13,30,89,31,142,31,142,30,73,31,73,30,46,31,46,30,71,31,253,31,17,31,19,31,19,30,175,31,7,31,7,30,187,31,195,31,195,30,8,31,234,31,59,31,237,31,249,31,223,31,202,31,115,31,115,30,189,31,189,30,2,31,2,30,105,31,105,30,2,31,210,31,214,31,102,31,119,31,250,31,5,31,115,31,34,31,246,31,245,31,244,31,219,31,10,31,10,30,225,31,145,31,137,31,123,31,248,31,224,31,2,31,167,31,167,30,203,31,255,31,255,30,163,31,177,31,2,31,2,30,79,31,82,31,238,31,127,31,176,31,237,31,108,31,25,31,76,31,152,31,66,31,182,31,182,30,182,29,18,31,235,31,48,31,77,31,25,31,89,31,200,31,200,30,222,31,18,31,127,31,81,31,168,31,168,30,166,31,166,30,218,31,122,31,165,31,53,31,173,31,90,31,173,31,195,31,113,31,113,30,113,29,108,31,170,31,165,31,165,30,50,31,170,31,170,30,52,31,25,31,172,31,109,31,185,31,157,31,223,31,13,31,66,31,243,31,211,31,109,31,109,30,185,31,204,31,27,31,98,31,248,31,248,30,246,31,246,30,179,31,154,31,154,30,209,31,96,31,96,30,51,31,51,30,166,31,166,30,130,31,49,31,136,31,45,31,129,31,58,31,244,31,25,31,56,31,56,30,99,31,232,31,159,31,195,31,148,31,148,30,35,31,35,30,233,31,20,31,35,31,167,31,214,31,94,31,198,31,35,31,96,31,4,31,90,31,90,30,90,29,44,31,19,31,191,31,218,31,241,31,178,31,178,30,178,29,99,31,181,31,109,31,109,30,217,31,18,31,143,31,38,31,38,30,179,31,122,31,208,31,136,31,136,30,28,31,8,31,52,31,185,31,185,30,211,31,76,31,162,31,160,31,241,31,72,31,164,31,152,31,224,31,82,31,192,31,192,30,170,31,200,31,158,31,129,31,76,31,145,31,138,31,138,30,186,31,186,30,100,31,154,31,154,30,44,31,65,31,93,31,93,30,93,29,93,28,52,31,254,31,254,30,232,31,80,31,157,31,186,31,162,31,192,31,138,31,73,31,73,30,234,31,14,31,89,31,89,30,92,31,161,31,220,31,253,31,253,30,107,31,166,31,180,31,180,30,99,31,119,31,106,31,106,30,211,31,198,31,8,31,196,31,65,31,39,31,62,31,142,31,42,31,90,31,109,31,109,30,109,29,222,31,126,31,15,31,179,31,190,31,239,31,254,31,208,31,208,30,208,29,218,31,255,31,224,31,96,31,58,31,127,31,124,31,87,31,87,30,53,31,13,31,237,31,39,31,20,31,123,31,187,31,54,31,146,31,146,31,128,31,141,31,141,30,122,31,122,30,24,31,24,30,97,31,6,31,190,31,26,31,34,31,34,30,228,31,129,31,159,31,64,31,16,31,16,31,142,31,221,31,102,31,28,31,28,30,244,31,6,31,169,31,11,31,11,30,252,31,84,31,3,31,40,31,170,31,170,30,102,31,46,31,118,31,252,31,54,31,108,31,172,31,119,31,119,30,80,31,163,31,196,31,42,31,151,31,115,31,164,31,155,31,184,31,138,31,197,31,138,31,73,31,69,31,69,30,55,31,13,31,98,31,98,30,98,29,98,28,26,31,152,31,179,31,25,31,25,30,25,29,25,28,25,27,110,31,110,30,110,29,78,31,78,30,39,31,97,31,73,31,223,31,176,31,7,31,118,31,240,31,240,30,141,31,141,30,141,29,12,31,12,30,12,29,115,31,206,31,222,31,222,30,91,31,166,31,53,31,220,31,112,31,112,31,112,30,160,31,160,30,132,31,6,31,6,30,24,31,24,30,155,31,96,31,252,31,252,30,13,31,109,31,80,31,80,30,22,31,37,31,255,31,216,31,38,31,85,31,61,31,165,31,165,30,165,29,165,28,220,31,101,31,124,31,170,31,135,31,240,31,234,31,234,30,234,29,144,31,134,31,64,31,64,30,184,31,243,31,188,31,132,31,191,31,191,30,125,31,1,31,112,31,239,31,72,31,208,31,114,31,249,31,67,31,67,30,44,31,193,31,185,31,140,31,159,31,159,30,6,31,24,31,6,31,111,31,29,31,202,31,202,30,38,31,169,31,169,30,203,31,247,31,247,30,20,31,89,31,69,31,53,31,83,31,83,30,36,31,90,31,90,30,55,31,94,31,193,31,189,31,189,30,239,31,45,31,27,31,144,31,51,31,132,31,20,31,206,31,206,31,206,30,83,31,14,31,157,31,162,31,102,31,203,31,103,31,103,30,103,29,103,31,122,31,176,31,248,31,220,31,220,30,37,31,200,31,200,30,78,31,18,31,109,31,210,31,210,30,72,31,237,31,223,31,151,31,29,31,197,31,172,31,172,30,57,31,222,31,14,31,123,31,101,31,237,31,19,31,19,30,19,29,33,31,33,30,230,31,194,31,47,31,134,31,46,31,46,30,77,31,37,31,24,31,33,31,20,31,213,31,175,31,175,30,166,31,166,30,51,31,51,30,68,31,68,30,158,31,224,31,133,31,133,30,21,31,121,31,121,30,104,31,104,30,104,29,162,31,223,31,252,31,174,31,6,31,180,31,180,30,178,31,178,30,149,31,43,31,148,31,148,30,60,31,114,31,168,31,168,30,59,31,59,30,84,31,241,31,167,31,147,31,109,31,252,31,59,31,72,31,220,31,220,30,173,31,222,31,97,31,240,31,150,31,73,31,49,31,183,31,229,31,229,30,229,29,179,31,220,31,204,31,240,31,35,31,35,31,82,31,200,31,236,31,93,31,25,31,173,31,173,30,255,31,255,30,255,29,172,31,110,31,204,31,204,30,22,31,89,31,209,31,54,31,235,31,161,31,90,31,62,31,95,31,36,31,4,31,28,31,209,31,27,31,116,31,129,31,146,31,46,31,223,31,223,30,223,29,223,28,252,31,30,31,108,31,108,30,57,31,253,31,160,31,248,31,248,30,49,31,125,31,41,31,175,31,175,30,134,31,231,31,62,31,38,31,69,31,157,31,196,31,6,31,58,31,104,31,73,31,73,30,16,31,80,31,13,31,222,31,241,31,56,31,200,31,119,31,161,31,182,31,132,31,193,31,210,31,210,30,129,31,129,30,244,31,219,31,226,31,229,31,40,31,40,30,14,31,14,30,14,29,164,31,164,30,92,31,170,31,138,31,138,30,96,31,23,31,23,30,100,31,100,30,98,31,106,31,165,31,116,31,228,31,215,31,98,31,24,31,24,30,24,29,90,31,237,31,103,31,252,31,179,31,246,31,98,31,148,31,186,31,186,30,10,31,21,31,77,31,53,31,148,31,25,31,185,31,185,30,185,29,114,31,219,31,165,31,65,31,65,30,29,31,12,31,195,31,172,31,14,31,90,31,204,31,68,31,118,31,118,30,150,31,150,30,22,31,131,31,178,31,28,31,28,30,28,29,81,31,81,30,141,31,74,31,173,31,173,30,65,31,100,31,18,31,141,31,56,31,161,31,11,31,240,31,205,31,47,31,63,31,161,31,59,31,172,31,249,31,253,31,181,31,173,31,56,31,224,31,246,31,203,31,203,30,60,31,64,31,70,31,68,31,143,31,251,31,248,31,90,31,152,31,115,31,115,30,251,31,251,30,68,31,68,30,97,31,169,31,169,30,114,31,78,31,26,31,26,30,205,31,158,31,127,31,19,31,209,31,70,31,255,31,47,31,103,31,176,31,255,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
