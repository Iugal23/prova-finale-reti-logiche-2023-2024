-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 447;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (8,0,19,0,113,0,210,0,153,0,136,0,44,0,191,0,203,0,214,0,175,0,237,0,0,0,69,0,151,0,31,0,0,0,0,0,75,0,0,0,0,0,17,0,254,0,7,0,0,0,211,0,132,0,66,0,0,0,15,0,45,0,207,0,149,0,102,0,216,0,176,0,53,0,0,0,0,0,233,0,33,0,95,0,66,0,165,0,116,0,0,0,122,0,91,0,206,0,0,0,18,0,205,0,218,0,92,0,220,0,178,0,62,0,39,0,167,0,28,0,47,0,233,0,0,0,48,0,149,0,0,0,105,0,120,0,141,0,64,0,14,0,236,0,175,0,72,0,254,0,84,0,239,0,200,0,131,0,127,0,0,0,106,0,216,0,30,0,0,0,85,0,142,0,23,0,25,0,215,0,0,0,0,0,186,0,177,0,0,0,118,0,22,0,17,0,143,0,0,0,160,0,167,0,0,0,31,0,0,0,232,0,0,0,171,0,19,0,6,0,32,0,116,0,0,0,108,0,98,0,166,0,142,0,0,0,74,0,171,0,161,0,0,0,181,0,220,0,38,0,8,0,84,0,1,0,221,0,134,0,0,0,162,0,170,0,216,0,253,0,0,0,254,0,121,0,62,0,201,0,0,0,0,0,181,0,49,0,0,0,214,0,73,0,59,0,165,0,202,0,249,0,81,0,0,0,140,0,0,0,0,0,215,0,232,0,55,0,13,0,203,0,210,0,71,0,0,0,200,0,19,0,154,0,13,0,111,0,158,0,93,0,231,0,207,0,0,0,173,0,58,0,172,0,0,0,0,0,32,0,0,0,150,0,161,0,4,0,0,0,0,0,160,0,0,0,0,0,230,0,0,0,146,0,236,0,240,0,104,0,147,0,79,0,0,0,93,0,134,0,0,0,108,0,246,0,56,0,68,0,39,0,54,0,25,0,239,0,205,0,253,0,211,0,67,0,39,0,15,0,139,0,0,0,44,0,1,0,184,0,20,0,5,0,0,0,0,0,138,0,0,0,243,0,186,0,197,0,18,0,0,0,169,0,247,0,195,0,84,0,184,0,248,0,68,0,203,0,220,0,0,0,0,0,230,0,127,0,0,0,228,0,213,0,76,0,71,0,150,0,202,0,124,0,0,0,234,0,87,0,156,0,160,0,65,0,114,0,0,0,140,0,4,0,0,0,0,0,115,0,231,0,54,0,75,0,0,0,0,0,0,0,119,0,51,0,0,0,217,0,44,0,60,0,124,0,230,0,198,0,240,0,82,0,84,0,175,0,125,0,118,0,213,0,0,0,171,0,199,0,167,0,108,0,50,0,102,0,86,0,159,0,0,0,27,0,90,0,0,0,163,0,150,0,41,0,72,0,100,0,147,0,5,0,143,0,109,0,167,0,250,0,44,0,200,0,166,0,82,0,122,0,0,0,0,0,25,0,0,0,0,0,0,0,150,0,17,0,32,0,0,0,0,0,117,0,215,0,11,0,171,0,0,0,120,0,66,0,99,0,255,0,93,0,33,0,177,0,221,0,254,0,0,0,89,0,155,0,0,0,143,0,216,0,188,0,0,0,0,0,108,0,0,0,104,0,95,0,0,0,184,0,81,0,114,0,137,0,130,0,19,0,129,0,0,0,0,0,123,0,132,0,0,0,69,0,81,0,106,0,247,0,77,0,0,0,241,0,77,0,145,0,25,0,119,0,208,0,131,0,0,0,43,0,0,0,8,0,0,0,2,0,0,0,0,0,41,0,1,0,180,0,0,0,221,0,243,0,196,0,201,0,26,0,135,0,110,0,43,0,247,0,186,0,130,0,0,0,20,0,84,0,109,0,4,0,148,0,228,0,219,0,0,0,8,0,176,0,148,0,0,0,154,0,146,0,0,0,89,0,253,0,108,0,175,0,0,0,102,0,200,0,56,0,61,0,241,0,37,0,186,0,0,0,192,0,248,0,32,0,93,0,140,0,203,0,192,0,220,0,5,0,112,0,170,0,165,0,31,0,205,0,228,0);
signal scenario_full  : scenario_type := (8,31,19,31,113,31,210,31,153,31,136,31,44,31,191,31,203,31,214,31,175,31,237,31,237,30,69,31,151,31,31,31,31,30,31,29,75,31,75,30,75,29,17,31,254,31,7,31,7,30,211,31,132,31,66,31,66,30,15,31,45,31,207,31,149,31,102,31,216,31,176,31,53,31,53,30,53,29,233,31,33,31,95,31,66,31,165,31,116,31,116,30,122,31,91,31,206,31,206,30,18,31,205,31,218,31,92,31,220,31,178,31,62,31,39,31,167,31,28,31,47,31,233,31,233,30,48,31,149,31,149,30,105,31,120,31,141,31,64,31,14,31,236,31,175,31,72,31,254,31,84,31,239,31,200,31,131,31,127,31,127,30,106,31,216,31,30,31,30,30,85,31,142,31,23,31,25,31,215,31,215,30,215,29,186,31,177,31,177,30,118,31,22,31,17,31,143,31,143,30,160,31,167,31,167,30,31,31,31,30,232,31,232,30,171,31,19,31,6,31,32,31,116,31,116,30,108,31,98,31,166,31,142,31,142,30,74,31,171,31,161,31,161,30,181,31,220,31,38,31,8,31,84,31,1,31,221,31,134,31,134,30,162,31,170,31,216,31,253,31,253,30,254,31,121,31,62,31,201,31,201,30,201,29,181,31,49,31,49,30,214,31,73,31,59,31,165,31,202,31,249,31,81,31,81,30,140,31,140,30,140,29,215,31,232,31,55,31,13,31,203,31,210,31,71,31,71,30,200,31,19,31,154,31,13,31,111,31,158,31,93,31,231,31,207,31,207,30,173,31,58,31,172,31,172,30,172,29,32,31,32,30,150,31,161,31,4,31,4,30,4,29,160,31,160,30,160,29,230,31,230,30,146,31,236,31,240,31,104,31,147,31,79,31,79,30,93,31,134,31,134,30,108,31,246,31,56,31,68,31,39,31,54,31,25,31,239,31,205,31,253,31,211,31,67,31,39,31,15,31,139,31,139,30,44,31,1,31,184,31,20,31,5,31,5,30,5,29,138,31,138,30,243,31,186,31,197,31,18,31,18,30,169,31,247,31,195,31,84,31,184,31,248,31,68,31,203,31,220,31,220,30,220,29,230,31,127,31,127,30,228,31,213,31,76,31,71,31,150,31,202,31,124,31,124,30,234,31,87,31,156,31,160,31,65,31,114,31,114,30,140,31,4,31,4,30,4,29,115,31,231,31,54,31,75,31,75,30,75,29,75,28,119,31,51,31,51,30,217,31,44,31,60,31,124,31,230,31,198,31,240,31,82,31,84,31,175,31,125,31,118,31,213,31,213,30,171,31,199,31,167,31,108,31,50,31,102,31,86,31,159,31,159,30,27,31,90,31,90,30,163,31,150,31,41,31,72,31,100,31,147,31,5,31,143,31,109,31,167,31,250,31,44,31,200,31,166,31,82,31,122,31,122,30,122,29,25,31,25,30,25,29,25,28,150,31,17,31,32,31,32,30,32,29,117,31,215,31,11,31,171,31,171,30,120,31,66,31,99,31,255,31,93,31,33,31,177,31,221,31,254,31,254,30,89,31,155,31,155,30,143,31,216,31,188,31,188,30,188,29,108,31,108,30,104,31,95,31,95,30,184,31,81,31,114,31,137,31,130,31,19,31,129,31,129,30,129,29,123,31,132,31,132,30,69,31,81,31,106,31,247,31,77,31,77,30,241,31,77,31,145,31,25,31,119,31,208,31,131,31,131,30,43,31,43,30,8,31,8,30,2,31,2,30,2,29,41,31,1,31,180,31,180,30,221,31,243,31,196,31,201,31,26,31,135,31,110,31,43,31,247,31,186,31,130,31,130,30,20,31,84,31,109,31,4,31,148,31,228,31,219,31,219,30,8,31,176,31,148,31,148,30,154,31,146,31,146,30,89,31,253,31,108,31,175,31,175,30,102,31,200,31,56,31,61,31,241,31,37,31,186,31,186,30,192,31,248,31,32,31,93,31,140,31,203,31,192,31,220,31,5,31,112,31,170,31,165,31,31,31,205,31,228,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
