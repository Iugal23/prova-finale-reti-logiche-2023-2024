-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 265;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (175,0,233,0,174,0,202,0,0,0,7,0,12,0,34,0,0,0,0,0,218,0,34,0,128,0,17,0,53,0,125,0,0,0,214,0,0,0,160,0,136,0,78,0,138,0,0,0,0,0,178,0,0,0,0,0,220,0,0,0,240,0,0,0,244,0,84,0,0,0,162,0,236,0,109,0,111,0,175,0,26,0,178,0,33,0,0,0,71,0,157,0,0,0,72,0,0,0,136,0,66,0,26,0,186,0,0,0,236,0,97,0,188,0,0,0,0,0,102,0,136,0,219,0,132,0,249,0,102,0,173,0,131,0,208,0,22,0,0,0,0,0,180,0,90,0,0,0,171,0,43,0,189,0,142,0,94,0,70,0,154,0,0,0,169,0,0,0,186,0,252,0,17,0,125,0,160,0,0,0,77,0,209,0,0,0,153,0,0,0,35,0,0,0,23,0,162,0,0,0,189,0,235,0,117,0,189,0,116,0,52,0,86,0,94,0,18,0,248,0,246,0,119,0,249,0,152,0,0,0,160,0,222,0,0,0,0,0,170,0,65,0,162,0,0,0,228,0,69,0,19,0,115,0,0,0,0,0,218,0,42,0,64,0,0,0,10,0,156,0,231,0,202,0,28,0,0,0,0,0,169,0,0,0,54,0,11,0,19,0,153,0,255,0,99,0,97,0,108,0,135,0,126,0,227,0,45,0,0,0,181,0,180,0,158,0,0,0,131,0,65,0,0,0,162,0,228,0,131,0,99,0,102,0,122,0,0,0,0,0,0,0,0,0,223,0,114,0,0,0,125,0,127,0,0,0,173,0,103,0,74,0,198,0,199,0,186,0,70,0,0,0,39,0,100,0,177,0,0,0,192,0,212,0,228,0,22,0,0,0,0,0,0,0,57,0,22,0,0,0,93,0,21,0,0,0,148,0,168,0,81,0,121,0,105,0,13,0,168,0,0,0,82,0,185,0,152,0,0,0,141,0,213,0,107,0,36,0,0,0,0,0,98,0,0,0,212,0,0,0,122,0,67,0,67,0,190,0,112,0,208,0,0,0,246,0,217,0,0,0,79,0,143,0,202,0,148,0,212,0,115,0,0,0,101,0,174,0,177,0,95,0,0,0,15,0,109,0,0,0,0,0,231,0,252,0,190,0,37,0,31,0,99,0,192,0,24,0,62,0,0,0,0,0,150,0,11,0,96,0);
signal scenario_full  : scenario_type := (175,31,233,31,174,31,202,31,202,30,7,31,12,31,34,31,34,30,34,29,218,31,34,31,128,31,17,31,53,31,125,31,125,30,214,31,214,30,160,31,136,31,78,31,138,31,138,30,138,29,178,31,178,30,178,29,220,31,220,30,240,31,240,30,244,31,84,31,84,30,162,31,236,31,109,31,111,31,175,31,26,31,178,31,33,31,33,30,71,31,157,31,157,30,72,31,72,30,136,31,66,31,26,31,186,31,186,30,236,31,97,31,188,31,188,30,188,29,102,31,136,31,219,31,132,31,249,31,102,31,173,31,131,31,208,31,22,31,22,30,22,29,180,31,90,31,90,30,171,31,43,31,189,31,142,31,94,31,70,31,154,31,154,30,169,31,169,30,186,31,252,31,17,31,125,31,160,31,160,30,77,31,209,31,209,30,153,31,153,30,35,31,35,30,23,31,162,31,162,30,189,31,235,31,117,31,189,31,116,31,52,31,86,31,94,31,18,31,248,31,246,31,119,31,249,31,152,31,152,30,160,31,222,31,222,30,222,29,170,31,65,31,162,31,162,30,228,31,69,31,19,31,115,31,115,30,115,29,218,31,42,31,64,31,64,30,10,31,156,31,231,31,202,31,28,31,28,30,28,29,169,31,169,30,54,31,11,31,19,31,153,31,255,31,99,31,97,31,108,31,135,31,126,31,227,31,45,31,45,30,181,31,180,31,158,31,158,30,131,31,65,31,65,30,162,31,228,31,131,31,99,31,102,31,122,31,122,30,122,29,122,28,122,27,223,31,114,31,114,30,125,31,127,31,127,30,173,31,103,31,74,31,198,31,199,31,186,31,70,31,70,30,39,31,100,31,177,31,177,30,192,31,212,31,228,31,22,31,22,30,22,29,22,28,57,31,22,31,22,30,93,31,21,31,21,30,148,31,168,31,81,31,121,31,105,31,13,31,168,31,168,30,82,31,185,31,152,31,152,30,141,31,213,31,107,31,36,31,36,30,36,29,98,31,98,30,212,31,212,30,122,31,67,31,67,31,190,31,112,31,208,31,208,30,246,31,217,31,217,30,79,31,143,31,202,31,148,31,212,31,115,31,115,30,101,31,174,31,177,31,95,31,95,30,15,31,109,31,109,30,109,29,231,31,252,31,190,31,37,31,31,31,99,31,192,31,24,31,62,31,62,30,62,29,150,31,11,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
