-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 352;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,155,0,11,0,131,0,91,0,197,0,110,0,0,0,0,0,192,0,143,0,0,0,152,0,147,0,0,0,234,0,0,0,196,0,103,0,0,0,149,0,241,0,38,0,183,0,5,0,224,0,232,0,0,0,0,0,175,0,0,0,76,0,205,0,117,0,191,0,60,0,45,0,142,0,29,0,101,0,0,0,0,0,237,0,112,0,182,0,0,0,156,0,0,0,0,0,0,0,43,0,106,0,28,0,109,0,139,0,183,0,28,0,140,0,111,0,2,0,99,0,0,0,224,0,0,0,229,0,63,0,52,0,229,0,116,0,252,0,0,0,227,0,192,0,230,0,90,0,222,0,49,0,193,0,37,0,88,0,0,0,133,0,248,0,104,0,213,0,29,0,0,0,196,0,233,0,148,0,0,0,0,0,135,0,209,0,143,0,0,0,67,0,191,0,243,0,0,0,53,0,10,0,54,0,0,0,241,0,40,0,174,0,110,0,78,0,238,0,0,0,239,0,0,0,95,0,81,0,133,0,254,0,0,0,39,0,147,0,182,0,167,0,165,0,180,0,0,0,204,0,156,0,67,0,68,0,184,0,70,0,99,0,248,0,255,0,115,0,205,0,0,0,206,0,47,0,164,0,0,0,229,0,112,0,172,0,106,0,0,0,0,0,246,0,232,0,0,0,127,0,70,0,0,0,223,0,13,0,238,0,84,0,38,0,147,0,0,0,140,0,172,0,126,0,4,0,69,0,179,0,0,0,17,0,0,0,71,0,62,0,139,0,213,0,226,0,172,0,0,0,234,0,106,0,78,0,79,0,56,0,43,0,0,0,135,0,148,0,197,0,0,0,243,0,6,0,0,0,222,0,2,0,129,0,138,0,104,0,168,0,189,0,102,0,0,0,49,0,91,0,144,0,0,0,32,0,108,0,0,0,86,0,0,0,44,0,0,0,241,0,0,0,66,0,185,0,166,0,181,0,0,0,43,0,64,0,146,0,49,0,119,0,207,0,193,0,63,0,0,0,0,0,231,0,14,0,108,0,131,0,248,0,0,0,60,0,105,0,0,0,212,0,163,0,162,0,31,0,0,0,18,0,0,0,103,0,123,0,253,0,23,0,98,0,0,0,205,0,0,0,230,0,212,0,186,0,116,0,220,0,101,0,140,0,181,0,188,0,220,0,200,0,107,0,115,0,0,0,227,0,0,0,54,0,39,0,18,0,38,0,0,0,67,0,38,0,117,0,61,0,194,0,0,0,36,0,60,0,252,0,193,0,53,0,117,0,181,0,0,0,153,0,234,0,106,0,207,0,0,0,250,0,0,0,26,0,52,0,0,0,0,0,0,0,35,0,251,0,50,0,12,0,141,0,25,0,0,0,166,0,0,0,76,0,28,0,117,0,4,0,176,0,224,0,2,0,0,0,137,0,27,0,0,0,54,0,68,0,135,0,0,0,187,0,243,0,220,0,116,0,168,0,0,0,116,0,0,0,2,0,115,0,0,0,13,0,213,0,76,0,0,0,128,0,0,0,213,0,239,0,0,0,86,0,224,0,211,0,83,0,180,0,138,0,219,0,234,0,154,0,28,0);
signal scenario_full  : scenario_type := (136,31,155,31,11,31,131,31,91,31,197,31,110,31,110,30,110,29,192,31,143,31,143,30,152,31,147,31,147,30,234,31,234,30,196,31,103,31,103,30,149,31,241,31,38,31,183,31,5,31,224,31,232,31,232,30,232,29,175,31,175,30,76,31,205,31,117,31,191,31,60,31,45,31,142,31,29,31,101,31,101,30,101,29,237,31,112,31,182,31,182,30,156,31,156,30,156,29,156,28,43,31,106,31,28,31,109,31,139,31,183,31,28,31,140,31,111,31,2,31,99,31,99,30,224,31,224,30,229,31,63,31,52,31,229,31,116,31,252,31,252,30,227,31,192,31,230,31,90,31,222,31,49,31,193,31,37,31,88,31,88,30,133,31,248,31,104,31,213,31,29,31,29,30,196,31,233,31,148,31,148,30,148,29,135,31,209,31,143,31,143,30,67,31,191,31,243,31,243,30,53,31,10,31,54,31,54,30,241,31,40,31,174,31,110,31,78,31,238,31,238,30,239,31,239,30,95,31,81,31,133,31,254,31,254,30,39,31,147,31,182,31,167,31,165,31,180,31,180,30,204,31,156,31,67,31,68,31,184,31,70,31,99,31,248,31,255,31,115,31,205,31,205,30,206,31,47,31,164,31,164,30,229,31,112,31,172,31,106,31,106,30,106,29,246,31,232,31,232,30,127,31,70,31,70,30,223,31,13,31,238,31,84,31,38,31,147,31,147,30,140,31,172,31,126,31,4,31,69,31,179,31,179,30,17,31,17,30,71,31,62,31,139,31,213,31,226,31,172,31,172,30,234,31,106,31,78,31,79,31,56,31,43,31,43,30,135,31,148,31,197,31,197,30,243,31,6,31,6,30,222,31,2,31,129,31,138,31,104,31,168,31,189,31,102,31,102,30,49,31,91,31,144,31,144,30,32,31,108,31,108,30,86,31,86,30,44,31,44,30,241,31,241,30,66,31,185,31,166,31,181,31,181,30,43,31,64,31,146,31,49,31,119,31,207,31,193,31,63,31,63,30,63,29,231,31,14,31,108,31,131,31,248,31,248,30,60,31,105,31,105,30,212,31,163,31,162,31,31,31,31,30,18,31,18,30,103,31,123,31,253,31,23,31,98,31,98,30,205,31,205,30,230,31,212,31,186,31,116,31,220,31,101,31,140,31,181,31,188,31,220,31,200,31,107,31,115,31,115,30,227,31,227,30,54,31,39,31,18,31,38,31,38,30,67,31,38,31,117,31,61,31,194,31,194,30,36,31,60,31,252,31,193,31,53,31,117,31,181,31,181,30,153,31,234,31,106,31,207,31,207,30,250,31,250,30,26,31,52,31,52,30,52,29,52,28,35,31,251,31,50,31,12,31,141,31,25,31,25,30,166,31,166,30,76,31,28,31,117,31,4,31,176,31,224,31,2,31,2,30,137,31,27,31,27,30,54,31,68,31,135,31,135,30,187,31,243,31,220,31,116,31,168,31,168,30,116,31,116,30,2,31,115,31,115,30,13,31,213,31,76,31,76,30,128,31,128,30,213,31,239,31,239,30,86,31,224,31,211,31,83,31,180,31,138,31,219,31,234,31,154,31,28,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
