-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 542;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (235,0,107,0,118,0,113,0,3,0,0,0,185,0,157,0,101,0,0,0,94,0,181,0,246,0,202,0,141,0,196,0,227,0,30,0,0,0,0,0,116,0,193,0,239,0,73,0,0,0,146,0,7,0,248,0,3,0,243,0,199,0,0,0,208,0,37,0,32,0,167,0,45,0,104,0,0,0,205,0,52,0,141,0,47,0,0,0,206,0,74,0,68,0,214,0,138,0,142,0,0,0,0,0,147,0,250,0,68,0,246,0,141,0,204,0,225,0,237,0,16,0,25,0,186,0,0,0,237,0,0,0,252,0,88,0,152,0,239,0,244,0,45,0,0,0,76,0,225,0,153,0,174,0,41,0,109,0,110,0,2,0,178,0,149,0,18,0,0,0,125,0,184,0,127,0,175,0,0,0,18,0,0,0,56,0,0,0,148,0,65,0,0,0,89,0,106,0,0,0,222,0,0,0,120,0,63,0,255,0,100,0,105,0,145,0,101,0,201,0,98,0,117,0,179,0,132,0,127,0,0,0,61,0,131,0,45,0,176,0,100,0,50,0,145,0,246,0,142,0,0,0,170,0,125,0,79,0,219,0,0,0,39,0,0,0,205,0,220,0,0,0,105,0,62,0,0,0,188,0,19,0,98,0,84,0,244,0,103,0,14,0,194,0,128,0,166,0,0,0,184,0,0,0,124,0,238,0,198,0,0,0,77,0,212,0,0,0,247,0,78,0,90,0,121,0,9,0,64,0,0,0,58,0,114,0,7,0,65,0,47,0,42,0,222,0,254,0,164,0,54,0,198,0,199,0,35,0,190,0,44,0,215,0,0,0,70,0,9,0,0,0,254,0,122,0,0,0,175,0,51,0,106,0,244,0,190,0,141,0,0,0,41,0,15,0,39,0,216,0,87,0,137,0,233,0,0,0,34,0,154,0,81,0,34,0,214,0,44,0,0,0,74,0,6,0,0,0,240,0,85,0,116,0,192,0,30,0,224,0,56,0,136,0,172,0,219,0,29,0,194,0,0,0,54,0,43,0,133,0,0,0,123,0,0,0,0,0,235,0,0,0,0,0,201,0,5,0,211,0,28,0,153,0,128,0,20,0,37,0,0,0,2,0,34,0,23,0,222,0,0,0,241,0,102,0,194,0,0,0,0,0,32,0,0,0,14,0,107,0,0,0,0,0,88,0,78,0,27,0,202,0,0,0,252,0,229,0,211,0,37,0,0,0,0,0,112,0,72,0,60,0,229,0,108,0,145,0,129,0,164,0,8,0,0,0,234,0,183,0,110,0,20,0,0,0,0,0,193,0,223,0,190,0,76,0,117,0,0,0,140,0,0,0,0,0,181,0,104,0,125,0,254,0,197,0,140,0,0,0,203,0,19,0,0,0,0,0,149,0,0,0,83,0,236,0,0,0,64,0,164,0,61,0,0,0,168,0,0,0,186,0,45,0,36,0,234,0,160,0,91,0,0,0,0,0,22,0,118,0,107,0,255,0,18,0,0,0,233,0,0,0,149,0,92,0,230,0,188,0,23,0,40,0,190,0,98,0,168,0,0,0,151,0,87,0,110,0,0,0,113,0,24,0,127,0,35,0,118,0,0,0,146,0,190,0,116,0,215,0,0,0,104,0,0,0,137,0,2,0,0,0,239,0,56,0,87,0,93,0,60,0,248,0,54,0,34,0,0,0,211,0,189,0,1,0,131,0,128,0,91,0,191,0,76,0,143,0,211,0,0,0,82,0,146,0,0,0,175,0,130,0,182,0,38,0,119,0,56,0,10,0,78,0,20,0,0,0,251,0,52,0,214,0,0,0,63,0,67,0,5,0,81,0,170,0,0,0,8,0,174,0,97,0,247,0,93,0,137,0,0,0,1,0,81,0,0,0,112,0,34,0,210,0,130,0,0,0,52,0,129,0,244,0,104,0,0,0,115,0,172,0,42,0,47,0,241,0,150,0,0,0,152,0,243,0,225,0,113,0,101,0,0,0,60,0,68,0,0,0,0,0,41,0,8,0,171,0,137,0,50,0,52,0,26,0,168,0,22,0,209,0,0,0,143,0,203,0,168,0,188,0,249,0,190,0,95,0,0,0,222,0,9,0,93,0,2,0,182,0,0,0,65,0,78,0,0,0,57,0,138,0,225,0,167,0,145,0,134,0,54,0,242,0,202,0,5,0,166,0,21,0,0,0,237,0,0,0,82,0,81,0,217,0,0,0,221,0,185,0,109,0,0,0,9,0,0,0,0,0,222,0,156,0,162,0,3,0,183,0,17,0,148,0,0,0,28,0,147,0,189,0,0,0,169,0,162,0,0,0,115,0,124,0,130,0,98,0,60,0,53,0,0,0,205,0,0,0,230,0,159,0,48,0,0,0,149,0,98,0,133,0,0,0,48,0,140,0,99,0,255,0,106,0,0,0,242,0,2,0,192,0,67,0);
signal scenario_full  : scenario_type := (235,31,107,31,118,31,113,31,3,31,3,30,185,31,157,31,101,31,101,30,94,31,181,31,246,31,202,31,141,31,196,31,227,31,30,31,30,30,30,29,116,31,193,31,239,31,73,31,73,30,146,31,7,31,248,31,3,31,243,31,199,31,199,30,208,31,37,31,32,31,167,31,45,31,104,31,104,30,205,31,52,31,141,31,47,31,47,30,206,31,74,31,68,31,214,31,138,31,142,31,142,30,142,29,147,31,250,31,68,31,246,31,141,31,204,31,225,31,237,31,16,31,25,31,186,31,186,30,237,31,237,30,252,31,88,31,152,31,239,31,244,31,45,31,45,30,76,31,225,31,153,31,174,31,41,31,109,31,110,31,2,31,178,31,149,31,18,31,18,30,125,31,184,31,127,31,175,31,175,30,18,31,18,30,56,31,56,30,148,31,65,31,65,30,89,31,106,31,106,30,222,31,222,30,120,31,63,31,255,31,100,31,105,31,145,31,101,31,201,31,98,31,117,31,179,31,132,31,127,31,127,30,61,31,131,31,45,31,176,31,100,31,50,31,145,31,246,31,142,31,142,30,170,31,125,31,79,31,219,31,219,30,39,31,39,30,205,31,220,31,220,30,105,31,62,31,62,30,188,31,19,31,98,31,84,31,244,31,103,31,14,31,194,31,128,31,166,31,166,30,184,31,184,30,124,31,238,31,198,31,198,30,77,31,212,31,212,30,247,31,78,31,90,31,121,31,9,31,64,31,64,30,58,31,114,31,7,31,65,31,47,31,42,31,222,31,254,31,164,31,54,31,198,31,199,31,35,31,190,31,44,31,215,31,215,30,70,31,9,31,9,30,254,31,122,31,122,30,175,31,51,31,106,31,244,31,190,31,141,31,141,30,41,31,15,31,39,31,216,31,87,31,137,31,233,31,233,30,34,31,154,31,81,31,34,31,214,31,44,31,44,30,74,31,6,31,6,30,240,31,85,31,116,31,192,31,30,31,224,31,56,31,136,31,172,31,219,31,29,31,194,31,194,30,54,31,43,31,133,31,133,30,123,31,123,30,123,29,235,31,235,30,235,29,201,31,5,31,211,31,28,31,153,31,128,31,20,31,37,31,37,30,2,31,34,31,23,31,222,31,222,30,241,31,102,31,194,31,194,30,194,29,32,31,32,30,14,31,107,31,107,30,107,29,88,31,78,31,27,31,202,31,202,30,252,31,229,31,211,31,37,31,37,30,37,29,112,31,72,31,60,31,229,31,108,31,145,31,129,31,164,31,8,31,8,30,234,31,183,31,110,31,20,31,20,30,20,29,193,31,223,31,190,31,76,31,117,31,117,30,140,31,140,30,140,29,181,31,104,31,125,31,254,31,197,31,140,31,140,30,203,31,19,31,19,30,19,29,149,31,149,30,83,31,236,31,236,30,64,31,164,31,61,31,61,30,168,31,168,30,186,31,45,31,36,31,234,31,160,31,91,31,91,30,91,29,22,31,118,31,107,31,255,31,18,31,18,30,233,31,233,30,149,31,92,31,230,31,188,31,23,31,40,31,190,31,98,31,168,31,168,30,151,31,87,31,110,31,110,30,113,31,24,31,127,31,35,31,118,31,118,30,146,31,190,31,116,31,215,31,215,30,104,31,104,30,137,31,2,31,2,30,239,31,56,31,87,31,93,31,60,31,248,31,54,31,34,31,34,30,211,31,189,31,1,31,131,31,128,31,91,31,191,31,76,31,143,31,211,31,211,30,82,31,146,31,146,30,175,31,130,31,182,31,38,31,119,31,56,31,10,31,78,31,20,31,20,30,251,31,52,31,214,31,214,30,63,31,67,31,5,31,81,31,170,31,170,30,8,31,174,31,97,31,247,31,93,31,137,31,137,30,1,31,81,31,81,30,112,31,34,31,210,31,130,31,130,30,52,31,129,31,244,31,104,31,104,30,115,31,172,31,42,31,47,31,241,31,150,31,150,30,152,31,243,31,225,31,113,31,101,31,101,30,60,31,68,31,68,30,68,29,41,31,8,31,171,31,137,31,50,31,52,31,26,31,168,31,22,31,209,31,209,30,143,31,203,31,168,31,188,31,249,31,190,31,95,31,95,30,222,31,9,31,93,31,2,31,182,31,182,30,65,31,78,31,78,30,57,31,138,31,225,31,167,31,145,31,134,31,54,31,242,31,202,31,5,31,166,31,21,31,21,30,237,31,237,30,82,31,81,31,217,31,217,30,221,31,185,31,109,31,109,30,9,31,9,30,9,29,222,31,156,31,162,31,3,31,183,31,17,31,148,31,148,30,28,31,147,31,189,31,189,30,169,31,162,31,162,30,115,31,124,31,130,31,98,31,60,31,53,31,53,30,205,31,205,30,230,31,159,31,48,31,48,30,149,31,98,31,133,31,133,30,48,31,140,31,99,31,255,31,106,31,106,30,242,31,2,31,192,31,67,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
