-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_206 is
end project_tb_206;

architecture project_tb_arch_206 of project_tb_206 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 417;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (123,0,170,0,0,0,241,0,178,0,117,0,174,0,172,0,101,0,89,0,245,0,36,0,143,0,100,0,38,0,94,0,182,0,196,0,0,0,49,0,1,0,61,0,134,0,154,0,13,0,209,0,193,0,105,0,205,0,0,0,89,0,0,0,148,0,185,0,119,0,27,0,54,0,0,0,37,0,169,0,23,0,19,0,163,0,0,0,0,0,0,0,86,0,111,0,142,0,0,0,0,0,140,0,169,0,14,0,0,0,0,0,137,0,99,0,246,0,210,0,0,0,78,0,147,0,53,0,115,0,224,0,124,0,28,0,0,0,168,0,191,0,235,0,161,0,71,0,128,0,71,0,0,0,189,0,209,0,164,0,0,0,93,0,238,0,146,0,0,0,234,0,164,0,23,0,0,0,0,0,0,0,7,0,0,0,179,0,113,0,233,0,159,0,61,0,159,0,0,0,139,0,10,0,0,0,123,0,42,0,234,0,204,0,105,0,167,0,185,0,118,0,10,0,245,0,49,0,247,0,179,0,0,0,125,0,0,0,167,0,23,0,203,0,87,0,207,0,86,0,200,0,185,0,37,0,29,0,213,0,72,0,228,0,82,0,142,0,25,0,254,0,103,0,99,0,0,0,63,0,45,0,12,0,118,0,0,0,36,0,0,0,5,0,242,0,102,0,170,0,109,0,0,0,197,0,140,0,100,0,103,0,0,0,69,0,161,0,84,0,253,0,123,0,1,0,3,0,177,0,22,0,43,0,94,0,228,0,38,0,61,0,164,0,56,0,183,0,175,0,14,0,0,0,243,0,236,0,124,0,0,0,134,0,29,0,83,0,0,0,122,0,0,0,0,0,0,0,148,0,0,0,132,0,119,0,96,0,131,0,154,0,222,0,135,0,217,0,0,0,79,0,142,0,226,0,28,0,196,0,201,0,154,0,24,0,181,0,10,0,32,0,6,0,125,0,71,0,223,0,122,0,202,0,53,0,64,0,29,0,29,0,123,0,189,0,156,0,31,0,237,0,238,0,6,0,189,0,195,0,86,0,0,0,96,0,135,0,233,0,146,0,34,0,231,0,0,0,100,0,254,0,194,0,0,0,155,0,243,0,184,0,0,0,119,0,184,0,142,0,0,0,0,0,105,0,8,0,184,0,186,0,146,0,51,0,109,0,236,0,98,0,145,0,123,0,12,0,193,0,242,0,142,0,0,0,70,0,0,0,231,0,212,0,214,0,254,0,0,0,0,0,180,0,58,0,36,0,0,0,192,0,188,0,155,0,0,0,192,0,0,0,7,0,45,0,220,0,0,0,3,0,0,0,18,0,194,0,36,0,249,0,0,0,193,0,0,0,43,0,0,0,40,0,219,0,65,0,148,0,120,0,118,0,122,0,84,0,0,0,0,0,160,0,58,0,105,0,61,0,91,0,142,0,106,0,85,0,143,0,0,0,178,0,0,0,243,0,117,0,31,0,102,0,12,0,216,0,11,0,55,0,106,0,125,0,0,0,91,0,101,0,137,0,47,0,32,0,219,0,215,0,0,0,0,0,0,0,114,0,19,0,108,0,34,0,31,0,0,0,200,0,96,0,21,0,132,0,33,0,139,0,0,0,85,0,38,0,71,0,113,0,232,0,250,0,138,0,196,0,204,0,37,0,167,0,163,0,188,0,207,0,0,0,147,0,117,0,62,0,236,0,0,0,112,0,153,0,39,0,0,0,150,0,0,0,162,0,234,0,191,0,255,0,88,0,70,0,168,0,53,0,247,0,50,0,40,0,0,0,37,0,196,0,129,0,151,0,7,0,234,0,0,0,0,0,240,0,0,0,202,0,128,0,27,0,0,0,0,0,0,0,0,0,17,0,0,0,221,0,0,0,0,0);
signal scenario_full  : scenario_type := (123,31,170,31,170,30,241,31,178,31,117,31,174,31,172,31,101,31,89,31,245,31,36,31,143,31,100,31,38,31,94,31,182,31,196,31,196,30,49,31,1,31,61,31,134,31,154,31,13,31,209,31,193,31,105,31,205,31,205,30,89,31,89,30,148,31,185,31,119,31,27,31,54,31,54,30,37,31,169,31,23,31,19,31,163,31,163,30,163,29,163,28,86,31,111,31,142,31,142,30,142,29,140,31,169,31,14,31,14,30,14,29,137,31,99,31,246,31,210,31,210,30,78,31,147,31,53,31,115,31,224,31,124,31,28,31,28,30,168,31,191,31,235,31,161,31,71,31,128,31,71,31,71,30,189,31,209,31,164,31,164,30,93,31,238,31,146,31,146,30,234,31,164,31,23,31,23,30,23,29,23,28,7,31,7,30,179,31,113,31,233,31,159,31,61,31,159,31,159,30,139,31,10,31,10,30,123,31,42,31,234,31,204,31,105,31,167,31,185,31,118,31,10,31,245,31,49,31,247,31,179,31,179,30,125,31,125,30,167,31,23,31,203,31,87,31,207,31,86,31,200,31,185,31,37,31,29,31,213,31,72,31,228,31,82,31,142,31,25,31,254,31,103,31,99,31,99,30,63,31,45,31,12,31,118,31,118,30,36,31,36,30,5,31,242,31,102,31,170,31,109,31,109,30,197,31,140,31,100,31,103,31,103,30,69,31,161,31,84,31,253,31,123,31,1,31,3,31,177,31,22,31,43,31,94,31,228,31,38,31,61,31,164,31,56,31,183,31,175,31,14,31,14,30,243,31,236,31,124,31,124,30,134,31,29,31,83,31,83,30,122,31,122,30,122,29,122,28,148,31,148,30,132,31,119,31,96,31,131,31,154,31,222,31,135,31,217,31,217,30,79,31,142,31,226,31,28,31,196,31,201,31,154,31,24,31,181,31,10,31,32,31,6,31,125,31,71,31,223,31,122,31,202,31,53,31,64,31,29,31,29,31,123,31,189,31,156,31,31,31,237,31,238,31,6,31,189,31,195,31,86,31,86,30,96,31,135,31,233,31,146,31,34,31,231,31,231,30,100,31,254,31,194,31,194,30,155,31,243,31,184,31,184,30,119,31,184,31,142,31,142,30,142,29,105,31,8,31,184,31,186,31,146,31,51,31,109,31,236,31,98,31,145,31,123,31,12,31,193,31,242,31,142,31,142,30,70,31,70,30,231,31,212,31,214,31,254,31,254,30,254,29,180,31,58,31,36,31,36,30,192,31,188,31,155,31,155,30,192,31,192,30,7,31,45,31,220,31,220,30,3,31,3,30,18,31,194,31,36,31,249,31,249,30,193,31,193,30,43,31,43,30,40,31,219,31,65,31,148,31,120,31,118,31,122,31,84,31,84,30,84,29,160,31,58,31,105,31,61,31,91,31,142,31,106,31,85,31,143,31,143,30,178,31,178,30,243,31,117,31,31,31,102,31,12,31,216,31,11,31,55,31,106,31,125,31,125,30,91,31,101,31,137,31,47,31,32,31,219,31,215,31,215,30,215,29,215,28,114,31,19,31,108,31,34,31,31,31,31,30,200,31,96,31,21,31,132,31,33,31,139,31,139,30,85,31,38,31,71,31,113,31,232,31,250,31,138,31,196,31,204,31,37,31,167,31,163,31,188,31,207,31,207,30,147,31,117,31,62,31,236,31,236,30,112,31,153,31,39,31,39,30,150,31,150,30,162,31,234,31,191,31,255,31,88,31,70,31,168,31,53,31,247,31,50,31,40,31,40,30,37,31,196,31,129,31,151,31,7,31,234,31,234,30,234,29,240,31,240,30,202,31,128,31,27,31,27,30,27,29,27,28,27,27,17,31,17,30,221,31,221,30,221,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
