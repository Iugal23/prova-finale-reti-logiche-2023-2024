-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 490;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,158,0,84,0,0,0,230,0,75,0,0,0,185,0,106,0,254,0,57,0,171,0,171,0,166,0,0,0,0,0,77,0,104,0,55,0,161,0,53,0,230,0,72,0,248,0,240,0,104,0,0,0,219,0,214,0,218,0,213,0,0,0,9,0,112,0,78,0,248,0,69,0,117,0,0,0,55,0,0,0,79,0,77,0,20,0,0,0,189,0,250,0,85,0,232,0,242,0,207,0,105,0,190,0,141,0,0,0,11,0,0,0,64,0,116,0,146,0,0,0,210,0,169,0,0,0,0,0,40,0,242,0,22,0,207,0,206,0,177,0,131,0,132,0,228,0,50,0,243,0,0,0,153,0,83,0,94,0,83,0,231,0,178,0,75,0,176,0,93,0,0,0,223,0,203,0,154,0,49,0,0,0,222,0,150,0,239,0,96,0,170,0,7,0,32,0,180,0,14,0,32,0,156,0,0,0,178,0,243,0,222,0,236,0,17,0,16,0,90,0,18,0,35,0,0,0,80,0,154,0,88,0,17,0,31,0,64,0,38,0,0,0,157,0,85,0,193,0,104,0,87,0,173,0,20,0,22,0,227,0,219,0,0,0,99,0,0,0,0,0,80,0,190,0,68,0,7,0,112,0,38,0,33,0,0,0,217,0,28,0,39,0,195,0,245,0,96,0,102,0,100,0,86,0,0,0,63,0,108,0,100,0,89,0,168,0,126,0,118,0,247,0,105,0,244,0,28,0,112,0,90,0,0,0,35,0,145,0,112,0,26,0,0,0,216,0,0,0,202,0,232,0,89,0,217,0,174,0,15,0,37,0,0,0,38,0,36,0,196,0,87,0,111,0,128,0,0,0,175,0,61,0,154,0,244,0,231,0,116,0,121,0,197,0,132,0,13,0,65,0,0,0,0,0,40,0,85,0,0,0,0,0,150,0,109,0,105,0,0,0,129,0,185,0,27,0,26,0,47,0,0,0,158,0,180,0,26,0,0,0,86,0,69,0,111,0,0,0,0,0,227,0,6,0,216,0,0,0,0,0,0,0,218,0,239,0,37,0,201,0,178,0,14,0,0,0,182,0,148,0,19,0,242,0,88,0,51,0,0,0,56,0,0,0,5,0,161,0,234,0,102,0,59,0,230,0,0,0,219,0,0,0,166,0,113,0,248,0,97,0,0,0,101,0,225,0,0,0,252,0,151,0,108,0,110,0,22,0,77,0,65,0,0,0,94,0,112,0,102,0,17,0,191,0,0,0,236,0,211,0,118,0,0,0,86,0,54,0,156,0,0,0,0,0,57,0,166,0,0,0,62,0,0,0,100,0,167,0,0,0,45,0,166,0,245,0,171,0,196,0,238,0,250,0,0,0,235,0,0,0,153,0,110,0,167,0,0,0,116,0,203,0,158,0,98,0,0,0,0,0,153,0,103,0,246,0,76,0,175,0,214,0,99,0,233,0,18,0,177,0,32,0,241,0,0,0,36,0,137,0,233,0,118,0,60,0,73,0,137,0,30,0,0,0,124,0,43,0,240,0,39,0,238,0,39,0,66,0,0,0,242,0,88,0,126,0,14,0,17,0,49,0,132,0,0,0,37,0,0,0,0,0,117,0,69,0,0,0,26,0,195,0,23,0,169,0,176,0,175,0,44,0,208,0,247,0,196,0,45,0,0,0,123,0,54,0,199,0,188,0,118,0,210,0,30,0,85,0,83,0,174,0,219,0,232,0,4,0,178,0,0,0,30,0,133,0,56,0,0,0,0,0,58,0,66,0,1,0,0,0,0,0,180,0,0,0,0,0,199,0,169,0,231,0,115,0,107,0,148,0,0,0,109,0,0,0,86,0,17,0,251,0,36,0,46,0,158,0,0,0,186,0,0,0,0,0,81,0,16,0,73,0,45,0,93,0,158,0,241,0,0,0,22,0,195,0,0,0,137,0,76,0,103,0,185,0,114,0,23,0,0,0,89,0,191,0,16,0,0,0,88,0,218,0,162,0,168,0,126,0,0,0,27,0,0,0,0,0,30,0,211,0,0,0,236,0,174,0,74,0,50,0,45,0,0,0,254,0,0,0,0,0,102,0,27,0,0,0,162,0,14,0,0,0,0,0,10,0,53,0,194,0,21,0,0,0,41,0,31,0,56,0,105,0,99,0,236,0,85,0,188,0,0,0,3,0,35,0,0,0,60,0,75,0,148,0,161,0);
signal scenario_full  : scenario_type := (95,31,158,31,84,31,84,30,230,31,75,31,75,30,185,31,106,31,254,31,57,31,171,31,171,31,166,31,166,30,166,29,77,31,104,31,55,31,161,31,53,31,230,31,72,31,248,31,240,31,104,31,104,30,219,31,214,31,218,31,213,31,213,30,9,31,112,31,78,31,248,31,69,31,117,31,117,30,55,31,55,30,79,31,77,31,20,31,20,30,189,31,250,31,85,31,232,31,242,31,207,31,105,31,190,31,141,31,141,30,11,31,11,30,64,31,116,31,146,31,146,30,210,31,169,31,169,30,169,29,40,31,242,31,22,31,207,31,206,31,177,31,131,31,132,31,228,31,50,31,243,31,243,30,153,31,83,31,94,31,83,31,231,31,178,31,75,31,176,31,93,31,93,30,223,31,203,31,154,31,49,31,49,30,222,31,150,31,239,31,96,31,170,31,7,31,32,31,180,31,14,31,32,31,156,31,156,30,178,31,243,31,222,31,236,31,17,31,16,31,90,31,18,31,35,31,35,30,80,31,154,31,88,31,17,31,31,31,64,31,38,31,38,30,157,31,85,31,193,31,104,31,87,31,173,31,20,31,22,31,227,31,219,31,219,30,99,31,99,30,99,29,80,31,190,31,68,31,7,31,112,31,38,31,33,31,33,30,217,31,28,31,39,31,195,31,245,31,96,31,102,31,100,31,86,31,86,30,63,31,108,31,100,31,89,31,168,31,126,31,118,31,247,31,105,31,244,31,28,31,112,31,90,31,90,30,35,31,145,31,112,31,26,31,26,30,216,31,216,30,202,31,232,31,89,31,217,31,174,31,15,31,37,31,37,30,38,31,36,31,196,31,87,31,111,31,128,31,128,30,175,31,61,31,154,31,244,31,231,31,116,31,121,31,197,31,132,31,13,31,65,31,65,30,65,29,40,31,85,31,85,30,85,29,150,31,109,31,105,31,105,30,129,31,185,31,27,31,26,31,47,31,47,30,158,31,180,31,26,31,26,30,86,31,69,31,111,31,111,30,111,29,227,31,6,31,216,31,216,30,216,29,216,28,218,31,239,31,37,31,201,31,178,31,14,31,14,30,182,31,148,31,19,31,242,31,88,31,51,31,51,30,56,31,56,30,5,31,161,31,234,31,102,31,59,31,230,31,230,30,219,31,219,30,166,31,113,31,248,31,97,31,97,30,101,31,225,31,225,30,252,31,151,31,108,31,110,31,22,31,77,31,65,31,65,30,94,31,112,31,102,31,17,31,191,31,191,30,236,31,211,31,118,31,118,30,86,31,54,31,156,31,156,30,156,29,57,31,166,31,166,30,62,31,62,30,100,31,167,31,167,30,45,31,166,31,245,31,171,31,196,31,238,31,250,31,250,30,235,31,235,30,153,31,110,31,167,31,167,30,116,31,203,31,158,31,98,31,98,30,98,29,153,31,103,31,246,31,76,31,175,31,214,31,99,31,233,31,18,31,177,31,32,31,241,31,241,30,36,31,137,31,233,31,118,31,60,31,73,31,137,31,30,31,30,30,124,31,43,31,240,31,39,31,238,31,39,31,66,31,66,30,242,31,88,31,126,31,14,31,17,31,49,31,132,31,132,30,37,31,37,30,37,29,117,31,69,31,69,30,26,31,195,31,23,31,169,31,176,31,175,31,44,31,208,31,247,31,196,31,45,31,45,30,123,31,54,31,199,31,188,31,118,31,210,31,30,31,85,31,83,31,174,31,219,31,232,31,4,31,178,31,178,30,30,31,133,31,56,31,56,30,56,29,58,31,66,31,1,31,1,30,1,29,180,31,180,30,180,29,199,31,169,31,231,31,115,31,107,31,148,31,148,30,109,31,109,30,86,31,17,31,251,31,36,31,46,31,158,31,158,30,186,31,186,30,186,29,81,31,16,31,73,31,45,31,93,31,158,31,241,31,241,30,22,31,195,31,195,30,137,31,76,31,103,31,185,31,114,31,23,31,23,30,89,31,191,31,16,31,16,30,88,31,218,31,162,31,168,31,126,31,126,30,27,31,27,30,27,29,30,31,211,31,211,30,236,31,174,31,74,31,50,31,45,31,45,30,254,31,254,30,254,29,102,31,27,31,27,30,162,31,14,31,14,30,14,29,10,31,53,31,194,31,21,31,21,30,41,31,31,31,56,31,105,31,99,31,236,31,85,31,188,31,188,30,3,31,35,31,35,30,60,31,75,31,148,31,161,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
