-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 911;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,118,0,0,0,91,0,196,0,0,0,182,0,0,0,199,0,177,0,181,0,76,0,26,0,48,0,0,0,57,0,224,0,87,0,0,0,4,0,0,0,188,0,230,0,204,0,0,0,143,0,139,0,54,0,235,0,165,0,204,0,197,0,236,0,83,0,128,0,11,0,88,0,154,0,242,0,124,0,0,0,204,0,205,0,0,0,26,0,36,0,86,0,129,0,213,0,0,0,0,0,167,0,69,0,0,0,94,0,32,0,6,0,75,0,85,0,224,0,144,0,136,0,241,0,13,0,43,0,84,0,231,0,158,0,0,0,191,0,171,0,72,0,240,0,233,0,165,0,0,0,125,0,157,0,54,0,102,0,247,0,193,0,0,0,221,0,0,0,205,0,193,0,245,0,142,0,125,0,108,0,215,0,182,0,0,0,216,0,42,0,209,0,186,0,104,0,25,0,103,0,55,0,77,0,233,0,228,0,46,0,115,0,0,0,0,0,0,0,141,0,92,0,134,0,132,0,0,0,40,0,200,0,0,0,20,0,102,0,110,0,129,0,227,0,25,0,0,0,93,0,17,0,209,0,180,0,244,0,110,0,0,0,13,0,28,0,219,0,7,0,210,0,182,0,0,0,191,0,47,0,235,0,0,0,30,0,169,0,0,0,61,0,96,0,171,0,221,0,143,0,110,0,206,0,48,0,0,0,242,0,235,0,117,0,0,0,255,0,68,0,54,0,138,0,197,0,0,0,38,0,155,0,246,0,246,0,237,0,131,0,0,0,0,0,177,0,28,0,4,0,212,0,81,0,71,0,190,0,183,0,0,0,171,0,125,0,64,0,28,0,0,0,0,0,0,0,134,0,159,0,240,0,69,0,212,0,95,0,151,0,236,0,181,0,136,0,170,0,188,0,36,0,159,0,137,0,35,0,44,0,35,0,10,0,203,0,173,0,230,0,241,0,0,0,190,0,83,0,189,0,87,0,138,0,224,0,41,0,208,0,50,0,178,0,0,0,105,0,167,0,88,0,0,0,95,0,0,0,202,0,0,0,44,0,0,0,116,0,115,0,0,0,73,0,0,0,0,0,173,0,202,0,95,0,144,0,0,0,94,0,0,0,254,0,93,0,204,0,65,0,192,0,156,0,0,0,65,0,211,0,30,0,223,0,249,0,235,0,0,0,194,0,96,0,218,0,109,0,222,0,98,0,140,0,183,0,113,0,32,0,169,0,26,0,59,0,105,0,106,0,106,0,77,0,240,0,7,0,0,0,146,0,0,0,206,0,64,0,68,0,15,0,175,0,0,0,58,0,163,0,14,0,0,0,0,0,239,0,18,0,49,0,133,0,74,0,142,0,190,0,0,0,183,0,222,0,113,0,0,0,175,0,228,0,3,0,1,0,102,0,119,0,20,0,0,0,226,0,134,0,95,0,0,0,0,0,30,0,254,0,0,0,147,0,169,0,0,0,130,0,190,0,76,0,57,0,89,0,180,0,0,0,151,0,117,0,42,0,151,0,3,0,34,0,43,0,36,0,116,0,193,0,207,0,237,0,240,0,196,0,221,0,60,0,214,0,58,0,203,0,186,0,188,0,115,0,103,0,223,0,241,0,122,0,150,0,8,0,123,0,198,0,230,0,67,0,242,0,24,0,1,0,159,0,151,0,22,0,29,0,0,0,253,0,86,0,55,0,154,0,81,0,80,0,37,0,0,0,0,0,111,0,203,0,121,0,253,0,228,0,151,0,0,0,33,0,223,0,126,0,189,0,203,0,56,0,242,0,202,0,250,0,0,0,253,0,76,0,192,0,55,0,64,0,228,0,0,0,166,0,31,0,255,0,0,0,69,0,241,0,103,0,69,0,0,0,0,0,24,0,0,0,245,0,0,0,147,0,76,0,0,0,178,0,96,0,0,0,18,0,50,0,0,0,160,0,131,0,0,0,172,0,0,0,0,0,0,0,0,0,139,0,247,0,105,0,250,0,223,0,253,0,242,0,132,0,0,0,39,0,141,0,0,0,249,0,46,0,88,0,192,0,147,0,93,0,143,0,50,0,0,0,106,0,149,0,0,0,0,0,239,0,214,0,47,0,224,0,0,0,0,0,32,0,221,0,125,0,34,0,0,0,206,0,198,0,184,0,114,0,0,0,4,0,0,0,246,0,88,0,198,0,19,0,23,0,254,0,228,0,102,0,0,0,70,0,0,0,0,0,0,0,193,0,0,0,159,0,220,0,29,0,0,0,63,0,152,0,0,0,167,0,204,0,0,0,111,0,37,0,0,0,210,0,0,0,0,0,242,0,149,0,157,0,0,0,148,0,3,0,147,0,145,0,204,0,219,0,0,0,0,0,0,0,230,0,58,0,197,0,0,0,252,0,100,0,136,0,209,0,48,0,27,0,109,0,123,0,87,0,140,0,0,0,164,0,112,0,87,0,229,0,64,0,0,0,0,0,67,0,236,0,0,0,56,0,13,0,27,0,210,0,170,0,0,0,99,0,157,0,100,0,0,0,0,0,205,0,96,0,83,0,0,0,225,0,0,0,185,0,160,0,255,0,177,0,179,0,133,0,79,0,230,0,88,0,132,0,103,0,210,0,218,0,186,0,220,0,38,0,97,0,0,0,0,0,116,0,239,0,181,0,226,0,0,0,139,0,33,0,154,0,0,0,230,0,0,0,79,0,0,0,187,0,0,0,42,0,210,0,18,0,158,0,95,0,66,0,179,0,189,0,29,0,210,0,0,0,0,0,179,0,64,0,0,0,156,0,0,0,203,0,5,0,169,0,51,0,17,0,118,0,0,0,73,0,0,0,156,0,100,0,0,0,55,0,21,0,219,0,86,0,201,0,0,0,122,0,88,0,0,0,0,0,142,0,207,0,238,0,0,0,115,0,123,0,0,0,0,0,0,0,100,0,0,0,0,0,0,0,177,0,15,0,215,0,173,0,0,0,0,0,157,0,0,0,0,0,183,0,17,0,0,0,146,0,85,0,123,0,153,0,70,0,24,0,246,0,53,0,227,0,219,0,113,0,164,0,172,0,212,0,155,0,103,0,122,0,23,0,226,0,89,0,250,0,25,0,34,0,216,0,126,0,0,0,225,0,19,0,61,0,32,0,58,0,199,0,56,0,0,0,0,0,144,0,32,0,193,0,213,0,22,0,57,0,0,0,0,0,77,0,225,0,142,0,188,0,85,0,82,0,0,0,198,0,243,0,177,0,0,0,93,0,53,0,112,0,0,0,138,0,0,0,203,0,144,0,0,0,0,0,22,0,153,0,0,0,195,0,0,0,125,0,0,0,183,0,145,0,158,0,115,0,0,0,107,0,124,0,85,0,26,0,27,0,39,0,0,0,202,0,213,0,184,0,141,0,0,0,50,0,231,0,0,0,76,0,0,0,54,0,141,0,0,0,230,0,0,0,52,0,86,0,39,0,117,0,98,0,224,0,119,0,0,0,92,0,0,0,152,0,212,0,198,0,118,0,60,0,124,0,35,0,0,0,104,0,73,0,65,0,121,0,0,0,129,0,71,0,0,0,19,0,0,0,240,0,160,0,0,0,39,0,104,0,0,0,0,0,115,0,171,0,248,0,207,0,0,0,195,0,15,0,75,0,94,0,119,0,0,0,80,0,241,0,0,0,0,0,129,0,27,0,252,0,121,0,51,0,0,0,163,0,70,0,50,0,59,0,197,0,169,0,161,0,172,0,178,0,160,0,79,0,90,0,143,0,248,0,138,0,166,0,247,0,11,0,0,0,166,0,0,0,21,0,38,0,175,0,0,0,75,0,192,0,116,0,146,0,0,0,62,0,0,0,167,0,222,0,238,0,162,0,0,0,193,0,217,0,0,0,0,0,0,0,185,0,34,0,201,0,166,0,123,0,0,0,0,0,67,0,229,0,239,0,0,0,97,0,32,0,221,0,85,0,0,0,103,0,158,0,95,0,202,0,246,0,34,0,100,0,161,0,120,0,128,0,145,0,181,0,54,0,171,0,215,0,0,0,121,0,15,0,158,0,131,0,70,0,46,0,93,0,255,0,0,0,116,0,233,0,4,0,38,0,0,0,235,0,226,0,0,0,0,0,75,0,8,0);
signal scenario_full  : scenario_type := (0,0,118,31,118,30,91,31,196,31,196,30,182,31,182,30,199,31,177,31,181,31,76,31,26,31,48,31,48,30,57,31,224,31,87,31,87,30,4,31,4,30,188,31,230,31,204,31,204,30,143,31,139,31,54,31,235,31,165,31,204,31,197,31,236,31,83,31,128,31,11,31,88,31,154,31,242,31,124,31,124,30,204,31,205,31,205,30,26,31,36,31,86,31,129,31,213,31,213,30,213,29,167,31,69,31,69,30,94,31,32,31,6,31,75,31,85,31,224,31,144,31,136,31,241,31,13,31,43,31,84,31,231,31,158,31,158,30,191,31,171,31,72,31,240,31,233,31,165,31,165,30,125,31,157,31,54,31,102,31,247,31,193,31,193,30,221,31,221,30,205,31,193,31,245,31,142,31,125,31,108,31,215,31,182,31,182,30,216,31,42,31,209,31,186,31,104,31,25,31,103,31,55,31,77,31,233,31,228,31,46,31,115,31,115,30,115,29,115,28,141,31,92,31,134,31,132,31,132,30,40,31,200,31,200,30,20,31,102,31,110,31,129,31,227,31,25,31,25,30,93,31,17,31,209,31,180,31,244,31,110,31,110,30,13,31,28,31,219,31,7,31,210,31,182,31,182,30,191,31,47,31,235,31,235,30,30,31,169,31,169,30,61,31,96,31,171,31,221,31,143,31,110,31,206,31,48,31,48,30,242,31,235,31,117,31,117,30,255,31,68,31,54,31,138,31,197,31,197,30,38,31,155,31,246,31,246,31,237,31,131,31,131,30,131,29,177,31,28,31,4,31,212,31,81,31,71,31,190,31,183,31,183,30,171,31,125,31,64,31,28,31,28,30,28,29,28,28,134,31,159,31,240,31,69,31,212,31,95,31,151,31,236,31,181,31,136,31,170,31,188,31,36,31,159,31,137,31,35,31,44,31,35,31,10,31,203,31,173,31,230,31,241,31,241,30,190,31,83,31,189,31,87,31,138,31,224,31,41,31,208,31,50,31,178,31,178,30,105,31,167,31,88,31,88,30,95,31,95,30,202,31,202,30,44,31,44,30,116,31,115,31,115,30,73,31,73,30,73,29,173,31,202,31,95,31,144,31,144,30,94,31,94,30,254,31,93,31,204,31,65,31,192,31,156,31,156,30,65,31,211,31,30,31,223,31,249,31,235,31,235,30,194,31,96,31,218,31,109,31,222,31,98,31,140,31,183,31,113,31,32,31,169,31,26,31,59,31,105,31,106,31,106,31,77,31,240,31,7,31,7,30,146,31,146,30,206,31,64,31,68,31,15,31,175,31,175,30,58,31,163,31,14,31,14,30,14,29,239,31,18,31,49,31,133,31,74,31,142,31,190,31,190,30,183,31,222,31,113,31,113,30,175,31,228,31,3,31,1,31,102,31,119,31,20,31,20,30,226,31,134,31,95,31,95,30,95,29,30,31,254,31,254,30,147,31,169,31,169,30,130,31,190,31,76,31,57,31,89,31,180,31,180,30,151,31,117,31,42,31,151,31,3,31,34,31,43,31,36,31,116,31,193,31,207,31,237,31,240,31,196,31,221,31,60,31,214,31,58,31,203,31,186,31,188,31,115,31,103,31,223,31,241,31,122,31,150,31,8,31,123,31,198,31,230,31,67,31,242,31,24,31,1,31,159,31,151,31,22,31,29,31,29,30,253,31,86,31,55,31,154,31,81,31,80,31,37,31,37,30,37,29,111,31,203,31,121,31,253,31,228,31,151,31,151,30,33,31,223,31,126,31,189,31,203,31,56,31,242,31,202,31,250,31,250,30,253,31,76,31,192,31,55,31,64,31,228,31,228,30,166,31,31,31,255,31,255,30,69,31,241,31,103,31,69,31,69,30,69,29,24,31,24,30,245,31,245,30,147,31,76,31,76,30,178,31,96,31,96,30,18,31,50,31,50,30,160,31,131,31,131,30,172,31,172,30,172,29,172,28,172,27,139,31,247,31,105,31,250,31,223,31,253,31,242,31,132,31,132,30,39,31,141,31,141,30,249,31,46,31,88,31,192,31,147,31,93,31,143,31,50,31,50,30,106,31,149,31,149,30,149,29,239,31,214,31,47,31,224,31,224,30,224,29,32,31,221,31,125,31,34,31,34,30,206,31,198,31,184,31,114,31,114,30,4,31,4,30,246,31,88,31,198,31,19,31,23,31,254,31,228,31,102,31,102,30,70,31,70,30,70,29,70,28,193,31,193,30,159,31,220,31,29,31,29,30,63,31,152,31,152,30,167,31,204,31,204,30,111,31,37,31,37,30,210,31,210,30,210,29,242,31,149,31,157,31,157,30,148,31,3,31,147,31,145,31,204,31,219,31,219,30,219,29,219,28,230,31,58,31,197,31,197,30,252,31,100,31,136,31,209,31,48,31,27,31,109,31,123,31,87,31,140,31,140,30,164,31,112,31,87,31,229,31,64,31,64,30,64,29,67,31,236,31,236,30,56,31,13,31,27,31,210,31,170,31,170,30,99,31,157,31,100,31,100,30,100,29,205,31,96,31,83,31,83,30,225,31,225,30,185,31,160,31,255,31,177,31,179,31,133,31,79,31,230,31,88,31,132,31,103,31,210,31,218,31,186,31,220,31,38,31,97,31,97,30,97,29,116,31,239,31,181,31,226,31,226,30,139,31,33,31,154,31,154,30,230,31,230,30,79,31,79,30,187,31,187,30,42,31,210,31,18,31,158,31,95,31,66,31,179,31,189,31,29,31,210,31,210,30,210,29,179,31,64,31,64,30,156,31,156,30,203,31,5,31,169,31,51,31,17,31,118,31,118,30,73,31,73,30,156,31,100,31,100,30,55,31,21,31,219,31,86,31,201,31,201,30,122,31,88,31,88,30,88,29,142,31,207,31,238,31,238,30,115,31,123,31,123,30,123,29,123,28,100,31,100,30,100,29,100,28,177,31,15,31,215,31,173,31,173,30,173,29,157,31,157,30,157,29,183,31,17,31,17,30,146,31,85,31,123,31,153,31,70,31,24,31,246,31,53,31,227,31,219,31,113,31,164,31,172,31,212,31,155,31,103,31,122,31,23,31,226,31,89,31,250,31,25,31,34,31,216,31,126,31,126,30,225,31,19,31,61,31,32,31,58,31,199,31,56,31,56,30,56,29,144,31,32,31,193,31,213,31,22,31,57,31,57,30,57,29,77,31,225,31,142,31,188,31,85,31,82,31,82,30,198,31,243,31,177,31,177,30,93,31,53,31,112,31,112,30,138,31,138,30,203,31,144,31,144,30,144,29,22,31,153,31,153,30,195,31,195,30,125,31,125,30,183,31,145,31,158,31,115,31,115,30,107,31,124,31,85,31,26,31,27,31,39,31,39,30,202,31,213,31,184,31,141,31,141,30,50,31,231,31,231,30,76,31,76,30,54,31,141,31,141,30,230,31,230,30,52,31,86,31,39,31,117,31,98,31,224,31,119,31,119,30,92,31,92,30,152,31,212,31,198,31,118,31,60,31,124,31,35,31,35,30,104,31,73,31,65,31,121,31,121,30,129,31,71,31,71,30,19,31,19,30,240,31,160,31,160,30,39,31,104,31,104,30,104,29,115,31,171,31,248,31,207,31,207,30,195,31,15,31,75,31,94,31,119,31,119,30,80,31,241,31,241,30,241,29,129,31,27,31,252,31,121,31,51,31,51,30,163,31,70,31,50,31,59,31,197,31,169,31,161,31,172,31,178,31,160,31,79,31,90,31,143,31,248,31,138,31,166,31,247,31,11,31,11,30,166,31,166,30,21,31,38,31,175,31,175,30,75,31,192,31,116,31,146,31,146,30,62,31,62,30,167,31,222,31,238,31,162,31,162,30,193,31,217,31,217,30,217,29,217,28,185,31,34,31,201,31,166,31,123,31,123,30,123,29,67,31,229,31,239,31,239,30,97,31,32,31,221,31,85,31,85,30,103,31,158,31,95,31,202,31,246,31,34,31,100,31,161,31,120,31,128,31,145,31,181,31,54,31,171,31,215,31,215,30,121,31,15,31,158,31,131,31,70,31,46,31,93,31,255,31,255,30,116,31,233,31,4,31,38,31,38,30,235,31,226,31,226,30,226,29,75,31,8,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
