-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_744 is
end project_tb_744;

architecture project_tb_arch_744 of project_tb_744 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 294;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,154,0,144,0,9,0,0,0,84,0,0,0,226,0,231,0,51,0,88,0,0,0,102,0,239,0,64,0,232,0,0,0,236,0,248,0,226,0,0,0,194,0,149,0,237,0,34,0,190,0,0,0,245,0,142,0,0,0,135,0,129,0,248,0,74,0,165,0,255,0,0,0,182,0,172,0,224,0,69,0,0,0,39,0,115,0,163,0,243,0,121,0,103,0,142,0,237,0,89,0,122,0,205,0,208,0,183,0,208,0,234,0,164,0,250,0,76,0,40,0,99,0,225,0,15,0,0,0,0,0,224,0,4,0,0,0,85,0,0,0,126,0,0,0,219,0,0,0,81,0,140,0,166,0,228,0,97,0,17,0,114,0,169,0,188,0,118,0,201,0,1,0,196,0,198,0,107,0,49,0,248,0,4,0,6,0,0,0,192,0,171,0,40,0,124,0,164,0,0,0,19,0,79,0,134,0,0,0,147,0,75,0,142,0,120,0,160,0,155,0,199,0,165,0,90,0,172,0,70,0,208,0,246,0,170,0,174,0,165,0,144,0,197,0,0,0,0,0,0,0,162,0,88,0,240,0,0,0,54,0,0,0,142,0,136,0,146,0,37,0,0,0,109,0,23,0,71,0,0,0,0,0,240,0,0,0,170,0,47,0,0,0,63,0,0,0,185,0,24,0,190,0,0,0,0,0,82,0,238,0,16,0,149,0,18,0,28,0,247,0,18,0,121,0,14,0,0,0,0,0,0,0,133,0,250,0,105,0,210,0,157,0,0,0,29,0,105,0,0,0,0,0,108,0,97,0,142,0,0,0,0,0,89,0,212,0,216,0,17,0,197,0,148,0,115,0,104,0,109,0,187,0,224,0,0,0,40,0,210,0,108,0,157,0,210,0,0,0,49,0,168,0,57,0,7,0,0,0,215,0,98,0,205,0,132,0,56,0,0,0,36,0,202,0,0,0,5,0,223,0,185,0,168,0,0,0,0,0,195,0,0,0,154,0,155,0,78,0,45,0,0,0,165,0,28,0,0,0,0,0,0,0,92,0,0,0,34,0,57,0,0,0,198,0,182,0,4,0,13,0,30,0,234,0,0,0,15,0,141,0,156,0,143,0,181,0,203,0,73,0,26,0,215,0,0,0,234,0,134,0,128,0,148,0,0,0,175,0,0,0,141,0,137,0,0,0,113,0,129,0,242,0,0,0,37,0,73,0,0,0,239,0,222,0,11,0,132,0,0,0,88,0,115,0,223,0,0,0,88,0,85,0,252,0,219,0,0,0,150,0,239,0,0,0,9,0,0,0,40,0,117,0,149,0,34,0);
signal scenario_full  : scenario_type := (0,0,154,31,144,31,9,31,9,30,84,31,84,30,226,31,231,31,51,31,88,31,88,30,102,31,239,31,64,31,232,31,232,30,236,31,248,31,226,31,226,30,194,31,149,31,237,31,34,31,190,31,190,30,245,31,142,31,142,30,135,31,129,31,248,31,74,31,165,31,255,31,255,30,182,31,172,31,224,31,69,31,69,30,39,31,115,31,163,31,243,31,121,31,103,31,142,31,237,31,89,31,122,31,205,31,208,31,183,31,208,31,234,31,164,31,250,31,76,31,40,31,99,31,225,31,15,31,15,30,15,29,224,31,4,31,4,30,85,31,85,30,126,31,126,30,219,31,219,30,81,31,140,31,166,31,228,31,97,31,17,31,114,31,169,31,188,31,118,31,201,31,1,31,196,31,198,31,107,31,49,31,248,31,4,31,6,31,6,30,192,31,171,31,40,31,124,31,164,31,164,30,19,31,79,31,134,31,134,30,147,31,75,31,142,31,120,31,160,31,155,31,199,31,165,31,90,31,172,31,70,31,208,31,246,31,170,31,174,31,165,31,144,31,197,31,197,30,197,29,197,28,162,31,88,31,240,31,240,30,54,31,54,30,142,31,136,31,146,31,37,31,37,30,109,31,23,31,71,31,71,30,71,29,240,31,240,30,170,31,47,31,47,30,63,31,63,30,185,31,24,31,190,31,190,30,190,29,82,31,238,31,16,31,149,31,18,31,28,31,247,31,18,31,121,31,14,31,14,30,14,29,14,28,133,31,250,31,105,31,210,31,157,31,157,30,29,31,105,31,105,30,105,29,108,31,97,31,142,31,142,30,142,29,89,31,212,31,216,31,17,31,197,31,148,31,115,31,104,31,109,31,187,31,224,31,224,30,40,31,210,31,108,31,157,31,210,31,210,30,49,31,168,31,57,31,7,31,7,30,215,31,98,31,205,31,132,31,56,31,56,30,36,31,202,31,202,30,5,31,223,31,185,31,168,31,168,30,168,29,195,31,195,30,154,31,155,31,78,31,45,31,45,30,165,31,28,31,28,30,28,29,28,28,92,31,92,30,34,31,57,31,57,30,198,31,182,31,4,31,13,31,30,31,234,31,234,30,15,31,141,31,156,31,143,31,181,31,203,31,73,31,26,31,215,31,215,30,234,31,134,31,128,31,148,31,148,30,175,31,175,30,141,31,137,31,137,30,113,31,129,31,242,31,242,30,37,31,73,31,73,30,239,31,222,31,11,31,132,31,132,30,88,31,115,31,223,31,223,30,88,31,85,31,252,31,219,31,219,30,150,31,239,31,239,30,9,31,9,30,40,31,117,31,149,31,34,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
