-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 295;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,9,0,0,0,12,0,0,0,86,0,165,0,30,0,0,0,54,0,0,0,32,0,131,0,200,0,11,0,237,0,133,0,60,0,219,0,207,0,14,0,0,0,0,0,0,0,243,0,247,0,216,0,204,0,106,0,247,0,0,0,152,0,127,0,116,0,105,0,0,0,145,0,94,0,96,0,88,0,181,0,82,0,0,0,0,0,0,0,76,0,89,0,58,0,16,0,76,0,131,0,117,0,236,0,14,0,0,0,109,0,0,0,36,0,68,0,6,0,83,0,2,0,249,0,104,0,0,0,183,0,0,0,0,0,199,0,0,0,138,0,137,0,142,0,0,0,151,0,147,0,0,0,159,0,191,0,0,0,0,0,179,0,3,0,92,0,0,0,209,0,53,0,255,0,0,0,102,0,153,0,53,0,92,0,6,0,0,0,0,0,214,0,0,0,30,0,78,0,24,0,100,0,101,0,144,0,216,0,53,0,12,0,211,0,0,0,35,0,49,0,139,0,133,0,77,0,16,0,41,0,51,0,115,0,149,0,188,0,160,0,220,0,198,0,0,0,214,0,159,0,210,0,144,0,142,0,80,0,0,0,245,0,217,0,188,0,148,0,173,0,135,0,237,0,3,0,0,0,158,0,104,0,235,0,89,0,0,0,197,0,118,0,59,0,148,0,0,0,141,0,0,0,177,0,98,0,0,0,45,0,235,0,120,0,144,0,30,0,0,0,76,0,0,0,217,0,237,0,0,0,143,0,199,0,0,0,211,0,168,0,97,0,198,0,127,0,0,0,0,0,199,0,244,0,211,0,181,0,197,0,214,0,239,0,63,0,89,0,99,0,247,0,0,0,165,0,73,0,235,0,58,0,115,0,66,0,59,0,102,0,0,0,36,0,0,0,0,0,171,0,112,0,0,0,92,0,66,0,156,0,101,0,184,0,116,0,202,0,75,0,176,0,184,0,143,0,87,0,0,0,216,0,0,0,123,0,0,0,163,0,11,0,71,0,253,0,138,0,231,0,20,0,0,0,0,0,0,0,220,0,146,0,0,0,249,0,140,0,9,0,116,0,9,0,201,0,0,0,152,0,136,0,225,0,67,0,135,0,162,0,0,0,95,0,124,0,11,0,131,0,203,0,118,0,165,0,0,0,0,0,0,0,167,0,0,0,234,0,142,0,98,0,228,0,148,0,8,0,8,0,0,0,0,0,26,0,0,0,0,0,40,0,82,0,0,0,0,0,251,0,220,0,29,0,13,0,89,0,248,0,75,0,0,0,193,0,13,0,0,0,31,0,43,0,158,0,38,0,0,0,134,0,172,0,0,0,72,0);
signal scenario_full  : scenario_type := (0,0,9,31,9,30,12,31,12,30,86,31,165,31,30,31,30,30,54,31,54,30,32,31,131,31,200,31,11,31,237,31,133,31,60,31,219,31,207,31,14,31,14,30,14,29,14,28,243,31,247,31,216,31,204,31,106,31,247,31,247,30,152,31,127,31,116,31,105,31,105,30,145,31,94,31,96,31,88,31,181,31,82,31,82,30,82,29,82,28,76,31,89,31,58,31,16,31,76,31,131,31,117,31,236,31,14,31,14,30,109,31,109,30,36,31,68,31,6,31,83,31,2,31,249,31,104,31,104,30,183,31,183,30,183,29,199,31,199,30,138,31,137,31,142,31,142,30,151,31,147,31,147,30,159,31,191,31,191,30,191,29,179,31,3,31,92,31,92,30,209,31,53,31,255,31,255,30,102,31,153,31,53,31,92,31,6,31,6,30,6,29,214,31,214,30,30,31,78,31,24,31,100,31,101,31,144,31,216,31,53,31,12,31,211,31,211,30,35,31,49,31,139,31,133,31,77,31,16,31,41,31,51,31,115,31,149,31,188,31,160,31,220,31,198,31,198,30,214,31,159,31,210,31,144,31,142,31,80,31,80,30,245,31,217,31,188,31,148,31,173,31,135,31,237,31,3,31,3,30,158,31,104,31,235,31,89,31,89,30,197,31,118,31,59,31,148,31,148,30,141,31,141,30,177,31,98,31,98,30,45,31,235,31,120,31,144,31,30,31,30,30,76,31,76,30,217,31,237,31,237,30,143,31,199,31,199,30,211,31,168,31,97,31,198,31,127,31,127,30,127,29,199,31,244,31,211,31,181,31,197,31,214,31,239,31,63,31,89,31,99,31,247,31,247,30,165,31,73,31,235,31,58,31,115,31,66,31,59,31,102,31,102,30,36,31,36,30,36,29,171,31,112,31,112,30,92,31,66,31,156,31,101,31,184,31,116,31,202,31,75,31,176,31,184,31,143,31,87,31,87,30,216,31,216,30,123,31,123,30,163,31,11,31,71,31,253,31,138,31,231,31,20,31,20,30,20,29,20,28,220,31,146,31,146,30,249,31,140,31,9,31,116,31,9,31,201,31,201,30,152,31,136,31,225,31,67,31,135,31,162,31,162,30,95,31,124,31,11,31,131,31,203,31,118,31,165,31,165,30,165,29,165,28,167,31,167,30,234,31,142,31,98,31,228,31,148,31,8,31,8,31,8,30,8,29,26,31,26,30,26,29,40,31,82,31,82,30,82,29,251,31,220,31,29,31,13,31,89,31,248,31,75,31,75,30,193,31,13,31,13,30,31,31,43,31,158,31,38,31,38,30,134,31,172,31,172,30,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
