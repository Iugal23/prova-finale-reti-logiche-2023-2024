-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_807 is
end project_tb_807;

architecture project_tb_arch_807 of project_tb_807 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 531;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (116,0,18,0,5,0,150,0,245,0,0,0,0,0,155,0,219,0,0,0,247,0,29,0,190,0,0,0,0,0,0,0,144,0,0,0,123,0,54,0,201,0,128,0,0,0,99,0,0,0,194,0,0,0,210,0,0,0,0,0,193,0,0,0,105,0,34,0,0,0,48,0,101,0,183,0,89,0,204,0,133,0,0,0,136,0,66,0,46,0,0,0,0,0,52,0,67,0,33,0,26,0,250,0,176,0,56,0,93,0,239,0,188,0,0,0,0,0,59,0,0,0,229,0,0,0,5,0,0,0,212,0,77,0,73,0,233,0,166,0,93,0,206,0,52,0,0,0,46,0,218,0,211,0,0,0,12,0,72,0,0,0,225,0,39,0,37,0,0,0,82,0,145,0,0,0,68,0,62,0,11,0,229,0,0,0,175,0,122,0,209,0,46,0,90,0,180,0,0,0,252,0,4,0,153,0,7,0,66,0,106,0,29,0,2,0,0,0,9,0,0,0,49,0,0,0,155,0,0,0,141,0,44,0,25,0,0,0,73,0,74,0,82,0,0,0,79,0,67,0,152,0,245,0,178,0,84,0,222,0,88,0,196,0,3,0,196,0,0,0,211,0,136,0,191,0,108,0,49,0,34,0,39,0,233,0,120,0,28,0,231,0,107,0,143,0,0,0,0,0,255,0,115,0,73,0,59,0,129,0,197,0,35,0,160,0,150,0,234,0,234,0,71,0,0,0,174,0,175,0,171,0,115,0,0,0,152,0,222,0,179,0,140,0,114,0,109,0,14,0,132,0,0,0,0,0,138,0,0,0,144,0,88,0,138,0,176,0,0,0,160,0,208,0,137,0,0,0,37,0,65,0,0,0,0,0,118,0,167,0,81,0,60,0,255,0,0,0,107,0,245,0,11,0,86,0,10,0,186,0,0,0,152,0,0,0,77,0,105,0,134,0,223,0,0,0,240,0,56,0,0,0,137,0,193,0,63,0,77,0,0,0,242,0,1,0,140,0,52,0,179,0,161,0,68,0,165,0,0,0,0,0,247,0,0,0,231,0,78,0,186,0,61,0,106,0,78,0,144,0,81,0,13,0,203,0,157,0,95,0,95,0,0,0,132,0,182,0,159,0,246,0,0,0,218,0,0,0,85,0,169,0,0,0,185,0,59,0,120,0,212,0,248,0,5,0,0,0,0,0,7,0,205,0,0,0,33,0,70,0,0,0,200,0,230,0,0,0,42,0,0,0,34,0,0,0,0,0,0,0,0,0,0,0,4,0,63,0,196,0,228,0,181,0,0,0,201,0,192,0,145,0,160,0,162,0,48,0,0,0,183,0,204,0,79,0,244,0,0,0,151,0,37,0,108,0,61,0,0,0,24,0,58,0,204,0,172,0,0,0,122,0,208,0,164,0,0,0,96,0,33,0,116,0,209,0,1,0,159,0,86,0,245,0,9,0,70,0,128,0,116,0,150,0,13,0,0,0,189,0,20,0,56,0,0,0,83,0,0,0,0,0,139,0,189,0,203,0,204,0,234,0,128,0,0,0,104,0,155,0,44,0,0,0,0,0,100,0,215,0,141,0,66,0,228,0,201,0,148,0,0,0,134,0,181,0,165,0,235,0,113,0,52,0,0,0,231,0,76,0,16,0,0,0,201,0,59,0,0,0,210,0,31,0,47,0,106,0,211,0,191,0,0,0,0,0,78,0,98,0,76,0,114,0,39,0,112,0,253,0,0,0,178,0,0,0,64,0,191,0,91,0,35,0,67,0,0,0,144,0,0,0,52,0,138,0,154,0,0,0,240,0,231,0,181,0,133,0,71,0,32,0,135,0,44,0,179,0,0,0,51,0,231,0,0,0,198,0,227,0,121,0,128,0,142,0,0,0,94,0,0,0,6,0,176,0,213,0,0,0,180,0,156,0,183,0,161,0,254,0,134,0,35,0,6,0,175,0,0,0,102,0,86,0,8,0,0,0,0,0,105,0,219,0,217,0,176,0,60,0,45,0,74,0,158,0,241,0,0,0,110,0,207,0,174,0,224,0,0,0,211,0,0,0,151,0,125,0,105,0,158,0,228,0,210,0,217,0,0,0,1,0,226,0,32,0,251,0,37,0,227,0,150,0,161,0,172,0,199,0,56,0,0,0,69,0,73,0,53,0,202,0,157,0,0,0,90,0,193,0,40,0,7,0,50,0,103,0,90,0,0,0,12,0,229,0,212,0,123,0,0,0,0,0,0,0,23,0,211,0,123,0,92,0,99,0,61,0,183,0,84,0,248,0,219,0,135,0,74,0,148,0,228,0,22,0,55,0,36,0,186,0,42,0,236,0,251,0,151,0,214,0,246,0,0,0,116,0,151,0,227,0,63,0,34,0,45,0,61,0,254,0);
signal scenario_full  : scenario_type := (116,31,18,31,5,31,150,31,245,31,245,30,245,29,155,31,219,31,219,30,247,31,29,31,190,31,190,30,190,29,190,28,144,31,144,30,123,31,54,31,201,31,128,31,128,30,99,31,99,30,194,31,194,30,210,31,210,30,210,29,193,31,193,30,105,31,34,31,34,30,48,31,101,31,183,31,89,31,204,31,133,31,133,30,136,31,66,31,46,31,46,30,46,29,52,31,67,31,33,31,26,31,250,31,176,31,56,31,93,31,239,31,188,31,188,30,188,29,59,31,59,30,229,31,229,30,5,31,5,30,212,31,77,31,73,31,233,31,166,31,93,31,206,31,52,31,52,30,46,31,218,31,211,31,211,30,12,31,72,31,72,30,225,31,39,31,37,31,37,30,82,31,145,31,145,30,68,31,62,31,11,31,229,31,229,30,175,31,122,31,209,31,46,31,90,31,180,31,180,30,252,31,4,31,153,31,7,31,66,31,106,31,29,31,2,31,2,30,9,31,9,30,49,31,49,30,155,31,155,30,141,31,44,31,25,31,25,30,73,31,74,31,82,31,82,30,79,31,67,31,152,31,245,31,178,31,84,31,222,31,88,31,196,31,3,31,196,31,196,30,211,31,136,31,191,31,108,31,49,31,34,31,39,31,233,31,120,31,28,31,231,31,107,31,143,31,143,30,143,29,255,31,115,31,73,31,59,31,129,31,197,31,35,31,160,31,150,31,234,31,234,31,71,31,71,30,174,31,175,31,171,31,115,31,115,30,152,31,222,31,179,31,140,31,114,31,109,31,14,31,132,31,132,30,132,29,138,31,138,30,144,31,88,31,138,31,176,31,176,30,160,31,208,31,137,31,137,30,37,31,65,31,65,30,65,29,118,31,167,31,81,31,60,31,255,31,255,30,107,31,245,31,11,31,86,31,10,31,186,31,186,30,152,31,152,30,77,31,105,31,134,31,223,31,223,30,240,31,56,31,56,30,137,31,193,31,63,31,77,31,77,30,242,31,1,31,140,31,52,31,179,31,161,31,68,31,165,31,165,30,165,29,247,31,247,30,231,31,78,31,186,31,61,31,106,31,78,31,144,31,81,31,13,31,203,31,157,31,95,31,95,31,95,30,132,31,182,31,159,31,246,31,246,30,218,31,218,30,85,31,169,31,169,30,185,31,59,31,120,31,212,31,248,31,5,31,5,30,5,29,7,31,205,31,205,30,33,31,70,31,70,30,200,31,230,31,230,30,42,31,42,30,34,31,34,30,34,29,34,28,34,27,34,26,4,31,63,31,196,31,228,31,181,31,181,30,201,31,192,31,145,31,160,31,162,31,48,31,48,30,183,31,204,31,79,31,244,31,244,30,151,31,37,31,108,31,61,31,61,30,24,31,58,31,204,31,172,31,172,30,122,31,208,31,164,31,164,30,96,31,33,31,116,31,209,31,1,31,159,31,86,31,245,31,9,31,70,31,128,31,116,31,150,31,13,31,13,30,189,31,20,31,56,31,56,30,83,31,83,30,83,29,139,31,189,31,203,31,204,31,234,31,128,31,128,30,104,31,155,31,44,31,44,30,44,29,100,31,215,31,141,31,66,31,228,31,201,31,148,31,148,30,134,31,181,31,165,31,235,31,113,31,52,31,52,30,231,31,76,31,16,31,16,30,201,31,59,31,59,30,210,31,31,31,47,31,106,31,211,31,191,31,191,30,191,29,78,31,98,31,76,31,114,31,39,31,112,31,253,31,253,30,178,31,178,30,64,31,191,31,91,31,35,31,67,31,67,30,144,31,144,30,52,31,138,31,154,31,154,30,240,31,231,31,181,31,133,31,71,31,32,31,135,31,44,31,179,31,179,30,51,31,231,31,231,30,198,31,227,31,121,31,128,31,142,31,142,30,94,31,94,30,6,31,176,31,213,31,213,30,180,31,156,31,183,31,161,31,254,31,134,31,35,31,6,31,175,31,175,30,102,31,86,31,8,31,8,30,8,29,105,31,219,31,217,31,176,31,60,31,45,31,74,31,158,31,241,31,241,30,110,31,207,31,174,31,224,31,224,30,211,31,211,30,151,31,125,31,105,31,158,31,228,31,210,31,217,31,217,30,1,31,226,31,32,31,251,31,37,31,227,31,150,31,161,31,172,31,199,31,56,31,56,30,69,31,73,31,53,31,202,31,157,31,157,30,90,31,193,31,40,31,7,31,50,31,103,31,90,31,90,30,12,31,229,31,212,31,123,31,123,30,123,29,123,28,23,31,211,31,123,31,92,31,99,31,61,31,183,31,84,31,248,31,219,31,135,31,74,31,148,31,228,31,22,31,55,31,36,31,186,31,42,31,236,31,251,31,151,31,214,31,246,31,246,30,116,31,151,31,227,31,63,31,34,31,45,31,61,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
