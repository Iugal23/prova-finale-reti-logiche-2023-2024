-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (103,0,238,0,22,0,218,0,227,0,59,0,78,0,89,0,178,0,9,0,231,0,172,0,124,0,186,0,244,0,20,0,0,0,65,0,178,0,209,0,55,0,202,0,194,0,70,0,18,0,0,0,95,0,0,0,72,0,254,0,1,0,0,0,19,0,0,0,68,0,15,0,220,0,0,0,5,0,75,0,18,0,154,0,54,0,153,0,4,0,75,0,119,0,110,0,185,0,117,0,10,0,12,0,14,0,197,0,6,0,195,0,188,0,114,0,77,0,242,0,138,0,176,0,7,0,207,0,158,0,63,0,124,0,217,0,158,0,113,0,52,0,0,0,0,0,21,0,127,0,3,0,74,0,217,0,1,0,41,0,242,0,79,0,166,0,54,0,0,0,0,0,0,0,189,0,0,0,0,0,102,0,195,0,174,0,3,0,16,0,192,0,0,0,0,0,170,0,130,0,100,0,11,0,120,0,207,0,234,0,112,0,232,0,103,0,193,0,170,0,98,0,28,0,0,0,0,0,240,0,144,0,17,0,0,0,0,0,0,0,166,0,0,0,0,0,0,0,45,0,36,0,251,0,151,0,0,0,0,0,190,0,197,0,137,0,224,0,124,0,200,0,68,0,155,0,91,0,255,0,221,0,10,0,0,0,62,0,88,0,0,0,191,0,137,0,234,0,52,0,61,0,176,0,0,0,189,0,235,0,248,0,59,0,241,0,166,0,167,0,233,0,0,0,223,0,197,0,50,0,174,0,109,0,0,0,174,0,23,0,207,0,142,0,206,0,79,0,168,0,0,0,136,0,0,0,0,0,219,0,0,0,140,0,15,0,183,0,255,0,26,0,0,0,0,0,23,0,184,0,211,0,0,0,186,0,0,0,100,0,131,0,189,0,181,0,57,0,112,0,135,0,0,0,0,0,208,0,82,0,0,0,70,0,213,0,220,0,215,0,230,0,0,0,0,0,0,0,84,0,0,0,131,0,0,0,135,0,0,0,146,0,209,0,0,0,193,0,207,0,245,0,217,0,73,0,48,0,204,0,251,0,136,0,0,0,58,0,0,0,192,0,210,0,28,0,0,0,34,0,26,0,127,0,122,0,2,0,163,0,197,0,0,0,0,0,188,0,169,0,19,0,53,0,0,0,137,0,35,0,48,0,232,0,23,0,9,0,0,0,187,0,0,0,247,0,147,0,0,0,66,0,211,0,234,0,9,0,135,0,73,0,0,0,244,0,106,0,75,0,231,0,100,0,134,0,84,0,101,0,98,0,0,0,184,0,54,0,149,0,0,0,191,0,169,0,10,0,0,0,181,0,0,0,201,0,192,0,116,0,189,0,41,0,0,0,93,0,130,0,97,0,113,0,0,0,68,0,59,0,15,0,19,0,32,0,0,0,122,0,14,0,242,0,146,0,0,0,45,0,4,0,228,0,190,0,0,0,133,0,0,0,19,0,13,0,19,0,222,0,89,0,11,0,116,0,61,0,212,0,0,0,0,0,242,0,196,0,0,0,244,0,0,0,0,0,55,0,153,0,120,0,17,0,94,0,253,0,76,0,251,0,0,0,0,0,0,0,65,0,174,0,245,0,237,0,50,0,0,0,207,0,196,0,231,0,209,0,50,0,170,0,2,0,0,0,175,0,206,0,0,0,234,0,234,0,135,0,58,0,0,0,0,0,205,0,162,0,0,0,0,0,92,0,0,0,0,0,129,0,2,0,0,0,88,0,31,0,167,0,0,0,0,0,221,0,125,0,0,0,130,0,134,0,152,0,250,0,16,0,232,0,0,0,0,0,163,0,0,0,220,0,29,0,83,0,0,0,155,0,138,0,157,0,151,0,0,0,0,0,45,0,205,0,28,0,9,0,70,0,220,0,0,0,27,0,213,0,106,0,0,0,81,0,112,0,15,0,209,0,0,0,160,0,14,0,20,0,157,0,191,0,0,0,248,0,173,0,200,0,50,0,231,0,238,0,188,0,20,0,235,0,0,0,239,0,16,0,252,0,0,0,0,0,161,0,21,0,135,0,113,0,0,0,188,0,245,0,42,0,0,0,58,0,151,0,128,0,218,0,144,0,253,0,25,0,186,0,181,0,164,0,121,0,78,0,201,0,75,0,231,0,111,0,250,0,178,0,62,0,0,0,0,0,30,0,202,0,178,0,61,0,33,0,0,0,135,0,0,0,199,0,54,0,237,0,42,0,11,0,12,0,205,0,67,0,135,0,103,0,0,0,126,0,219,0,123,0,79,0,0,0,0,0,217,0,227,0,4,0,113,0,22,0,46,0,0,0,46,0,0,0,166,0,204,0,115,0,29,0,0,0,244,0,252,0,192,0,0,0,222,0,165,0,71,0,189,0,0,0,174,0,194,0,190,0,94,0,197,0,238,0,95,0,125,0,189,0,255,0,0,0,45,0,90,0,254,0,0,0,69,0,84,0,136,0,60,0,121,0,161,0,66,0,189,0,101,0,211,0,0,0,247,0,230,0,0,0,17,0,1,0,53,0,185,0,90,0,14,0,150,0,177,0,48,0,196,0,69,0,220,0,77,0,10,0,0,0,96,0,157,0,0,0,69,0,147,0,207,0,0,0,0,0,159,0,174,0,0,0,53,0,81,0,151,0,11,0,235,0,198,0,254,0,79,0,255,0,194,0,60,0,0,0,69,0,253,0,69,0,14,0,28,0,14,0,36,0,73,0,0,0,0,0,223,0,144,0,125,0,0,0,0,0,113,0,0,0,233,0,44,0,156,0,1,0,184,0,2,0,204,0,40,0,230,0,0,0,117,0,241,0,0,0,0,0,207,0,124,0,59,0,132,0,138,0,127,0,0,0,0,0,253,0,214,0,47,0,14,0,136,0,88,0,147,0,248,0,143,0,221,0,0,0,158,0,148,0,0,0,138,0,79,0,10,0,190,0,242,0,106,0,63,0,12,0,154,0,38,0,111,0,63,0,49,0,0,0,58,0,225,0,241,0,8,0,94,0,0,0,0,0,124,0,244,0,173,0,0,0,22,0,251,0,215,0,86,0,140,0,54,0,170,0,137,0,3,0,0,0,46,0,0,0,205,0,84,0,0,0,180,0,78,0,30,0,68,0,135,0,33,0,0,0,76,0,233,0,26,0,58,0,67,0,0,0,225,0,55,0,79,0,3,0,58,0,218,0,143,0,242,0,178,0,0,0,84,0,57,0,213,0,181,0,53,0,0,0,183,0,80,0,125,0,106,0,113,0,76,0,0,0,124,0,231,0,237,0,180,0,136,0,68,0,0,0,107,0,108,0,63,0,123,0,31,0,13,0,131,0,210,0,53,0,230,0,113,0,23,0,0,0,245,0,18,0,155,0,0,0,232,0,66,0,0,0,0,0,45,0,79,0,33,0,254,0,239,0,0,0,0,0,60,0,37,0,88,0,29,0,251,0,151,0,214,0,170,0,209,0,22,0,154,0,121,0,0,0,177,0,93,0,0,0,119,0,240,0,162,0,109,0,65,0,20,0,189,0,0,0,0,0,55,0,229,0,0,0,36,0,44,0,0,0,24,0,126,0,115,0,198,0,36,0,151,0,61,0,64,0,0,0,150,0,0,0,0,0,128,0,4,0,6,0,0,0,200,0,97,0,6,0,247,0,146,0,80,0,197,0,196,0,0,0,174,0,195,0,234,0,20,0,175,0,35,0,245,0,164,0,48,0,37,0,172,0,0,0,207,0,248,0,16,0,195,0,0,0,0,0,0,0,113,0,225,0,0,0,0,0,0,0,190,0,192,0,113,0,0,0,0,0,45,0,234,0,5,0,0,0,237,0,111,0,217,0,0,0,87,0,57,0,174,0,0,0,0,0,217,0,147,0,224,0);
signal scenario_full  : scenario_type := (103,31,238,31,22,31,218,31,227,31,59,31,78,31,89,31,178,31,9,31,231,31,172,31,124,31,186,31,244,31,20,31,20,30,65,31,178,31,209,31,55,31,202,31,194,31,70,31,18,31,18,30,95,31,95,30,72,31,254,31,1,31,1,30,19,31,19,30,68,31,15,31,220,31,220,30,5,31,75,31,18,31,154,31,54,31,153,31,4,31,75,31,119,31,110,31,185,31,117,31,10,31,12,31,14,31,197,31,6,31,195,31,188,31,114,31,77,31,242,31,138,31,176,31,7,31,207,31,158,31,63,31,124,31,217,31,158,31,113,31,52,31,52,30,52,29,21,31,127,31,3,31,74,31,217,31,1,31,41,31,242,31,79,31,166,31,54,31,54,30,54,29,54,28,189,31,189,30,189,29,102,31,195,31,174,31,3,31,16,31,192,31,192,30,192,29,170,31,130,31,100,31,11,31,120,31,207,31,234,31,112,31,232,31,103,31,193,31,170,31,98,31,28,31,28,30,28,29,240,31,144,31,17,31,17,30,17,29,17,28,166,31,166,30,166,29,166,28,45,31,36,31,251,31,151,31,151,30,151,29,190,31,197,31,137,31,224,31,124,31,200,31,68,31,155,31,91,31,255,31,221,31,10,31,10,30,62,31,88,31,88,30,191,31,137,31,234,31,52,31,61,31,176,31,176,30,189,31,235,31,248,31,59,31,241,31,166,31,167,31,233,31,233,30,223,31,197,31,50,31,174,31,109,31,109,30,174,31,23,31,207,31,142,31,206,31,79,31,168,31,168,30,136,31,136,30,136,29,219,31,219,30,140,31,15,31,183,31,255,31,26,31,26,30,26,29,23,31,184,31,211,31,211,30,186,31,186,30,100,31,131,31,189,31,181,31,57,31,112,31,135,31,135,30,135,29,208,31,82,31,82,30,70,31,213,31,220,31,215,31,230,31,230,30,230,29,230,28,84,31,84,30,131,31,131,30,135,31,135,30,146,31,209,31,209,30,193,31,207,31,245,31,217,31,73,31,48,31,204,31,251,31,136,31,136,30,58,31,58,30,192,31,210,31,28,31,28,30,34,31,26,31,127,31,122,31,2,31,163,31,197,31,197,30,197,29,188,31,169,31,19,31,53,31,53,30,137,31,35,31,48,31,232,31,23,31,9,31,9,30,187,31,187,30,247,31,147,31,147,30,66,31,211,31,234,31,9,31,135,31,73,31,73,30,244,31,106,31,75,31,231,31,100,31,134,31,84,31,101,31,98,31,98,30,184,31,54,31,149,31,149,30,191,31,169,31,10,31,10,30,181,31,181,30,201,31,192,31,116,31,189,31,41,31,41,30,93,31,130,31,97,31,113,31,113,30,68,31,59,31,15,31,19,31,32,31,32,30,122,31,14,31,242,31,146,31,146,30,45,31,4,31,228,31,190,31,190,30,133,31,133,30,19,31,13,31,19,31,222,31,89,31,11,31,116,31,61,31,212,31,212,30,212,29,242,31,196,31,196,30,244,31,244,30,244,29,55,31,153,31,120,31,17,31,94,31,253,31,76,31,251,31,251,30,251,29,251,28,65,31,174,31,245,31,237,31,50,31,50,30,207,31,196,31,231,31,209,31,50,31,170,31,2,31,2,30,175,31,206,31,206,30,234,31,234,31,135,31,58,31,58,30,58,29,205,31,162,31,162,30,162,29,92,31,92,30,92,29,129,31,2,31,2,30,88,31,31,31,167,31,167,30,167,29,221,31,125,31,125,30,130,31,134,31,152,31,250,31,16,31,232,31,232,30,232,29,163,31,163,30,220,31,29,31,83,31,83,30,155,31,138,31,157,31,151,31,151,30,151,29,45,31,205,31,28,31,9,31,70,31,220,31,220,30,27,31,213,31,106,31,106,30,81,31,112,31,15,31,209,31,209,30,160,31,14,31,20,31,157,31,191,31,191,30,248,31,173,31,200,31,50,31,231,31,238,31,188,31,20,31,235,31,235,30,239,31,16,31,252,31,252,30,252,29,161,31,21,31,135,31,113,31,113,30,188,31,245,31,42,31,42,30,58,31,151,31,128,31,218,31,144,31,253,31,25,31,186,31,181,31,164,31,121,31,78,31,201,31,75,31,231,31,111,31,250,31,178,31,62,31,62,30,62,29,30,31,202,31,178,31,61,31,33,31,33,30,135,31,135,30,199,31,54,31,237,31,42,31,11,31,12,31,205,31,67,31,135,31,103,31,103,30,126,31,219,31,123,31,79,31,79,30,79,29,217,31,227,31,4,31,113,31,22,31,46,31,46,30,46,31,46,30,166,31,204,31,115,31,29,31,29,30,244,31,252,31,192,31,192,30,222,31,165,31,71,31,189,31,189,30,174,31,194,31,190,31,94,31,197,31,238,31,95,31,125,31,189,31,255,31,255,30,45,31,90,31,254,31,254,30,69,31,84,31,136,31,60,31,121,31,161,31,66,31,189,31,101,31,211,31,211,30,247,31,230,31,230,30,17,31,1,31,53,31,185,31,90,31,14,31,150,31,177,31,48,31,196,31,69,31,220,31,77,31,10,31,10,30,96,31,157,31,157,30,69,31,147,31,207,31,207,30,207,29,159,31,174,31,174,30,53,31,81,31,151,31,11,31,235,31,198,31,254,31,79,31,255,31,194,31,60,31,60,30,69,31,253,31,69,31,14,31,28,31,14,31,36,31,73,31,73,30,73,29,223,31,144,31,125,31,125,30,125,29,113,31,113,30,233,31,44,31,156,31,1,31,184,31,2,31,204,31,40,31,230,31,230,30,117,31,241,31,241,30,241,29,207,31,124,31,59,31,132,31,138,31,127,31,127,30,127,29,253,31,214,31,47,31,14,31,136,31,88,31,147,31,248,31,143,31,221,31,221,30,158,31,148,31,148,30,138,31,79,31,10,31,190,31,242,31,106,31,63,31,12,31,154,31,38,31,111,31,63,31,49,31,49,30,58,31,225,31,241,31,8,31,94,31,94,30,94,29,124,31,244,31,173,31,173,30,22,31,251,31,215,31,86,31,140,31,54,31,170,31,137,31,3,31,3,30,46,31,46,30,205,31,84,31,84,30,180,31,78,31,30,31,68,31,135,31,33,31,33,30,76,31,233,31,26,31,58,31,67,31,67,30,225,31,55,31,79,31,3,31,58,31,218,31,143,31,242,31,178,31,178,30,84,31,57,31,213,31,181,31,53,31,53,30,183,31,80,31,125,31,106,31,113,31,76,31,76,30,124,31,231,31,237,31,180,31,136,31,68,31,68,30,107,31,108,31,63,31,123,31,31,31,13,31,131,31,210,31,53,31,230,31,113,31,23,31,23,30,245,31,18,31,155,31,155,30,232,31,66,31,66,30,66,29,45,31,79,31,33,31,254,31,239,31,239,30,239,29,60,31,37,31,88,31,29,31,251,31,151,31,214,31,170,31,209,31,22,31,154,31,121,31,121,30,177,31,93,31,93,30,119,31,240,31,162,31,109,31,65,31,20,31,189,31,189,30,189,29,55,31,229,31,229,30,36,31,44,31,44,30,24,31,126,31,115,31,198,31,36,31,151,31,61,31,64,31,64,30,150,31,150,30,150,29,128,31,4,31,6,31,6,30,200,31,97,31,6,31,247,31,146,31,80,31,197,31,196,31,196,30,174,31,195,31,234,31,20,31,175,31,35,31,245,31,164,31,48,31,37,31,172,31,172,30,207,31,248,31,16,31,195,31,195,30,195,29,195,28,113,31,225,31,225,30,225,29,225,28,190,31,192,31,113,31,113,30,113,29,45,31,234,31,5,31,5,30,237,31,111,31,217,31,217,30,87,31,57,31,174,31,174,30,174,29,217,31,147,31,224,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
