-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_17 is
end project_tb_17;

architecture project_tb_arch_17 of project_tb_17 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 407;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,0,0,15,0,226,0,99,0,140,0,90,0,0,0,1,0,13,0,0,0,112,0,235,0,134,0,1,0,0,0,187,0,27,0,0,0,2,0,25,0,0,0,191,0,0,0,45,0,0,0,97,0,54,0,0,0,8,0,173,0,0,0,148,0,169,0,20,0,109,0,221,0,33,0,28,0,196,0,131,0,242,0,0,0,183,0,0,0,0,0,144,0,0,0,46,0,51,0,0,0,0,0,150,0,7,0,190,0,240,0,0,0,155,0,0,0,33,0,39,0,0,0,88,0,155,0,141,0,170,0,250,0,175,0,0,0,161,0,0,0,175,0,130,0,245,0,103,0,101,0,239,0,0,0,0,0,0,0,141,0,49,0,100,0,24,0,178,0,127,0,207,0,146,0,248,0,153,0,0,0,88,0,237,0,156,0,34,0,0,0,85,0,0,0,0,0,83,0,164,0,141,0,91,0,38,0,64,0,0,0,206,0,137,0,229,0,168,0,147,0,0,0,0,0,86,0,97,0,241,0,116,0,33,0,248,0,10,0,191,0,243,0,145,0,0,0,220,0,0,0,148,0,131,0,18,0,11,0,219,0,33,0,116,0,0,0,178,0,221,0,150,0,99,0,72,0,33,0,175,0,0,0,102,0,0,0,193,0,156,0,178,0,0,0,56,0,244,0,168,0,170,0,160,0,112,0,0,0,255,0,24,0,97,0,73,0,92,0,196,0,0,0,229,0,193,0,226,0,136,0,101,0,29,0,97,0,0,0,137,0,14,0,107,0,245,0,239,0,235,0,0,0,12,0,39,0,0,0,177,0,0,0,80,0,177,0,14,0,58,0,203,0,0,0,139,0,79,0,232,0,36,0,68,0,220,0,198,0,0,0,74,0,0,0,196,0,195,0,4,0,224,0,28,0,247,0,238,0,0,0,15,0,0,0,190,0,187,0,0,0,90,0,246,0,66,0,42,0,19,0,0,0,125,0,186,0,0,0,131,0,82,0,241,0,60,0,88,0,85,0,211,0,248,0,137,0,66,0,43,0,246,0,69,0,245,0,197,0,0,0,218,0,45,0,29,0,141,0,0,0,0,0,0,0,46,0,49,0,214,0,245,0,118,0,127,0,65,0,5,0,68,0,111,0,94,0,123,0,198,0,158,0,130,0,134,0,224,0,178,0,135,0,52,0,0,0,254,0,0,0,140,0,152,0,69,0,204,0,254,0,158,0,222,0,32,0,0,0,0,0,180,0,154,0,0,0,21,0,182,0,28,0,0,0,249,0,185,0,28,0,218,0,106,0,221,0,40,0,138,0,207,0,0,0,101,0,170,0,128,0,39,0,2,0,0,0,76,0,0,0,168,0,51,0,0,0,0,0,219,0,207,0,19,0,30,0,224,0,67,0,20,0,242,0,241,0,55,0,69,0,70,0,7,0,129,0,216,0,0,0,51,0,76,0,144,0,46,0,11,0,72,0,0,0,0,0,86,0,36,0,110,0,12,0,132,0,105,0,61,0,34,0,144,0,115,0,197,0,22,0,206,0,158,0,79,0,0,0,218,0,0,0,0,0,0,0,52,0,173,0,118,0,211,0,52,0,186,0,221,0,174,0,0,0,67,0,35,0,198,0,242,0,237,0,176,0,0,0,213,0,212,0,39,0,0,0,10,0,193,0,0,0,0,0,0,0,18,0,189,0,151,0,36,0,10,0,39,0,0,0,210,0,0,0,0,0,217,0,6,0,0,0,26,0,0,0,105,0,83,0,146,0,21,0,217,0,226,0,221,0,172,0,0,0,180,0,147,0,18,0,6,0,0,0,24,0,0,0,43,0,0,0);
signal scenario_full  : scenario_type := (56,31,56,30,15,31,226,31,99,31,140,31,90,31,90,30,1,31,13,31,13,30,112,31,235,31,134,31,1,31,1,30,187,31,27,31,27,30,2,31,25,31,25,30,191,31,191,30,45,31,45,30,97,31,54,31,54,30,8,31,173,31,173,30,148,31,169,31,20,31,109,31,221,31,33,31,28,31,196,31,131,31,242,31,242,30,183,31,183,30,183,29,144,31,144,30,46,31,51,31,51,30,51,29,150,31,7,31,190,31,240,31,240,30,155,31,155,30,33,31,39,31,39,30,88,31,155,31,141,31,170,31,250,31,175,31,175,30,161,31,161,30,175,31,130,31,245,31,103,31,101,31,239,31,239,30,239,29,239,28,141,31,49,31,100,31,24,31,178,31,127,31,207,31,146,31,248,31,153,31,153,30,88,31,237,31,156,31,34,31,34,30,85,31,85,30,85,29,83,31,164,31,141,31,91,31,38,31,64,31,64,30,206,31,137,31,229,31,168,31,147,31,147,30,147,29,86,31,97,31,241,31,116,31,33,31,248,31,10,31,191,31,243,31,145,31,145,30,220,31,220,30,148,31,131,31,18,31,11,31,219,31,33,31,116,31,116,30,178,31,221,31,150,31,99,31,72,31,33,31,175,31,175,30,102,31,102,30,193,31,156,31,178,31,178,30,56,31,244,31,168,31,170,31,160,31,112,31,112,30,255,31,24,31,97,31,73,31,92,31,196,31,196,30,229,31,193,31,226,31,136,31,101,31,29,31,97,31,97,30,137,31,14,31,107,31,245,31,239,31,235,31,235,30,12,31,39,31,39,30,177,31,177,30,80,31,177,31,14,31,58,31,203,31,203,30,139,31,79,31,232,31,36,31,68,31,220,31,198,31,198,30,74,31,74,30,196,31,195,31,4,31,224,31,28,31,247,31,238,31,238,30,15,31,15,30,190,31,187,31,187,30,90,31,246,31,66,31,42,31,19,31,19,30,125,31,186,31,186,30,131,31,82,31,241,31,60,31,88,31,85,31,211,31,248,31,137,31,66,31,43,31,246,31,69,31,245,31,197,31,197,30,218,31,45,31,29,31,141,31,141,30,141,29,141,28,46,31,49,31,214,31,245,31,118,31,127,31,65,31,5,31,68,31,111,31,94,31,123,31,198,31,158,31,130,31,134,31,224,31,178,31,135,31,52,31,52,30,254,31,254,30,140,31,152,31,69,31,204,31,254,31,158,31,222,31,32,31,32,30,32,29,180,31,154,31,154,30,21,31,182,31,28,31,28,30,249,31,185,31,28,31,218,31,106,31,221,31,40,31,138,31,207,31,207,30,101,31,170,31,128,31,39,31,2,31,2,30,76,31,76,30,168,31,51,31,51,30,51,29,219,31,207,31,19,31,30,31,224,31,67,31,20,31,242,31,241,31,55,31,69,31,70,31,7,31,129,31,216,31,216,30,51,31,76,31,144,31,46,31,11,31,72,31,72,30,72,29,86,31,36,31,110,31,12,31,132,31,105,31,61,31,34,31,144,31,115,31,197,31,22,31,206,31,158,31,79,31,79,30,218,31,218,30,218,29,218,28,52,31,173,31,118,31,211,31,52,31,186,31,221,31,174,31,174,30,67,31,35,31,198,31,242,31,237,31,176,31,176,30,213,31,212,31,39,31,39,30,10,31,193,31,193,30,193,29,193,28,18,31,189,31,151,31,36,31,10,31,39,31,39,30,210,31,210,30,210,29,217,31,6,31,6,30,26,31,26,30,105,31,83,31,146,31,21,31,217,31,226,31,221,31,172,31,172,30,180,31,147,31,18,31,6,31,6,30,24,31,24,30,43,31,43,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
