-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 296;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (161,0,0,0,6,0,110,0,46,0,190,0,0,0,0,0,108,0,158,0,0,0,192,0,0,0,123,0,53,0,0,0,97,0,153,0,247,0,178,0,0,0,124,0,233,0,0,0,69,0,112,0,79,0,0,0,88,0,73,0,37,0,0,0,211,0,182,0,189,0,195,0,131,0,149,0,86,0,125,0,167,0,188,0,61,0,236,0,0,0,0,0,223,0,100,0,218,0,12,0,205,0,43,0,83,0,201,0,0,0,0,0,146,0,43,0,80,0,92,0,33,0,60,0,89,0,250,0,255,0,131,0,55,0,135,0,0,0,251,0,146,0,245,0,57,0,29,0,58,0,255,0,198,0,166,0,3,0,185,0,217,0,24,0,0,0,107,0,77,0,204,0,128,0,60,0,100,0,0,0,0,0,55,0,0,0,12,0,67,0,151,0,192,0,54,0,125,0,77,0,196,0,211,0,172,0,0,0,223,0,150,0,143,0,90,0,241,0,81,0,103,0,45,0,196,0,0,0,110,0,224,0,247,0,93,0,42,0,5,0,229,0,0,0,169,0,234,0,0,0,0,0,93,0,204,0,243,0,112,0,0,0,66,0,213,0,0,0,0,0,204,0,146,0,90,0,57,0,139,0,226,0,0,0,110,0,46,0,52,0,186,0,0,0,5,0,107,0,93,0,0,0,0,0,137,0,224,0,189,0,84,0,222,0,92,0,74,0,241,0,40,0,79,0,0,0,44,0,207,0,194,0,93,0,24,0,154,0,42,0,100,0,94,0,45,0,17,0,41,0,207,0,71,0,140,0,140,0,0,0,5,0,195,0,0,0,1,0,185,0,250,0,189,0,92,0,254,0,222,0,31,0,121,0,0,0,210,0,149,0,74,0,136,0,79,0,88,0,141,0,188,0,48,0,162,0,0,0,123,0,0,0,243,0,166,0,93,0,218,0,197,0,0,0,254,0,100,0,0,0,232,0,132,0,227,0,79,0,63,0,68,0,19,0,167,0,0,0,75,0,101,0,245,0,0,0,0,0,0,0,0,0,124,0,82,0,116,0,42,0,0,0,203,0,51,0,250,0,121,0,18,0,14,0,0,0,2,0,1,0,206,0,10,0,0,0,0,0,42,0,75,0,226,0,98,0,52,0,0,0,148,0,147,0,4,0,0,0,167,0,29,0,234,0,125,0,52,0,200,0,67,0,4,0,232,0,13,0,210,0,153,0,0,0,0,0,0,0,133,0,45,0,23,0,140,0,129,0,222,0,81,0,29,0,0,0,10,0,34,0,144,0,0,0,218,0,198,0,231,0,97,0,0,0,69,0,0,0,226,0,0,0);
signal scenario_full  : scenario_type := (161,31,161,30,6,31,110,31,46,31,190,31,190,30,190,29,108,31,158,31,158,30,192,31,192,30,123,31,53,31,53,30,97,31,153,31,247,31,178,31,178,30,124,31,233,31,233,30,69,31,112,31,79,31,79,30,88,31,73,31,37,31,37,30,211,31,182,31,189,31,195,31,131,31,149,31,86,31,125,31,167,31,188,31,61,31,236,31,236,30,236,29,223,31,100,31,218,31,12,31,205,31,43,31,83,31,201,31,201,30,201,29,146,31,43,31,80,31,92,31,33,31,60,31,89,31,250,31,255,31,131,31,55,31,135,31,135,30,251,31,146,31,245,31,57,31,29,31,58,31,255,31,198,31,166,31,3,31,185,31,217,31,24,31,24,30,107,31,77,31,204,31,128,31,60,31,100,31,100,30,100,29,55,31,55,30,12,31,67,31,151,31,192,31,54,31,125,31,77,31,196,31,211,31,172,31,172,30,223,31,150,31,143,31,90,31,241,31,81,31,103,31,45,31,196,31,196,30,110,31,224,31,247,31,93,31,42,31,5,31,229,31,229,30,169,31,234,31,234,30,234,29,93,31,204,31,243,31,112,31,112,30,66,31,213,31,213,30,213,29,204,31,146,31,90,31,57,31,139,31,226,31,226,30,110,31,46,31,52,31,186,31,186,30,5,31,107,31,93,31,93,30,93,29,137,31,224,31,189,31,84,31,222,31,92,31,74,31,241,31,40,31,79,31,79,30,44,31,207,31,194,31,93,31,24,31,154,31,42,31,100,31,94,31,45,31,17,31,41,31,207,31,71,31,140,31,140,31,140,30,5,31,195,31,195,30,1,31,185,31,250,31,189,31,92,31,254,31,222,31,31,31,121,31,121,30,210,31,149,31,74,31,136,31,79,31,88,31,141,31,188,31,48,31,162,31,162,30,123,31,123,30,243,31,166,31,93,31,218,31,197,31,197,30,254,31,100,31,100,30,232,31,132,31,227,31,79,31,63,31,68,31,19,31,167,31,167,30,75,31,101,31,245,31,245,30,245,29,245,28,245,27,124,31,82,31,116,31,42,31,42,30,203,31,51,31,250,31,121,31,18,31,14,31,14,30,2,31,1,31,206,31,10,31,10,30,10,29,42,31,75,31,226,31,98,31,52,31,52,30,148,31,147,31,4,31,4,30,167,31,29,31,234,31,125,31,52,31,200,31,67,31,4,31,232,31,13,31,210,31,153,31,153,30,153,29,153,28,133,31,45,31,23,31,140,31,129,31,222,31,81,31,29,31,29,30,10,31,34,31,144,31,144,30,218,31,198,31,231,31,97,31,97,30,69,31,69,30,226,31,226,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
