-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 424;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,234,0,146,0,166,0,0,0,199,0,121,0,136,0,32,0,0,0,82,0,189,0,96,0,249,0,99,0,232,0,77,0,101,0,247,0,210,0,134,0,236,0,57,0,193,0,161,0,205,0,0,0,66,0,203,0,15,0,41,0,42,0,99,0,211,0,0,0,46,0,253,0,122,0,238,0,0,0,0,0,0,0,84,0,44,0,252,0,165,0,55,0,64,0,140,0,176,0,106,0,16,0,0,0,151,0,94,0,246,0,228,0,254,0,215,0,73,0,0,0,137,0,0,0,3,0,100,0,164,0,192,0,0,0,0,0,0,0,177,0,24,0,78,0,177,0,0,0,65,0,0,0,0,0,249,0,53,0,220,0,128,0,1,0,124,0,45,0,235,0,81,0,3,0,101,0,232,0,216,0,187,0,167,0,0,0,138,0,0,0,0,0,155,0,49,0,131,0,255,0,190,0,240,0,232,0,84,0,121,0,11,0,0,0,45,0,19,0,15,0,168,0,10,0,242,0,242,0,67,0,240,0,1,0,198,0,145,0,57,0,113,0,128,0,233,0,143,0,126,0,0,0,24,0,111,0,194,0,0,0,39,0,242,0,241,0,226,0,14,0,141,0,253,0,0,0,165,0,23,0,255,0,172,0,20,0,126,0,43,0,39,0,106,0,0,0,99,0,137,0,201,0,153,0,186,0,0,0,217,0,80,0,37,0,70,0,193,0,0,0,157,0,10,0,173,0,13,0,0,0,183,0,0,0,12,0,71,0,232,0,29,0,139,0,173,0,97,0,243,0,167,0,224,0,84,0,0,0,0,0,154,0,0,0,126,0,156,0,28,0,148,0,212,0,57,0,0,0,0,0,224,0,112,0,95,0,147,0,101,0,175,0,0,0,19,0,7,0,254,0,221,0,193,0,139,0,96,0,215,0,236,0,41,0,211,0,0,0,100,0,113,0,117,0,0,0,208,0,112,0,103,0,210,0,80,0,116,0,0,0,84,0,118,0,128,0,160,0,0,0,54,0,172,0,225,0,113,0,7,0,246,0,119,0,148,0,20,0,92,0,118,0,58,0,0,0,0,0,95,0,0,0,39,0,184,0,0,0,146,0,253,0,242,0,116,0,234,0,72,0,186,0,31,0,59,0,33,0,110,0,60,0,60,0,0,0,134,0,0,0,120,0,221,0,134,0,0,0,20,0,1,0,1,0,4,0,108,0,146,0,106,0,81,0,164,0,87,0,14,0,12,0,0,0,244,0,138,0,118,0,127,0,0,0,81,0,159,0,61,0,0,0,0,0,121,0,0,0,206,0,80,0,179,0,48,0,0,0,79,0,12,0,40,0,212,0,180,0,124,0,228,0,168,0,218,0,4,0,59,0,0,0,0,0,115,0,186,0,0,0,0,0,204,0,25,0,47,0,243,0,115,0,0,0,0,0,0,0,131,0,31,0,21,0,183,0,23,0,182,0,242,0,239,0,0,0,17,0,120,0,71,0,35,0,0,0,0,0,152,0,119,0,100,0,118,0,0,0,49,0,117,0,68,0,57,0,97,0,6,0,16,0,176,0,243,0,128,0,234,0,27,0,35,0,0,0,198,0,199,0,111,0,0,0,0,0,113,0,51,0,133,0,0,0,84,0,50,0,105,0,234,0,193,0,19,0,217,0,140,0,156,0,223,0,97,0,0,0,133,0,0,0,183,0,251,0,115,0,173,0,227,0,0,0,15,0,163,0,95,0,64,0,38,0,0,0,154,0,140,0,19,0,113,0,255,0,87,0,0,0,102,0,45,0,237,0,13,0,0,0,147,0,19,0,0,0,69,0,210,0,135,0,9,0,239,0,255,0,58,0,100,0,119,0,67,0,149,0,0,0,207,0,0,0,87,0,95,0,101,0,98,0,0,0,146,0);
signal scenario_full  : scenario_type := (0,0,234,31,146,31,166,31,166,30,199,31,121,31,136,31,32,31,32,30,82,31,189,31,96,31,249,31,99,31,232,31,77,31,101,31,247,31,210,31,134,31,236,31,57,31,193,31,161,31,205,31,205,30,66,31,203,31,15,31,41,31,42,31,99,31,211,31,211,30,46,31,253,31,122,31,238,31,238,30,238,29,238,28,84,31,44,31,252,31,165,31,55,31,64,31,140,31,176,31,106,31,16,31,16,30,151,31,94,31,246,31,228,31,254,31,215,31,73,31,73,30,137,31,137,30,3,31,100,31,164,31,192,31,192,30,192,29,192,28,177,31,24,31,78,31,177,31,177,30,65,31,65,30,65,29,249,31,53,31,220,31,128,31,1,31,124,31,45,31,235,31,81,31,3,31,101,31,232,31,216,31,187,31,167,31,167,30,138,31,138,30,138,29,155,31,49,31,131,31,255,31,190,31,240,31,232,31,84,31,121,31,11,31,11,30,45,31,19,31,15,31,168,31,10,31,242,31,242,31,67,31,240,31,1,31,198,31,145,31,57,31,113,31,128,31,233,31,143,31,126,31,126,30,24,31,111,31,194,31,194,30,39,31,242,31,241,31,226,31,14,31,141,31,253,31,253,30,165,31,23,31,255,31,172,31,20,31,126,31,43,31,39,31,106,31,106,30,99,31,137,31,201,31,153,31,186,31,186,30,217,31,80,31,37,31,70,31,193,31,193,30,157,31,10,31,173,31,13,31,13,30,183,31,183,30,12,31,71,31,232,31,29,31,139,31,173,31,97,31,243,31,167,31,224,31,84,31,84,30,84,29,154,31,154,30,126,31,156,31,28,31,148,31,212,31,57,31,57,30,57,29,224,31,112,31,95,31,147,31,101,31,175,31,175,30,19,31,7,31,254,31,221,31,193,31,139,31,96,31,215,31,236,31,41,31,211,31,211,30,100,31,113,31,117,31,117,30,208,31,112,31,103,31,210,31,80,31,116,31,116,30,84,31,118,31,128,31,160,31,160,30,54,31,172,31,225,31,113,31,7,31,246,31,119,31,148,31,20,31,92,31,118,31,58,31,58,30,58,29,95,31,95,30,39,31,184,31,184,30,146,31,253,31,242,31,116,31,234,31,72,31,186,31,31,31,59,31,33,31,110,31,60,31,60,31,60,30,134,31,134,30,120,31,221,31,134,31,134,30,20,31,1,31,1,31,4,31,108,31,146,31,106,31,81,31,164,31,87,31,14,31,12,31,12,30,244,31,138,31,118,31,127,31,127,30,81,31,159,31,61,31,61,30,61,29,121,31,121,30,206,31,80,31,179,31,48,31,48,30,79,31,12,31,40,31,212,31,180,31,124,31,228,31,168,31,218,31,4,31,59,31,59,30,59,29,115,31,186,31,186,30,186,29,204,31,25,31,47,31,243,31,115,31,115,30,115,29,115,28,131,31,31,31,21,31,183,31,23,31,182,31,242,31,239,31,239,30,17,31,120,31,71,31,35,31,35,30,35,29,152,31,119,31,100,31,118,31,118,30,49,31,117,31,68,31,57,31,97,31,6,31,16,31,176,31,243,31,128,31,234,31,27,31,35,31,35,30,198,31,199,31,111,31,111,30,111,29,113,31,51,31,133,31,133,30,84,31,50,31,105,31,234,31,193,31,19,31,217,31,140,31,156,31,223,31,97,31,97,30,133,31,133,30,183,31,251,31,115,31,173,31,227,31,227,30,15,31,163,31,95,31,64,31,38,31,38,30,154,31,140,31,19,31,113,31,255,31,87,31,87,30,102,31,45,31,237,31,13,31,13,30,147,31,19,31,19,30,69,31,210,31,135,31,9,31,239,31,255,31,58,31,100,31,119,31,67,31,149,31,149,30,207,31,207,30,87,31,95,31,101,31,98,31,98,30,146,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
