-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_883 is
end project_tb_883;

architecture project_tb_arch_883 of project_tb_883 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 671;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,94,0,0,0,11,0,134,0,0,0,232,0,56,0,219,0,187,0,196,0,12,0,0,0,23,0,145,0,199,0,33,0,185,0,102,0,110,0,67,0,163,0,179,0,185,0,153,0,0,0,0,0,108,0,57,0,247,0,92,0,234,0,0,0,200,0,233,0,121,0,68,0,16,0,168,0,72,0,0,0,0,0,30,0,103,0,105,0,8,0,0,0,235,0,7,0,9,0,179,0,123,0,25,0,0,0,168,0,211,0,0,0,160,0,210,0,221,0,0,0,0,0,142,0,241,0,161,0,87,0,0,0,0,0,17,0,231,0,226,0,0,0,0,0,131,0,51,0,25,0,130,0,229,0,9,0,60,0,182,0,222,0,223,0,165,0,0,0,0,0,103,0,201,0,242,0,252,0,193,0,195,0,11,0,220,0,152,0,215,0,15,0,24,0,153,0,49,0,90,0,227,0,0,0,172,0,198,0,253,0,99,0,34,0,0,0,220,0,112,0,240,0,208,0,64,0,246,0,218,0,0,0,48,0,249,0,166,0,0,0,224,0,146,0,251,0,185,0,6,0,214,0,147,0,0,0,115,0,18,0,13,0,142,0,100,0,46,0,237,0,127,0,241,0,186,0,113,0,79,0,194,0,165,0,140,0,87,0,171,0,22,0,161,0,59,0,33,0,0,0,206,0,56,0,175,0,0,0,6,0,72,0,39,0,45,0,113,0,62,0,15,0,68,0,199,0,0,0,108,0,134,0,246,0,28,0,0,0,93,0,139,0,0,0,188,0,0,0,189,0,6,0,186,0,231,0,190,0,212,0,98,0,229,0,254,0,0,0,168,0,203,0,153,0,0,0,195,0,193,0,0,0,0,0,0,0,235,0,24,0,220,0,7,0,76,0,138,0,0,0,0,0,26,0,223,0,119,0,71,0,117,0,1,0,100,0,37,0,225,0,0,0,0,0,111,0,0,0,122,0,73,0,66,0,188,0,151,0,204,0,36,0,171,0,215,0,168,0,133,0,120,0,184,0,0,0,20,0,231,0,169,0,0,0,0,0,38,0,61,0,69,0,195,0,0,0,0,0,32,0,0,0,0,0,155,0,75,0,0,0,175,0,0,0,1,0,255,0,0,0,172,0,133,0,180,0,194,0,0,0,164,0,95,0,236,0,236,0,218,0,0,0,156,0,198,0,14,0,197,0,146,0,115,0,220,0,144,0,222,0,116,0,6,0,0,0,248,0,205,0,252,0,139,0,13,0,104,0,96,0,21,0,141,0,51,0,212,0,119,0,231,0,0,0,232,0,0,0,104,0,120,0,5,0,141,0,213,0,88,0,0,0,0,0,24,0,0,0,0,0,0,0,34,0,95,0,0,0,0,0,128,0,36,0,111,0,134,0,46,0,53,0,101,0,143,0,235,0,34,0,103,0,0,0,0,0,228,0,215,0,255,0,0,0,50,0,245,0,194,0,179,0,141,0,186,0,77,0,174,0,210,0,224,0,31,0,123,0,223,0,151,0,119,0,33,0,130,0,132,0,0,0,58,0,11,0,214,0,85,0,0,0,219,0,153,0,0,0,0,0,84,0,167,0,162,0,236,0,217,0,106,0,55,0,159,0,25,0,105,0,24,0,62,0,179,0,103,0,0,0,0,0,78,0,0,0,244,0,234,0,104,0,121,0,0,0,29,0,0,0,143,0,168,0,135,0,122,0,83,0,0,0,207,0,0,0,104,0,0,0,0,0,44,0,58,0,131,0,36,0,0,0,212,0,242,0,177,0,230,0,172,0,0,0,198,0,198,0,113,0,116,0,206,0,163,0,14,0,118,0,188,0,93,0,0,0,0,0,0,0,196,0,232,0,76,0,0,0,0,0,0,0,61,0,107,0,210,0,25,0,199,0,115,0,143,0,0,0,112,0,34,0,15,0,230,0,24,0,133,0,41,0,0,0,0,0,0,0,125,0,223,0,0,0,112,0,176,0,45,0,114,0,195,0,0,0,60,0,252,0,124,0,195,0,76,0,14,0,222,0,172,0,227,0,0,0,0,0,24,0,248,0,134,0,172,0,107,0,119,0,0,0,242,0,81,0,166,0,218,0,197,0,143,0,144,0,25,0,224,0,169,0,51,0,0,0,94,0,234,0,136,0,241,0,58,0,190,0,143,0,188,0,54,0,101,0,232,0,251,0,204,0,0,0,0,0,126,0,67,0,0,0,101,0,42,0,0,0,0,0,164,0,126,0,215,0,157,0,0,0,2,0,126,0,0,0,65,0,35,0,0,0,0,0,0,0,118,0,137,0,58,0,250,0,163,0,233,0,31,0,0,0,179,0,0,0,0,0,24,0,231,0,214,0,255,0,35,0,75,0,233,0,25,0,0,0,55,0,0,0,0,0,0,0,16,0,78,0,0,0,149,0,101,0,54,0,212,0,158,0,91,0,217,0,252,0,212,0,124,0,0,0,19,0,208,0,183,0,30,0,0,0,0,0,140,0,19,0,141,0,0,0,46,0,0,0,0,0,11,0,38,0,0,0,77,0,132,0,46,0,3,0,46,0,209,0,0,0,0,0,109,0,0,0,82,0,154,0,0,0,143,0,209,0,37,0,165,0,255,0,0,0,0,0,176,0,0,0,198,0,3,0,82,0,114,0,20,0,190,0,253,0,102,0,151,0,245,0,0,0,65,0,225,0,128,0,0,0,60,0,0,0,176,0,43,0,220,0,0,0,236,0,73,0,192,0,187,0,187,0,0,0,191,0,0,0,141,0,196,0,0,0,12,0,0,0,18,0,195,0,229,0,81,0,60,0,83,0,208,0,0,0,206,0,37,0,0,0,132,0,0,0,57,0,136,0,145,0,244,0,221,0,44,0,219,0,73,0,0,0,66,0,0,0,81,0,93,0,28,0,88,0,0,0,103,0,234,0,39,0,80,0,18,0,158,0,0,0,192,0,14,0,113,0,0,0,163,0,158,0,82,0,216,0,214,0,213,0,250,0,60,0,230,0,0,0,24,0,28,0);
signal scenario_full  : scenario_type := (0,0,94,31,94,30,11,31,134,31,134,30,232,31,56,31,219,31,187,31,196,31,12,31,12,30,23,31,145,31,199,31,33,31,185,31,102,31,110,31,67,31,163,31,179,31,185,31,153,31,153,30,153,29,108,31,57,31,247,31,92,31,234,31,234,30,200,31,233,31,121,31,68,31,16,31,168,31,72,31,72,30,72,29,30,31,103,31,105,31,8,31,8,30,235,31,7,31,9,31,179,31,123,31,25,31,25,30,168,31,211,31,211,30,160,31,210,31,221,31,221,30,221,29,142,31,241,31,161,31,87,31,87,30,87,29,17,31,231,31,226,31,226,30,226,29,131,31,51,31,25,31,130,31,229,31,9,31,60,31,182,31,222,31,223,31,165,31,165,30,165,29,103,31,201,31,242,31,252,31,193,31,195,31,11,31,220,31,152,31,215,31,15,31,24,31,153,31,49,31,90,31,227,31,227,30,172,31,198,31,253,31,99,31,34,31,34,30,220,31,112,31,240,31,208,31,64,31,246,31,218,31,218,30,48,31,249,31,166,31,166,30,224,31,146,31,251,31,185,31,6,31,214,31,147,31,147,30,115,31,18,31,13,31,142,31,100,31,46,31,237,31,127,31,241,31,186,31,113,31,79,31,194,31,165,31,140,31,87,31,171,31,22,31,161,31,59,31,33,31,33,30,206,31,56,31,175,31,175,30,6,31,72,31,39,31,45,31,113,31,62,31,15,31,68,31,199,31,199,30,108,31,134,31,246,31,28,31,28,30,93,31,139,31,139,30,188,31,188,30,189,31,6,31,186,31,231,31,190,31,212,31,98,31,229,31,254,31,254,30,168,31,203,31,153,31,153,30,195,31,193,31,193,30,193,29,193,28,235,31,24,31,220,31,7,31,76,31,138,31,138,30,138,29,26,31,223,31,119,31,71,31,117,31,1,31,100,31,37,31,225,31,225,30,225,29,111,31,111,30,122,31,73,31,66,31,188,31,151,31,204,31,36,31,171,31,215,31,168,31,133,31,120,31,184,31,184,30,20,31,231,31,169,31,169,30,169,29,38,31,61,31,69,31,195,31,195,30,195,29,32,31,32,30,32,29,155,31,75,31,75,30,175,31,175,30,1,31,255,31,255,30,172,31,133,31,180,31,194,31,194,30,164,31,95,31,236,31,236,31,218,31,218,30,156,31,198,31,14,31,197,31,146,31,115,31,220,31,144,31,222,31,116,31,6,31,6,30,248,31,205,31,252,31,139,31,13,31,104,31,96,31,21,31,141,31,51,31,212,31,119,31,231,31,231,30,232,31,232,30,104,31,120,31,5,31,141,31,213,31,88,31,88,30,88,29,24,31,24,30,24,29,24,28,34,31,95,31,95,30,95,29,128,31,36,31,111,31,134,31,46,31,53,31,101,31,143,31,235,31,34,31,103,31,103,30,103,29,228,31,215,31,255,31,255,30,50,31,245,31,194,31,179,31,141,31,186,31,77,31,174,31,210,31,224,31,31,31,123,31,223,31,151,31,119,31,33,31,130,31,132,31,132,30,58,31,11,31,214,31,85,31,85,30,219,31,153,31,153,30,153,29,84,31,167,31,162,31,236,31,217,31,106,31,55,31,159,31,25,31,105,31,24,31,62,31,179,31,103,31,103,30,103,29,78,31,78,30,244,31,234,31,104,31,121,31,121,30,29,31,29,30,143,31,168,31,135,31,122,31,83,31,83,30,207,31,207,30,104,31,104,30,104,29,44,31,58,31,131,31,36,31,36,30,212,31,242,31,177,31,230,31,172,31,172,30,198,31,198,31,113,31,116,31,206,31,163,31,14,31,118,31,188,31,93,31,93,30,93,29,93,28,196,31,232,31,76,31,76,30,76,29,76,28,61,31,107,31,210,31,25,31,199,31,115,31,143,31,143,30,112,31,34,31,15,31,230,31,24,31,133,31,41,31,41,30,41,29,41,28,125,31,223,31,223,30,112,31,176,31,45,31,114,31,195,31,195,30,60,31,252,31,124,31,195,31,76,31,14,31,222,31,172,31,227,31,227,30,227,29,24,31,248,31,134,31,172,31,107,31,119,31,119,30,242,31,81,31,166,31,218,31,197,31,143,31,144,31,25,31,224,31,169,31,51,31,51,30,94,31,234,31,136,31,241,31,58,31,190,31,143,31,188,31,54,31,101,31,232,31,251,31,204,31,204,30,204,29,126,31,67,31,67,30,101,31,42,31,42,30,42,29,164,31,126,31,215,31,157,31,157,30,2,31,126,31,126,30,65,31,35,31,35,30,35,29,35,28,118,31,137,31,58,31,250,31,163,31,233,31,31,31,31,30,179,31,179,30,179,29,24,31,231,31,214,31,255,31,35,31,75,31,233,31,25,31,25,30,55,31,55,30,55,29,55,28,16,31,78,31,78,30,149,31,101,31,54,31,212,31,158,31,91,31,217,31,252,31,212,31,124,31,124,30,19,31,208,31,183,31,30,31,30,30,30,29,140,31,19,31,141,31,141,30,46,31,46,30,46,29,11,31,38,31,38,30,77,31,132,31,46,31,3,31,46,31,209,31,209,30,209,29,109,31,109,30,82,31,154,31,154,30,143,31,209,31,37,31,165,31,255,31,255,30,255,29,176,31,176,30,198,31,3,31,82,31,114,31,20,31,190,31,253,31,102,31,151,31,245,31,245,30,65,31,225,31,128,31,128,30,60,31,60,30,176,31,43,31,220,31,220,30,236,31,73,31,192,31,187,31,187,31,187,30,191,31,191,30,141,31,196,31,196,30,12,31,12,30,18,31,195,31,229,31,81,31,60,31,83,31,208,31,208,30,206,31,37,31,37,30,132,31,132,30,57,31,136,31,145,31,244,31,221,31,44,31,219,31,73,31,73,30,66,31,66,30,81,31,93,31,28,31,88,31,88,30,103,31,234,31,39,31,80,31,18,31,158,31,158,30,192,31,14,31,113,31,113,30,163,31,158,31,82,31,216,31,214,31,213,31,250,31,60,31,230,31,230,30,24,31,28,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
