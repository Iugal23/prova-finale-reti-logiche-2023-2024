-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 752;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (227,0,152,0,0,0,0,0,25,0,144,0,40,0,34,0,0,0,230,0,0,0,3,0,0,0,149,0,0,0,24,0,0,0,156,0,0,0,0,0,0,0,0,0,65,0,0,0,86,0,235,0,179,0,62,0,111,0,0,0,234,0,0,0,62,0,127,0,117,0,115,0,241,0,228,0,186,0,173,0,190,0,13,0,85,0,13,0,168,0,19,0,249,0,114,0,0,0,11,0,51,0,135,0,237,0,249,0,230,0,26,0,3,0,19,0,0,0,31,0,116,0,0,0,0,0,68,0,0,0,113,0,198,0,0,0,148,0,0,0,40,0,0,0,88,0,20,0,153,0,157,0,217,0,198,0,156,0,10,0,120,0,37,0,227,0,1,0,181,0,239,0,190,0,201,0,82,0,3,0,146,0,57,0,26,0,231,0,61,0,0,0,0,0,172,0,178,0,158,0,197,0,0,0,0,0,130,0,45,0,53,0,184,0,246,0,0,0,151,0,51,0,186,0,0,0,0,0,196,0,173,0,0,0,253,0,177,0,237,0,91,0,46,0,62,0,0,0,220,0,153,0,9,0,169,0,0,0,195,0,68,0,211,0,0,0,144,0,188,0,190,0,239,0,201,0,0,0,0,0,153,0,225,0,9,0,243,0,0,0,213,0,0,0,0,0,0,0,0,0,116,0,148,0,207,0,38,0,83,0,186,0,210,0,109,0,163,0,91,0,0,0,50,0,48,0,27,0,15,0,232,0,148,0,88,0,79,0,12,0,119,0,159,0,226,0,0,0,62,0,123,0,218,0,242,0,185,0,161,0,124,0,212,0,5,0,0,0,0,0,172,0,33,0,0,0,146,0,182,0,1,0,32,0,0,0,21,0,155,0,65,0,134,0,154,0,243,0,45,0,17,0,139,0,217,0,128,0,232,0,222,0,0,0,97,0,0,0,0,0,0,0,0,0,193,0,217,0,131,0,178,0,214,0,62,0,242,0,104,0,0,0,58,0,247,0,33,0,0,0,0,0,163,0,130,0,61,0,139,0,171,0,0,0,121,0,8,0,42,0,0,0,176,0,2,0,200,0,0,0,121,0,228,0,0,0,7,0,55,0,237,0,69,0,173,0,247,0,149,0,226,0,107,0,186,0,237,0,0,0,150,0,44,0,227,0,0,0,231,0,154,0,0,0,0,0,176,0,238,0,68,0,0,0,203,0,93,0,254,0,77,0,0,0,0,0,228,0,5,0,45,0,130,0,0,0,47,0,218,0,96,0,85,0,0,0,148,0,72,0,130,0,168,0,7,0,240,0,134,0,83,0,100,0,142,0,21,0,23,0,12,0,108,0,71,0,153,0,0,0,243,0,242,0,203,0,0,0,77,0,0,0,18,0,232,0,122,0,147,0,60,0,0,0,108,0,0,0,105,0,225,0,0,0,62,0,139,0,156,0,213,0,5,0,0,0,248,0,84,0,92,0,0,0,0,0,141,0,206,0,181,0,128,0,0,0,239,0,30,0,45,0,0,0,0,0,42,0,208,0,142,0,7,0,223,0,173,0,122,0,208,0,0,0,255,0,228,0,26,0,195,0,0,0,218,0,52,0,143,0,14,0,166,0,134,0,226,0,0,0,0,0,233,0,153,0,180,0,0,0,0,0,115,0,92,0,153,0,248,0,0,0,132,0,171,0,165,0,224,0,239,0,74,0,0,0,177,0,221,0,154,0,140,0,0,0,153,0,194,0,86,0,230,0,4,0,121,0,196,0,204,0,14,0,0,0,234,0,11,0,0,0,133,0,0,0,236,0,34,0,166,0,143,0,0,0,190,0,189,0,13,0,120,0,15,0,183,0,159,0,208,0,236,0,124,0,17,0,25,0,187,0,128,0,71,0,216,0,209,0,45,0,0,0,33,0,14,0,7,0,0,0,216,0,229,0,0,0,0,0,146,0,217,0,108,0,0,0,99,0,0,0,254,0,195,0,187,0,34,0,0,0,0,0,239,0,0,0,63,0,208,0,0,0,81,0,0,0,107,0,131,0,33,0,164,0,190,0,70,0,0,0,9,0,0,0,141,0,239,0,134,0,55,0,237,0,234,0,173,0,59,0,181,0,240,0,0,0,191,0,198,0,145,0,81,0,184,0,28,0,157,0,183,0,99,0,156,0,116,0,248,0,224,0,143,0,190,0,237,0,0,0,43,0,32,0,170,0,46,0,141,0,91,0,0,0,0,0,0,0,142,0,60,0,190,0,42,0,0,0,94,0,174,0,209,0,127,0,1,0,0,0,62,0,0,0,117,0,32,0,35,0,158,0,224,0,154,0,86,0,41,0,197,0,158,0,63,0,0,0,0,0,176,0,243,0,43,0,100,0,173,0,173,0,0,0,72,0,120,0,57,0,0,0,64,0,154,0,0,0,54,0,247,0,93,0,135,0,108,0,0,0,170,0,0,0,206,0,244,0,160,0,189,0,0,0,161,0,254,0,158,0,0,0,122,0,84,0,66,0,147,0,231,0,248,0,0,0,51,0,29,0,0,0,106,0,21,0,0,0,146,0,79,0,7,0,0,0,36,0,0,0,0,0,204,0,111,0,132,0,236,0,182,0,206,0,230,0,0,0,254,0,133,0,0,0,70,0,4,0,131,0,33,0,42,0,115,0,195,0,178,0,130,0,143,0,87,0,0,0,0,0,0,0,128,0,94,0,88,0,35,0,5,0,174,0,51,0,0,0,18,0,54,0,56,0,137,0,0,0,0,0,0,0,24,0,0,0,30,0,99,0,130,0,192,0,41,0,179,0,211,0,0,0,91,0,112,0,155,0,244,0,0,0,244,0,115,0,235,0,32,0,222,0,97,0,98,0,114,0,14,0,210,0,0,0,86,0,170,0,19,0,0,0,95,0,3,0,0,0,123,0,86,0,154,0,217,0,130,0,0,0,178,0,147,0,59,0,245,0,198,0,23,0,242,0,231,0,14,0,0,0,7,0,176,0,63,0,43,0,0,0,235,0,3,0,0,0,178,0,238,0,195,0,192,0,64,0,171,0,10,0,111,0,23,0,78,0,36,0,240,0,196,0,199,0,19,0,62,0,147,0,62,0,35,0,203,0,194,0,0,0,44,0,204,0,43,0,248,0,70,0,35,0,171,0,0,0,53,0,252,0,0,0,252,0,13,0,144,0,115,0,54,0,189,0,59,0,5,0,133,0,12,0,0,0,0,0,125,0,78,0,15,0,0,0,197,0,0,0,16,0,153,0,197,0,35,0,143,0,0,0,0,0,163,0,212,0,0,0,0,0,255,0,0,0,0,0,96,0,225,0,246,0,0,0,166,0,25,0,103,0,36,0,153,0,135,0,129,0,31,0,182,0,229,0,138,0,176,0,222,0,0,0);
signal scenario_full  : scenario_type := (227,31,152,31,152,30,152,29,25,31,144,31,40,31,34,31,34,30,230,31,230,30,3,31,3,30,149,31,149,30,24,31,24,30,156,31,156,30,156,29,156,28,156,27,65,31,65,30,86,31,235,31,179,31,62,31,111,31,111,30,234,31,234,30,62,31,127,31,117,31,115,31,241,31,228,31,186,31,173,31,190,31,13,31,85,31,13,31,168,31,19,31,249,31,114,31,114,30,11,31,51,31,135,31,237,31,249,31,230,31,26,31,3,31,19,31,19,30,31,31,116,31,116,30,116,29,68,31,68,30,113,31,198,31,198,30,148,31,148,30,40,31,40,30,88,31,20,31,153,31,157,31,217,31,198,31,156,31,10,31,120,31,37,31,227,31,1,31,181,31,239,31,190,31,201,31,82,31,3,31,146,31,57,31,26,31,231,31,61,31,61,30,61,29,172,31,178,31,158,31,197,31,197,30,197,29,130,31,45,31,53,31,184,31,246,31,246,30,151,31,51,31,186,31,186,30,186,29,196,31,173,31,173,30,253,31,177,31,237,31,91,31,46,31,62,31,62,30,220,31,153,31,9,31,169,31,169,30,195,31,68,31,211,31,211,30,144,31,188,31,190,31,239,31,201,31,201,30,201,29,153,31,225,31,9,31,243,31,243,30,213,31,213,30,213,29,213,28,213,27,116,31,148,31,207,31,38,31,83,31,186,31,210,31,109,31,163,31,91,31,91,30,50,31,48,31,27,31,15,31,232,31,148,31,88,31,79,31,12,31,119,31,159,31,226,31,226,30,62,31,123,31,218,31,242,31,185,31,161,31,124,31,212,31,5,31,5,30,5,29,172,31,33,31,33,30,146,31,182,31,1,31,32,31,32,30,21,31,155,31,65,31,134,31,154,31,243,31,45,31,17,31,139,31,217,31,128,31,232,31,222,31,222,30,97,31,97,30,97,29,97,28,97,27,193,31,217,31,131,31,178,31,214,31,62,31,242,31,104,31,104,30,58,31,247,31,33,31,33,30,33,29,163,31,130,31,61,31,139,31,171,31,171,30,121,31,8,31,42,31,42,30,176,31,2,31,200,31,200,30,121,31,228,31,228,30,7,31,55,31,237,31,69,31,173,31,247,31,149,31,226,31,107,31,186,31,237,31,237,30,150,31,44,31,227,31,227,30,231,31,154,31,154,30,154,29,176,31,238,31,68,31,68,30,203,31,93,31,254,31,77,31,77,30,77,29,228,31,5,31,45,31,130,31,130,30,47,31,218,31,96,31,85,31,85,30,148,31,72,31,130,31,168,31,7,31,240,31,134,31,83,31,100,31,142,31,21,31,23,31,12,31,108,31,71,31,153,31,153,30,243,31,242,31,203,31,203,30,77,31,77,30,18,31,232,31,122,31,147,31,60,31,60,30,108,31,108,30,105,31,225,31,225,30,62,31,139,31,156,31,213,31,5,31,5,30,248,31,84,31,92,31,92,30,92,29,141,31,206,31,181,31,128,31,128,30,239,31,30,31,45,31,45,30,45,29,42,31,208,31,142,31,7,31,223,31,173,31,122,31,208,31,208,30,255,31,228,31,26,31,195,31,195,30,218,31,52,31,143,31,14,31,166,31,134,31,226,31,226,30,226,29,233,31,153,31,180,31,180,30,180,29,115,31,92,31,153,31,248,31,248,30,132,31,171,31,165,31,224,31,239,31,74,31,74,30,177,31,221,31,154,31,140,31,140,30,153,31,194,31,86,31,230,31,4,31,121,31,196,31,204,31,14,31,14,30,234,31,11,31,11,30,133,31,133,30,236,31,34,31,166,31,143,31,143,30,190,31,189,31,13,31,120,31,15,31,183,31,159,31,208,31,236,31,124,31,17,31,25,31,187,31,128,31,71,31,216,31,209,31,45,31,45,30,33,31,14,31,7,31,7,30,216,31,229,31,229,30,229,29,146,31,217,31,108,31,108,30,99,31,99,30,254,31,195,31,187,31,34,31,34,30,34,29,239,31,239,30,63,31,208,31,208,30,81,31,81,30,107,31,131,31,33,31,164,31,190,31,70,31,70,30,9,31,9,30,141,31,239,31,134,31,55,31,237,31,234,31,173,31,59,31,181,31,240,31,240,30,191,31,198,31,145,31,81,31,184,31,28,31,157,31,183,31,99,31,156,31,116,31,248,31,224,31,143,31,190,31,237,31,237,30,43,31,32,31,170,31,46,31,141,31,91,31,91,30,91,29,91,28,142,31,60,31,190,31,42,31,42,30,94,31,174,31,209,31,127,31,1,31,1,30,62,31,62,30,117,31,32,31,35,31,158,31,224,31,154,31,86,31,41,31,197,31,158,31,63,31,63,30,63,29,176,31,243,31,43,31,100,31,173,31,173,31,173,30,72,31,120,31,57,31,57,30,64,31,154,31,154,30,54,31,247,31,93,31,135,31,108,31,108,30,170,31,170,30,206,31,244,31,160,31,189,31,189,30,161,31,254,31,158,31,158,30,122,31,84,31,66,31,147,31,231,31,248,31,248,30,51,31,29,31,29,30,106,31,21,31,21,30,146,31,79,31,7,31,7,30,36,31,36,30,36,29,204,31,111,31,132,31,236,31,182,31,206,31,230,31,230,30,254,31,133,31,133,30,70,31,4,31,131,31,33,31,42,31,115,31,195,31,178,31,130,31,143,31,87,31,87,30,87,29,87,28,128,31,94,31,88,31,35,31,5,31,174,31,51,31,51,30,18,31,54,31,56,31,137,31,137,30,137,29,137,28,24,31,24,30,30,31,99,31,130,31,192,31,41,31,179,31,211,31,211,30,91,31,112,31,155,31,244,31,244,30,244,31,115,31,235,31,32,31,222,31,97,31,98,31,114,31,14,31,210,31,210,30,86,31,170,31,19,31,19,30,95,31,3,31,3,30,123,31,86,31,154,31,217,31,130,31,130,30,178,31,147,31,59,31,245,31,198,31,23,31,242,31,231,31,14,31,14,30,7,31,176,31,63,31,43,31,43,30,235,31,3,31,3,30,178,31,238,31,195,31,192,31,64,31,171,31,10,31,111,31,23,31,78,31,36,31,240,31,196,31,199,31,19,31,62,31,147,31,62,31,35,31,203,31,194,31,194,30,44,31,204,31,43,31,248,31,70,31,35,31,171,31,171,30,53,31,252,31,252,30,252,31,13,31,144,31,115,31,54,31,189,31,59,31,5,31,133,31,12,31,12,30,12,29,125,31,78,31,15,31,15,30,197,31,197,30,16,31,153,31,197,31,35,31,143,31,143,30,143,29,163,31,212,31,212,30,212,29,255,31,255,30,255,29,96,31,225,31,246,31,246,30,166,31,25,31,103,31,36,31,153,31,135,31,129,31,31,31,182,31,229,31,138,31,176,31,222,31,222,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
