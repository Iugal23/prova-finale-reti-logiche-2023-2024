-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 986;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,223,0,0,0,111,0,98,0,121,0,105,0,178,0,84,0,120,0,210,0,41,0,10,0,178,0,115,0,19,0,196,0,241,0,65,0,42,0,255,0,0,0,0,0,189,0,107,0,4,0,2,0,95,0,9,0,179,0,120,0,130,0,58,0,5,0,208,0,101,0,124,0,139,0,186,0,167,0,199,0,196,0,119,0,0,0,147,0,246,0,0,0,53,0,77,0,89,0,38,0,81,0,33,0,0,0,0,0,92,0,5,0,61,0,24,0,170,0,69,0,135,0,0,0,32,0,66,0,194,0,136,0,72,0,13,0,0,0,33,0,210,0,233,0,0,0,169,0,52,0,158,0,0,0,121,0,225,0,127,0,46,0,154,0,0,0,218,0,148,0,0,0,148,0,249,0,215,0,170,0,139,0,103,0,0,0,146,0,51,0,208,0,140,0,110,0,73,0,5,0,12,0,0,0,0,0,180,0,22,0,113,0,103,0,0,0,51,0,249,0,0,0,111,0,224,0,229,0,184,0,165,0,0,0,98,0,140,0,165,0,114,0,78,0,210,0,115,0,172,0,189,0,76,0,46,0,138,0,1,0,8,0,0,0,218,0,189,0,38,0,10,0,185,0,0,0,213,0,69,0,134,0,77,0,229,0,0,0,54,0,3,0,0,0,203,0,111,0,39,0,120,0,95,0,182,0,0,0,79,0,53,0,215,0,39,0,254,0,109,0,41,0,64,0,149,0,0,0,223,0,0,0,118,0,92,0,253,0,0,0,170,0,232,0,18,0,112,0,221,0,0,0,0,0,92,0,128,0,0,0,236,0,0,0,164,0,166,0,80,0,0,0,172,0,83,0,19,0,0,0,0,0,214,0,133,0,76,0,66,0,206,0,124,0,170,0,0,0,183,0,0,0,0,0,46,0,39,0,80,0,0,0,0,0,0,0,85,0,103,0,0,0,246,0,7,0,176,0,243,0,79,0,42,0,30,0,0,0,133,0,0,0,0,0,22,0,56,0,193,0,224,0,0,0,156,0,75,0,255,0,0,0,132,0,0,0,237,0,221,0,158,0,0,0,235,0,234,0,183,0,40,0,0,0,61,0,0,0,6,0,0,0,197,0,81,0,26,0,221,0,67,0,189,0,0,0,108,0,104,0,252,0,234,0,55,0,112,0,216,0,66,0,203,0,62,0,134,0,10,0,0,0,24,0,94,0,122,0,197,0,67,0,0,0,0,0,0,0,121,0,119,0,0,0,213,0,125,0,93,0,0,0,49,0,0,0,0,0,80,0,212,0,0,0,5,0,112,0,254,0,0,0,0,0,186,0,191,0,68,0,75,0,233,0,190,0,0,0,177,0,34,0,118,0,0,0,64,0,168,0,35,0,0,0,205,0,217,0,217,0,185,0,113,0,43,0,91,0,150,0,42,0,191,0,0,0,217,0,201,0,234,0,0,0,0,0,0,0,89,0,11,0,244,0,168,0,0,0,18,0,134,0,196,0,14,0,80,0,0,0,172,0,184,0,93,0,215,0,0,0,29,0,157,0,90,0,29,0,163,0,167,0,0,0,0,0,194,0,0,0,166,0,118,0,139,0,0,0,243,0,132,0,110,0,174,0,105,0,0,0,167,0,231,0,249,0,133,0,87,0,47,0,175,0,59,0,21,0,140,0,193,0,0,0,185,0,82,0,97,0,235,0,166,0,75,0,218,0,39,0,100,0,184,0,193,0,245,0,209,0,113,0,218,0,132,0,100,0,0,0,50,0,0,0,163,0,0,0,165,0,154,0,210,0,167,0,0,0,0,0,174,0,40,0,0,0,118,0,52,0,72,0,167,0,0,0,146,0,28,0,70,0,0,0,107,0,176,0,233,0,0,0,106,0,4,0,203,0,137,0,162,0,148,0,44,0,188,0,0,0,0,0,0,0,191,0,33,0,79,0,85,0,0,0,204,0,11,0,30,0,14,0,226,0,195,0,206,0,148,0,54,0,118,0,230,0,122,0,120,0,0,0,103,0,106,0,101,0,6,0,0,0,79,0,111,0,99,0,63,0,0,0,25,0,77,0,0,0,128,0,0,0,186,0,166,0,53,0,0,0,137,0,125,0,0,0,237,0,78,0,148,0,0,0,244,0,167,0,42,0,235,0,126,0,70,0,56,0,233,0,237,0,132,0,0,0,0,0,246,0,173,0,53,0,0,0,189,0,108,0,161,0,241,0,238,0,76,0,181,0,77,0,249,0,195,0,0,0,54,0,155,0,87,0,45,0,204,0,233,0,0,0,105,0,175,0,154,0,0,0,179,0,126,0,0,0,59,0,21,0,125,0,108,0,117,0,229,0,163,0,0,0,63,0,0,0,18,0,0,0,80,0,134,0,80,0,198,0,250,0,235,0,132,0,39,0,63,0,250,0,11,0,0,0,10,0,63,0,211,0,200,0,115,0,143,0,198,0,0,0,179,0,249,0,197,0,41,0,126,0,189,0,0,0,0,0,241,0,237,0,150,0,178,0,0,0,0,0,202,0,195,0,241,0,200,0,196,0,0,0,0,0,162,0,220,0,124,0,65,0,60,0,126,0,89,0,230,0,0,0,16,0,0,0,90,0,89,0,210,0,0,0,170,0,74,0,71,0,0,0,117,0,108,0,73,0,255,0,35,0,112,0,0,0,171,0,215,0,45,0,57,0,0,0,61,0,38,0,177,0,235,0,129,0,49,0,221,0,194,0,199,0,127,0,10,0,78,0,0,0,183,0,218,0,154,0,207,0,250,0,166,0,250,0,132,0,252,0,60,0,0,0,248,0,222,0,238,0,0,0,73,0,188,0,0,0,45,0,211,0,250,0,121,0,242,0,129,0,186,0,146,0,23,0,59,0,94,0,50,0,32,0,35,0,9,0,135,0,0,0,0,0,133,0,0,0,164,0,0,0,105,0,38,0,0,0,58,0,137,0,170,0,0,0,78,0,196,0,85,0,0,0,116,0,0,0,4,0,0,0,78,0,185,0,0,0,0,0,211,0,89,0,222,0,0,0,185,0,0,0,12,0,48,0,57,0,56,0,0,0,52,0,160,0,133,0,236,0,159,0,4,0,0,0,86,0,0,0,70,0,162,0,189,0,90,0,32,0,127,0,140,0,69,0,235,0,188,0,57,0,0,0,138,0,0,0,108,0,84,0,0,0,0,0,16,0,11,0,53,0,24,0,23,0,213,0,0,0,31,0,253,0,138,0,134,0,87,0,51,0,0,0,0,0,109,0,0,0,149,0,164,0,187,0,67,0,0,0,161,0,77,0,15,0,214,0,0,0,0,0,0,0,225,0,212,0,241,0,0,0,112,0,71,0,117,0,223,0,133,0,0,0,81,0,166,0,48,0,140,0,0,0,182,0,253,0,28,0,29,0,68,0,0,0,115,0,143,0,17,0,25,0,27,0,0,0,0,0,253,0,0,0,71,0,91,0,189,0,0,0,243,0,177,0,2,0,0,0,89,0,0,0,166,0,18,0,138,0,188,0,243,0,149,0,80,0,0,0,67,0,62,0,150,0,0,0,249,0,0,0,104,0,100,0,153,0,78,0,181,0,229,0,0,0,123,0,66,0,213,0,17,0,125,0,39,0,118,0,20,0,189,0,0,0,157,0,0,0,0,0,75,0,253,0,0,0,238,0,145,0,0,0,102,0,0,0,89,0,244,0,0,0,242,0,0,0,97,0,180,0,0,0,250,0,0,0,227,0,24,0,85,0,115,0,126,0,175,0,232,0,211,0,0,0,103,0,57,0,208,0,0,0,63,0,191,0,197,0,204,0,0,0,114,0,135,0,0,0,225,0,39,0,39,0,8,0,168,0,239,0,161,0,88,0,146,0,87,0,107,0,205,0,150,0,5,0,0,0,198,0,165,0,140,0,5,0,124,0,32,0,109,0,0,0,67,0,0,0,114,0,199,0,208,0,64,0,0,0,0,0,162,0,161,0,0,0,0,0,170,0,200,0,0,0,206,0,0,0,144,0,50,0,229,0,205,0,216,0,0,0,17,0,241,0,174,0,0,0,254,0,241,0,170,0,184,0,77,0,15,0,32,0,237,0,0,0,136,0,240,0,237,0,0,0,132,0,245,0,0,0,0,0,98,0,125,0,170,0,79,0,178,0,73,0,0,0,70,0,0,0,158,0,106,0,235,0,189,0,129,0,146,0,67,0,188,0,253,0,0,0,103,0,40,0,0,0,0,0,70,0,225,0,49,0,148,0,0,0,169,0,91,0,37,0,0,0,163,0,0,0,129,0,220,0,0,0,163,0,111,0,65,0,244,0,222,0,104,0,122,0,198,0,243,0,76,0,242,0,0,0,114,0,129,0,79,0,0,0,71,0,99,0,0,0,0,0,172,0,0,0,229,0,66,0,0,0,80,0,160,0,153,0,228,0,19,0,0,0,220,0);
signal scenario_full  : scenario_type := (71,31,223,31,223,30,111,31,98,31,121,31,105,31,178,31,84,31,120,31,210,31,41,31,10,31,178,31,115,31,19,31,196,31,241,31,65,31,42,31,255,31,255,30,255,29,189,31,107,31,4,31,2,31,95,31,9,31,179,31,120,31,130,31,58,31,5,31,208,31,101,31,124,31,139,31,186,31,167,31,199,31,196,31,119,31,119,30,147,31,246,31,246,30,53,31,77,31,89,31,38,31,81,31,33,31,33,30,33,29,92,31,5,31,61,31,24,31,170,31,69,31,135,31,135,30,32,31,66,31,194,31,136,31,72,31,13,31,13,30,33,31,210,31,233,31,233,30,169,31,52,31,158,31,158,30,121,31,225,31,127,31,46,31,154,31,154,30,218,31,148,31,148,30,148,31,249,31,215,31,170,31,139,31,103,31,103,30,146,31,51,31,208,31,140,31,110,31,73,31,5,31,12,31,12,30,12,29,180,31,22,31,113,31,103,31,103,30,51,31,249,31,249,30,111,31,224,31,229,31,184,31,165,31,165,30,98,31,140,31,165,31,114,31,78,31,210,31,115,31,172,31,189,31,76,31,46,31,138,31,1,31,8,31,8,30,218,31,189,31,38,31,10,31,185,31,185,30,213,31,69,31,134,31,77,31,229,31,229,30,54,31,3,31,3,30,203,31,111,31,39,31,120,31,95,31,182,31,182,30,79,31,53,31,215,31,39,31,254,31,109,31,41,31,64,31,149,31,149,30,223,31,223,30,118,31,92,31,253,31,253,30,170,31,232,31,18,31,112,31,221,31,221,30,221,29,92,31,128,31,128,30,236,31,236,30,164,31,166,31,80,31,80,30,172,31,83,31,19,31,19,30,19,29,214,31,133,31,76,31,66,31,206,31,124,31,170,31,170,30,183,31,183,30,183,29,46,31,39,31,80,31,80,30,80,29,80,28,85,31,103,31,103,30,246,31,7,31,176,31,243,31,79,31,42,31,30,31,30,30,133,31,133,30,133,29,22,31,56,31,193,31,224,31,224,30,156,31,75,31,255,31,255,30,132,31,132,30,237,31,221,31,158,31,158,30,235,31,234,31,183,31,40,31,40,30,61,31,61,30,6,31,6,30,197,31,81,31,26,31,221,31,67,31,189,31,189,30,108,31,104,31,252,31,234,31,55,31,112,31,216,31,66,31,203,31,62,31,134,31,10,31,10,30,24,31,94,31,122,31,197,31,67,31,67,30,67,29,67,28,121,31,119,31,119,30,213,31,125,31,93,31,93,30,49,31,49,30,49,29,80,31,212,31,212,30,5,31,112,31,254,31,254,30,254,29,186,31,191,31,68,31,75,31,233,31,190,31,190,30,177,31,34,31,118,31,118,30,64,31,168,31,35,31,35,30,205,31,217,31,217,31,185,31,113,31,43,31,91,31,150,31,42,31,191,31,191,30,217,31,201,31,234,31,234,30,234,29,234,28,89,31,11,31,244,31,168,31,168,30,18,31,134,31,196,31,14,31,80,31,80,30,172,31,184,31,93,31,215,31,215,30,29,31,157,31,90,31,29,31,163,31,167,31,167,30,167,29,194,31,194,30,166,31,118,31,139,31,139,30,243,31,132,31,110,31,174,31,105,31,105,30,167,31,231,31,249,31,133,31,87,31,47,31,175,31,59,31,21,31,140,31,193,31,193,30,185,31,82,31,97,31,235,31,166,31,75,31,218,31,39,31,100,31,184,31,193,31,245,31,209,31,113,31,218,31,132,31,100,31,100,30,50,31,50,30,163,31,163,30,165,31,154,31,210,31,167,31,167,30,167,29,174,31,40,31,40,30,118,31,52,31,72,31,167,31,167,30,146,31,28,31,70,31,70,30,107,31,176,31,233,31,233,30,106,31,4,31,203,31,137,31,162,31,148,31,44,31,188,31,188,30,188,29,188,28,191,31,33,31,79,31,85,31,85,30,204,31,11,31,30,31,14,31,226,31,195,31,206,31,148,31,54,31,118,31,230,31,122,31,120,31,120,30,103,31,106,31,101,31,6,31,6,30,79,31,111,31,99,31,63,31,63,30,25,31,77,31,77,30,128,31,128,30,186,31,166,31,53,31,53,30,137,31,125,31,125,30,237,31,78,31,148,31,148,30,244,31,167,31,42,31,235,31,126,31,70,31,56,31,233,31,237,31,132,31,132,30,132,29,246,31,173,31,53,31,53,30,189,31,108,31,161,31,241,31,238,31,76,31,181,31,77,31,249,31,195,31,195,30,54,31,155,31,87,31,45,31,204,31,233,31,233,30,105,31,175,31,154,31,154,30,179,31,126,31,126,30,59,31,21,31,125,31,108,31,117,31,229,31,163,31,163,30,63,31,63,30,18,31,18,30,80,31,134,31,80,31,198,31,250,31,235,31,132,31,39,31,63,31,250,31,11,31,11,30,10,31,63,31,211,31,200,31,115,31,143,31,198,31,198,30,179,31,249,31,197,31,41,31,126,31,189,31,189,30,189,29,241,31,237,31,150,31,178,31,178,30,178,29,202,31,195,31,241,31,200,31,196,31,196,30,196,29,162,31,220,31,124,31,65,31,60,31,126,31,89,31,230,31,230,30,16,31,16,30,90,31,89,31,210,31,210,30,170,31,74,31,71,31,71,30,117,31,108,31,73,31,255,31,35,31,112,31,112,30,171,31,215,31,45,31,57,31,57,30,61,31,38,31,177,31,235,31,129,31,49,31,221,31,194,31,199,31,127,31,10,31,78,31,78,30,183,31,218,31,154,31,207,31,250,31,166,31,250,31,132,31,252,31,60,31,60,30,248,31,222,31,238,31,238,30,73,31,188,31,188,30,45,31,211,31,250,31,121,31,242,31,129,31,186,31,146,31,23,31,59,31,94,31,50,31,32,31,35,31,9,31,135,31,135,30,135,29,133,31,133,30,164,31,164,30,105,31,38,31,38,30,58,31,137,31,170,31,170,30,78,31,196,31,85,31,85,30,116,31,116,30,4,31,4,30,78,31,185,31,185,30,185,29,211,31,89,31,222,31,222,30,185,31,185,30,12,31,48,31,57,31,56,31,56,30,52,31,160,31,133,31,236,31,159,31,4,31,4,30,86,31,86,30,70,31,162,31,189,31,90,31,32,31,127,31,140,31,69,31,235,31,188,31,57,31,57,30,138,31,138,30,108,31,84,31,84,30,84,29,16,31,11,31,53,31,24,31,23,31,213,31,213,30,31,31,253,31,138,31,134,31,87,31,51,31,51,30,51,29,109,31,109,30,149,31,164,31,187,31,67,31,67,30,161,31,77,31,15,31,214,31,214,30,214,29,214,28,225,31,212,31,241,31,241,30,112,31,71,31,117,31,223,31,133,31,133,30,81,31,166,31,48,31,140,31,140,30,182,31,253,31,28,31,29,31,68,31,68,30,115,31,143,31,17,31,25,31,27,31,27,30,27,29,253,31,253,30,71,31,91,31,189,31,189,30,243,31,177,31,2,31,2,30,89,31,89,30,166,31,18,31,138,31,188,31,243,31,149,31,80,31,80,30,67,31,62,31,150,31,150,30,249,31,249,30,104,31,100,31,153,31,78,31,181,31,229,31,229,30,123,31,66,31,213,31,17,31,125,31,39,31,118,31,20,31,189,31,189,30,157,31,157,30,157,29,75,31,253,31,253,30,238,31,145,31,145,30,102,31,102,30,89,31,244,31,244,30,242,31,242,30,97,31,180,31,180,30,250,31,250,30,227,31,24,31,85,31,115,31,126,31,175,31,232,31,211,31,211,30,103,31,57,31,208,31,208,30,63,31,191,31,197,31,204,31,204,30,114,31,135,31,135,30,225,31,39,31,39,31,8,31,168,31,239,31,161,31,88,31,146,31,87,31,107,31,205,31,150,31,5,31,5,30,198,31,165,31,140,31,5,31,124,31,32,31,109,31,109,30,67,31,67,30,114,31,199,31,208,31,64,31,64,30,64,29,162,31,161,31,161,30,161,29,170,31,200,31,200,30,206,31,206,30,144,31,50,31,229,31,205,31,216,31,216,30,17,31,241,31,174,31,174,30,254,31,241,31,170,31,184,31,77,31,15,31,32,31,237,31,237,30,136,31,240,31,237,31,237,30,132,31,245,31,245,30,245,29,98,31,125,31,170,31,79,31,178,31,73,31,73,30,70,31,70,30,158,31,106,31,235,31,189,31,129,31,146,31,67,31,188,31,253,31,253,30,103,31,40,31,40,30,40,29,70,31,225,31,49,31,148,31,148,30,169,31,91,31,37,31,37,30,163,31,163,30,129,31,220,31,220,30,163,31,111,31,65,31,244,31,222,31,104,31,122,31,198,31,243,31,76,31,242,31,242,30,114,31,129,31,79,31,79,30,71,31,99,31,99,30,99,29,172,31,172,30,229,31,66,31,66,30,80,31,160,31,153,31,228,31,19,31,19,30,220,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
