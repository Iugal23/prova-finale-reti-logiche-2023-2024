-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_126 is
end project_tb_126;

architecture project_tb_arch_126 of project_tb_126 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 791;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (163,0,24,0,151,0,0,0,0,0,25,0,120,0,233,0,223,0,118,0,174,0,209,0,0,0,91,0,70,0,43,0,0,0,224,0,0,0,144,0,178,0,0,0,0,0,16,0,194,0,128,0,12,0,159,0,254,0,165,0,55,0,204,0,95,0,163,0,63,0,201,0,0,0,97,0,183,0,133,0,231,0,15,0,0,0,0,0,197,0,0,0,42,0,60,0,82,0,0,0,236,0,198,0,180,0,58,0,140,0,76,0,10,0,14,0,87,0,183,0,170,0,0,0,0,0,0,0,242,0,19,0,92,0,171,0,115,0,246,0,49,0,0,0,148,0,13,0,159,0,89,0,0,0,0,0,17,0,180,0,0,0,130,0,64,0,0,0,33,0,0,0,44,0,254,0,184,0,0,0,98,0,182,0,152,0,98,0,77,0,0,0,0,0,0,0,150,0,0,0,56,0,158,0,198,0,158,0,224,0,69,0,45,0,99,0,7,0,0,0,0,0,0,0,67,0,0,0,142,0,97,0,37,0,167,0,184,0,106,0,169,0,186,0,14,0,211,0,177,0,163,0,227,0,0,0,209,0,168,0,0,0,110,0,180,0,179,0,192,0,95,0,163,0,0,0,107,0,2,0,3,0,0,0,252,0,0,0,7,0,53,0,0,0,117,0,191,0,119,0,0,0,6,0,160,0,252,0,0,0,30,0,28,0,90,0,217,0,244,0,22,0,229,0,222,0,5,0,0,0,197,0,61,0,0,0,0,0,0,0,181,0,0,0,93,0,156,0,47,0,94,0,137,0,138,0,0,0,10,0,105,0,0,0,0,0,249,0,185,0,111,0,130,0,110,0,107,0,0,0,0,0,0,0,219,0,108,0,160,0,127,0,220,0,3,0,17,0,20,0,202,0,151,0,56,0,75,0,102,0,219,0,0,0,0,0,166,0,229,0,16,0,82,0,210,0,104,0,13,0,67,0,112,0,253,0,155,0,117,0,88,0,177,0,17,0,18,0,245,0,205,0,0,0,141,0,0,0,58,0,0,0,214,0,44,0,31,0,108,0,241,0,14,0,100,0,110,0,137,0,0,0,114,0,0,0,215,0,5,0,1,0,139,0,0,0,195,0,21,0,227,0,76,0,63,0,0,0,0,0,227,0,104,0,199,0,39,0,0,0,77,0,0,0,97,0,141,0,208,0,226,0,32,0,158,0,229,0,0,0,2,0,183,0,217,0,173,0,162,0,49,0,27,0,201,0,30,0,0,0,169,0,233,0,157,0,82,0,0,0,157,0,8,0,87,0,204,0,74,0,234,0,0,0,250,0,0,0,145,0,53,0,197,0,22,0,66,0,198,0,18,0,211,0,61,0,0,0,192,0,0,0,0,0,44,0,143,0,56,0,0,0,54,0,0,0,200,0,0,0,231,0,0,0,39,0,191,0,0,0,76,0,209,0,56,0,152,0,186,0,42,0,198,0,192,0,64,0,22,0,193,0,0,0,107,0,189,0,203,0,150,0,0,0,221,0,131,0,196,0,66,0,159,0,0,0,76,0,128,0,75,0,187,0,233,0,254,0,162,0,127,0,171,0,60,0,133,0,142,0,0,0,42,0,201,0,43,0,94,0,203,0,0,0,156,0,54,0,148,0,180,0,213,0,201,0,109,0,0,0,184,0,61,0,33,0,175,0,35,0,80,0,251,0,0,0,82,0,122,0,167,0,64,0,142,0,155,0,34,0,155,0,158,0,0,0,0,0,95,0,29,0,107,0,246,0,175,0,0,0,68,0,128,0,76,0,76,0,142,0,59,0,0,0,111,0,106,0,65,0,138,0,2,0,43,0,143,0,0,0,2,0,39,0,218,0,180,0,87,0,221,0,2,0,0,0,223,0,205,0,227,0,190,0,59,0,199,0,27,0,54,0,18,0,246,0,0,0,166,0,167,0,48,0,165,0,0,0,155,0,22,0,7,0,216,0,0,0,137,0,151,0,38,0,0,0,89,0,249,0,0,0,12,0,197,0,21,0,0,0,136,0,0,0,0,0,145,0,77,0,68,0,143,0,133,0,0,0,211,0,59,0,0,0,232,0,224,0,126,0,163,0,0,0,29,0,134,0,9,0,179,0,134,0,42,0,164,0,0,0,29,0,0,0,76,0,249,0,232,0,205,0,252,0,0,0,0,0,81,0,81,0,25,0,233,0,108,0,88,0,253,0,158,0,233,0,0,0,0,0,72,0,108,0,0,0,0,0,174,0,69,0,0,0,19,0,0,0,160,0,214,0,88,0,168,0,213,0,180,0,13,0,212,0,0,0,96,0,43,0,23,0,149,0,33,0,165,0,193,0,178,0,0,0,0,0,0,0,64,0,167,0,75,0,12,0,228,0,195,0,80,0,197,0,0,0,219,0,9,0,208,0,146,0,44,0,0,0,17,0,160,0,136,0,61,0,132,0,54,0,94,0,0,0,161,0,0,0,215,0,97,0,0,0,13,0,0,0,33,0,0,0,37,0,58,0,76,0,219,0,6,0,0,0,81,0,180,0,0,0,211,0,166,0,188,0,24,0,104,0,0,0,0,0,252,0,85,0,170,0,0,0,213,0,100,0,0,0,244,0,102,0,56,0,196,0,132,0,254,0,0,0,34,0,212,0,46,0,119,0,244,0,224,0,0,0,0,0,176,0,58,0,185,0,118,0,57,0,150,0,255,0,17,0,0,0,3,0,205,0,36,0,186,0,0,0,154,0,214,0,133,0,16,0,47,0,185,0,161,0,0,0,203,0,75,0,219,0,189,0,64,0,169,0,249,0,125,0,0,0,0,0,31,0,0,0,22,0,169,0,219,0,133,0,118,0,141,0,0,0,78,0,8,0,187,0,248,0,64,0,161,0,23,0,109,0,170,0,65,0,0,0,31,0,57,0,19,0,111,0,123,0,251,0,171,0,24,0,197,0,218,0,46,0,117,0,59,0,0,0,0,0,203,0,0,0,251,0,208,0,161,0,36,0,123,0,245,0,0,0,172,0,243,0,97,0,114,0,0,0,246,0,66,0,18,0,3,0,0,0,165,0,127,0,87,0,195,0,0,0,41,0,214,0,238,0,0,0,175,0,221,0,0,0,159,0,79,0,56,0,0,0,0,0,45,0,0,0,144,0,20,0,0,0,97,0,115,0,139,0,0,0,18,0,137,0,233,0,254,0,255,0,139,0,43,0,120,0,190,0,19,0,139,0,123,0,46,0,103,0,150,0,8,0,39,0,0,0,0,0,77,0,119,0,184,0,147,0,84,0,0,0,22,0,61,0,0,0,148,0,216,0,0,0,76,0,117,0,134,0,0,0,0,0,43,0,71,0,73,0,0,0,240,0,0,0,154,0,203,0,47,0,119,0,148,0,0,0,129,0,24,0,214,0,115,0,129,0,25,0,0,0,0,0,125,0,231,0,100,0,99,0,153,0,120,0,0,0,56,0,17,0,249,0,37,0,9,0,148,0,182,0,194,0,150,0,136,0,38,0,0,0,0,0,181,0,150,0,88,0,20,0,17,0,124,0,253,0,38,0,0,0);
signal scenario_full  : scenario_type := (163,31,24,31,151,31,151,30,151,29,25,31,120,31,233,31,223,31,118,31,174,31,209,31,209,30,91,31,70,31,43,31,43,30,224,31,224,30,144,31,178,31,178,30,178,29,16,31,194,31,128,31,12,31,159,31,254,31,165,31,55,31,204,31,95,31,163,31,63,31,201,31,201,30,97,31,183,31,133,31,231,31,15,31,15,30,15,29,197,31,197,30,42,31,60,31,82,31,82,30,236,31,198,31,180,31,58,31,140,31,76,31,10,31,14,31,87,31,183,31,170,31,170,30,170,29,170,28,242,31,19,31,92,31,171,31,115,31,246,31,49,31,49,30,148,31,13,31,159,31,89,31,89,30,89,29,17,31,180,31,180,30,130,31,64,31,64,30,33,31,33,30,44,31,254,31,184,31,184,30,98,31,182,31,152,31,98,31,77,31,77,30,77,29,77,28,150,31,150,30,56,31,158,31,198,31,158,31,224,31,69,31,45,31,99,31,7,31,7,30,7,29,7,28,67,31,67,30,142,31,97,31,37,31,167,31,184,31,106,31,169,31,186,31,14,31,211,31,177,31,163,31,227,31,227,30,209,31,168,31,168,30,110,31,180,31,179,31,192,31,95,31,163,31,163,30,107,31,2,31,3,31,3,30,252,31,252,30,7,31,53,31,53,30,117,31,191,31,119,31,119,30,6,31,160,31,252,31,252,30,30,31,28,31,90,31,217,31,244,31,22,31,229,31,222,31,5,31,5,30,197,31,61,31,61,30,61,29,61,28,181,31,181,30,93,31,156,31,47,31,94,31,137,31,138,31,138,30,10,31,105,31,105,30,105,29,249,31,185,31,111,31,130,31,110,31,107,31,107,30,107,29,107,28,219,31,108,31,160,31,127,31,220,31,3,31,17,31,20,31,202,31,151,31,56,31,75,31,102,31,219,31,219,30,219,29,166,31,229,31,16,31,82,31,210,31,104,31,13,31,67,31,112,31,253,31,155,31,117,31,88,31,177,31,17,31,18,31,245,31,205,31,205,30,141,31,141,30,58,31,58,30,214,31,44,31,31,31,108,31,241,31,14,31,100,31,110,31,137,31,137,30,114,31,114,30,215,31,5,31,1,31,139,31,139,30,195,31,21,31,227,31,76,31,63,31,63,30,63,29,227,31,104,31,199,31,39,31,39,30,77,31,77,30,97,31,141,31,208,31,226,31,32,31,158,31,229,31,229,30,2,31,183,31,217,31,173,31,162,31,49,31,27,31,201,31,30,31,30,30,169,31,233,31,157,31,82,31,82,30,157,31,8,31,87,31,204,31,74,31,234,31,234,30,250,31,250,30,145,31,53,31,197,31,22,31,66,31,198,31,18,31,211,31,61,31,61,30,192,31,192,30,192,29,44,31,143,31,56,31,56,30,54,31,54,30,200,31,200,30,231,31,231,30,39,31,191,31,191,30,76,31,209,31,56,31,152,31,186,31,42,31,198,31,192,31,64,31,22,31,193,31,193,30,107,31,189,31,203,31,150,31,150,30,221,31,131,31,196,31,66,31,159,31,159,30,76,31,128,31,75,31,187,31,233,31,254,31,162,31,127,31,171,31,60,31,133,31,142,31,142,30,42,31,201,31,43,31,94,31,203,31,203,30,156,31,54,31,148,31,180,31,213,31,201,31,109,31,109,30,184,31,61,31,33,31,175,31,35,31,80,31,251,31,251,30,82,31,122,31,167,31,64,31,142,31,155,31,34,31,155,31,158,31,158,30,158,29,95,31,29,31,107,31,246,31,175,31,175,30,68,31,128,31,76,31,76,31,142,31,59,31,59,30,111,31,106,31,65,31,138,31,2,31,43,31,143,31,143,30,2,31,39,31,218,31,180,31,87,31,221,31,2,31,2,30,223,31,205,31,227,31,190,31,59,31,199,31,27,31,54,31,18,31,246,31,246,30,166,31,167,31,48,31,165,31,165,30,155,31,22,31,7,31,216,31,216,30,137,31,151,31,38,31,38,30,89,31,249,31,249,30,12,31,197,31,21,31,21,30,136,31,136,30,136,29,145,31,77,31,68,31,143,31,133,31,133,30,211,31,59,31,59,30,232,31,224,31,126,31,163,31,163,30,29,31,134,31,9,31,179,31,134,31,42,31,164,31,164,30,29,31,29,30,76,31,249,31,232,31,205,31,252,31,252,30,252,29,81,31,81,31,25,31,233,31,108,31,88,31,253,31,158,31,233,31,233,30,233,29,72,31,108,31,108,30,108,29,174,31,69,31,69,30,19,31,19,30,160,31,214,31,88,31,168,31,213,31,180,31,13,31,212,31,212,30,96,31,43,31,23,31,149,31,33,31,165,31,193,31,178,31,178,30,178,29,178,28,64,31,167,31,75,31,12,31,228,31,195,31,80,31,197,31,197,30,219,31,9,31,208,31,146,31,44,31,44,30,17,31,160,31,136,31,61,31,132,31,54,31,94,31,94,30,161,31,161,30,215,31,97,31,97,30,13,31,13,30,33,31,33,30,37,31,58,31,76,31,219,31,6,31,6,30,81,31,180,31,180,30,211,31,166,31,188,31,24,31,104,31,104,30,104,29,252,31,85,31,170,31,170,30,213,31,100,31,100,30,244,31,102,31,56,31,196,31,132,31,254,31,254,30,34,31,212,31,46,31,119,31,244,31,224,31,224,30,224,29,176,31,58,31,185,31,118,31,57,31,150,31,255,31,17,31,17,30,3,31,205,31,36,31,186,31,186,30,154,31,214,31,133,31,16,31,47,31,185,31,161,31,161,30,203,31,75,31,219,31,189,31,64,31,169,31,249,31,125,31,125,30,125,29,31,31,31,30,22,31,169,31,219,31,133,31,118,31,141,31,141,30,78,31,8,31,187,31,248,31,64,31,161,31,23,31,109,31,170,31,65,31,65,30,31,31,57,31,19,31,111,31,123,31,251,31,171,31,24,31,197,31,218,31,46,31,117,31,59,31,59,30,59,29,203,31,203,30,251,31,208,31,161,31,36,31,123,31,245,31,245,30,172,31,243,31,97,31,114,31,114,30,246,31,66,31,18,31,3,31,3,30,165,31,127,31,87,31,195,31,195,30,41,31,214,31,238,31,238,30,175,31,221,31,221,30,159,31,79,31,56,31,56,30,56,29,45,31,45,30,144,31,20,31,20,30,97,31,115,31,139,31,139,30,18,31,137,31,233,31,254,31,255,31,139,31,43,31,120,31,190,31,19,31,139,31,123,31,46,31,103,31,150,31,8,31,39,31,39,30,39,29,77,31,119,31,184,31,147,31,84,31,84,30,22,31,61,31,61,30,148,31,216,31,216,30,76,31,117,31,134,31,134,30,134,29,43,31,71,31,73,31,73,30,240,31,240,30,154,31,203,31,47,31,119,31,148,31,148,30,129,31,24,31,214,31,115,31,129,31,25,31,25,30,25,29,125,31,231,31,100,31,99,31,153,31,120,31,120,30,56,31,17,31,249,31,37,31,9,31,148,31,182,31,194,31,150,31,136,31,38,31,38,30,38,29,181,31,150,31,88,31,20,31,17,31,124,31,253,31,38,31,38,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
