-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 921;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,0,0,69,0,164,0,193,0,116,0,82,0,128,0,186,0,0,0,240,0,39,0,76,0,227,0,255,0,77,0,63,0,199,0,180,0,99,0,160,0,90,0,246,0,58,0,68,0,212,0,97,0,137,0,0,0,121,0,35,0,0,0,121,0,38,0,111,0,120,0,222,0,200,0,181,0,98,0,0,0,0,0,180,0,0,0,0,0,0,0,56,0,128,0,122,0,61,0,69,0,0,0,74,0,222,0,229,0,0,0,13,0,110,0,218,0,23,0,194,0,5,0,0,0,0,0,0,0,204,0,217,0,0,0,102,0,83,0,185,0,34,0,11,0,109,0,0,0,50,0,0,0,224,0,84,0,26,0,113,0,159,0,0,0,224,0,239,0,54,0,75,0,0,0,0,0,0,0,235,0,94,0,0,0,251,0,126,0,30,0,19,0,203,0,191,0,139,0,154,0,52,0,64,0,69,0,0,0,227,0,86,0,177,0,185,0,51,0,181,0,54,0,1,0,1,0,79,0,0,0,93,0,178,0,170,0,63,0,113,0,0,0,231,0,59,0,130,0,116,0,0,0,169,0,95,0,18,0,253,0,0,0,197,0,11,0,51,0,0,0,92,0,132,0,150,0,157,0,186,0,0,0,0,0,212,0,241,0,39,0,128,0,99,0,0,0,2,0,7,0,95,0,29,0,121,0,0,0,249,0,130,0,86,0,0,0,41,0,89,0,148,0,254,0,148,0,46,0,0,0,180,0,228,0,191,0,239,0,226,0,0,0,0,0,83,0,0,0,87,0,73,0,159,0,60,0,0,0,246,0,108,0,0,0,184,0,56,0,3,0,212,0,67,0,162,0,229,0,0,0,0,0,0,0,0,0,100,0,10,0,123,0,106,0,99,0,43,0,110,0,250,0,90,0,151,0,234,0,46,0,54,0,0,0,66,0,95,0,221,0,94,0,0,0,0,0,0,0,81,0,221,0,216,0,0,0,200,0,215,0,12,0,0,0,0,0,0,0,212,0,18,0,0,0,0,0,225,0,0,0,0,0,138,0,244,0,10,0,20,0,0,0,127,0,203,0,30,0,21,0,0,0,254,0,205,0,0,0,173,0,81,0,50,0,0,0,100,0,162,0,0,0,122,0,4,0,131,0,219,0,0,0,150,0,228,0,0,0,19,0,0,0,60,0,18,0,0,0,0,0,0,0,37,0,23,0,7,0,19,0,110,0,32,0,245,0,194,0,180,0,121,0,137,0,198,0,0,0,174,0,0,0,160,0,83,0,55,0,0,0,222,0,187,0,203,0,219,0,196,0,0,0,0,0,249,0,0,0,65,0,0,0,27,0,0,0,0,0,0,0,14,0,210,0,0,0,100,0,0,0,38,0,121,0,42,0,101,0,0,0,88,0,253,0,142,0,186,0,147,0,59,0,0,0,127,0,0,0,0,0,158,0,0,0,0,0,95,0,198,0,90,0,0,0,84,0,0,0,10,0,194,0,104,0,0,0,197,0,216,0,124,0,169,0,0,0,125,0,49,0,145,0,0,0,64,0,0,0,59,0,231,0,221,0,137,0,252,0,129,0,211,0,116,0,235,0,104,0,99,0,40,0,215,0,12,0,0,0,209,0,162,0,0,0,0,0,142,0,61,0,0,0,0,0,15,0,186,0,67,0,66,0,0,0,46,0,174,0,210,0,0,0,54,0,140,0,80,0,70,0,30,0,117,0,0,0,216,0,162,0,50,0,0,0,246,0,136,0,158,0,173,0,215,0,57,0,134,0,0,0,40,0,113,0,83,0,0,0,0,0,218,0,52,0,199,0,254,0,24,0,92,0,0,0,126,0,0,0,86,0,149,0,241,0,20,0,32,0,177,0,146,0,230,0,25,0,5,0,178,0,163,0,6,0,53,0,191,0,0,0,186,0,0,0,0,0,231,0,98,0,122,0,0,0,255,0,212,0,0,0,0,0,230,0,62,0,0,0,171,0,228,0,151,0,151,0,180,0,75,0,204,0,134,0,75,0,201,0,98,0,148,0,39,0,0,0,123,0,61,0,155,0,108,0,42,0,148,0,0,0,108,0,172,0,113,0,127,0,122,0,0,0,91,0,0,0,0,0,168,0,165,0,65,0,219,0,253,0,105,0,0,0,56,0,8,0,235,0,6,0,0,0,68,0,98,0,201,0,13,0,4,0,198,0,58,0,100,0,0,0,131,0,0,0,31,0,79,0,74,0,110,0,57,0,0,0,142,0,0,0,62,0,95,0,65,0,115,0,58,0,241,0,0,0,157,0,208,0,26,0,225,0,230,0,135,0,0,0,184,0,106,0,0,0,0,0,83,0,106,0,0,0,0,0,20,0,147,0,10,0,120,0,142,0,74,0,189,0,178,0,3,0,39,0,0,0,150,0,126,0,68,0,6,0,0,0,144,0,115,0,170,0,187,0,10,0,0,0,58,0,116,0,112,0,0,0,171,0,242,0,230,0,55,0,143,0,185,0,0,0,4,0,40,0,169,0,33,0,119,0,5,0,0,0,0,0,86,0,0,0,17,0,92,0,187,0,0,0,0,0,96,0,170,0,0,0,246,0,241,0,0,0,161,0,166,0,0,0,0,0,172,0,100,0,183,0,2,0,184,0,0,0,221,0,68,0,252,0,0,0,255,0,174,0,89,0,234,0,183,0,83,0,0,0,93,0,196,0,26,0,142,0,50,0,163,0,208,0,189,0,207,0,99,0,144,0,120,0,0,0,14,0,110,0,89,0,122,0,22,0,0,0,210,0,241,0,0,0,173,0,0,0,8,0,131,0,145,0,235,0,226,0,232,0,0,0,72,0,167,0,141,0,215,0,57,0,19,0,0,0,75,0,253,0,169,0,221,0,0,0,72,0,129,0,0,0,26,0,100,0,168,0,251,0,0,0,0,0,0,0,0,0,0,0,169,0,0,0,0,0,184,0,128,0,150,0,156,0,92,0,201,0,125,0,91,0,111,0,0,0,76,0,138,0,0,0,116,0,214,0,225,0,248,0,90,0,241,0,221,0,87,0,123,0,218,0,74,0,88,0,168,0,0,0,226,0,150,0,230,0,204,0,161,0,0,0,68,0,223,0,154,0,76,0,12,0,0,0,116,0,246,0,104,0,134,0,20,0,11,0,0,0,29,0,168,0,0,0,0,0,145,0,1,0,183,0,140,0,0,0,153,0,62,0,252,0,5,0,132,0,216,0,85,0,123,0,76,0,33,0,64,0,23,0,26,0,103,0,209,0,0,0,40,0,122,0,0,0,178,0,183,0,131,0,52,0,226,0,0,0,246,0,91,0,217,0,0,0,152,0,237,0,0,0,3,0,134,0,207,0,239,0,153,0,115,0,0,0,112,0,3,0,72,0,197,0,162,0,93,0,0,0,213,0,206,0,6,0,0,0,188,0,46,0,17,0,167,0,61,0,171,0,118,0,0,0,199,0,126,0,211,0,102,0,0,0,226,0,0,0,77,0,15,0,206,0,14,0,252,0,87,0,59,0,0,0,0,0,147,0,223,0,11,0,0,0,207,0,1,0,52,0,0,0,0,0,28,0,161,0,238,0,0,0,165,0,241,0,77,0,38,0,195,0,142,0,158,0,124,0,0,0,9,0,0,0,36,0,28,0,141,0,0,0,0,0,204,0,0,0,73,0,104,0,0,0,0,0,32,0,250,0,186,0,38,0,240,0,216,0,68,0,174,0,110,0,125,0,233,0,114,0,34,0,221,0,0,0,252,0,127,0,155,0,0,0,137,0,68,0,158,0,10,0,153,0,94,0,0,0,237,0,231,0,215,0,112,0,16,0,117,0,0,0,98,0,191,0,0,0,159,0,236,0,0,0,208,0,0,0,0,0,143,0,117,0,117,0,0,0,0,0,91,0,238,0,29,0,138,0,198,0,84,0,130,0,0,0,219,0,71,0,52,0,66,0,141,0,181,0,150,0,134,0,0,0,198,0,0,0,65,0,113,0,74,0,219,0,105,0,0,0,0,0,173,0,0,0,0,0,41,0,91,0,14,0,0,0,0,0,128,0,126,0,0,0,192,0,70,0,170,0,202,0,160,0,225,0,45,0,0,0,209,0,246,0,0,0,115,0,60,0,0,0,229,0,0,0,0,0);
signal scenario_full  : scenario_type := (201,31,201,30,69,31,164,31,193,31,116,31,82,31,128,31,186,31,186,30,240,31,39,31,76,31,227,31,255,31,77,31,63,31,199,31,180,31,99,31,160,31,90,31,246,31,58,31,68,31,212,31,97,31,137,31,137,30,121,31,35,31,35,30,121,31,38,31,111,31,120,31,222,31,200,31,181,31,98,31,98,30,98,29,180,31,180,30,180,29,180,28,56,31,128,31,122,31,61,31,69,31,69,30,74,31,222,31,229,31,229,30,13,31,110,31,218,31,23,31,194,31,5,31,5,30,5,29,5,28,204,31,217,31,217,30,102,31,83,31,185,31,34,31,11,31,109,31,109,30,50,31,50,30,224,31,84,31,26,31,113,31,159,31,159,30,224,31,239,31,54,31,75,31,75,30,75,29,75,28,235,31,94,31,94,30,251,31,126,31,30,31,19,31,203,31,191,31,139,31,154,31,52,31,64,31,69,31,69,30,227,31,86,31,177,31,185,31,51,31,181,31,54,31,1,31,1,31,79,31,79,30,93,31,178,31,170,31,63,31,113,31,113,30,231,31,59,31,130,31,116,31,116,30,169,31,95,31,18,31,253,31,253,30,197,31,11,31,51,31,51,30,92,31,132,31,150,31,157,31,186,31,186,30,186,29,212,31,241,31,39,31,128,31,99,31,99,30,2,31,7,31,95,31,29,31,121,31,121,30,249,31,130,31,86,31,86,30,41,31,89,31,148,31,254,31,148,31,46,31,46,30,180,31,228,31,191,31,239,31,226,31,226,30,226,29,83,31,83,30,87,31,73,31,159,31,60,31,60,30,246,31,108,31,108,30,184,31,56,31,3,31,212,31,67,31,162,31,229,31,229,30,229,29,229,28,229,27,100,31,10,31,123,31,106,31,99,31,43,31,110,31,250,31,90,31,151,31,234,31,46,31,54,31,54,30,66,31,95,31,221,31,94,31,94,30,94,29,94,28,81,31,221,31,216,31,216,30,200,31,215,31,12,31,12,30,12,29,12,28,212,31,18,31,18,30,18,29,225,31,225,30,225,29,138,31,244,31,10,31,20,31,20,30,127,31,203,31,30,31,21,31,21,30,254,31,205,31,205,30,173,31,81,31,50,31,50,30,100,31,162,31,162,30,122,31,4,31,131,31,219,31,219,30,150,31,228,31,228,30,19,31,19,30,60,31,18,31,18,30,18,29,18,28,37,31,23,31,7,31,19,31,110,31,32,31,245,31,194,31,180,31,121,31,137,31,198,31,198,30,174,31,174,30,160,31,83,31,55,31,55,30,222,31,187,31,203,31,219,31,196,31,196,30,196,29,249,31,249,30,65,31,65,30,27,31,27,30,27,29,27,28,14,31,210,31,210,30,100,31,100,30,38,31,121,31,42,31,101,31,101,30,88,31,253,31,142,31,186,31,147,31,59,31,59,30,127,31,127,30,127,29,158,31,158,30,158,29,95,31,198,31,90,31,90,30,84,31,84,30,10,31,194,31,104,31,104,30,197,31,216,31,124,31,169,31,169,30,125,31,49,31,145,31,145,30,64,31,64,30,59,31,231,31,221,31,137,31,252,31,129,31,211,31,116,31,235,31,104,31,99,31,40,31,215,31,12,31,12,30,209,31,162,31,162,30,162,29,142,31,61,31,61,30,61,29,15,31,186,31,67,31,66,31,66,30,46,31,174,31,210,31,210,30,54,31,140,31,80,31,70,31,30,31,117,31,117,30,216,31,162,31,50,31,50,30,246,31,136,31,158,31,173,31,215,31,57,31,134,31,134,30,40,31,113,31,83,31,83,30,83,29,218,31,52,31,199,31,254,31,24,31,92,31,92,30,126,31,126,30,86,31,149,31,241,31,20,31,32,31,177,31,146,31,230,31,25,31,5,31,178,31,163,31,6,31,53,31,191,31,191,30,186,31,186,30,186,29,231,31,98,31,122,31,122,30,255,31,212,31,212,30,212,29,230,31,62,31,62,30,171,31,228,31,151,31,151,31,180,31,75,31,204,31,134,31,75,31,201,31,98,31,148,31,39,31,39,30,123,31,61,31,155,31,108,31,42,31,148,31,148,30,108,31,172,31,113,31,127,31,122,31,122,30,91,31,91,30,91,29,168,31,165,31,65,31,219,31,253,31,105,31,105,30,56,31,8,31,235,31,6,31,6,30,68,31,98,31,201,31,13,31,4,31,198,31,58,31,100,31,100,30,131,31,131,30,31,31,79,31,74,31,110,31,57,31,57,30,142,31,142,30,62,31,95,31,65,31,115,31,58,31,241,31,241,30,157,31,208,31,26,31,225,31,230,31,135,31,135,30,184,31,106,31,106,30,106,29,83,31,106,31,106,30,106,29,20,31,147,31,10,31,120,31,142,31,74,31,189,31,178,31,3,31,39,31,39,30,150,31,126,31,68,31,6,31,6,30,144,31,115,31,170,31,187,31,10,31,10,30,58,31,116,31,112,31,112,30,171,31,242,31,230,31,55,31,143,31,185,31,185,30,4,31,40,31,169,31,33,31,119,31,5,31,5,30,5,29,86,31,86,30,17,31,92,31,187,31,187,30,187,29,96,31,170,31,170,30,246,31,241,31,241,30,161,31,166,31,166,30,166,29,172,31,100,31,183,31,2,31,184,31,184,30,221,31,68,31,252,31,252,30,255,31,174,31,89,31,234,31,183,31,83,31,83,30,93,31,196,31,26,31,142,31,50,31,163,31,208,31,189,31,207,31,99,31,144,31,120,31,120,30,14,31,110,31,89,31,122,31,22,31,22,30,210,31,241,31,241,30,173,31,173,30,8,31,131,31,145,31,235,31,226,31,232,31,232,30,72,31,167,31,141,31,215,31,57,31,19,31,19,30,75,31,253,31,169,31,221,31,221,30,72,31,129,31,129,30,26,31,100,31,168,31,251,31,251,30,251,29,251,28,251,27,251,26,169,31,169,30,169,29,184,31,128,31,150,31,156,31,92,31,201,31,125,31,91,31,111,31,111,30,76,31,138,31,138,30,116,31,214,31,225,31,248,31,90,31,241,31,221,31,87,31,123,31,218,31,74,31,88,31,168,31,168,30,226,31,150,31,230,31,204,31,161,31,161,30,68,31,223,31,154,31,76,31,12,31,12,30,116,31,246,31,104,31,134,31,20,31,11,31,11,30,29,31,168,31,168,30,168,29,145,31,1,31,183,31,140,31,140,30,153,31,62,31,252,31,5,31,132,31,216,31,85,31,123,31,76,31,33,31,64,31,23,31,26,31,103,31,209,31,209,30,40,31,122,31,122,30,178,31,183,31,131,31,52,31,226,31,226,30,246,31,91,31,217,31,217,30,152,31,237,31,237,30,3,31,134,31,207,31,239,31,153,31,115,31,115,30,112,31,3,31,72,31,197,31,162,31,93,31,93,30,213,31,206,31,6,31,6,30,188,31,46,31,17,31,167,31,61,31,171,31,118,31,118,30,199,31,126,31,211,31,102,31,102,30,226,31,226,30,77,31,15,31,206,31,14,31,252,31,87,31,59,31,59,30,59,29,147,31,223,31,11,31,11,30,207,31,1,31,52,31,52,30,52,29,28,31,161,31,238,31,238,30,165,31,241,31,77,31,38,31,195,31,142,31,158,31,124,31,124,30,9,31,9,30,36,31,28,31,141,31,141,30,141,29,204,31,204,30,73,31,104,31,104,30,104,29,32,31,250,31,186,31,38,31,240,31,216,31,68,31,174,31,110,31,125,31,233,31,114,31,34,31,221,31,221,30,252,31,127,31,155,31,155,30,137,31,68,31,158,31,10,31,153,31,94,31,94,30,237,31,231,31,215,31,112,31,16,31,117,31,117,30,98,31,191,31,191,30,159,31,236,31,236,30,208,31,208,30,208,29,143,31,117,31,117,31,117,30,117,29,91,31,238,31,29,31,138,31,198,31,84,31,130,31,130,30,219,31,71,31,52,31,66,31,141,31,181,31,150,31,134,31,134,30,198,31,198,30,65,31,113,31,74,31,219,31,105,31,105,30,105,29,173,31,173,30,173,29,41,31,91,31,14,31,14,30,14,29,128,31,126,31,126,30,192,31,70,31,170,31,202,31,160,31,225,31,45,31,45,30,209,31,246,31,246,30,115,31,60,31,60,30,229,31,229,30,229,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
