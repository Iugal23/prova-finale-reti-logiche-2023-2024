-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 295;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,33,0,182,0,90,0,163,0,0,0,0,0,0,0,177,0,0,0,190,0,185,0,111,0,134,0,96,0,81,0,0,0,148,0,124,0,193,0,232,0,197,0,208,0,105,0,197,0,221,0,114,0,218,0,235,0,0,0,175,0,126,0,85,0,1,0,177,0,0,0,0,0,218,0,39,0,36,0,143,0,0,0,162,0,176,0,11,0,123,0,243,0,145,0,201,0,0,0,157,0,103,0,0,0,64,0,125,0,190,0,4,0,43,0,7,0,241,0,0,0,194,0,144,0,183,0,223,0,24,0,80,0,0,0,219,0,195,0,73,0,226,0,0,0,26,0,74,0,0,0,14,0,46,0,14,0,216,0,0,0,239,0,110,0,138,0,141,0,41,0,194,0,114,0,113,0,150,0,113,0,110,0,0,0,0,0,178,0,189,0,215,0,192,0,241,0,31,0,38,0,65,0,116,0,185,0,172,0,93,0,0,0,70,0,104,0,146,0,245,0,82,0,0,0,254,0,0,0,18,0,51,0,33,0,209,0,88,0,168,0,105,0,0,0,0,0,146,0,145,0,153,0,0,0,207,0,48,0,225,0,44,0,63,0,188,0,51,0,48,0,186,0,16,0,119,0,0,0,28,0,23,0,34,0,0,0,10,0,52,0,157,0,0,0,0,0,10,0,208,0,1,0,20,0,128,0,133,0,0,0,0,0,187,0,0,0,0,0,0,0,245,0,204,0,147,0,166,0,189,0,109,0,133,0,84,0,0,0,240,0,0,0,12,0,219,0,98,0,0,0,61,0,243,0,245,0,56,0,130,0,0,0,160,0,151,0,191,0,0,0,0,0,106,0,208,0,74,0,254,0,5,0,77,0,0,0,0,0,47,0,126,0,27,0,9,0,0,0,156,0,230,0,166,0,124,0,0,0,0,0,0,0,169,0,2,0,0,0,55,0,21,0,78,0,247,0,104,0,50,0,202,0,0,0,105,0,188,0,150,0,223,0,0,0,0,0,21,0,17,0,130,0,121,0,0,0,93,0,0,0,231,0,193,0,0,0,137,0,52,0,23,0,116,0,159,0,200,0,230,0,175,0,82,0,186,0,0,0,9,0,89,0,139,0,248,0,226,0,0,0,185,0,30,0,34,0,0,0,151,0,0,0,0,0,146,0,113,0,47,0,76,0,202,0,49,0,127,0,0,0,101,0,174,0,93,0,111,0,123,0,102,0,187,0,156,0,194,0,0,0,75,0,151,0,147,0,191,0,59,0,0,0,199,0,202,0,148,0,245,0,186,0,78,0,229,0,247,0,199,0,55,0,0,0,162,0,0,0);
signal scenario_full  : scenario_type := (0,0,33,31,182,31,90,31,163,31,163,30,163,29,163,28,177,31,177,30,190,31,185,31,111,31,134,31,96,31,81,31,81,30,148,31,124,31,193,31,232,31,197,31,208,31,105,31,197,31,221,31,114,31,218,31,235,31,235,30,175,31,126,31,85,31,1,31,177,31,177,30,177,29,218,31,39,31,36,31,143,31,143,30,162,31,176,31,11,31,123,31,243,31,145,31,201,31,201,30,157,31,103,31,103,30,64,31,125,31,190,31,4,31,43,31,7,31,241,31,241,30,194,31,144,31,183,31,223,31,24,31,80,31,80,30,219,31,195,31,73,31,226,31,226,30,26,31,74,31,74,30,14,31,46,31,14,31,216,31,216,30,239,31,110,31,138,31,141,31,41,31,194,31,114,31,113,31,150,31,113,31,110,31,110,30,110,29,178,31,189,31,215,31,192,31,241,31,31,31,38,31,65,31,116,31,185,31,172,31,93,31,93,30,70,31,104,31,146,31,245,31,82,31,82,30,254,31,254,30,18,31,51,31,33,31,209,31,88,31,168,31,105,31,105,30,105,29,146,31,145,31,153,31,153,30,207,31,48,31,225,31,44,31,63,31,188,31,51,31,48,31,186,31,16,31,119,31,119,30,28,31,23,31,34,31,34,30,10,31,52,31,157,31,157,30,157,29,10,31,208,31,1,31,20,31,128,31,133,31,133,30,133,29,187,31,187,30,187,29,187,28,245,31,204,31,147,31,166,31,189,31,109,31,133,31,84,31,84,30,240,31,240,30,12,31,219,31,98,31,98,30,61,31,243,31,245,31,56,31,130,31,130,30,160,31,151,31,191,31,191,30,191,29,106,31,208,31,74,31,254,31,5,31,77,31,77,30,77,29,47,31,126,31,27,31,9,31,9,30,156,31,230,31,166,31,124,31,124,30,124,29,124,28,169,31,2,31,2,30,55,31,21,31,78,31,247,31,104,31,50,31,202,31,202,30,105,31,188,31,150,31,223,31,223,30,223,29,21,31,17,31,130,31,121,31,121,30,93,31,93,30,231,31,193,31,193,30,137,31,52,31,23,31,116,31,159,31,200,31,230,31,175,31,82,31,186,31,186,30,9,31,89,31,139,31,248,31,226,31,226,30,185,31,30,31,34,31,34,30,151,31,151,30,151,29,146,31,113,31,47,31,76,31,202,31,49,31,127,31,127,30,101,31,174,31,93,31,111,31,123,31,102,31,187,31,156,31,194,31,194,30,75,31,151,31,147,31,191,31,59,31,59,30,199,31,202,31,148,31,245,31,186,31,78,31,229,31,247,31,199,31,55,31,55,30,162,31,162,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
