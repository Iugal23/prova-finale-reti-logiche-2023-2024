-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_204 is
end project_tb_204;

architecture project_tb_arch_204 of project_tb_204 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 932;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,71,0,225,0,54,0,154,0,0,0,197,0,172,0,6,0,208,0,0,0,93,0,0,0,57,0,150,0,230,0,189,0,83,0,199,0,225,0,24,0,0,0,0,0,7,0,142,0,39,0,150,0,80,0,236,0,177,0,99,0,64,0,0,0,145,0,0,0,136,0,0,0,197,0,0,0,226,0,108,0,112,0,101,0,72,0,209,0,0,0,0,0,244,0,57,0,0,0,202,0,181,0,10,0,196,0,18,0,0,0,85,0,0,0,232,0,0,0,136,0,242,0,117,0,66,0,169,0,41,0,80,0,119,0,0,0,217,0,236,0,161,0,0,0,0,0,230,0,212,0,231,0,125,0,247,0,114,0,192,0,94,0,0,0,214,0,235,0,246,0,0,0,32,0,170,0,130,0,158,0,210,0,97,0,80,0,191,0,9,0,0,0,201,0,171,0,52,0,99,0,239,0,160,0,67,0,8,0,158,0,0,0,168,0,114,0,68,0,51,0,213,0,0,0,71,0,47,0,10,0,85,0,141,0,164,0,181,0,180,0,143,0,0,0,2,0,186,0,159,0,204,0,222,0,220,0,2,0,216,0,228,0,0,0,191,0,125,0,248,0,0,0,0,0,10,0,34,0,82,0,0,0,151,0,207,0,245,0,1,0,180,0,38,0,0,0,140,0,0,0,182,0,35,0,121,0,53,0,27,0,227,0,0,0,0,0,0,0,28,0,0,0,12,0,6,0,223,0,210,0,129,0,196,0,86,0,183,0,31,0,0,0,161,0,127,0,120,0,1,0,208,0,195,0,7,0,120,0,62,0,126,0,144,0,0,0,0,0,0,0,46,0,200,0,239,0,38,0,109,0,111,0,127,0,59,0,0,0,0,0,192,0,153,0,19,0,240,0,99,0,189,0,75,0,159,0,0,0,0,0,48,0,0,0,0,0,0,0,247,0,206,0,125,0,170,0,107,0,89,0,30,0,43,0,0,0,123,0,64,0,186,0,66,0,223,0,195,0,76,0,187,0,74,0,0,0,219,0,202,0,54,0,0,0,47,0,117,0,159,0,223,0,230,0,249,0,0,0,0,0,145,0,143,0,55,0,0,0,0,0,0,0,123,0,122,0,23,0,87,0,102,0,163,0,175,0,246,0,188,0,0,0,27,0,216,0,117,0,99,0,13,0,165,0,238,0,22,0,107,0,126,0,91,0,0,0,199,0,230,0,177,0,30,0,29,0,53,0,0,0,99,0,0,0,146,0,143,0,56,0,67,0,147,0,60,0,35,0,43,0,16,0,250,0,0,0,88,0,157,0,184,0,0,0,0,0,0,0,94,0,136,0,121,0,184,0,68,0,140,0,50,0,54,0,0,0,126,0,206,0,192,0,0,0,127,0,0,0,169,0,120,0,220,0,4,0,0,0,0,0,206,0,0,0,167,0,47,0,119,0,180,0,57,0,142,0,66,0,0,0,175,0,204,0,229,0,0,0,0,0,8,0,37,0,0,0,0,0,127,0,228,0,155,0,158,0,0,0,160,0,94,0,112,0,195,0,73,0,23,0,0,0,0,0,123,0,44,0,51,0,126,0,22,0,205,0,145,0,0,0,218,0,162,0,94,0,0,0,90,0,250,0,209,0,56,0,155,0,127,0,0,0,105,0,187,0,93,0,169,0,124,0,0,0,0,0,146,0,224,0,131,0,233,0,126,0,223,0,102,0,0,0,210,0,121,0,152,0,0,0,229,0,75,0,225,0,233,0,75,0,0,0,154,0,0,0,232,0,199,0,244,0,162,0,0,0,3,0,22,0,52,0,0,0,220,0,74,0,26,0,54,0,176,0,154,0,125,0,105,0,196,0,162,0,101,0,56,0,0,0,52,0,46,0,179,0,0,0,17,0,0,0,32,0,7,0,234,0,40,0,64,0,223,0,171,0,53,0,248,0,181,0,111,0,154,0,0,0,0,0,200,0,124,0,103,0,42,0,241,0,122,0,12,0,0,0,233,0,168,0,87,0,218,0,0,0,0,0,67,0,39,0,0,0,170,0,0,0,89,0,111,0,184,0,0,0,0,0,98,0,74,0,163,0,93,0,19,0,137,0,0,0,128,0,240,0,116,0,57,0,30,0,130,0,0,0,116,0,115,0,0,0,206,0,224,0,103,0,63,0,240,0,0,0,0,0,131,0,151,0,0,0,64,0,157,0,83,0,86,0,28,0,53,0,223,0,29,0,107,0,0,0,0,0,71,0,0,0,95,0,144,0,27,0,191,0,51,0,132,0,241,0,89,0,68,0,167,0,113,0,0,0,0,0,0,0,156,0,0,0,94,0,254,0,221,0,0,0,0,0,232,0,78,0,250,0,0,0,0,0,27,0,163,0,10,0,167,0,0,0,100,0,143,0,22,0,29,0,159,0,147,0,0,0,83,0,106,0,32,0,158,0,143,0,197,0,178,0,119,0,75,0,0,0,0,0,0,0,2,0,133,0,208,0,132,0,11,0,198,0,11,0,53,0,155,0,194,0,169,0,57,0,0,0,224,0,123,0,197,0,64,0,199,0,185,0,189,0,177,0,50,0,57,0,150,0,0,0,71,0,79,0,89,0,73,0,103,0,145,0,90,0,73,0,49,0,226,0,106,0,140,0,202,0,0,0,231,0,216,0,139,0,0,0,42,0,95,0,114,0,111,0,74,0,72,0,125,0,152,0,146,0,0,0,174,0,119,0,93,0,0,0,102,0,128,0,79,0,198,0,7,0,138,0,0,0,3,0,0,0,200,0,249,0,23,0,102,0,0,0,0,0,0,0,87,0,64,0,36,0,127,0,0,0,104,0,94,0,150,0,199,0,118,0,0,0,22,0,27,0,68,0,142,0,29,0,1,0,0,0,125,0,162,0,0,0,73,0,149,0,85,0,157,0,205,0,106,0,204,0,76,0,167,0,51,0,253,0,252,0,50,0,124,0,154,0,175,0,0,0,9,0,0,0,148,0,86,0,0,0,114,0,182,0,171,0,254,0,115,0,6,0,223,0,6,0,81,0,52,0,0,0,0,0,198,0,20,0,213,0,0,0,125,0,105,0,0,0,228,0,167,0,42,0,212,0,203,0,32,0,6,0,220,0,135,0,188,0,218,0,10,0,89,0,58,0,70,0,0,0,155,0,62,0,65,0,123,0,0,0,0,0,17,0,191,0,0,0,252,0,232,0,181,0,0,0,252,0,141,0,63,0,138,0,196,0,64,0,218,0,120,0,244,0,126,0,35,0,0,0,190,0,156,0,218,0,196,0,218,0,216,0,0,0,162,0,115,0,70,0,175,0,0,0,0,0,0,0,239,0,203,0,234,0,127,0,224,0,202,0,24,0,213,0,200,0,20,0,57,0,0,0,206,0,0,0,222,0,108,0,20,0,223,0,77,0,227,0,0,0,7,0,191,0,220,0,174,0,160,0,207,0,123,0,13,0,242,0,0,0,223,0,99,0,0,0,164,0,32,0,0,0,67,0,123,0,0,0,230,0,38,0,197,0,66,0,36,0,0,0,54,0,121,0,78,0,115,0,188,0,148,0,128,0,173,0,0,0,123,0,4,0,189,0,106,0,40,0,83,0,24,0,156,0,174,0,250,0,0,0,185,0,228,0,69,0,0,0,180,0,0,0,63,0,0,0,202,0,221,0,151,0,42,0,0,0,58,0,0,0,248,0,230,0,201,0,60,0,217,0,0,0,238,0,48,0,9,0,0,0,92,0,23,0,122,0,70,0,174,0,252,0,177,0,1,0,0,0,0,0,0,0,101,0,0,0,0,0,116,0,186,0,174,0,239,0,224,0,106,0,175,0,0,0,80,0,62,0,56,0,1,0,6,0,0,0,35,0,200,0,46,0,142,0,0,0,0,0,183,0,0,0,141,0,211,0,0,0,24,0,94,0,185,0,0,0,68,0,236,0,190,0,195,0,0,0,192,0,216,0,186,0,229,0,240,0,72,0,53,0,0,0,0,0,214,0,5,0,175,0,58,0,0,0,0,0,125,0,209,0,0,0,0,0,0,0,0,0,68,0,168,0,38,0,175,0,118,0,227,0,39,0,54,0,142,0,0,0,98,0,23,0,143,0,104,0,66,0,80,0,150,0,250,0,21,0,177,0,24,0,176,0,101,0,31,0,209,0,0,0,61,0,54,0,147,0,99,0,32,0,249,0);
signal scenario_full  : scenario_type := (49,31,71,31,225,31,54,31,154,31,154,30,197,31,172,31,6,31,208,31,208,30,93,31,93,30,57,31,150,31,230,31,189,31,83,31,199,31,225,31,24,31,24,30,24,29,7,31,142,31,39,31,150,31,80,31,236,31,177,31,99,31,64,31,64,30,145,31,145,30,136,31,136,30,197,31,197,30,226,31,108,31,112,31,101,31,72,31,209,31,209,30,209,29,244,31,57,31,57,30,202,31,181,31,10,31,196,31,18,31,18,30,85,31,85,30,232,31,232,30,136,31,242,31,117,31,66,31,169,31,41,31,80,31,119,31,119,30,217,31,236,31,161,31,161,30,161,29,230,31,212,31,231,31,125,31,247,31,114,31,192,31,94,31,94,30,214,31,235,31,246,31,246,30,32,31,170,31,130,31,158,31,210,31,97,31,80,31,191,31,9,31,9,30,201,31,171,31,52,31,99,31,239,31,160,31,67,31,8,31,158,31,158,30,168,31,114,31,68,31,51,31,213,31,213,30,71,31,47,31,10,31,85,31,141,31,164,31,181,31,180,31,143,31,143,30,2,31,186,31,159,31,204,31,222,31,220,31,2,31,216,31,228,31,228,30,191,31,125,31,248,31,248,30,248,29,10,31,34,31,82,31,82,30,151,31,207,31,245,31,1,31,180,31,38,31,38,30,140,31,140,30,182,31,35,31,121,31,53,31,27,31,227,31,227,30,227,29,227,28,28,31,28,30,12,31,6,31,223,31,210,31,129,31,196,31,86,31,183,31,31,31,31,30,161,31,127,31,120,31,1,31,208,31,195,31,7,31,120,31,62,31,126,31,144,31,144,30,144,29,144,28,46,31,200,31,239,31,38,31,109,31,111,31,127,31,59,31,59,30,59,29,192,31,153,31,19,31,240,31,99,31,189,31,75,31,159,31,159,30,159,29,48,31,48,30,48,29,48,28,247,31,206,31,125,31,170,31,107,31,89,31,30,31,43,31,43,30,123,31,64,31,186,31,66,31,223,31,195,31,76,31,187,31,74,31,74,30,219,31,202,31,54,31,54,30,47,31,117,31,159,31,223,31,230,31,249,31,249,30,249,29,145,31,143,31,55,31,55,30,55,29,55,28,123,31,122,31,23,31,87,31,102,31,163,31,175,31,246,31,188,31,188,30,27,31,216,31,117,31,99,31,13,31,165,31,238,31,22,31,107,31,126,31,91,31,91,30,199,31,230,31,177,31,30,31,29,31,53,31,53,30,99,31,99,30,146,31,143,31,56,31,67,31,147,31,60,31,35,31,43,31,16,31,250,31,250,30,88,31,157,31,184,31,184,30,184,29,184,28,94,31,136,31,121,31,184,31,68,31,140,31,50,31,54,31,54,30,126,31,206,31,192,31,192,30,127,31,127,30,169,31,120,31,220,31,4,31,4,30,4,29,206,31,206,30,167,31,47,31,119,31,180,31,57,31,142,31,66,31,66,30,175,31,204,31,229,31,229,30,229,29,8,31,37,31,37,30,37,29,127,31,228,31,155,31,158,31,158,30,160,31,94,31,112,31,195,31,73,31,23,31,23,30,23,29,123,31,44,31,51,31,126,31,22,31,205,31,145,31,145,30,218,31,162,31,94,31,94,30,90,31,250,31,209,31,56,31,155,31,127,31,127,30,105,31,187,31,93,31,169,31,124,31,124,30,124,29,146,31,224,31,131,31,233,31,126,31,223,31,102,31,102,30,210,31,121,31,152,31,152,30,229,31,75,31,225,31,233,31,75,31,75,30,154,31,154,30,232,31,199,31,244,31,162,31,162,30,3,31,22,31,52,31,52,30,220,31,74,31,26,31,54,31,176,31,154,31,125,31,105,31,196,31,162,31,101,31,56,31,56,30,52,31,46,31,179,31,179,30,17,31,17,30,32,31,7,31,234,31,40,31,64,31,223,31,171,31,53,31,248,31,181,31,111,31,154,31,154,30,154,29,200,31,124,31,103,31,42,31,241,31,122,31,12,31,12,30,233,31,168,31,87,31,218,31,218,30,218,29,67,31,39,31,39,30,170,31,170,30,89,31,111,31,184,31,184,30,184,29,98,31,74,31,163,31,93,31,19,31,137,31,137,30,128,31,240,31,116,31,57,31,30,31,130,31,130,30,116,31,115,31,115,30,206,31,224,31,103,31,63,31,240,31,240,30,240,29,131,31,151,31,151,30,64,31,157,31,83,31,86,31,28,31,53,31,223,31,29,31,107,31,107,30,107,29,71,31,71,30,95,31,144,31,27,31,191,31,51,31,132,31,241,31,89,31,68,31,167,31,113,31,113,30,113,29,113,28,156,31,156,30,94,31,254,31,221,31,221,30,221,29,232,31,78,31,250,31,250,30,250,29,27,31,163,31,10,31,167,31,167,30,100,31,143,31,22,31,29,31,159,31,147,31,147,30,83,31,106,31,32,31,158,31,143,31,197,31,178,31,119,31,75,31,75,30,75,29,75,28,2,31,133,31,208,31,132,31,11,31,198,31,11,31,53,31,155,31,194,31,169,31,57,31,57,30,224,31,123,31,197,31,64,31,199,31,185,31,189,31,177,31,50,31,57,31,150,31,150,30,71,31,79,31,89,31,73,31,103,31,145,31,90,31,73,31,49,31,226,31,106,31,140,31,202,31,202,30,231,31,216,31,139,31,139,30,42,31,95,31,114,31,111,31,74,31,72,31,125,31,152,31,146,31,146,30,174,31,119,31,93,31,93,30,102,31,128,31,79,31,198,31,7,31,138,31,138,30,3,31,3,30,200,31,249,31,23,31,102,31,102,30,102,29,102,28,87,31,64,31,36,31,127,31,127,30,104,31,94,31,150,31,199,31,118,31,118,30,22,31,27,31,68,31,142,31,29,31,1,31,1,30,125,31,162,31,162,30,73,31,149,31,85,31,157,31,205,31,106,31,204,31,76,31,167,31,51,31,253,31,252,31,50,31,124,31,154,31,175,31,175,30,9,31,9,30,148,31,86,31,86,30,114,31,182,31,171,31,254,31,115,31,6,31,223,31,6,31,81,31,52,31,52,30,52,29,198,31,20,31,213,31,213,30,125,31,105,31,105,30,228,31,167,31,42,31,212,31,203,31,32,31,6,31,220,31,135,31,188,31,218,31,10,31,89,31,58,31,70,31,70,30,155,31,62,31,65,31,123,31,123,30,123,29,17,31,191,31,191,30,252,31,232,31,181,31,181,30,252,31,141,31,63,31,138,31,196,31,64,31,218,31,120,31,244,31,126,31,35,31,35,30,190,31,156,31,218,31,196,31,218,31,216,31,216,30,162,31,115,31,70,31,175,31,175,30,175,29,175,28,239,31,203,31,234,31,127,31,224,31,202,31,24,31,213,31,200,31,20,31,57,31,57,30,206,31,206,30,222,31,108,31,20,31,223,31,77,31,227,31,227,30,7,31,191,31,220,31,174,31,160,31,207,31,123,31,13,31,242,31,242,30,223,31,99,31,99,30,164,31,32,31,32,30,67,31,123,31,123,30,230,31,38,31,197,31,66,31,36,31,36,30,54,31,121,31,78,31,115,31,188,31,148,31,128,31,173,31,173,30,123,31,4,31,189,31,106,31,40,31,83,31,24,31,156,31,174,31,250,31,250,30,185,31,228,31,69,31,69,30,180,31,180,30,63,31,63,30,202,31,221,31,151,31,42,31,42,30,58,31,58,30,248,31,230,31,201,31,60,31,217,31,217,30,238,31,48,31,9,31,9,30,92,31,23,31,122,31,70,31,174,31,252,31,177,31,1,31,1,30,1,29,1,28,101,31,101,30,101,29,116,31,186,31,174,31,239,31,224,31,106,31,175,31,175,30,80,31,62,31,56,31,1,31,6,31,6,30,35,31,200,31,46,31,142,31,142,30,142,29,183,31,183,30,141,31,211,31,211,30,24,31,94,31,185,31,185,30,68,31,236,31,190,31,195,31,195,30,192,31,216,31,186,31,229,31,240,31,72,31,53,31,53,30,53,29,214,31,5,31,175,31,58,31,58,30,58,29,125,31,209,31,209,30,209,29,209,28,209,27,68,31,168,31,38,31,175,31,118,31,227,31,39,31,54,31,142,31,142,30,98,31,23,31,143,31,104,31,66,31,80,31,150,31,250,31,21,31,177,31,24,31,176,31,101,31,31,31,209,31,209,30,61,31,54,31,147,31,99,31,32,31,249,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
