-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_450 is
end project_tb_450;

architecture project_tb_arch_450 of project_tb_450 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 716;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,189,0,211,0,218,0,129,0,43,0,215,0,185,0,20,0,164,0,11,0,0,0,0,0,89,0,24,0,48,0,160,0,0,0,105,0,127,0,203,0,0,0,19,0,0,0,57,0,150,0,7,0,132,0,170,0,31,0,0,0,185,0,136,0,165,0,7,0,14,0,61,0,94,0,0,0,0,0,147,0,105,0,88,0,41,0,145,0,107,0,213,0,0,0,255,0,239,0,0,0,0,0,96,0,153,0,163,0,109,0,119,0,175,0,164,0,182,0,15,0,159,0,224,0,70,0,0,0,43,0,0,0,0,0,244,0,176,0,240,0,149,0,255,0,181,0,127,0,0,0,0,0,181,0,115,0,174,0,220,0,9,0,163,0,128,0,21,0,223,0,50,0,14,0,58,0,35,0,3,0,42,0,48,0,119,0,155,0,231,0,241,0,71,0,37,0,40,0,38,0,0,0,204,0,164,0,41,0,239,0,226,0,31,0,204,0,66,0,0,0,220,0,181,0,0,0,147,0,0,0,142,0,0,0,161,0,234,0,152,0,0,0,0,0,0,0,103,0,192,0,177,0,105,0,188,0,38,0,234,0,201,0,138,0,239,0,0,0,0,0,2,0,0,0,37,0,75,0,183,0,175,0,177,0,5,0,105,0,0,0,248,0,225,0,152,0,205,0,103,0,235,0,217,0,81,0,0,0,157,0,52,0,250,0,7,0,0,0,0,0,0,0,102,0,63,0,230,0,120,0,216,0,0,0,0,0,18,0,93,0,144,0,182,0,80,0,205,0,186,0,0,0,0,0,171,0,0,0,167,0,239,0,0,0,0,0,160,0,239,0,0,0,62,0,180,0,59,0,20,0,0,0,48,0,0,0,123,0,34,0,242,0,87,0,37,0,49,0,0,0,175,0,126,0,132,0,154,0,60,0,108,0,215,0,150,0,187,0,164,0,157,0,65,0,90,0,0,0,16,0,139,0,24,0,77,0,197,0,147,0,247,0,188,0,218,0,164,0,42,0,25,0,143,0,89,0,103,0,0,0,19,0,0,0,78,0,12,0,0,0,20,0,180,0,0,0,223,0,29,0,34,0,0,0,179,0,29,0,0,0,73,0,103,0,4,0,226,0,0,0,17,0,76,0,29,0,225,0,63,0,106,0,78,0,194,0,153,0,14,0,58,0,175,0,161,0,224,0,0,0,180,0,105,0,227,0,180,0,97,0,202,0,134,0,192,0,83,0,191,0,233,0,77,0,194,0,175,0,0,0,55,0,157,0,29,0,0,0,71,0,116,0,0,0,147,0,127,0,187,0,207,0,64,0,171,0,183,0,237,0,0,0,213,0,202,0,92,0,0,0,235,0,40,0,210,0,194,0,108,0,79,0,248,0,230,0,126,0,60,0,54,0,207,0,226,0,201,0,13,0,32,0,44,0,49,0,22,0,110,0,0,0,244,0,77,0,80,0,21,0,5,0,196,0,54,0,42,0,0,0,99,0,51,0,108,0,0,0,0,0,145,0,224,0,209,0,65,0,84,0,166,0,245,0,114,0,30,0,115,0,228,0,114,0,135,0,16,0,244,0,140,0,95,0,235,0,78,0,181,0,89,0,0,0,198,0,98,0,0,0,181,0,153,0,13,0,36,0,45,0,156,0,5,0,15,0,0,0,75,0,150,0,97,0,189,0,155,0,105,0,133,0,0,0,153,0,204,0,59,0,0,0,193,0,209,0,150,0,175,0,218,0,166,0,0,0,41,0,252,0,107,0,0,0,141,0,15,0,21,0,0,0,198,0,43,0,226,0,44,0,165,0,0,0,192,0,0,0,0,0,0,0,213,0,158,0,14,0,0,0,2,0,28,0,204,0,200,0,0,0,199,0,0,0,144,0,186,0,97,0,76,0,32,0,191,0,0,0,10,0,203,0,24,0,232,0,132,0,204,0,0,0,114,0,37,0,145,0,42,0,233,0,4,0,158,0,150,0,62,0,32,0,97,0,132,0,128,0,157,0,0,0,39,0,139,0,0,0,56,0,0,0,21,0,108,0,123,0,49,0,0,0,5,0,24,0,18,0,38,0,162,0,55,0,241,0,0,0,221,0,9,0,0,0,206,0,96,0,199,0,172,0,246,0,178,0,203,0,78,0,0,0,76,0,204,0,0,0,0,0,126,0,142,0,100,0,145,0,219,0,187,0,132,0,125,0,174,0,2,0,14,0,122,0,209,0,0,0,111,0,0,0,100,0,126,0,197,0,228,0,207,0,0,0,186,0,78,0,89,0,0,0,251,0,159,0,0,0,231,0,253,0,134,0,59,0,0,0,146,0,18,0,0,0,209,0,78,0,172,0,69,0,0,0,67,0,231,0,0,0,0,0,234,0,27,0,186,0,178,0,22,0,35,0,0,0,226,0,229,0,245,0,10,0,0,0,20,0,130,0,250,0,43,0,140,0,0,0,241,0,238,0,230,0,22,0,115,0,175,0,133,0,0,0,6,0,85,0,168,0,0,0,179,0,157,0,71,0,188,0,0,0,20,0,0,0,204,0,69,0,3,0,19,0,170,0,145,0,107,0,116,0,224,0,6,0,184,0,104,0,101,0,243,0,215,0,60,0,202,0,0,0,113,0,239,0,0,0,223,0,14,0,0,0,155,0,214,0,178,0,0,0,35,0,117,0,0,0,65,0,0,0,213,0,0,0,0,0,190,0,65,0,235,0,228,0,14,0,92,0,0,0,187,0,92,0,252,0,209,0,226,0,0,0,0,0,125,0,133,0,135,0,201,0,0,0,0,0,0,0,233,0,134,0,67,0,245,0,109,0,0,0,215,0,0,0,200,0,118,0,0,0,230,0,0,0,121,0,250,0,103,0,118,0,255,0,76,0,192,0,0,0,202,0,0,0,116,0,0,0,13,0,195,0,33,0,0,0,123,0,85,0,0,0,173,0,238,0,190,0,81,0,0,0,56,0,230,0,89,0,186,0,0,0,42,0,0,0,186,0,25,0,213,0,0,0,114,0,0,0,0,0,132,0,117,0,246,0,95,0,128,0,149,0,170,0,41,0,131,0,17,0,92,0,34,0,0,0,45,0,168,0,4,0,193,0,9,0,0,0,76,0,172,0,0,0,106,0,236,0,0,0,44,0,176,0,160,0,193,0,0,0,252,0,0,0,197,0,139,0,44,0,35,0,0,0,127,0,60,0,51,0,0,0,59,0,253,0,123,0);
signal scenario_full  : scenario_type := (133,31,189,31,211,31,218,31,129,31,43,31,215,31,185,31,20,31,164,31,11,31,11,30,11,29,89,31,24,31,48,31,160,31,160,30,105,31,127,31,203,31,203,30,19,31,19,30,57,31,150,31,7,31,132,31,170,31,31,31,31,30,185,31,136,31,165,31,7,31,14,31,61,31,94,31,94,30,94,29,147,31,105,31,88,31,41,31,145,31,107,31,213,31,213,30,255,31,239,31,239,30,239,29,96,31,153,31,163,31,109,31,119,31,175,31,164,31,182,31,15,31,159,31,224,31,70,31,70,30,43,31,43,30,43,29,244,31,176,31,240,31,149,31,255,31,181,31,127,31,127,30,127,29,181,31,115,31,174,31,220,31,9,31,163,31,128,31,21,31,223,31,50,31,14,31,58,31,35,31,3,31,42,31,48,31,119,31,155,31,231,31,241,31,71,31,37,31,40,31,38,31,38,30,204,31,164,31,41,31,239,31,226,31,31,31,204,31,66,31,66,30,220,31,181,31,181,30,147,31,147,30,142,31,142,30,161,31,234,31,152,31,152,30,152,29,152,28,103,31,192,31,177,31,105,31,188,31,38,31,234,31,201,31,138,31,239,31,239,30,239,29,2,31,2,30,37,31,75,31,183,31,175,31,177,31,5,31,105,31,105,30,248,31,225,31,152,31,205,31,103,31,235,31,217,31,81,31,81,30,157,31,52,31,250,31,7,31,7,30,7,29,7,28,102,31,63,31,230,31,120,31,216,31,216,30,216,29,18,31,93,31,144,31,182,31,80,31,205,31,186,31,186,30,186,29,171,31,171,30,167,31,239,31,239,30,239,29,160,31,239,31,239,30,62,31,180,31,59,31,20,31,20,30,48,31,48,30,123,31,34,31,242,31,87,31,37,31,49,31,49,30,175,31,126,31,132,31,154,31,60,31,108,31,215,31,150,31,187,31,164,31,157,31,65,31,90,31,90,30,16,31,139,31,24,31,77,31,197,31,147,31,247,31,188,31,218,31,164,31,42,31,25,31,143,31,89,31,103,31,103,30,19,31,19,30,78,31,12,31,12,30,20,31,180,31,180,30,223,31,29,31,34,31,34,30,179,31,29,31,29,30,73,31,103,31,4,31,226,31,226,30,17,31,76,31,29,31,225,31,63,31,106,31,78,31,194,31,153,31,14,31,58,31,175,31,161,31,224,31,224,30,180,31,105,31,227,31,180,31,97,31,202,31,134,31,192,31,83,31,191,31,233,31,77,31,194,31,175,31,175,30,55,31,157,31,29,31,29,30,71,31,116,31,116,30,147,31,127,31,187,31,207,31,64,31,171,31,183,31,237,31,237,30,213,31,202,31,92,31,92,30,235,31,40,31,210,31,194,31,108,31,79,31,248,31,230,31,126,31,60,31,54,31,207,31,226,31,201,31,13,31,32,31,44,31,49,31,22,31,110,31,110,30,244,31,77,31,80,31,21,31,5,31,196,31,54,31,42,31,42,30,99,31,51,31,108,31,108,30,108,29,145,31,224,31,209,31,65,31,84,31,166,31,245,31,114,31,30,31,115,31,228,31,114,31,135,31,16,31,244,31,140,31,95,31,235,31,78,31,181,31,89,31,89,30,198,31,98,31,98,30,181,31,153,31,13,31,36,31,45,31,156,31,5,31,15,31,15,30,75,31,150,31,97,31,189,31,155,31,105,31,133,31,133,30,153,31,204,31,59,31,59,30,193,31,209,31,150,31,175,31,218,31,166,31,166,30,41,31,252,31,107,31,107,30,141,31,15,31,21,31,21,30,198,31,43,31,226,31,44,31,165,31,165,30,192,31,192,30,192,29,192,28,213,31,158,31,14,31,14,30,2,31,28,31,204,31,200,31,200,30,199,31,199,30,144,31,186,31,97,31,76,31,32,31,191,31,191,30,10,31,203,31,24,31,232,31,132,31,204,31,204,30,114,31,37,31,145,31,42,31,233,31,4,31,158,31,150,31,62,31,32,31,97,31,132,31,128,31,157,31,157,30,39,31,139,31,139,30,56,31,56,30,21,31,108,31,123,31,49,31,49,30,5,31,24,31,18,31,38,31,162,31,55,31,241,31,241,30,221,31,9,31,9,30,206,31,96,31,199,31,172,31,246,31,178,31,203,31,78,31,78,30,76,31,204,31,204,30,204,29,126,31,142,31,100,31,145,31,219,31,187,31,132,31,125,31,174,31,2,31,14,31,122,31,209,31,209,30,111,31,111,30,100,31,126,31,197,31,228,31,207,31,207,30,186,31,78,31,89,31,89,30,251,31,159,31,159,30,231,31,253,31,134,31,59,31,59,30,146,31,18,31,18,30,209,31,78,31,172,31,69,31,69,30,67,31,231,31,231,30,231,29,234,31,27,31,186,31,178,31,22,31,35,31,35,30,226,31,229,31,245,31,10,31,10,30,20,31,130,31,250,31,43,31,140,31,140,30,241,31,238,31,230,31,22,31,115,31,175,31,133,31,133,30,6,31,85,31,168,31,168,30,179,31,157,31,71,31,188,31,188,30,20,31,20,30,204,31,69,31,3,31,19,31,170,31,145,31,107,31,116,31,224,31,6,31,184,31,104,31,101,31,243,31,215,31,60,31,202,31,202,30,113,31,239,31,239,30,223,31,14,31,14,30,155,31,214,31,178,31,178,30,35,31,117,31,117,30,65,31,65,30,213,31,213,30,213,29,190,31,65,31,235,31,228,31,14,31,92,31,92,30,187,31,92,31,252,31,209,31,226,31,226,30,226,29,125,31,133,31,135,31,201,31,201,30,201,29,201,28,233,31,134,31,67,31,245,31,109,31,109,30,215,31,215,30,200,31,118,31,118,30,230,31,230,30,121,31,250,31,103,31,118,31,255,31,76,31,192,31,192,30,202,31,202,30,116,31,116,30,13,31,195,31,33,31,33,30,123,31,85,31,85,30,173,31,238,31,190,31,81,31,81,30,56,31,230,31,89,31,186,31,186,30,42,31,42,30,186,31,25,31,213,31,213,30,114,31,114,30,114,29,132,31,117,31,246,31,95,31,128,31,149,31,170,31,41,31,131,31,17,31,92,31,34,31,34,30,45,31,168,31,4,31,193,31,9,31,9,30,76,31,172,31,172,30,106,31,236,31,236,30,44,31,176,31,160,31,193,31,193,30,252,31,252,30,197,31,139,31,44,31,35,31,35,30,127,31,60,31,51,31,51,30,59,31,253,31,123,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
