-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 564;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (123,0,248,0,209,0,252,0,174,0,0,0,0,0,0,0,197,0,49,0,195,0,5,0,9,0,231,0,0,0,125,0,41,0,0,0,1,0,222,0,196,0,157,0,142,0,95,0,123,0,154,0,230,0,13,0,212,0,17,0,116,0,0,0,57,0,70,0,42,0,148,0,30,0,0,0,0,0,14,0,192,0,89,0,104,0,0,0,248,0,216,0,69,0,0,0,144,0,242,0,35,0,250,0,148,0,162,0,246,0,74,0,179,0,193,0,0,0,246,0,59,0,136,0,244,0,60,0,0,0,0,0,85,0,107,0,26,0,120,0,143,0,89,0,62,0,115,0,186,0,78,0,0,0,248,0,200,0,143,0,52,0,14,0,66,0,92,0,154,0,51,0,0,0,249,0,166,0,15,0,152,0,159,0,155,0,0,0,163,0,249,0,140,0,25,0,0,0,165,0,73,0,184,0,21,0,0,0,39,0,212,0,0,0,3,0,243,0,0,0,189,0,0,0,74,0,200,0,17,0,0,0,12,0,24,0,165,0,162,0,136,0,0,0,58,0,148,0,0,0,0,0,182,0,0,0,0,0,72,0,12,0,66,0,14,0,230,0,169,0,0,0,190,0,157,0,0,0,98,0,195,0,135,0,14,0,147,0,12,0,247,0,20,0,252,0,108,0,0,0,228,0,0,0,43,0,126,0,182,0,236,0,60,0,0,0,0,0,45,0,119,0,86,0,123,0,148,0,163,0,107,0,20,0,16,0,153,0,197,0,234,0,148,0,148,0,0,0,190,0,108,0,0,0,163,0,130,0,182,0,31,0,136,0,19,0,158,0,163,0,18,0,0,0,0,0,126,0,227,0,48,0,29,0,0,0,0,0,13,0,170,0,3,0,9,0,127,0,0,0,0,0,211,0,0,0,105,0,219,0,49,0,153,0,0,0,109,0,73,0,170,0,128,0,0,0,140,0,45,0,129,0,0,0,231,0,183,0,57,0,119,0,69,0,199,0,211,0,107,0,39,0,136,0,128,0,211,0,148,0,37,0,254,0,0,0,0,0,255,0,0,0,30,0,170,0,201,0,1,0,176,0,154,0,181,0,249,0,50,0,228,0,95,0,72,0,28,0,4,0,0,0,124,0,219,0,214,0,65,0,60,0,140,0,3,0,99,0,56,0,0,0,65,0,0,0,52,0,17,0,67,0,104,0,45,0,146,0,122,0,62,0,0,0,109,0,23,0,118,0,171,0,94,0,1,0,0,0,232,0,0,0,72,0,0,0,149,0,0,0,78,0,0,0,136,0,137,0,190,0,0,0,49,0,0,0,85,0,62,0,65,0,191,0,71,0,245,0,127,0,196,0,69,0,0,0,219,0,109,0,183,0,235,0,0,0,224,0,126,0,0,0,0,0,184,0,68,0,211,0,227,0,218,0,88,0,191,0,0,0,13,0,188,0,94,0,148,0,231,0,223,0,188,0,9,0,46,0,4,0,45,0,6,0,0,0,0,0,0,0,74,0,0,0,0,0,129,0,1,0,20,0,166,0,206,0,29,0,91,0,214,0,217,0,0,0,0,0,0,0,117,0,24,0,0,0,78,0,229,0,180,0,67,0,23,0,0,0,47,0,46,0,228,0,65,0,0,0,0,0,0,0,239,0,225,0,49,0,50,0,30,0,230,0,104,0,0,0,239,0,131,0,0,0,18,0,58,0,0,0,20,0,0,0,202,0,60,0,64,0,0,0,0,0,246,0,99,0,229,0,41,0,46,0,123,0,0,0,0,0,0,0,78,0,0,0,15,0,209,0,181,0,81,0,120,0,198,0,39,0,47,0,0,0,70,0,0,0,7,0,144,0,52,0,0,0,180,0,124,0,9,0,232,0,31,0,68,0,0,0,0,0,115,0,42,0,90,0,129,0,180,0,45,0,27,0,0,0,100,0,194,0,0,0,215,0,3,0,1,0,114,0,0,0,0,0,147,0,145,0,155,0,226,0,130,0,231,0,198,0,187,0,115,0,50,0,62,0,51,0,17,0,53,0,24,0,222,0,2,0,69,0,208,0,20,0,139,0,194,0,233,0,43,0,253,0,42,0,176,0,126,0,80,0,80,0,229,0,0,0,191,0,235,0,18,0,209,0,253,0,0,0,240,0,147,0,129,0,67,0,94,0,77,0,0,0,232,0,0,0,172,0,9,0,238,0,168,0,0,0,68,0,0,0,55,0,170,0,113,0,150,0,0,0,226,0,242,0,97,0,115,0,232,0,0,0,83,0,4,0,165,0,0,0,249,0,0,0,70,0,0,0,71,0,99,0,222,0,148,0,0,0,31,0,236,0,0,0,0,0,0,0,11,0,73,0,0,0,196,0,202,0,116,0,15,0,0,0,199,0,0,0,147,0,148,0,27,0,152,0,206,0,50,0,28,0,23,0,102,0,122,0,152,0,138,0,187,0,83,0,209,0,251,0,111,0,36,0,116,0,130,0,0,0,4,0,0,0,111,0,238,0,0,0,79,0,0,0,26,0,25,0,45,0,0,0,0,0);
signal scenario_full  : scenario_type := (123,31,248,31,209,31,252,31,174,31,174,30,174,29,174,28,197,31,49,31,195,31,5,31,9,31,231,31,231,30,125,31,41,31,41,30,1,31,222,31,196,31,157,31,142,31,95,31,123,31,154,31,230,31,13,31,212,31,17,31,116,31,116,30,57,31,70,31,42,31,148,31,30,31,30,30,30,29,14,31,192,31,89,31,104,31,104,30,248,31,216,31,69,31,69,30,144,31,242,31,35,31,250,31,148,31,162,31,246,31,74,31,179,31,193,31,193,30,246,31,59,31,136,31,244,31,60,31,60,30,60,29,85,31,107,31,26,31,120,31,143,31,89,31,62,31,115,31,186,31,78,31,78,30,248,31,200,31,143,31,52,31,14,31,66,31,92,31,154,31,51,31,51,30,249,31,166,31,15,31,152,31,159,31,155,31,155,30,163,31,249,31,140,31,25,31,25,30,165,31,73,31,184,31,21,31,21,30,39,31,212,31,212,30,3,31,243,31,243,30,189,31,189,30,74,31,200,31,17,31,17,30,12,31,24,31,165,31,162,31,136,31,136,30,58,31,148,31,148,30,148,29,182,31,182,30,182,29,72,31,12,31,66,31,14,31,230,31,169,31,169,30,190,31,157,31,157,30,98,31,195,31,135,31,14,31,147,31,12,31,247,31,20,31,252,31,108,31,108,30,228,31,228,30,43,31,126,31,182,31,236,31,60,31,60,30,60,29,45,31,119,31,86,31,123,31,148,31,163,31,107,31,20,31,16,31,153,31,197,31,234,31,148,31,148,31,148,30,190,31,108,31,108,30,163,31,130,31,182,31,31,31,136,31,19,31,158,31,163,31,18,31,18,30,18,29,126,31,227,31,48,31,29,31,29,30,29,29,13,31,170,31,3,31,9,31,127,31,127,30,127,29,211,31,211,30,105,31,219,31,49,31,153,31,153,30,109,31,73,31,170,31,128,31,128,30,140,31,45,31,129,31,129,30,231,31,183,31,57,31,119,31,69,31,199,31,211,31,107,31,39,31,136,31,128,31,211,31,148,31,37,31,254,31,254,30,254,29,255,31,255,30,30,31,170,31,201,31,1,31,176,31,154,31,181,31,249,31,50,31,228,31,95,31,72,31,28,31,4,31,4,30,124,31,219,31,214,31,65,31,60,31,140,31,3,31,99,31,56,31,56,30,65,31,65,30,52,31,17,31,67,31,104,31,45,31,146,31,122,31,62,31,62,30,109,31,23,31,118,31,171,31,94,31,1,31,1,30,232,31,232,30,72,31,72,30,149,31,149,30,78,31,78,30,136,31,137,31,190,31,190,30,49,31,49,30,85,31,62,31,65,31,191,31,71,31,245,31,127,31,196,31,69,31,69,30,219,31,109,31,183,31,235,31,235,30,224,31,126,31,126,30,126,29,184,31,68,31,211,31,227,31,218,31,88,31,191,31,191,30,13,31,188,31,94,31,148,31,231,31,223,31,188,31,9,31,46,31,4,31,45,31,6,31,6,30,6,29,6,28,74,31,74,30,74,29,129,31,1,31,20,31,166,31,206,31,29,31,91,31,214,31,217,31,217,30,217,29,217,28,117,31,24,31,24,30,78,31,229,31,180,31,67,31,23,31,23,30,47,31,46,31,228,31,65,31,65,30,65,29,65,28,239,31,225,31,49,31,50,31,30,31,230,31,104,31,104,30,239,31,131,31,131,30,18,31,58,31,58,30,20,31,20,30,202,31,60,31,64,31,64,30,64,29,246,31,99,31,229,31,41,31,46,31,123,31,123,30,123,29,123,28,78,31,78,30,15,31,209,31,181,31,81,31,120,31,198,31,39,31,47,31,47,30,70,31,70,30,7,31,144,31,52,31,52,30,180,31,124,31,9,31,232,31,31,31,68,31,68,30,68,29,115,31,42,31,90,31,129,31,180,31,45,31,27,31,27,30,100,31,194,31,194,30,215,31,3,31,1,31,114,31,114,30,114,29,147,31,145,31,155,31,226,31,130,31,231,31,198,31,187,31,115,31,50,31,62,31,51,31,17,31,53,31,24,31,222,31,2,31,69,31,208,31,20,31,139,31,194,31,233,31,43,31,253,31,42,31,176,31,126,31,80,31,80,31,229,31,229,30,191,31,235,31,18,31,209,31,253,31,253,30,240,31,147,31,129,31,67,31,94,31,77,31,77,30,232,31,232,30,172,31,9,31,238,31,168,31,168,30,68,31,68,30,55,31,170,31,113,31,150,31,150,30,226,31,242,31,97,31,115,31,232,31,232,30,83,31,4,31,165,31,165,30,249,31,249,30,70,31,70,30,71,31,99,31,222,31,148,31,148,30,31,31,236,31,236,30,236,29,236,28,11,31,73,31,73,30,196,31,202,31,116,31,15,31,15,30,199,31,199,30,147,31,148,31,27,31,152,31,206,31,50,31,28,31,23,31,102,31,122,31,152,31,138,31,187,31,83,31,209,31,251,31,111,31,36,31,116,31,130,31,130,30,4,31,4,30,111,31,238,31,238,30,79,31,79,30,26,31,25,31,45,31,45,30,45,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
