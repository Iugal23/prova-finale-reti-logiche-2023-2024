-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 982;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (110,0,102,0,196,0,165,0,116,0,17,0,19,0,11,0,0,0,155,0,0,0,82,0,112,0,0,0,0,0,161,0,54,0,89,0,0,0,252,0,212,0,17,0,132,0,11,0,244,0,183,0,154,0,236,0,3,0,101,0,88,0,177,0,41,0,88,0,180,0,10,0,118,0,135,0,64,0,110,0,64,0,105,0,97,0,7,0,24,0,205,0,192,0,209,0,0,0,228,0,0,0,135,0,214,0,0,0,40,0,0,0,155,0,0,0,230,0,92,0,0,0,117,0,122,0,86,0,185,0,129,0,23,0,41,0,0,0,116,0,147,0,55,0,0,0,145,0,0,0,203,0,72,0,0,0,86,0,11,0,13,0,241,0,0,0,225,0,42,0,84,0,118,0,48,0,91,0,120,0,82,0,195,0,225,0,0,0,249,0,48,0,124,0,26,0,25,0,89,0,135,0,194,0,237,0,47,0,123,0,171,0,198,0,47,0,234,0,86,0,0,0,12,0,197,0,125,0,178,0,0,0,21,0,38,0,52,0,116,0,27,0,12,0,107,0,200,0,42,0,128,0,155,0,195,0,193,0,155,0,221,0,188,0,0,0,119,0,92,0,54,0,252,0,245,0,136,0,220,0,39,0,224,0,206,0,232,0,74,0,125,0,104,0,84,0,223,0,71,0,236,0,0,0,0,0,114,0,0,0,0,0,222,0,0,0,0,0,33,0,0,0,29,0,20,0,67,0,173,0,122,0,139,0,206,0,143,0,0,0,37,0,0,0,0,0,61,0,0,0,0,0,41,0,0,0,233,0,239,0,111,0,0,0,0,0,78,0,0,0,155,0,61,0,94,0,135,0,14,0,125,0,12,0,113,0,234,0,102,0,244,0,0,0,74,0,99,0,44,0,54,0,158,0,252,0,129,0,64,0,0,0,174,0,205,0,33,0,167,0,0,0,0,0,16,0,191,0,1,0,63,0,239,0,220,0,116,0,22,0,236,0,0,0,106,0,103,0,0,0,0,0,17,0,213,0,68,0,246,0,157,0,111,0,29,0,93,0,252,0,0,0,87,0,70,0,133,0,206,0,0,0,30,0,81,0,152,0,0,0,11,0,191,0,126,0,244,0,121,0,72,0,244,0,20,0,47,0,26,0,120,0,0,0,0,0,82,0,228,0,0,0,83,0,90,0,0,0,108,0,179,0,0,0,2,0,181,0,245,0,68,0,31,0,0,0,24,0,0,0,74,0,91,0,176,0,64,0,0,0,0,0,0,0,124,0,82,0,207,0,201,0,120,0,108,0,46,0,89,0,58,0,103,0,69,0,0,0,37,0,0,0,36,0,186,0,2,0,37,0,50,0,53,0,147,0,185,0,39,0,111,0,238,0,0,0,154,0,222,0,0,0,53,0,247,0,0,0,191,0,95,0,94,0,113,0,155,0,78,0,81,0,48,0,172,0,10,0,172,0,2,0,10,0,16,0,167,0,114,0,109,0,0,0,43,0,95,0,6,0,90,0,162,0,111,0,146,0,4,0,0,0,138,0,0,0,9,0,74,0,112,0,12,0,0,0,254,0,48,0,6,0,41,0,0,0,95,0,226,0,13,0,76,0,236,0,173,0,0,0,26,0,36,0,170,0,18,0,0,0,141,0,72,0,0,0,0,0,244,0,0,0,153,0,191,0,47,0,6,0,0,0,55,0,43,0,107,0,50,0,0,0,20,0,0,0,245,0,132,0,255,0,197,0,0,0,10,0,24,0,131,0,205,0,0,0,136,0,50,0,0,0,53,0,62,0,0,0,101,0,183,0,184,0,165,0,52,0,79,0,241,0,0,0,71,0,117,0,31,0,247,0,19,0,156,0,187,0,213,0,244,0,111,0,46,0,24,0,197,0,171,0,100,0,75,0,113,0,112,0,0,0,89,0,60,0,11,0,223,0,65,0,178,0,54,0,245,0,93,0,13,0,14,0,64,0,158,0,0,0,143,0,217,0,58,0,105,0,98,0,76,0,0,0,0,0,203,0,19,0,0,0,7,0,0,0,181,0,0,0,213,0,0,0,65,0,230,0,0,0,0,0,9,0,248,0,211,0,0,0,95,0,174,0,211,0,90,0,172,0,106,0,27,0,0,0,184,0,198,0,149,0,180,0,105,0,156,0,0,0,186,0,56,0,245,0,0,0,130,0,0,0,16,0,0,0,1,0,94,0,166,0,245,0,210,0,174,0,84,0,111,0,95,0,9,0,30,0,249,0,229,0,198,0,26,0,127,0,59,0,18,0,250,0,86,0,183,0,229,0,242,0,0,0,144,0,65,0,115,0,0,0,18,0,0,0,95,0,56,0,106,0,19,0,132,0,59,0,92,0,173,0,0,0,13,0,150,0,58,0,4,0,168,0,211,0,123,0,222,0,240,0,0,0,101,0,0,0,15,0,222,0,50,0,182,0,214,0,17,0,0,0,189,0,160,0,201,0,155,0,97,0,161,0,221,0,149,0,196,0,163,0,36,0,241,0,201,0,110,0,46,0,0,0,15,0,165,0,173,0,82,0,39,0,67,0,255,0,240,0,146,0,86,0,0,0,221,0,0,0,211,0,104,0,0,0,188,0,234,0,36,0,0,0,156,0,141,0,206,0,0,0,206,0,152,0,225,0,201,0,136,0,95,0,0,0,165,0,111,0,33,0,225,0,0,0,222,0,24,0,63,0,34,0,16,0,4,0,232,0,0,0,0,0,227,0,173,0,40,0,47,0,177,0,241,0,0,0,27,0,109,0,24,0,156,0,216,0,51,0,0,0,144,0,130,0,226,0,176,0,94,0,68,0,143,0,177,0,52,0,62,0,233,0,199,0,0,0,0,0,211,0,205,0,38,0,0,0,0,0,173,0,0,0,30,0,45,0,96,0,131,0,7,0,171,0,222,0,142,0,15,0,39,0,129,0,14,0,47,0,35,0,102,0,76,0,59,0,154,0,215,0,79,0,240,0,132,0,206,0,33,0,77,0,46,0,221,0,47,0,0,0,219,0,253,0,170,0,219,0,177,0,0,0,51,0,207,0,0,0,119,0,97,0,198,0,174,0,79,0,169,0,0,0,0,0,133,0,248,0,105,0,134,0,87,0,36,0,0,0,0,0,102,0,163,0,220,0,159,0,0,0,0,0,25,0,0,0,179,0,188,0,194,0,232,0,132,0,69,0,0,0,201,0,119,0,141,0,0,0,0,0,0,0,76,0,224,0,0,0,223,0,106,0,145,0,243,0,122,0,180,0,72,0,122,0,0,0,201,0,155,0,45,0,242,0,0,0,155,0,200,0,172,0,0,0,67,0,165,0,0,0,106,0,93,0,10,0,31,0,30,0,0,0,134,0,26,0,213,0,186,0,179,0,169,0,234,0,154,0,101,0,0,0,55,0,0,0,9,0,176,0,2,0,180,0,120,0,173,0,24,0,96,0,218,0,75,0,0,0,199,0,45,0,221,0,170,0,20,0,0,0,107,0,133,0,122,0,222,0,55,0,94,0,192,0,0,0,169,0,33,0,37,0,151,0,0,0,49,0,0,0,177,0,250,0,125,0,110,0,176,0,0,0,208,0,136,0,70,0,204,0,36,0,116,0,136,0,0,0,88,0,0,0,0,0,7,0,0,0,0,0,18,0,0,0,225,0,0,0,157,0,41,0,237,0,225,0,157,0,66,0,102,0,0,0,156,0,161,0,0,0,82,0,191,0,28,0,183,0,125,0,9,0,6,0,181,0,0,0,104,0,152,0,0,0,183,0,0,0,248,0,167,0,93,0,0,0,199,0,159,0,34,0,60,0,73,0,96,0,103,0,120,0,66,0,199,0,0,0,0,0,204,0,27,0,173,0,74,0,245,0,201,0,0,0,0,0,82,0,74,0,37,0,98,0,235,0,154,0,215,0,201,0,29,0,0,0,212,0,244,0,17,0,196,0,0,0,115,0,112,0,0,0,100,0,254,0,106,0,226,0,51,0,186,0,76,0,130,0,0,0,223,0,0,0,40,0,7,0,70,0,0,0,16,0,235,0,33,0,88,0,31,0,0,0,236,0,0,0,29,0,28,0,0,0,127,0,44,0,219,0,0,0,155,0,0,0,251,0,67,0,160,0,152,0,0,0,13,0,91,0,18,0,150,0,26,0,0,0,88,0,0,0,0,0,147,0,0,0,34,0,140,0,213,0,118,0,0,0,81,0,0,0,0,0,0,0,53,0,73,0,216,0,0,0,189,0,2,0,185,0,21,0,0,0,3,0,0,0,5,0,203,0,2,0,9,0,68,0,93,0,170,0,91,0,0,0,47,0,166,0,255,0,44,0,23,0,238,0,242,0,79,0,3,0,46,0,125,0,141,0,16,0,199,0,167,0,125,0,60,0,93,0,0,0,227,0,3,0,75,0,60,0);
signal scenario_full  : scenario_type := (110,31,102,31,196,31,165,31,116,31,17,31,19,31,11,31,11,30,155,31,155,30,82,31,112,31,112,30,112,29,161,31,54,31,89,31,89,30,252,31,212,31,17,31,132,31,11,31,244,31,183,31,154,31,236,31,3,31,101,31,88,31,177,31,41,31,88,31,180,31,10,31,118,31,135,31,64,31,110,31,64,31,105,31,97,31,7,31,24,31,205,31,192,31,209,31,209,30,228,31,228,30,135,31,214,31,214,30,40,31,40,30,155,31,155,30,230,31,92,31,92,30,117,31,122,31,86,31,185,31,129,31,23,31,41,31,41,30,116,31,147,31,55,31,55,30,145,31,145,30,203,31,72,31,72,30,86,31,11,31,13,31,241,31,241,30,225,31,42,31,84,31,118,31,48,31,91,31,120,31,82,31,195,31,225,31,225,30,249,31,48,31,124,31,26,31,25,31,89,31,135,31,194,31,237,31,47,31,123,31,171,31,198,31,47,31,234,31,86,31,86,30,12,31,197,31,125,31,178,31,178,30,21,31,38,31,52,31,116,31,27,31,12,31,107,31,200,31,42,31,128,31,155,31,195,31,193,31,155,31,221,31,188,31,188,30,119,31,92,31,54,31,252,31,245,31,136,31,220,31,39,31,224,31,206,31,232,31,74,31,125,31,104,31,84,31,223,31,71,31,236,31,236,30,236,29,114,31,114,30,114,29,222,31,222,30,222,29,33,31,33,30,29,31,20,31,67,31,173,31,122,31,139,31,206,31,143,31,143,30,37,31,37,30,37,29,61,31,61,30,61,29,41,31,41,30,233,31,239,31,111,31,111,30,111,29,78,31,78,30,155,31,61,31,94,31,135,31,14,31,125,31,12,31,113,31,234,31,102,31,244,31,244,30,74,31,99,31,44,31,54,31,158,31,252,31,129,31,64,31,64,30,174,31,205,31,33,31,167,31,167,30,167,29,16,31,191,31,1,31,63,31,239,31,220,31,116,31,22,31,236,31,236,30,106,31,103,31,103,30,103,29,17,31,213,31,68,31,246,31,157,31,111,31,29,31,93,31,252,31,252,30,87,31,70,31,133,31,206,31,206,30,30,31,81,31,152,31,152,30,11,31,191,31,126,31,244,31,121,31,72,31,244,31,20,31,47,31,26,31,120,31,120,30,120,29,82,31,228,31,228,30,83,31,90,31,90,30,108,31,179,31,179,30,2,31,181,31,245,31,68,31,31,31,31,30,24,31,24,30,74,31,91,31,176,31,64,31,64,30,64,29,64,28,124,31,82,31,207,31,201,31,120,31,108,31,46,31,89,31,58,31,103,31,69,31,69,30,37,31,37,30,36,31,186,31,2,31,37,31,50,31,53,31,147,31,185,31,39,31,111,31,238,31,238,30,154,31,222,31,222,30,53,31,247,31,247,30,191,31,95,31,94,31,113,31,155,31,78,31,81,31,48,31,172,31,10,31,172,31,2,31,10,31,16,31,167,31,114,31,109,31,109,30,43,31,95,31,6,31,90,31,162,31,111,31,146,31,4,31,4,30,138,31,138,30,9,31,74,31,112,31,12,31,12,30,254,31,48,31,6,31,41,31,41,30,95,31,226,31,13,31,76,31,236,31,173,31,173,30,26,31,36,31,170,31,18,31,18,30,141,31,72,31,72,30,72,29,244,31,244,30,153,31,191,31,47,31,6,31,6,30,55,31,43,31,107,31,50,31,50,30,20,31,20,30,245,31,132,31,255,31,197,31,197,30,10,31,24,31,131,31,205,31,205,30,136,31,50,31,50,30,53,31,62,31,62,30,101,31,183,31,184,31,165,31,52,31,79,31,241,31,241,30,71,31,117,31,31,31,247,31,19,31,156,31,187,31,213,31,244,31,111,31,46,31,24,31,197,31,171,31,100,31,75,31,113,31,112,31,112,30,89,31,60,31,11,31,223,31,65,31,178,31,54,31,245,31,93,31,13,31,14,31,64,31,158,31,158,30,143,31,217,31,58,31,105,31,98,31,76,31,76,30,76,29,203,31,19,31,19,30,7,31,7,30,181,31,181,30,213,31,213,30,65,31,230,31,230,30,230,29,9,31,248,31,211,31,211,30,95,31,174,31,211,31,90,31,172,31,106,31,27,31,27,30,184,31,198,31,149,31,180,31,105,31,156,31,156,30,186,31,56,31,245,31,245,30,130,31,130,30,16,31,16,30,1,31,94,31,166,31,245,31,210,31,174,31,84,31,111,31,95,31,9,31,30,31,249,31,229,31,198,31,26,31,127,31,59,31,18,31,250,31,86,31,183,31,229,31,242,31,242,30,144,31,65,31,115,31,115,30,18,31,18,30,95,31,56,31,106,31,19,31,132,31,59,31,92,31,173,31,173,30,13,31,150,31,58,31,4,31,168,31,211,31,123,31,222,31,240,31,240,30,101,31,101,30,15,31,222,31,50,31,182,31,214,31,17,31,17,30,189,31,160,31,201,31,155,31,97,31,161,31,221,31,149,31,196,31,163,31,36,31,241,31,201,31,110,31,46,31,46,30,15,31,165,31,173,31,82,31,39,31,67,31,255,31,240,31,146,31,86,31,86,30,221,31,221,30,211,31,104,31,104,30,188,31,234,31,36,31,36,30,156,31,141,31,206,31,206,30,206,31,152,31,225,31,201,31,136,31,95,31,95,30,165,31,111,31,33,31,225,31,225,30,222,31,24,31,63,31,34,31,16,31,4,31,232,31,232,30,232,29,227,31,173,31,40,31,47,31,177,31,241,31,241,30,27,31,109,31,24,31,156,31,216,31,51,31,51,30,144,31,130,31,226,31,176,31,94,31,68,31,143,31,177,31,52,31,62,31,233,31,199,31,199,30,199,29,211,31,205,31,38,31,38,30,38,29,173,31,173,30,30,31,45,31,96,31,131,31,7,31,171,31,222,31,142,31,15,31,39,31,129,31,14,31,47,31,35,31,102,31,76,31,59,31,154,31,215,31,79,31,240,31,132,31,206,31,33,31,77,31,46,31,221,31,47,31,47,30,219,31,253,31,170,31,219,31,177,31,177,30,51,31,207,31,207,30,119,31,97,31,198,31,174,31,79,31,169,31,169,30,169,29,133,31,248,31,105,31,134,31,87,31,36,31,36,30,36,29,102,31,163,31,220,31,159,31,159,30,159,29,25,31,25,30,179,31,188,31,194,31,232,31,132,31,69,31,69,30,201,31,119,31,141,31,141,30,141,29,141,28,76,31,224,31,224,30,223,31,106,31,145,31,243,31,122,31,180,31,72,31,122,31,122,30,201,31,155,31,45,31,242,31,242,30,155,31,200,31,172,31,172,30,67,31,165,31,165,30,106,31,93,31,10,31,31,31,30,31,30,30,134,31,26,31,213,31,186,31,179,31,169,31,234,31,154,31,101,31,101,30,55,31,55,30,9,31,176,31,2,31,180,31,120,31,173,31,24,31,96,31,218,31,75,31,75,30,199,31,45,31,221,31,170,31,20,31,20,30,107,31,133,31,122,31,222,31,55,31,94,31,192,31,192,30,169,31,33,31,37,31,151,31,151,30,49,31,49,30,177,31,250,31,125,31,110,31,176,31,176,30,208,31,136,31,70,31,204,31,36,31,116,31,136,31,136,30,88,31,88,30,88,29,7,31,7,30,7,29,18,31,18,30,225,31,225,30,157,31,41,31,237,31,225,31,157,31,66,31,102,31,102,30,156,31,161,31,161,30,82,31,191,31,28,31,183,31,125,31,9,31,6,31,181,31,181,30,104,31,152,31,152,30,183,31,183,30,248,31,167,31,93,31,93,30,199,31,159,31,34,31,60,31,73,31,96,31,103,31,120,31,66,31,199,31,199,30,199,29,204,31,27,31,173,31,74,31,245,31,201,31,201,30,201,29,82,31,74,31,37,31,98,31,235,31,154,31,215,31,201,31,29,31,29,30,212,31,244,31,17,31,196,31,196,30,115,31,112,31,112,30,100,31,254,31,106,31,226,31,51,31,186,31,76,31,130,31,130,30,223,31,223,30,40,31,7,31,70,31,70,30,16,31,235,31,33,31,88,31,31,31,31,30,236,31,236,30,29,31,28,31,28,30,127,31,44,31,219,31,219,30,155,31,155,30,251,31,67,31,160,31,152,31,152,30,13,31,91,31,18,31,150,31,26,31,26,30,88,31,88,30,88,29,147,31,147,30,34,31,140,31,213,31,118,31,118,30,81,31,81,30,81,29,81,28,53,31,73,31,216,31,216,30,189,31,2,31,185,31,21,31,21,30,3,31,3,30,5,31,203,31,2,31,9,31,68,31,93,31,170,31,91,31,91,30,47,31,166,31,255,31,44,31,23,31,238,31,242,31,79,31,3,31,46,31,125,31,141,31,16,31,199,31,167,31,125,31,60,31,93,31,93,30,227,31,3,31,75,31,60,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
