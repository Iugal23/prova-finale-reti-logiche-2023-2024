-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_615 is
end project_tb_615;

architecture project_tb_arch_615 of project_tb_615 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 171;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,117,0,138,0,103,0,102,0,189,0,252,0,4,0,130,0,194,0,176,0,198,0,243,0,254,0,7,0,76,0,0,0,187,0,0,0,42,0,222,0,209,0,156,0,19,0,0,0,0,0,169,0,20,0,171,0,134,0,155,0,0,0,57,0,39,0,193,0,181,0,0,0,46,0,62,0,182,0,142,0,234,0,124,0,0,0,97,0,210,0,0,0,171,0,87,0,207,0,24,0,57,0,0,0,86,0,14,0,75,0,222,0,182,0,220,0,99,0,0,0,112,0,88,0,252,0,128,0,165,0,191,0,194,0,114,0,29,0,229,0,98,0,0,0,122,0,26,0,193,0,0,0,97,0,65,0,22,0,0,0,62,0,0,0,138,0,15,0,81,0,29,0,132,0,0,0,246,0,187,0,20,0,228,0,174,0,235,0,211,0,0,0,0,0,233,0,133,0,217,0,161,0,229,0,103,0,9,0,45,0,39,0,0,0,24,0,228,0,221,0,11,0,112,0,0,0,38,0,127,0,143,0,252,0,83,0,0,0,86,0,0,0,240,0,81,0,0,0,19,0,0,0,6,0,18,0,92,0,8,0,0,0,239,0,0,0,115,0,227,0,100,0,8,0,0,0,219,0,103,0,0,0,179,0,0,0,51,0,0,0,123,0,95,0,0,0,47,0,88,0,0,0,219,0,137,0,232,0,214,0,0,0,170,0,93,0,221,0,111,0,22,0,210,0,255,0,0,0,10,0,117,0,38,0,121,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,117,31,138,31,103,31,102,31,189,31,252,31,4,31,130,31,194,31,176,31,198,31,243,31,254,31,7,31,76,31,76,30,187,31,187,30,42,31,222,31,209,31,156,31,19,31,19,30,19,29,169,31,20,31,171,31,134,31,155,31,155,30,57,31,39,31,193,31,181,31,181,30,46,31,62,31,182,31,142,31,234,31,124,31,124,30,97,31,210,31,210,30,171,31,87,31,207,31,24,31,57,31,57,30,86,31,14,31,75,31,222,31,182,31,220,31,99,31,99,30,112,31,88,31,252,31,128,31,165,31,191,31,194,31,114,31,29,31,229,31,98,31,98,30,122,31,26,31,193,31,193,30,97,31,65,31,22,31,22,30,62,31,62,30,138,31,15,31,81,31,29,31,132,31,132,30,246,31,187,31,20,31,228,31,174,31,235,31,211,31,211,30,211,29,233,31,133,31,217,31,161,31,229,31,103,31,9,31,45,31,39,31,39,30,24,31,228,31,221,31,11,31,112,31,112,30,38,31,127,31,143,31,252,31,83,31,83,30,86,31,86,30,240,31,81,31,81,30,19,31,19,30,6,31,18,31,92,31,8,31,8,30,239,31,239,30,115,31,227,31,100,31,8,31,8,30,219,31,103,31,103,30,179,31,179,30,51,31,51,30,123,31,95,31,95,30,47,31,88,31,88,30,219,31,137,31,232,31,214,31,214,30,170,31,93,31,221,31,111,31,22,31,210,31,255,31,255,30,10,31,117,31,38,31,121,31,121,30,121,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
