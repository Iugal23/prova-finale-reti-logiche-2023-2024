-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 249;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,0,0,54,0,242,0,39,0,0,0,240,0,169,0,162,0,111,0,124,0,183,0,37,0,247,0,115,0,129,0,237,0,0,0,66,0,212,0,43,0,37,0,43,0,0,0,0,0,215,0,234,0,65,0,60,0,0,0,232,0,200,0,49,0,192,0,0,0,249,0,35,0,90,0,23,0,18,0,0,0,12,0,122,0,182,0,211,0,0,0,129,0,105,0,186,0,0,0,0,0,111,0,94,0,80,0,112,0,0,0,0,0,226,0,243,0,253,0,212,0,169,0,81,0,249,0,164,0,236,0,226,0,65,0,0,0,232,0,231,0,120,0,194,0,155,0,196,0,183,0,34,0,243,0,204,0,254,0,242,0,158,0,86,0,78,0,133,0,0,0,253,0,1,0,249,0,9,0,135,0,0,0,0,0,0,0,239,0,117,0,18,0,0,0,80,0,49,0,167,0,141,0,0,0,108,0,0,0,0,0,76,0,87,0,199,0,207,0,255,0,188,0,53,0,180,0,250,0,0,0,112,0,0,0,0,0,45,0,244,0,102,0,75,0,76,0,173,0,254,0,255,0,204,0,60,0,84,0,121,0,0,0,236,0,37,0,74,0,0,0,42,0,153,0,221,0,0,0,30,0,255,0,148,0,216,0,105,0,194,0,63,0,108,0,205,0,225,0,231,0,178,0,0,0,99,0,0,0,116,0,212,0,16,0,172,0,157,0,240,0,32,0,144,0,139,0,0,0,223,0,191,0,241,0,0,0,77,0,230,0,230,0,88,0,55,0,188,0,181,0,149,0,175,0,48,0,21,0,31,0,90,0,217,0,240,0,0,0,209,0,11,0,126,0,0,0,0,0,194,0,51,0,154,0,163,0,46,0,195,0,215,0,26,0,190,0,76,0,179,0,156,0,64,0,29,0,125,0,254,0,30,0,165,0,197,0,134,0,24,0,0,0,186,0,144,0,138,0,67,0,159,0,42,0,0,0,0,0,201,0,142,0,123,0,116,0,0,0,70,0,4,0,121,0,224,0,214,0,0,0,35,0,235,0,0,0,216,0,66,0,57,0,21,0,147,0,71,0,60,0,9,0,0,0,114,0,0,0,144,0,143,0,115,0,85,0);
signal scenario_full  : scenario_type := (135,31,135,30,54,31,242,31,39,31,39,30,240,31,169,31,162,31,111,31,124,31,183,31,37,31,247,31,115,31,129,31,237,31,237,30,66,31,212,31,43,31,37,31,43,31,43,30,43,29,215,31,234,31,65,31,60,31,60,30,232,31,200,31,49,31,192,31,192,30,249,31,35,31,90,31,23,31,18,31,18,30,12,31,122,31,182,31,211,31,211,30,129,31,105,31,186,31,186,30,186,29,111,31,94,31,80,31,112,31,112,30,112,29,226,31,243,31,253,31,212,31,169,31,81,31,249,31,164,31,236,31,226,31,65,31,65,30,232,31,231,31,120,31,194,31,155,31,196,31,183,31,34,31,243,31,204,31,254,31,242,31,158,31,86,31,78,31,133,31,133,30,253,31,1,31,249,31,9,31,135,31,135,30,135,29,135,28,239,31,117,31,18,31,18,30,80,31,49,31,167,31,141,31,141,30,108,31,108,30,108,29,76,31,87,31,199,31,207,31,255,31,188,31,53,31,180,31,250,31,250,30,112,31,112,30,112,29,45,31,244,31,102,31,75,31,76,31,173,31,254,31,255,31,204,31,60,31,84,31,121,31,121,30,236,31,37,31,74,31,74,30,42,31,153,31,221,31,221,30,30,31,255,31,148,31,216,31,105,31,194,31,63,31,108,31,205,31,225,31,231,31,178,31,178,30,99,31,99,30,116,31,212,31,16,31,172,31,157,31,240,31,32,31,144,31,139,31,139,30,223,31,191,31,241,31,241,30,77,31,230,31,230,31,88,31,55,31,188,31,181,31,149,31,175,31,48,31,21,31,31,31,90,31,217,31,240,31,240,30,209,31,11,31,126,31,126,30,126,29,194,31,51,31,154,31,163,31,46,31,195,31,215,31,26,31,190,31,76,31,179,31,156,31,64,31,29,31,125,31,254,31,30,31,165,31,197,31,134,31,24,31,24,30,186,31,144,31,138,31,67,31,159,31,42,31,42,30,42,29,201,31,142,31,123,31,116,31,116,30,70,31,4,31,121,31,224,31,214,31,214,30,35,31,235,31,235,30,216,31,66,31,57,31,21,31,147,31,71,31,60,31,9,31,9,30,114,31,114,30,144,31,143,31,115,31,85,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
