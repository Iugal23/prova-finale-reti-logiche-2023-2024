-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 357;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (246,0,0,0,0,0,0,0,61,0,153,0,0,0,36,0,0,0,34,0,103,0,51,0,37,0,193,0,121,0,206,0,4,0,126,0,123,0,200,0,235,0,0,0,40,0,57,0,0,0,101,0,27,0,229,0,160,0,170,0,161,0,104,0,188,0,0,0,89,0,100,0,8,0,80,0,86,0,18,0,0,0,248,0,42,0,0,0,67,0,171,0,0,0,128,0,83,0,95,0,0,0,161,0,199,0,0,0,50,0,28,0,151,0,0,0,251,0,49,0,194,0,87,0,113,0,224,0,110,0,10,0,199,0,0,0,127,0,0,0,191,0,10,0,0,0,244,0,97,0,52,0,132,0,0,0,5,0,0,0,92,0,0,0,0,0,175,0,232,0,254,0,0,0,97,0,5,0,33,0,231,0,95,0,199,0,0,0,0,0,167,0,82,0,63,0,68,0,0,0,0,0,30,0,0,0,98,0,191,0,42,0,0,0,130,0,35,0,114,0,74,0,97,0,180,0,0,0,0,0,246,0,225,0,44,0,14,0,221,0,184,0,183,0,0,0,164,0,0,0,229,0,107,0,0,0,157,0,205,0,0,0,65,0,0,0,0,0,102,0,80,0,0,0,204,0,117,0,0,0,0,0,232,0,0,0,193,0,107,0,186,0,0,0,8,0,0,0,187,0,160,0,0,0,25,0,19,0,34,0,0,0,37,0,39,0,74,0,31,0,55,0,137,0,181,0,54,0,109,0,2,0,0,0,35,0,116,0,127,0,79,0,155,0,48,0,2,0,131,0,225,0,255,0,34,0,132,0,0,0,0,0,13,0,154,0,142,0,53,0,79,0,34,0,72,0,145,0,131,0,0,0,28,0,26,0,82,0,229,0,142,0,45,0,10,0,244,0,201,0,39,0,76,0,124,0,216,0,104,0,30,0,139,0,105,0,0,0,22,0,216,0,180,0,238,0,0,0,10,0,228,0,0,0,126,0,7,0,163,0,214,0,106,0,180,0,6,0,89,0,199,0,163,0,0,0,62,0,207,0,0,0,160,0,244,0,158,0,73,0,0,0,0,0,0,0,170,0,132,0,212,0,78,0,21,0,208,0,35,0,42,0,191,0,0,0,12,0,66,0,68,0,114,0,110,0,143,0,0,0,137,0,0,0,119,0,72,0,0,0,190,0,149,0,36,0,40,0,178,0,226,0,142,0,0,0,90,0,147,0,0,0,7,0,0,0,176,0,92,0,0,0,142,0,81,0,44,0,162,0,137,0,79,0,44,0,0,0,146,0,146,0,229,0,63,0,84,0,223,0,244,0,145,0,48,0,90,0,160,0,0,0,40,0,12,0,0,0,165,0,0,0,0,0,33,0,152,0,0,0,2,0,51,0,147,0,70,0,0,0,71,0,102,0,137,0,160,0,211,0,0,0,44,0,206,0,0,0,222,0,158,0,205,0,52,0,157,0,231,0,0,0,170,0,0,0,133,0,4,0,96,0,0,0,72,0,152,0,0,0,196,0,174,0,0,0,75,0,234,0,80,0,142,0,31,0,207,0,166,0,0,0,0,0,243,0,174,0,0,0,82,0,56,0,0,0,20,0,141,0,249,0,124,0);
signal scenario_full  : scenario_type := (246,31,246,30,246,29,246,28,61,31,153,31,153,30,36,31,36,30,34,31,103,31,51,31,37,31,193,31,121,31,206,31,4,31,126,31,123,31,200,31,235,31,235,30,40,31,57,31,57,30,101,31,27,31,229,31,160,31,170,31,161,31,104,31,188,31,188,30,89,31,100,31,8,31,80,31,86,31,18,31,18,30,248,31,42,31,42,30,67,31,171,31,171,30,128,31,83,31,95,31,95,30,161,31,199,31,199,30,50,31,28,31,151,31,151,30,251,31,49,31,194,31,87,31,113,31,224,31,110,31,10,31,199,31,199,30,127,31,127,30,191,31,10,31,10,30,244,31,97,31,52,31,132,31,132,30,5,31,5,30,92,31,92,30,92,29,175,31,232,31,254,31,254,30,97,31,5,31,33,31,231,31,95,31,199,31,199,30,199,29,167,31,82,31,63,31,68,31,68,30,68,29,30,31,30,30,98,31,191,31,42,31,42,30,130,31,35,31,114,31,74,31,97,31,180,31,180,30,180,29,246,31,225,31,44,31,14,31,221,31,184,31,183,31,183,30,164,31,164,30,229,31,107,31,107,30,157,31,205,31,205,30,65,31,65,30,65,29,102,31,80,31,80,30,204,31,117,31,117,30,117,29,232,31,232,30,193,31,107,31,186,31,186,30,8,31,8,30,187,31,160,31,160,30,25,31,19,31,34,31,34,30,37,31,39,31,74,31,31,31,55,31,137,31,181,31,54,31,109,31,2,31,2,30,35,31,116,31,127,31,79,31,155,31,48,31,2,31,131,31,225,31,255,31,34,31,132,31,132,30,132,29,13,31,154,31,142,31,53,31,79,31,34,31,72,31,145,31,131,31,131,30,28,31,26,31,82,31,229,31,142,31,45,31,10,31,244,31,201,31,39,31,76,31,124,31,216,31,104,31,30,31,139,31,105,31,105,30,22,31,216,31,180,31,238,31,238,30,10,31,228,31,228,30,126,31,7,31,163,31,214,31,106,31,180,31,6,31,89,31,199,31,163,31,163,30,62,31,207,31,207,30,160,31,244,31,158,31,73,31,73,30,73,29,73,28,170,31,132,31,212,31,78,31,21,31,208,31,35,31,42,31,191,31,191,30,12,31,66,31,68,31,114,31,110,31,143,31,143,30,137,31,137,30,119,31,72,31,72,30,190,31,149,31,36,31,40,31,178,31,226,31,142,31,142,30,90,31,147,31,147,30,7,31,7,30,176,31,92,31,92,30,142,31,81,31,44,31,162,31,137,31,79,31,44,31,44,30,146,31,146,31,229,31,63,31,84,31,223,31,244,31,145,31,48,31,90,31,160,31,160,30,40,31,12,31,12,30,165,31,165,30,165,29,33,31,152,31,152,30,2,31,51,31,147,31,70,31,70,30,71,31,102,31,137,31,160,31,211,31,211,30,44,31,206,31,206,30,222,31,158,31,205,31,52,31,157,31,231,31,231,30,170,31,170,30,133,31,4,31,96,31,96,30,72,31,152,31,152,30,196,31,174,31,174,30,75,31,234,31,80,31,142,31,31,31,207,31,166,31,166,30,166,29,243,31,174,31,174,30,82,31,56,31,56,30,20,31,141,31,249,31,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
