-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_222 is
end project_tb_222;

architecture project_tb_arch_222 of project_tb_222 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 704;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (231,0,4,0,94,0,123,0,70,0,152,0,0,0,0,0,211,0,53,0,123,0,106,0,6,0,88,0,56,0,62,0,0,0,26,0,199,0,0,0,187,0,69,0,204,0,143,0,22,0,116,0,160,0,178,0,0,0,222,0,156,0,0,0,98,0,0,0,24,0,126,0,162,0,210,0,237,0,0,0,92,0,123,0,252,0,0,0,148,0,88,0,0,0,243,0,148,0,233,0,0,0,252,0,10,0,0,0,242,0,129,0,250,0,72,0,0,0,54,0,33,0,65,0,178,0,216,0,0,0,0,0,161,0,26,0,215,0,0,0,0,0,187,0,194,0,31,0,71,0,247,0,225,0,145,0,36,0,81,0,126,0,0,0,217,0,18,0,36,0,71,0,0,0,208,0,111,0,0,0,13,0,78,0,135,0,82,0,108,0,194,0,193,0,255,0,112,0,252,0,198,0,0,0,86,0,205,0,26,0,238,0,183,0,0,0,66,0,99,0,77,0,112,0,255,0,211,0,0,0,0,0,231,0,159,0,241,0,0,0,119,0,0,0,85,0,74,0,184,0,76,0,0,0,0,0,140,0,122,0,0,0,0,0,0,0,251,0,61,0,76,0,0,0,44,0,0,0,240,0,195,0,164,0,249,0,0,0,0,0,32,0,65,0,190,0,9,0,0,0,0,0,234,0,168,0,43,0,172,0,136,0,0,0,98,0,111,0,221,0,66,0,47,0,49,0,94,0,129,0,0,0,15,0,0,0,2,0,19,0,175,0,21,0,148,0,241,0,36,0,91,0,0,0,249,0,51,0,201,0,143,0,194,0,190,0,220,0,37,0,217,0,234,0,123,0,0,0,225,0,0,0,160,0,171,0,84,0,168,0,0,0,251,0,108,0,193,0,202,0,126,0,0,0,107,0,178,0,189,0,99,0,209,0,221,0,220,0,125,0,113,0,78,0,14,0,0,0,59,0,0,0,140,0,122,0,0,0,0,0,110,0,58,0,226,0,150,0,208,0,0,0,0,0,186,0,244,0,19,0,18,0,109,0,0,0,20,0,189,0,234,0,0,0,75,0,239,0,139,0,0,0,192,0,94,0,35,0,0,0,103,0,0,0,222,0,0,0,116,0,55,0,137,0,165,0,0,0,209,0,154,0,173,0,188,0,0,0,255,0,137,0,204,0,150,0,241,0,74,0,24,0,0,0,181,0,164,0,38,0,117,0,154,0,9,0,8,0,163,0,154,0,229,0,146,0,168,0,179,0,135,0,9,0,0,0,249,0,2,0,0,0,77,0,242,0,126,0,0,0,0,0,13,0,204,0,56,0,137,0,85,0,136,0,0,0,161,0,95,0,225,0,99,0,158,0,181,0,0,0,179,0,99,0,228,0,0,0,160,0,241,0,145,0,212,0,76,0,0,0,18,0,115,0,254,0,62,0,231,0,0,0,182,0,88,0,152,0,0,0,252,0,164,0,231,0,131,0,164,0,78,0,0,0,139,0,210,0,46,0,153,0,42,0,0,0,11,0,190,0,171,0,50,0,148,0,135,0,162,0,17,0,170,0,39,0,206,0,82,0,30,0,66,0,193,0,254,0,121,0,205,0,176,0,194,0,118,0,131,0,181,0,102,0,9,0,141,0,103,0,0,0,0,0,76,0,224,0,215,0,0,0,0,0,233,0,0,0,183,0,124,0,207,0,141,0,142,0,0,0,53,0,119,0,221,0,166,0,0,0,0,0,27,0,48,0,0,0,12,0,101,0,144,0,0,0,0,0,30,0,244,0,227,0,157,0,0,0,72,0,77,0,223,0,140,0,150,0,0,0,164,0,0,0,0,0,77,0,18,0,0,0,249,0,74,0,117,0,91,0,144,0,211,0,109,0,0,0,155,0,214,0,185,0,162,0,149,0,188,0,14,0,36,0,81,0,37,0,155,0,218,0,186,0,189,0,0,0,112,0,0,0,205,0,152,0,109,0,211,0,4,0,26,0,41,0,118,0,203,0,63,0,0,0,124,0,198,0,59,0,0,0,149,0,0,0,2,0,234,0,178,0,23,0,90,0,211,0,0,0,230,0,123,0,36,0,131,0,173,0,0,0,45,0,77,0,111,0,214,0,238,0,177,0,184,0,62,0,194,0,99,0,188,0,162,0,9,0,102,0,0,0,26,0,84,0,219,0,0,0,102,0,0,0,89,0,48,0,241,0,41,0,59,0,86,0,125,0,110,0,213,0,95,0,53,0,65,0,219,0,63,0,68,0,191,0,89,0,0,0,153,0,0,0,5,0,237,0,15,0,146,0,239,0,145,0,158,0,0,0,170,0,203,0,0,0,239,0,254,0,0,0,53,0,46,0,123,0,189,0,200,0,63,0,193,0,162,0,248,0,93,0,183,0,136,0,13,0,249,0,0,0,127,0,0,0,0,0,44,0,22,0,0,0,179,0,97,0,187,0,206,0,51,0,94,0,26,0,34,0,140,0,60,0,105,0,152,0,155,0,170,0,98,0,138,0,208,0,108,0,11,0,88,0,0,0,140,0,71,0,36,0,240,0,0,0,140,0,26,0,203,0,0,0,43,0,167,0,193,0,208,0,0,0,0,0,31,0,76,0,11,0,0,0,39,0,30,0,162,0,227,0,234,0,211,0,0,0,185,0,245,0,84,0,140,0,121,0,29,0,199,0,33,0,106,0,185,0,98,0,10,0,0,0,190,0,198,0,45,0,198,0,0,0,153,0,53,0,0,0,89,0,246,0,0,0,123,0,17,0,0,0,166,0,0,0,98,0,6,0,4,0,43,0,203,0,0,0,0,0,177,0,0,0,121,0,246,0,0,0,192,0,227,0,56,0,0,0,81,0,102,0,124,0,195,0,189,0,148,0,120,0,67,0,2,0,113,0,20,0,61,0,0,0,233,0,66,0,19,0,254,0,0,0,92,0,68,0,170,0,207,0,203,0,54,0,74,0,27,0,224,0,0,0,34,0,44,0,130,0,185,0,179,0,66,0,0,0,210,0,103,0,115,0,0,0,184,0,66,0,80,0,0,0,203,0,2,0,144,0,62,0,206,0,212,0,210,0,0,0,17,0,239,0,125,0,142,0,78,0,0,0,238,0,26,0,56,0,68,0,185,0,135,0,0,0,43,0,95,0,166,0,149,0,164,0,28,0);
signal scenario_full  : scenario_type := (231,31,4,31,94,31,123,31,70,31,152,31,152,30,152,29,211,31,53,31,123,31,106,31,6,31,88,31,56,31,62,31,62,30,26,31,199,31,199,30,187,31,69,31,204,31,143,31,22,31,116,31,160,31,178,31,178,30,222,31,156,31,156,30,98,31,98,30,24,31,126,31,162,31,210,31,237,31,237,30,92,31,123,31,252,31,252,30,148,31,88,31,88,30,243,31,148,31,233,31,233,30,252,31,10,31,10,30,242,31,129,31,250,31,72,31,72,30,54,31,33,31,65,31,178,31,216,31,216,30,216,29,161,31,26,31,215,31,215,30,215,29,187,31,194,31,31,31,71,31,247,31,225,31,145,31,36,31,81,31,126,31,126,30,217,31,18,31,36,31,71,31,71,30,208,31,111,31,111,30,13,31,78,31,135,31,82,31,108,31,194,31,193,31,255,31,112,31,252,31,198,31,198,30,86,31,205,31,26,31,238,31,183,31,183,30,66,31,99,31,77,31,112,31,255,31,211,31,211,30,211,29,231,31,159,31,241,31,241,30,119,31,119,30,85,31,74,31,184,31,76,31,76,30,76,29,140,31,122,31,122,30,122,29,122,28,251,31,61,31,76,31,76,30,44,31,44,30,240,31,195,31,164,31,249,31,249,30,249,29,32,31,65,31,190,31,9,31,9,30,9,29,234,31,168,31,43,31,172,31,136,31,136,30,98,31,111,31,221,31,66,31,47,31,49,31,94,31,129,31,129,30,15,31,15,30,2,31,19,31,175,31,21,31,148,31,241,31,36,31,91,31,91,30,249,31,51,31,201,31,143,31,194,31,190,31,220,31,37,31,217,31,234,31,123,31,123,30,225,31,225,30,160,31,171,31,84,31,168,31,168,30,251,31,108,31,193,31,202,31,126,31,126,30,107,31,178,31,189,31,99,31,209,31,221,31,220,31,125,31,113,31,78,31,14,31,14,30,59,31,59,30,140,31,122,31,122,30,122,29,110,31,58,31,226,31,150,31,208,31,208,30,208,29,186,31,244,31,19,31,18,31,109,31,109,30,20,31,189,31,234,31,234,30,75,31,239,31,139,31,139,30,192,31,94,31,35,31,35,30,103,31,103,30,222,31,222,30,116,31,55,31,137,31,165,31,165,30,209,31,154,31,173,31,188,31,188,30,255,31,137,31,204,31,150,31,241,31,74,31,24,31,24,30,181,31,164,31,38,31,117,31,154,31,9,31,8,31,163,31,154,31,229,31,146,31,168,31,179,31,135,31,9,31,9,30,249,31,2,31,2,30,77,31,242,31,126,31,126,30,126,29,13,31,204,31,56,31,137,31,85,31,136,31,136,30,161,31,95,31,225,31,99,31,158,31,181,31,181,30,179,31,99,31,228,31,228,30,160,31,241,31,145,31,212,31,76,31,76,30,18,31,115,31,254,31,62,31,231,31,231,30,182,31,88,31,152,31,152,30,252,31,164,31,231,31,131,31,164,31,78,31,78,30,139,31,210,31,46,31,153,31,42,31,42,30,11,31,190,31,171,31,50,31,148,31,135,31,162,31,17,31,170,31,39,31,206,31,82,31,30,31,66,31,193,31,254,31,121,31,205,31,176,31,194,31,118,31,131,31,181,31,102,31,9,31,141,31,103,31,103,30,103,29,76,31,224,31,215,31,215,30,215,29,233,31,233,30,183,31,124,31,207,31,141,31,142,31,142,30,53,31,119,31,221,31,166,31,166,30,166,29,27,31,48,31,48,30,12,31,101,31,144,31,144,30,144,29,30,31,244,31,227,31,157,31,157,30,72,31,77,31,223,31,140,31,150,31,150,30,164,31,164,30,164,29,77,31,18,31,18,30,249,31,74,31,117,31,91,31,144,31,211,31,109,31,109,30,155,31,214,31,185,31,162,31,149,31,188,31,14,31,36,31,81,31,37,31,155,31,218,31,186,31,189,31,189,30,112,31,112,30,205,31,152,31,109,31,211,31,4,31,26,31,41,31,118,31,203,31,63,31,63,30,124,31,198,31,59,31,59,30,149,31,149,30,2,31,234,31,178,31,23,31,90,31,211,31,211,30,230,31,123,31,36,31,131,31,173,31,173,30,45,31,77,31,111,31,214,31,238,31,177,31,184,31,62,31,194,31,99,31,188,31,162,31,9,31,102,31,102,30,26,31,84,31,219,31,219,30,102,31,102,30,89,31,48,31,241,31,41,31,59,31,86,31,125,31,110,31,213,31,95,31,53,31,65,31,219,31,63,31,68,31,191,31,89,31,89,30,153,31,153,30,5,31,237,31,15,31,146,31,239,31,145,31,158,31,158,30,170,31,203,31,203,30,239,31,254,31,254,30,53,31,46,31,123,31,189,31,200,31,63,31,193,31,162,31,248,31,93,31,183,31,136,31,13,31,249,31,249,30,127,31,127,30,127,29,44,31,22,31,22,30,179,31,97,31,187,31,206,31,51,31,94,31,26,31,34,31,140,31,60,31,105,31,152,31,155,31,170,31,98,31,138,31,208,31,108,31,11,31,88,31,88,30,140,31,71,31,36,31,240,31,240,30,140,31,26,31,203,31,203,30,43,31,167,31,193,31,208,31,208,30,208,29,31,31,76,31,11,31,11,30,39,31,30,31,162,31,227,31,234,31,211,31,211,30,185,31,245,31,84,31,140,31,121,31,29,31,199,31,33,31,106,31,185,31,98,31,10,31,10,30,190,31,198,31,45,31,198,31,198,30,153,31,53,31,53,30,89,31,246,31,246,30,123,31,17,31,17,30,166,31,166,30,98,31,6,31,4,31,43,31,203,31,203,30,203,29,177,31,177,30,121,31,246,31,246,30,192,31,227,31,56,31,56,30,81,31,102,31,124,31,195,31,189,31,148,31,120,31,67,31,2,31,113,31,20,31,61,31,61,30,233,31,66,31,19,31,254,31,254,30,92,31,68,31,170,31,207,31,203,31,54,31,74,31,27,31,224,31,224,30,34,31,44,31,130,31,185,31,179,31,66,31,66,30,210,31,103,31,115,31,115,30,184,31,66,31,80,31,80,30,203,31,2,31,144,31,62,31,206,31,212,31,210,31,210,30,17,31,239,31,125,31,142,31,78,31,78,30,238,31,26,31,56,31,68,31,185,31,135,31,135,30,43,31,95,31,166,31,149,31,164,31,28,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
