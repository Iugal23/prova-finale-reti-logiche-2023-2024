-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 825;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,64,0,92,0,0,0,153,0,170,0,252,0,130,0,13,0,16,0,27,0,161,0,153,0,0,0,0,0,208,0,31,0,234,0,0,0,21,0,119,0,41,0,167,0,96,0,83,0,166,0,0,0,0,0,159,0,0,0,146,0,51,0,20,0,0,0,223,0,12,0,64,0,0,0,100,0,71,0,209,0,87,0,68,0,235,0,0,0,121,0,130,0,132,0,16,0,120,0,148,0,99,0,218,0,191,0,0,0,161,0,82,0,46,0,0,0,114,0,182,0,101,0,247,0,60,0,0,0,0,0,0,0,0,0,75,0,63,0,209,0,242,0,134,0,0,0,92,0,248,0,141,0,44,0,30,0,0,0,0,0,196,0,144,0,41,0,159,0,246,0,0,0,175,0,91,0,0,0,0,0,0,0,106,0,40,0,142,0,227,0,0,0,0,0,0,0,0,0,0,0,0,0,9,0,138,0,109,0,0,0,145,0,0,0,232,0,115,0,50,0,49,0,0,0,148,0,213,0,20,0,105,0,228,0,212,0,0,0,0,0,93,0,0,0,122,0,103,0,166,0,0,0,20,0,60,0,163,0,98,0,198,0,191,0,124,0,139,0,222,0,165,0,242,0,186,0,13,0,0,0,137,0,86,0,233,0,165,0,0,0,0,0,233,0,0,0,137,0,0,0,46,0,0,0,0,0,0,0,111,0,250,0,0,0,204,0,97,0,164,0,72,0,0,0,79,0,190,0,155,0,102,0,202,0,173,0,0,0,71,0,92,0,112,0,100,0,52,0,9,0,0,0,36,0,0,0,230,0,204,0,232,0,241,0,0,0,205,0,50,0,8,0,65,0,222,0,0,0,187,0,159,0,77,0,138,0,254,0,0,0,130,0,189,0,0,0,97,0,168,0,3,0,193,0,85,0,246,0,25,0,74,0,21,0,65,0,0,0,67,0,72,0,94,0,109,0,84,0,77,0,12,0,198,0,27,0,0,0,237,0,166,0,90,0,234,0,9,0,211,0,246,0,192,0,52,0,162,0,54,0,0,0,22,0,119,0,153,0,68,0,149,0,181,0,134,0,235,0,135,0,0,0,105,0,50,0,172,0,25,0,0,0,13,0,0,0,216,0,108,0,24,0,76,0,233,0,249,0,17,0,58,0,77,0,98,0,152,0,225,0,81,0,67,0,0,0,197,0,47,0,72,0,193,0,161,0,84,0,0,0,21,0,35,0,4,0,0,0,173,0,0,0,244,0,57,0,185,0,54,0,249,0,248,0,228,0,240,0,160,0,0,0,217,0,50,0,214,0,0,0,85,0,242,0,0,0,128,0,37,0,176,0,26,0,150,0,114,0,136,0,205,0,105,0,245,0,199,0,0,0,0,0,195,0,0,0,23,0,71,0,240,0,132,0,159,0,102,0,38,0,143,0,61,0,0,0,146,0,119,0,118,0,107,0,57,0,0,0,114,0,17,0,249,0,87,0,250,0,198,0,0,0,165,0,0,0,33,0,232,0,0,0,0,0,155,0,0,0,40,0,0,0,69,0,0,0,252,0,0,0,158,0,38,0,172,0,56,0,35,0,40,0,84,0,21,0,169,0,67,0,0,0,95,0,0,0,108,0,141,0,223,0,155,0,162,0,0,0,45,0,32,0,140,0,29,0,216,0,234,0,68,0,0,0,0,0,183,0,22,0,105,0,196,0,253,0,174,0,0,0,246,0,76,0,0,0,109,0,90,0,0,0,163,0,246,0,0,0,90,0,225,0,83,0,0,0,0,0,78,0,0,0,0,0,9,0,0,0,149,0,60,0,47,0,47,0,0,0,73,0,53,0,81,0,41,0,187,0,17,0,181,0,128,0,213,0,151,0,168,0,0,0,0,0,0,0,2,0,0,0,18,0,112,0,228,0,0,0,233,0,102,0,244,0,215,0,0,0,0,0,0,0,85,0,219,0,77,0,74,0,0,0,58,0,175,0,146,0,162,0,101,0,176,0,160,0,14,0,0,0,0,0,120,0,119,0,46,0,0,0,19,0,98,0,0,0,203,0,0,0,0,0,0,0,253,0,0,0,157,0,0,0,0,0,236,0,0,0,107,0,196,0,0,0,71,0,10,0,172,0,92,0,159,0,224,0,0,0,151,0,188,0,254,0,94,0,233,0,0,0,124,0,27,0,140,0,135,0,183,0,93,0,132,0,0,0,106,0,7,0,0,0,0,0,239,0,32,0,190,0,4,0,17,0,138,0,0,0,221,0,0,0,231,0,6,0,231,0,13,0,118,0,0,0,0,0,130,0,0,0,0,0,44,0,243,0,69,0,221,0,58,0,68,0,63,0,0,0,37,0,247,0,0,0,105,0,142,0,133,0,218,0,0,0,68,0,0,0,179,0,18,0,81,0,155,0,120,0,0,0,162,0,224,0,172,0,112,0,194,0,203,0,71,0,0,0,12,0,0,0,62,0,212,0,180,0,94,0,161,0,0,0,68,0,50,0,0,0,73,0,0,0,92,0,0,0,88,0,0,0,192,0,249,0,48,0,0,0,118,0,225,0,151,0,161,0,192,0,0,0,204,0,98,0,83,0,221,0,0,0,2,0,83,0,146,0,137,0,165,0,191,0,191,0,60,0,197,0,186,0,111,0,28,0,236,0,73,0,89,0,79,0,149,0,159,0,227,0,52,0,244,0,120,0,121,0,0,0,6,0,55,0,237,0,101,0,155,0,165,0,101,0,0,0,114,0,142,0,178,0,157,0,66,0,66,0,185,0,0,0,24,0,166,0,210,0,60,0,209,0,0,0,152,0,14,0,0,0,150,0,0,0,202,0,133,0,0,0,0,0,15,0,0,0,223,0,182,0,0,0,173,0,140,0,78,0,0,0,55,0,151,0,0,0,58,0,18,0,27,0,170,0,0,0,0,0,152,0,166,0,20,0,143,0,183,0,247,0,222,0,0,0,165,0,236,0,155,0,249,0,122,0,0,0,167,0,0,0,62,0,0,0,0,0,0,0,47,0,0,0,159,0,16,0,0,0,176,0,0,0,245,0,0,0,0,0,143,0,136,0,25,0,7,0,0,0,57,0,220,0,241,0,111,0,198,0,234,0,191,0,0,0,243,0,174,0,29,0,182,0,142,0,227,0,223,0,74,0,147,0,175,0,0,0,0,0,0,0,246,0,219,0,124,0,171,0,0,0,142,0,129,0,128,0,157,0,98,0,241,0,117,0,147,0,0,0,4,0,183,0,0,0,92,0,118,0,42,0,27,0,0,0,0,0,58,0,255,0,110,0,119,0,102,0,186,0,6,0,207,0,78,0,187,0,145,0,6,0,0,0,39,0,175,0,209,0,0,0,69,0,92,0,235,0,25,0,50,0,0,0,0,0,10,0,120,0,0,0,35,0,252,0,72,0,59,0,224,0,230,0,81,0,185,0,214,0,211,0,77,0,201,0,227,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,179,0,167,0,131,0,4,0,82,0,0,0,131,0,178,0,202,0,0,0,127,0,152,0,242,0,6,0,75,0,154,0,249,0,228,0,157,0,174,0,49,0,197,0,236,0,21,0,33,0,75,0,153,0,86,0,99,0,209,0,220,0,14,0,129,0,194,0,0,0,133,0,22,0,35,0,134,0,155,0,65,0,85,0,228,0,94,0,51,0,195,0,171,0,0,0,249,0,209,0);
signal scenario_full  : scenario_type := (56,31,64,31,92,31,92,30,153,31,170,31,252,31,130,31,13,31,16,31,27,31,161,31,153,31,153,30,153,29,208,31,31,31,234,31,234,30,21,31,119,31,41,31,167,31,96,31,83,31,166,31,166,30,166,29,159,31,159,30,146,31,51,31,20,31,20,30,223,31,12,31,64,31,64,30,100,31,71,31,209,31,87,31,68,31,235,31,235,30,121,31,130,31,132,31,16,31,120,31,148,31,99,31,218,31,191,31,191,30,161,31,82,31,46,31,46,30,114,31,182,31,101,31,247,31,60,31,60,30,60,29,60,28,60,27,75,31,63,31,209,31,242,31,134,31,134,30,92,31,248,31,141,31,44,31,30,31,30,30,30,29,196,31,144,31,41,31,159,31,246,31,246,30,175,31,91,31,91,30,91,29,91,28,106,31,40,31,142,31,227,31,227,30,227,29,227,28,227,27,227,26,227,25,9,31,138,31,109,31,109,30,145,31,145,30,232,31,115,31,50,31,49,31,49,30,148,31,213,31,20,31,105,31,228,31,212,31,212,30,212,29,93,31,93,30,122,31,103,31,166,31,166,30,20,31,60,31,163,31,98,31,198,31,191,31,124,31,139,31,222,31,165,31,242,31,186,31,13,31,13,30,137,31,86,31,233,31,165,31,165,30,165,29,233,31,233,30,137,31,137,30,46,31,46,30,46,29,46,28,111,31,250,31,250,30,204,31,97,31,164,31,72,31,72,30,79,31,190,31,155,31,102,31,202,31,173,31,173,30,71,31,92,31,112,31,100,31,52,31,9,31,9,30,36,31,36,30,230,31,204,31,232,31,241,31,241,30,205,31,50,31,8,31,65,31,222,31,222,30,187,31,159,31,77,31,138,31,254,31,254,30,130,31,189,31,189,30,97,31,168,31,3,31,193,31,85,31,246,31,25,31,74,31,21,31,65,31,65,30,67,31,72,31,94,31,109,31,84,31,77,31,12,31,198,31,27,31,27,30,237,31,166,31,90,31,234,31,9,31,211,31,246,31,192,31,52,31,162,31,54,31,54,30,22,31,119,31,153,31,68,31,149,31,181,31,134,31,235,31,135,31,135,30,105,31,50,31,172,31,25,31,25,30,13,31,13,30,216,31,108,31,24,31,76,31,233,31,249,31,17,31,58,31,77,31,98,31,152,31,225,31,81,31,67,31,67,30,197,31,47,31,72,31,193,31,161,31,84,31,84,30,21,31,35,31,4,31,4,30,173,31,173,30,244,31,57,31,185,31,54,31,249,31,248,31,228,31,240,31,160,31,160,30,217,31,50,31,214,31,214,30,85,31,242,31,242,30,128,31,37,31,176,31,26,31,150,31,114,31,136,31,205,31,105,31,245,31,199,31,199,30,199,29,195,31,195,30,23,31,71,31,240,31,132,31,159,31,102,31,38,31,143,31,61,31,61,30,146,31,119,31,118,31,107,31,57,31,57,30,114,31,17,31,249,31,87,31,250,31,198,31,198,30,165,31,165,30,33,31,232,31,232,30,232,29,155,31,155,30,40,31,40,30,69,31,69,30,252,31,252,30,158,31,38,31,172,31,56,31,35,31,40,31,84,31,21,31,169,31,67,31,67,30,95,31,95,30,108,31,141,31,223,31,155,31,162,31,162,30,45,31,32,31,140,31,29,31,216,31,234,31,68,31,68,30,68,29,183,31,22,31,105,31,196,31,253,31,174,31,174,30,246,31,76,31,76,30,109,31,90,31,90,30,163,31,246,31,246,30,90,31,225,31,83,31,83,30,83,29,78,31,78,30,78,29,9,31,9,30,149,31,60,31,47,31,47,31,47,30,73,31,53,31,81,31,41,31,187,31,17,31,181,31,128,31,213,31,151,31,168,31,168,30,168,29,168,28,2,31,2,30,18,31,112,31,228,31,228,30,233,31,102,31,244,31,215,31,215,30,215,29,215,28,85,31,219,31,77,31,74,31,74,30,58,31,175,31,146,31,162,31,101,31,176,31,160,31,14,31,14,30,14,29,120,31,119,31,46,31,46,30,19,31,98,31,98,30,203,31,203,30,203,29,203,28,253,31,253,30,157,31,157,30,157,29,236,31,236,30,107,31,196,31,196,30,71,31,10,31,172,31,92,31,159,31,224,31,224,30,151,31,188,31,254,31,94,31,233,31,233,30,124,31,27,31,140,31,135,31,183,31,93,31,132,31,132,30,106,31,7,31,7,30,7,29,239,31,32,31,190,31,4,31,17,31,138,31,138,30,221,31,221,30,231,31,6,31,231,31,13,31,118,31,118,30,118,29,130,31,130,30,130,29,44,31,243,31,69,31,221,31,58,31,68,31,63,31,63,30,37,31,247,31,247,30,105,31,142,31,133,31,218,31,218,30,68,31,68,30,179,31,18,31,81,31,155,31,120,31,120,30,162,31,224,31,172,31,112,31,194,31,203,31,71,31,71,30,12,31,12,30,62,31,212,31,180,31,94,31,161,31,161,30,68,31,50,31,50,30,73,31,73,30,92,31,92,30,88,31,88,30,192,31,249,31,48,31,48,30,118,31,225,31,151,31,161,31,192,31,192,30,204,31,98,31,83,31,221,31,221,30,2,31,83,31,146,31,137,31,165,31,191,31,191,31,60,31,197,31,186,31,111,31,28,31,236,31,73,31,89,31,79,31,149,31,159,31,227,31,52,31,244,31,120,31,121,31,121,30,6,31,55,31,237,31,101,31,155,31,165,31,101,31,101,30,114,31,142,31,178,31,157,31,66,31,66,31,185,31,185,30,24,31,166,31,210,31,60,31,209,31,209,30,152,31,14,31,14,30,150,31,150,30,202,31,133,31,133,30,133,29,15,31,15,30,223,31,182,31,182,30,173,31,140,31,78,31,78,30,55,31,151,31,151,30,58,31,18,31,27,31,170,31,170,30,170,29,152,31,166,31,20,31,143,31,183,31,247,31,222,31,222,30,165,31,236,31,155,31,249,31,122,31,122,30,167,31,167,30,62,31,62,30,62,29,62,28,47,31,47,30,159,31,16,31,16,30,176,31,176,30,245,31,245,30,245,29,143,31,136,31,25,31,7,31,7,30,57,31,220,31,241,31,111,31,198,31,234,31,191,31,191,30,243,31,174,31,29,31,182,31,142,31,227,31,223,31,74,31,147,31,175,31,175,30,175,29,175,28,246,31,219,31,124,31,171,31,171,30,142,31,129,31,128,31,157,31,98,31,241,31,117,31,147,31,147,30,4,31,183,31,183,30,92,31,118,31,42,31,27,31,27,30,27,29,58,31,255,31,110,31,119,31,102,31,186,31,6,31,207,31,78,31,187,31,145,31,6,31,6,30,39,31,175,31,209,31,209,30,69,31,92,31,235,31,25,31,50,31,50,30,50,29,10,31,120,31,120,30,35,31,252,31,72,31,59,31,224,31,230,31,81,31,185,31,214,31,211,31,77,31,201,31,227,31,227,30,227,29,227,28,227,27,227,26,227,25,227,24,179,31,167,31,131,31,4,31,82,31,82,30,131,31,178,31,202,31,202,30,127,31,152,31,242,31,6,31,75,31,154,31,249,31,228,31,157,31,174,31,49,31,197,31,236,31,21,31,33,31,75,31,153,31,86,31,99,31,209,31,220,31,14,31,129,31,194,31,194,30,133,31,22,31,35,31,134,31,155,31,65,31,85,31,228,31,94,31,51,31,195,31,171,31,171,30,249,31,209,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
