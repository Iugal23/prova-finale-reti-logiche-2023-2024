-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_779 is
end project_tb_779;

architecture project_tb_arch_779 of project_tb_779 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 561;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (78,0,188,0,151,0,73,0,229,0,0,0,187,0,234,0,238,0,144,0,0,0,31,0,0,0,164,0,0,0,0,0,0,0,160,0,7,0,0,0,51,0,49,0,181,0,37,0,109,0,132,0,92,0,0,0,96,0,66,0,0,0,251,0,44,0,60,0,1,0,161,0,191,0,218,0,0,0,187,0,0,0,3,0,97,0,41,0,144,0,214,0,205,0,0,0,59,0,141,0,151,0,225,0,83,0,0,0,0,0,151,0,44,0,149,0,185,0,193,0,126,0,237,0,28,0,0,0,0,0,43,0,212,0,28,0,233,0,15,0,165,0,165,0,0,0,190,0,80,0,0,0,64,0,42,0,212,0,16,0,87,0,19,0,147,0,0,0,25,0,189,0,244,0,109,0,203,0,165,0,175,0,233,0,236,0,0,0,95,0,222,0,38,0,0,0,53,0,146,0,34,0,117,0,57,0,0,0,136,0,200,0,110,0,71,0,1,0,144,0,0,0,75,0,61,0,125,0,193,0,226,0,204,0,237,0,78,0,78,0,96,0,4,0,253,0,34,0,4,0,0,0,0,0,160,0,76,0,9,0,182,0,10,0,65,0,127,0,57,0,191,0,231,0,140,0,185,0,44,0,0,0,0,0,185,0,251,0,18,0,140,0,239,0,188,0,135,0,135,0,146,0,188,0,183,0,116,0,17,0,74,0,37,0,0,0,101,0,180,0,0,0,0,0,60,0,0,0,228,0,0,0,63,0,0,0,42,0,110,0,191,0,137,0,160,0,160,0,44,0,101,0,0,0,135,0,83,0,234,0,244,0,80,0,98,0,119,0,136,0,0,0,0,0,105,0,0,0,92,0,38,0,0,0,0,0,65,0,88,0,139,0,25,0,96,0,143,0,104,0,71,0,189,0,192,0,0,0,167,0,0,0,0,0,0,0,251,0,207,0,83,0,20,0,191,0,178,0,147,0,215,0,29,0,178,0,0,0,236,0,69,0,236,0,235,0,227,0,176,0,0,0,0,0,11,0,46,0,19,0,88,0,207,0,189,0,0,0,200,0,0,0,4,0,0,0,0,0,205,0,218,0,0,0,156,0,0,0,115,0,8,0,244,0,53,0,209,0,59,0,16,0,0,0,67,0,8,0,123,0,132,0,0,0,133,0,248,0,87,0,157,0,109,0,54,0,235,0,20,0,234,0,203,0,0,0,193,0,29,0,0,0,63,0,19,0,235,0,4,0,218,0,20,0,166,0,0,0,168,0,162,0,56,0,159,0,91,0,0,0,200,0,210,0,108,0,58,0,0,0,90,0,0,0,0,0,228,0,0,0,98,0,122,0,0,0,232,0,96,0,203,0,0,0,210,0,60,0,252,0,124,0,127,0,73,0,204,0,153,0,91,0,0,0,0,0,134,0,0,0,0,0,194,0,69,0,0,0,0,0,50,0,170,0,202,0,58,0,104,0,145,0,85,0,215,0,59,0,117,0,157,0,158,0,230,0,247,0,149,0,0,0,0,0,247,0,185,0,176,0,13,0,180,0,66,0,0,0,56,0,46,0,159,0,244,0,82,0,243,0,224,0,178,0,75,0,157,0,133,0,63,0,34,0,183,0,160,0,103,0,216,0,130,0,0,0,32,0,0,0,159,0,149,0,215,0,87,0,81,0,0,0,0,0,174,0,151,0,209,0,11,0,254,0,229,0,128,0,81,0,249,0,87,0,249,0,28,0,101,0,16,0,0,0,44,0,0,0,121,0,0,0,0,0,0,0,101,0,97,0,230,0,241,0,0,0,18,0,212,0,197,0,247,0,162,0,68,0,0,0,223,0,198,0,203,0,40,0,5,0,210,0,199,0,49,0,129,0,206,0,43,0,54,0,150,0,168,0,228,0,128,0,138,0,216,0,13,0,115,0,169,0,79,0,252,0,252,0,64,0,83,0,138,0,58,0,171,0,88,0,225,0,103,0,203,0,247,0,15,0,184,0,65,0,0,0,137,0,0,0,155,0,164,0,61,0,22,0,129,0,0,0,46,0,32,0,127,0,0,0,0,0,0,0,50,0,187,0,19,0,112,0,0,0,58,0,32,0,206,0,0,0,89,0,36,0,209,0,56,0,52,0,210,0,0,0,190,0,0,0,117,0,0,0,0,0,223,0,137,0,0,0,95,0,147,0,129,0,46,0,0,0,202,0,185,0,99,0,154,0,89,0,81,0,162,0,131,0,142,0,0,0,0,0,10,0,134,0,0,0,0,0,0,0,60,0,0,0,0,0,34,0,135,0,18,0,26,0,101,0,171,0,133,0,126,0,109,0,237,0,89,0,140,0,147,0,0,0,14,0,0,0,12,0,174,0,89,0,0,0,0,0,196,0,0,0,110,0,71,0,20,0,149,0,217,0,102,0,99,0,138,0,0,0,140,0,0,0,66,0,18,0,180,0,138,0,254,0,225,0,222,0,118,0,159,0,20,0,215,0,75,0,211,0,0,0,0,0,0,0,118,0,187,0,254,0,69,0,140,0,64,0);
signal scenario_full  : scenario_type := (78,31,188,31,151,31,73,31,229,31,229,30,187,31,234,31,238,31,144,31,144,30,31,31,31,30,164,31,164,30,164,29,164,28,160,31,7,31,7,30,51,31,49,31,181,31,37,31,109,31,132,31,92,31,92,30,96,31,66,31,66,30,251,31,44,31,60,31,1,31,161,31,191,31,218,31,218,30,187,31,187,30,3,31,97,31,41,31,144,31,214,31,205,31,205,30,59,31,141,31,151,31,225,31,83,31,83,30,83,29,151,31,44,31,149,31,185,31,193,31,126,31,237,31,28,31,28,30,28,29,43,31,212,31,28,31,233,31,15,31,165,31,165,31,165,30,190,31,80,31,80,30,64,31,42,31,212,31,16,31,87,31,19,31,147,31,147,30,25,31,189,31,244,31,109,31,203,31,165,31,175,31,233,31,236,31,236,30,95,31,222,31,38,31,38,30,53,31,146,31,34,31,117,31,57,31,57,30,136,31,200,31,110,31,71,31,1,31,144,31,144,30,75,31,61,31,125,31,193,31,226,31,204,31,237,31,78,31,78,31,96,31,4,31,253,31,34,31,4,31,4,30,4,29,160,31,76,31,9,31,182,31,10,31,65,31,127,31,57,31,191,31,231,31,140,31,185,31,44,31,44,30,44,29,185,31,251,31,18,31,140,31,239,31,188,31,135,31,135,31,146,31,188,31,183,31,116,31,17,31,74,31,37,31,37,30,101,31,180,31,180,30,180,29,60,31,60,30,228,31,228,30,63,31,63,30,42,31,110,31,191,31,137,31,160,31,160,31,44,31,101,31,101,30,135,31,83,31,234,31,244,31,80,31,98,31,119,31,136,31,136,30,136,29,105,31,105,30,92,31,38,31,38,30,38,29,65,31,88,31,139,31,25,31,96,31,143,31,104,31,71,31,189,31,192,31,192,30,167,31,167,30,167,29,167,28,251,31,207,31,83,31,20,31,191,31,178,31,147,31,215,31,29,31,178,31,178,30,236,31,69,31,236,31,235,31,227,31,176,31,176,30,176,29,11,31,46,31,19,31,88,31,207,31,189,31,189,30,200,31,200,30,4,31,4,30,4,29,205,31,218,31,218,30,156,31,156,30,115,31,8,31,244,31,53,31,209,31,59,31,16,31,16,30,67,31,8,31,123,31,132,31,132,30,133,31,248,31,87,31,157,31,109,31,54,31,235,31,20,31,234,31,203,31,203,30,193,31,29,31,29,30,63,31,19,31,235,31,4,31,218,31,20,31,166,31,166,30,168,31,162,31,56,31,159,31,91,31,91,30,200,31,210,31,108,31,58,31,58,30,90,31,90,30,90,29,228,31,228,30,98,31,122,31,122,30,232,31,96,31,203,31,203,30,210,31,60,31,252,31,124,31,127,31,73,31,204,31,153,31,91,31,91,30,91,29,134,31,134,30,134,29,194,31,69,31,69,30,69,29,50,31,170,31,202,31,58,31,104,31,145,31,85,31,215,31,59,31,117,31,157,31,158,31,230,31,247,31,149,31,149,30,149,29,247,31,185,31,176,31,13,31,180,31,66,31,66,30,56,31,46,31,159,31,244,31,82,31,243,31,224,31,178,31,75,31,157,31,133,31,63,31,34,31,183,31,160,31,103,31,216,31,130,31,130,30,32,31,32,30,159,31,149,31,215,31,87,31,81,31,81,30,81,29,174,31,151,31,209,31,11,31,254,31,229,31,128,31,81,31,249,31,87,31,249,31,28,31,101,31,16,31,16,30,44,31,44,30,121,31,121,30,121,29,121,28,101,31,97,31,230,31,241,31,241,30,18,31,212,31,197,31,247,31,162,31,68,31,68,30,223,31,198,31,203,31,40,31,5,31,210,31,199,31,49,31,129,31,206,31,43,31,54,31,150,31,168,31,228,31,128,31,138,31,216,31,13,31,115,31,169,31,79,31,252,31,252,31,64,31,83,31,138,31,58,31,171,31,88,31,225,31,103,31,203,31,247,31,15,31,184,31,65,31,65,30,137,31,137,30,155,31,164,31,61,31,22,31,129,31,129,30,46,31,32,31,127,31,127,30,127,29,127,28,50,31,187,31,19,31,112,31,112,30,58,31,32,31,206,31,206,30,89,31,36,31,209,31,56,31,52,31,210,31,210,30,190,31,190,30,117,31,117,30,117,29,223,31,137,31,137,30,95,31,147,31,129,31,46,31,46,30,202,31,185,31,99,31,154,31,89,31,81,31,162,31,131,31,142,31,142,30,142,29,10,31,134,31,134,30,134,29,134,28,60,31,60,30,60,29,34,31,135,31,18,31,26,31,101,31,171,31,133,31,126,31,109,31,237,31,89,31,140,31,147,31,147,30,14,31,14,30,12,31,174,31,89,31,89,30,89,29,196,31,196,30,110,31,71,31,20,31,149,31,217,31,102,31,99,31,138,31,138,30,140,31,140,30,66,31,18,31,180,31,138,31,254,31,225,31,222,31,118,31,159,31,20,31,215,31,75,31,211,31,211,30,211,29,211,28,118,31,187,31,254,31,69,31,140,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
