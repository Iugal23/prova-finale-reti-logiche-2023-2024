-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_441 is
end project_tb_441;

architecture project_tb_arch_441 of project_tb_441 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 851;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,121,0,0,0,62,0,134,0,102,0,128,0,36,0,75,0,191,0,60,0,195,0,0,0,27,0,0,0,255,0,175,0,222,0,0,0,0,0,4,0,0,0,135,0,76,0,6,0,169,0,40,0,155,0,0,0,81,0,203,0,64,0,197,0,0,0,248,0,0,0,212,0,7,0,44,0,124,0,0,0,41,0,2,0,255,0,185,0,119,0,0,0,207,0,32,0,216,0,61,0,204,0,71,0,123,0,240,0,98,0,243,0,175,0,0,0,123,0,107,0,169,0,4,0,0,0,84,0,127,0,73,0,0,0,195,0,0,0,19,0,89,0,0,0,179,0,151,0,218,0,221,0,0,0,245,0,119,0,0,0,213,0,114,0,0,0,174,0,0,0,0,0,33,0,249,0,227,0,0,0,225,0,0,0,111,0,0,0,143,0,140,0,207,0,101,0,183,0,131,0,102,0,89,0,75,0,0,0,162,0,177,0,41,0,134,0,201,0,13,0,0,0,145,0,177,0,230,0,49,0,0,0,30,0,0,0,235,0,245,0,85,0,0,0,0,0,117,0,109,0,226,0,66,0,208,0,119,0,87,0,0,0,131,0,141,0,0,0,47,0,0,0,186,0,105,0,0,0,0,0,99,0,161,0,0,0,231,0,144,0,0,0,0,0,159,0,60,0,128,0,0,0,5,0,13,0,58,0,25,0,0,0,251,0,194,0,149,0,207,0,236,0,33,0,114,0,130,0,41,0,187,0,0,0,91,0,174,0,134,0,190,0,81,0,8,0,207,0,186,0,119,0,163,0,159,0,44,0,0,0,41,0,54,0,107,0,28,0,219,0,166,0,106,0,110,0,0,0,97,0,73,0,0,0,197,0,185,0,0,0,52,0,141,0,150,0,194,0,40,0,200,0,10,0,56,0,0,0,0,0,130,0,178,0,143,0,0,0,0,0,0,0,144,0,90,0,250,0,186,0,185,0,0,0,0,0,34,0,26,0,10,0,11,0,253,0,0,0,8,0,137,0,119,0,114,0,197,0,32,0,185,0,239,0,165,0,216,0,158,0,186,0,14,0,43,0,225,0,121,0,0,0,56,0,0,0,168,0,0,0,72,0,154,0,0,0,182,0,25,0,31,0,0,0,230,0,0,0,204,0,175,0,146,0,119,0,185,0,161,0,111,0,0,0,0,0,0,0,52,0,3,0,0,0,73,0,54,0,71,0,252,0,21,0,229,0,179,0,0,0,84,0,18,0,107,0,12,0,154,0,141,0,68,0,81,0,37,0,212,0,168,0,130,0,220,0,0,0,7,0,170,0,43,0,188,0,122,0,239,0,0,0,4,0,0,0,248,0,225,0,146,0,38,0,109,0,201,0,65,0,39,0,141,0,196,0,5,0,0,0,0,0,160,0,125,0,176,0,106,0,103,0,93,0,66,0,198,0,132,0,194,0,0,0,244,0,149,0,16,0,137,0,114,0,0,0,214,0,0,0,113,0,0,0,0,0,4,0,215,0,79,0,0,0,101,0,135,0,46,0,98,0,19,0,212,0,31,0,28,0,154,0,0,0,171,0,247,0,151,0,0,0,149,0,97,0,248,0,51,0,38,0,0,0,47,0,48,0,250,0,91,0,36,0,196,0,108,0,0,0,250,0,63,0,235,0,71,0,82,0,237,0,1,0,248,0,235,0,118,0,221,0,59,0,77,0,128,0,0,0,136,0,234,0,103,0,236,0,103,0,0,0,25,0,0,0,210,0,50,0,158,0,104,0,92,0,58,0,138,0,203,0,254,0,0,0,134,0,217,0,240,0,202,0,0,0,143,0,153,0,164,0,76,0,0,0,0,0,182,0,167,0,43,0,101,0,218,0,164,0,0,0,156,0,61,0,0,0,0,0,239,0,213,0,123,0,49,0,119,0,73,0,51,0,0,0,86,0,0,0,15,0,33,0,97,0,47,0,99,0,10,0,158,0,213,0,235,0,17,0,11,0,253,0,27,0,82,0,241,0,162,0,211,0,120,0,44,0,113,0,227,0,228,0,224,0,42,0,0,0,79,0,59,0,166,0,111,0,0,0,74,0,59,0,254,0,206,0,232,0,0,0,216,0,167,0,190,0,249,0,90,0,244,0,0,0,140,0,154,0,122,0,137,0,0,0,0,0,0,0,188,0,105,0,105,0,174,0,143,0,31,0,152,0,62,0,226,0,140,0,0,0,0,0,255,0,145,0,192,0,82,0,174,0,206,0,0,0,0,0,67,0,0,0,49,0,175,0,70,0,0,0,255,0,167,0,81,0,216,0,136,0,61,0,119,0,0,0,38,0,212,0,232,0,219,0,223,0,161,0,163,0,46,0,230,0,193,0,133,0,58,0,126,0,106,0,114,0,0,0,205,0,181,0,225,0,0,0,128,0,0,0,237,0,187,0,107,0,0,0,67,0,157,0,179,0,182,0,239,0,42,0,31,0,0,0,221,0,15,0,0,0,0,0,128,0,163,0,162,0,164,0,193,0,72,0,25,0,243,0,79,0,164,0,73,0,120,0,2,0,0,0,132,0,177,0,36,0,0,0,212,0,222,0,199,0,96,0,0,0,49,0,130,0,89,0,13,0,21,0,0,0,253,0,187,0,229,0,221,0,209,0,162,0,0,0,9,0,79,0,39,0,0,0,26,0,230,0,93,0,0,0,173,0,0,0,90,0,0,0,115,0,197,0,153,0,237,0,0,0,204,0,0,0,0,0,192,0,53,0,200,0,154,0,0,0,201,0,25,0,68,0,154,0,0,0,0,0,26,0,10,0,16,0,149,0,192,0,0,0,235,0,246,0,0,0,221,0,111,0,164,0,0,0,155,0,0,0,0,0,74,0,246,0,251,0,0,0,0,0,0,0,76,0,220,0,182,0,91,0,86,0,0,0,184,0,210,0,198,0,23,0,6,0,100,0,144,0,49,0,233,0,0,0,166,0,104,0,0,0,26,0,152,0,160,0,0,0,179,0,18,0,180,0,54,0,112,0,0,0,137,0,210,0,4,0,229,0,89,0,215,0,21,0,132,0,87,0,235,0,113,0,254,0,164,0,0,0,159,0,85,0,242,0,246,0,170,0,0,0,111,0,59,0,0,0,0,0,0,0,116,0,139,0,0,0,19,0,13,0,107,0,51,0,246,0,103,0,63,0,238,0,203,0,224,0,110,0,232,0,240,0,0,0,227,0,253,0,187,0,0,0,137,0,129,0,154,0,85,0,193,0,77,0,211,0,19,0,0,0,0,0,114,0,120,0,149,0,215,0,82,0,132,0,70,0,249,0,0,0,201,0,173,0,159,0,0,0,14,0,7,0,96,0,35,0,195,0,161,0,79,0,164,0,0,0,72,0,139,0,35,0,198,0,236,0,130,0,55,0,32,0,224,0,56,0,20,0,254,0,108,0,79,0,41,0,230,0,248,0,35,0,197,0,224,0,158,0,0,0,0,0,141,0,187,0,0,0,0,0,247,0,50,0,0,0,173,0,190,0,196,0,95,0,0,0,150,0,29,0,251,0,44,0,0,0,214,0,245,0,57,0,204,0,117,0,0,0,232,0,117,0,117,0,0,0,0,0,0,0,172,0,159,0,102,0,0,0,120,0,216,0,22,0,87,0,159,0,7,0,0,0,70,0,19,0,5,0,0,0,0,0,127,0,45,0,0,0,15,0,65,0,196,0,133,0,119,0,1,0,34,0,162,0,87,0,134,0,68,0,151,0,22,0,148,0,52,0,140,0,0,0,101,0,163,0,63,0,99,0,8,0,0,0,223,0,217,0,12,0,6,0,0,0,178,0,90,0,0,0);
signal scenario_full  : scenario_type := (0,0,121,31,121,30,62,31,134,31,102,31,128,31,36,31,75,31,191,31,60,31,195,31,195,30,27,31,27,30,255,31,175,31,222,31,222,30,222,29,4,31,4,30,135,31,76,31,6,31,169,31,40,31,155,31,155,30,81,31,203,31,64,31,197,31,197,30,248,31,248,30,212,31,7,31,44,31,124,31,124,30,41,31,2,31,255,31,185,31,119,31,119,30,207,31,32,31,216,31,61,31,204,31,71,31,123,31,240,31,98,31,243,31,175,31,175,30,123,31,107,31,169,31,4,31,4,30,84,31,127,31,73,31,73,30,195,31,195,30,19,31,89,31,89,30,179,31,151,31,218,31,221,31,221,30,245,31,119,31,119,30,213,31,114,31,114,30,174,31,174,30,174,29,33,31,249,31,227,31,227,30,225,31,225,30,111,31,111,30,143,31,140,31,207,31,101,31,183,31,131,31,102,31,89,31,75,31,75,30,162,31,177,31,41,31,134,31,201,31,13,31,13,30,145,31,177,31,230,31,49,31,49,30,30,31,30,30,235,31,245,31,85,31,85,30,85,29,117,31,109,31,226,31,66,31,208,31,119,31,87,31,87,30,131,31,141,31,141,30,47,31,47,30,186,31,105,31,105,30,105,29,99,31,161,31,161,30,231,31,144,31,144,30,144,29,159,31,60,31,128,31,128,30,5,31,13,31,58,31,25,31,25,30,251,31,194,31,149,31,207,31,236,31,33,31,114,31,130,31,41,31,187,31,187,30,91,31,174,31,134,31,190,31,81,31,8,31,207,31,186,31,119,31,163,31,159,31,44,31,44,30,41,31,54,31,107,31,28,31,219,31,166,31,106,31,110,31,110,30,97,31,73,31,73,30,197,31,185,31,185,30,52,31,141,31,150,31,194,31,40,31,200,31,10,31,56,31,56,30,56,29,130,31,178,31,143,31,143,30,143,29,143,28,144,31,90,31,250,31,186,31,185,31,185,30,185,29,34,31,26,31,10,31,11,31,253,31,253,30,8,31,137,31,119,31,114,31,197,31,32,31,185,31,239,31,165,31,216,31,158,31,186,31,14,31,43,31,225,31,121,31,121,30,56,31,56,30,168,31,168,30,72,31,154,31,154,30,182,31,25,31,31,31,31,30,230,31,230,30,204,31,175,31,146,31,119,31,185,31,161,31,111,31,111,30,111,29,111,28,52,31,3,31,3,30,73,31,54,31,71,31,252,31,21,31,229,31,179,31,179,30,84,31,18,31,107,31,12,31,154,31,141,31,68,31,81,31,37,31,212,31,168,31,130,31,220,31,220,30,7,31,170,31,43,31,188,31,122,31,239,31,239,30,4,31,4,30,248,31,225,31,146,31,38,31,109,31,201,31,65,31,39,31,141,31,196,31,5,31,5,30,5,29,160,31,125,31,176,31,106,31,103,31,93,31,66,31,198,31,132,31,194,31,194,30,244,31,149,31,16,31,137,31,114,31,114,30,214,31,214,30,113,31,113,30,113,29,4,31,215,31,79,31,79,30,101,31,135,31,46,31,98,31,19,31,212,31,31,31,28,31,154,31,154,30,171,31,247,31,151,31,151,30,149,31,97,31,248,31,51,31,38,31,38,30,47,31,48,31,250,31,91,31,36,31,196,31,108,31,108,30,250,31,63,31,235,31,71,31,82,31,237,31,1,31,248,31,235,31,118,31,221,31,59,31,77,31,128,31,128,30,136,31,234,31,103,31,236,31,103,31,103,30,25,31,25,30,210,31,50,31,158,31,104,31,92,31,58,31,138,31,203,31,254,31,254,30,134,31,217,31,240,31,202,31,202,30,143,31,153,31,164,31,76,31,76,30,76,29,182,31,167,31,43,31,101,31,218,31,164,31,164,30,156,31,61,31,61,30,61,29,239,31,213,31,123,31,49,31,119,31,73,31,51,31,51,30,86,31,86,30,15,31,33,31,97,31,47,31,99,31,10,31,158,31,213,31,235,31,17,31,11,31,253,31,27,31,82,31,241,31,162,31,211,31,120,31,44,31,113,31,227,31,228,31,224,31,42,31,42,30,79,31,59,31,166,31,111,31,111,30,74,31,59,31,254,31,206,31,232,31,232,30,216,31,167,31,190,31,249,31,90,31,244,31,244,30,140,31,154,31,122,31,137,31,137,30,137,29,137,28,188,31,105,31,105,31,174,31,143,31,31,31,152,31,62,31,226,31,140,31,140,30,140,29,255,31,145,31,192,31,82,31,174,31,206,31,206,30,206,29,67,31,67,30,49,31,175,31,70,31,70,30,255,31,167,31,81,31,216,31,136,31,61,31,119,31,119,30,38,31,212,31,232,31,219,31,223,31,161,31,163,31,46,31,230,31,193,31,133,31,58,31,126,31,106,31,114,31,114,30,205,31,181,31,225,31,225,30,128,31,128,30,237,31,187,31,107,31,107,30,67,31,157,31,179,31,182,31,239,31,42,31,31,31,31,30,221,31,15,31,15,30,15,29,128,31,163,31,162,31,164,31,193,31,72,31,25,31,243,31,79,31,164,31,73,31,120,31,2,31,2,30,132,31,177,31,36,31,36,30,212,31,222,31,199,31,96,31,96,30,49,31,130,31,89,31,13,31,21,31,21,30,253,31,187,31,229,31,221,31,209,31,162,31,162,30,9,31,79,31,39,31,39,30,26,31,230,31,93,31,93,30,173,31,173,30,90,31,90,30,115,31,197,31,153,31,237,31,237,30,204,31,204,30,204,29,192,31,53,31,200,31,154,31,154,30,201,31,25,31,68,31,154,31,154,30,154,29,26,31,10,31,16,31,149,31,192,31,192,30,235,31,246,31,246,30,221,31,111,31,164,31,164,30,155,31,155,30,155,29,74,31,246,31,251,31,251,30,251,29,251,28,76,31,220,31,182,31,91,31,86,31,86,30,184,31,210,31,198,31,23,31,6,31,100,31,144,31,49,31,233,31,233,30,166,31,104,31,104,30,26,31,152,31,160,31,160,30,179,31,18,31,180,31,54,31,112,31,112,30,137,31,210,31,4,31,229,31,89,31,215,31,21,31,132,31,87,31,235,31,113,31,254,31,164,31,164,30,159,31,85,31,242,31,246,31,170,31,170,30,111,31,59,31,59,30,59,29,59,28,116,31,139,31,139,30,19,31,13,31,107,31,51,31,246,31,103,31,63,31,238,31,203,31,224,31,110,31,232,31,240,31,240,30,227,31,253,31,187,31,187,30,137,31,129,31,154,31,85,31,193,31,77,31,211,31,19,31,19,30,19,29,114,31,120,31,149,31,215,31,82,31,132,31,70,31,249,31,249,30,201,31,173,31,159,31,159,30,14,31,7,31,96,31,35,31,195,31,161,31,79,31,164,31,164,30,72,31,139,31,35,31,198,31,236,31,130,31,55,31,32,31,224,31,56,31,20,31,254,31,108,31,79,31,41,31,230,31,248,31,35,31,197,31,224,31,158,31,158,30,158,29,141,31,187,31,187,30,187,29,247,31,50,31,50,30,173,31,190,31,196,31,95,31,95,30,150,31,29,31,251,31,44,31,44,30,214,31,245,31,57,31,204,31,117,31,117,30,232,31,117,31,117,31,117,30,117,29,117,28,172,31,159,31,102,31,102,30,120,31,216,31,22,31,87,31,159,31,7,31,7,30,70,31,19,31,5,31,5,30,5,29,127,31,45,31,45,30,15,31,65,31,196,31,133,31,119,31,1,31,34,31,162,31,87,31,134,31,68,31,151,31,22,31,148,31,52,31,140,31,140,30,101,31,163,31,63,31,99,31,8,31,8,30,223,31,217,31,12,31,6,31,6,30,178,31,90,31,90,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
