-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 958;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,191,0,85,0,143,0,78,0,0,0,3,0,103,0,28,0,200,0,196,0,90,0,202,0,251,0,40,0,46,0,239,0,111,0,249,0,235,0,178,0,200,0,0,0,221,0,21,0,127,0,145,0,253,0,218,0,178,0,117,0,0,0,104,0,190,0,105,0,178,0,0,0,153,0,158,0,21,0,214,0,134,0,27,0,20,0,0,0,158,0,21,0,13,0,0,0,142,0,144,0,12,0,147,0,63,0,244,0,164,0,0,0,29,0,240,0,0,0,7,0,115,0,126,0,83,0,244,0,0,0,241,0,114,0,143,0,138,0,0,0,0,0,7,0,159,0,0,0,214,0,134,0,134,0,0,0,202,0,0,0,156,0,253,0,246,0,161,0,146,0,52,0,149,0,0,0,11,0,181,0,105,0,224,0,0,0,82,0,106,0,64,0,0,0,1,0,0,0,173,0,130,0,0,0,53,0,76,0,123,0,120,0,21,0,153,0,156,0,66,0,126,0,69,0,176,0,254,0,148,0,136,0,0,0,40,0,137,0,215,0,88,0,100,0,14,0,206,0,9,0,58,0,0,0,67,0,186,0,140,0,179,0,31,0,50,0,0,0,220,0,0,0,40,0,0,0,0,0,25,0,0,0,14,0,0,0,0,0,239,0,92,0,232,0,229,0,248,0,0,0,122,0,0,0,53,0,142,0,0,0,168,0,186,0,226,0,59,0,210,0,0,0,227,0,209,0,43,0,229,0,49,0,239,0,24,0,188,0,211,0,58,0,210,0,192,0,9,0,159,0,63,0,146,0,114,0,43,0,150,0,133,0,128,0,53,0,128,0,0,0,98,0,130,0,0,0,0,0,225,0,107,0,139,0,77,0,135,0,236,0,43,0,106,0,210,0,55,0,54,0,117,0,216,0,0,0,0,0,96,0,184,0,233,0,39,0,51,0,108,0,229,0,107,0,161,0,0,0,0,0,24,0,62,0,220,0,197,0,0,0,248,0,48,0,143,0,17,0,116,0,0,0,113,0,134,0,194,0,156,0,0,0,103,0,244,0,70,0,35,0,130,0,104,0,28,0,168,0,74,0,248,0,34,0,0,0,223,0,180,0,134,0,126,0,171,0,0,0,101,0,174,0,0,0,108,0,67,0,255,0,19,0,0,0,68,0,137,0,0,0,49,0,36,0,185,0,72,0,71,0,188,0,225,0,254,0,169,0,0,0,0,0,37,0,159,0,172,0,46,0,0,0,0,0,0,0,39,0,23,0,186,0,0,0,84,0,106,0,65,0,29,0,0,0,0,0,205,0,246,0,227,0,243,0,199,0,174,0,0,0,156,0,0,0,236,0,63,0,227,0,70,0,84,0,98,0,9,0,53,0,38,0,255,0,83,0,0,0,217,0,221,0,83,0,75,0,149,0,160,0,0,0,80,0,46,0,180,0,0,0,181,0,0,0,157,0,141,0,84,0,168,0,0,0,157,0,109,0,241,0,86,0,79,0,167,0,177,0,7,0,95,0,224,0,0,0,233,0,203,0,0,0,195,0,81,0,45,0,168,0,64,0,91,0,169,0,19,0,122,0,10,0,0,0,186,0,28,0,72,0,231,0,120,0,0,0,0,0,90,0,123,0,26,0,195,0,30,0,237,0,67,0,169,0,62,0,0,0,245,0,167,0,130,0,50,0,112,0,45,0,113,0,84,0,112,0,0,0,196,0,150,0,89,0,255,0,106,0,130,0,44,0,10,0,179,0,0,0,88,0,182,0,71,0,215,0,62,0,0,0,73,0,118,0,143,0,228,0,198,0,98,0,36,0,70,0,230,0,214,0,0,0,239,0,100,0,0,0,184,0,53,0,0,0,179,0,195,0,244,0,252,0,21,0,121,0,157,0,0,0,0,0,96,0,136,0,232,0,33,0,78,0,70,0,171,0,62,0,206,0,251,0,3,0,189,0,252,0,120,0,0,0,0,0,195,0,1,0,132,0,129,0,19,0,72,0,127,0,0,0,15,0,161,0,0,0,0,0,109,0,192,0,180,0,196,0,16,0,0,0,204,0,242,0,211,0,0,0,170,0,107,0,43,0,42,0,61,0,93,0,44,0,144,0,229,0,52,0,75,0,111,0,184,0,124,0,235,0,0,0,245,0,38,0,195,0,180,0,233,0,255,0,250,0,192,0,31,0,0,0,48,0,243,0,94,0,172,0,201,0,94,0,55,0,156,0,33,0,92,0,39,0,133,0,200,0,121,0,78,0,16,0,231,0,0,0,169,0,150,0,143,0,240,0,0,0,59,0,93,0,197,0,0,0,194,0,115,0,71,0,0,0,0,0,220,0,7,0,226,0,47,0,0,0,201,0,0,0,184,0,0,0,249,0,0,0,158,0,254,0,50,0,150,0,88,0,34,0,0,0,0,0,3,0,238,0,0,0,123,0,68,0,4,0,0,0,54,0,30,0,0,0,67,0,227,0,157,0,168,0,193,0,246,0,19,0,0,0,0,0,147,0,249,0,0,0,64,0,0,0,116,0,0,0,0,0,217,0,27,0,97,0,192,0,254,0,255,0,0,0,0,0,74,0,221,0,91,0,0,0,0,0,19,0,231,0,12,0,54,0,240,0,120,0,225,0,91,0,252,0,59,0,0,0,0,0,251,0,77,0,0,0,55,0,131,0,226,0,68,0,74,0,198,0,26,0,39,0,19,0,132,0,168,0,190,0,186,0,198,0,45,0,125,0,37,0,35,0,27,0,0,0,7,0,185,0,141,0,40,0,0,0,172,0,146,0,74,0,140,0,0,0,243,0,229,0,0,0,250,0,0,0,40,0,226,0,223,0,0,0,0,0,0,0,120,0,0,0,47,0,0,0,0,0,15,0,156,0,198,0,40,0,231,0,124,0,250,0,106,0,170,0,218,0,237,0,83,0,0,0,174,0,148,0,64,0,145,0,0,0,183,0,217,0,0,0,164,0,0,0,9,0,168,0,54,0,40,0,68,0,127,0,184,0,24,0,209,0,0,0,27,0,25,0,28,0,0,0,190,0,178,0,46,0,28,0,111,0,129,0,0,0,21,0,131,0,102,0,198,0,212,0,212,0,139,0,161,0,0,0,104,0,28,0,0,0,245,0,178,0,204,0,82,0,207,0,185,0,125,0,167,0,33,0,0,0,197,0,124,0,200,0,106,0,17,0,169,0,0,0,195,0,125,0,237,0,0,0,224,0,229,0,140,0,140,0,0,0,0,0,236,0,64,0,64,0,0,0,31,0,174,0,204,0,0,0,7,0,68,0,0,0,70,0,75,0,223,0,80,0,247,0,11,0,10,0,0,0,158,0,97,0,210,0,50,0,30,0,201,0,113,0,198,0,196,0,177,0,78,0,0,0,81,0,213,0,47,0,11,0,112,0,163,0,180,0,136,0,42,0,242,0,0,0,253,0,192,0,0,0,37,0,28,0,210,0,231,0,53,0,0,0,183,0,145,0,116,0,0,0,0,0,148,0,170,0,5,0,230,0,221,0,53,0,74,0,27,0,144,0,209,0,90,0,175,0,73,0,143,0,147,0,54,0,163,0,186,0,194,0,0,0,0,0,66,0,227,0,71,0,0,0,83,0,79,0,229,0,0,0,6,0,17,0,0,0,121,0,137,0,150,0,0,0,56,0,93,0,0,0,64,0,205,0,0,0,237,0,0,0,15,0,89,0,157,0,0,0,123,0,0,0,38,0,15,0,0,0,13,0,15,0,181,0,124,0,0,0,53,0,228,0,0,0,215,0,16,0,169,0,39,0,246,0,20,0,0,0,25,0,230,0,63,0,0,0,13,0,241,0,13,0,132,0,3,0,0,0,123,0,130,0,223,0,3,0,11,0,167,0,199,0,0,0,88,0,180,0,0,0,235,0,243,0,0,0,23,0,124,0,35,0,0,0,0,0,162,0,148,0,175,0,0,0,160,0,167,0,238,0,225,0,21,0,157,0,217,0,184,0,126,0,252,0,174,0,179,0,39,0,48,0,0,0,215,0,22,0,118,0,0,0,245,0,162,0,195,0,184,0,63,0,175,0,4,0,0,0,0,0,183,0,0,0,24,0,56,0,182,0,0,0,168,0,0,0,185,0,243,0,0,0,54,0,236,0,0,0,68,0,253,0,0,0,66,0,0,0,132,0,0,0,165,0,34,0,0,0,118,0,7,0,0,0,192,0,171,0,172,0,0,0,124,0,156,0,55,0,134,0,0,0,7,0,230,0,0,0,147,0,166,0,190,0,0,0,197,0,227,0,125,0,229,0,223,0,64,0,10,0,79,0,219,0);
signal scenario_full  : scenario_type := (56,31,191,31,85,31,143,31,78,31,78,30,3,31,103,31,28,31,200,31,196,31,90,31,202,31,251,31,40,31,46,31,239,31,111,31,249,31,235,31,178,31,200,31,200,30,221,31,21,31,127,31,145,31,253,31,218,31,178,31,117,31,117,30,104,31,190,31,105,31,178,31,178,30,153,31,158,31,21,31,214,31,134,31,27,31,20,31,20,30,158,31,21,31,13,31,13,30,142,31,144,31,12,31,147,31,63,31,244,31,164,31,164,30,29,31,240,31,240,30,7,31,115,31,126,31,83,31,244,31,244,30,241,31,114,31,143,31,138,31,138,30,138,29,7,31,159,31,159,30,214,31,134,31,134,31,134,30,202,31,202,30,156,31,253,31,246,31,161,31,146,31,52,31,149,31,149,30,11,31,181,31,105,31,224,31,224,30,82,31,106,31,64,31,64,30,1,31,1,30,173,31,130,31,130,30,53,31,76,31,123,31,120,31,21,31,153,31,156,31,66,31,126,31,69,31,176,31,254,31,148,31,136,31,136,30,40,31,137,31,215,31,88,31,100,31,14,31,206,31,9,31,58,31,58,30,67,31,186,31,140,31,179,31,31,31,50,31,50,30,220,31,220,30,40,31,40,30,40,29,25,31,25,30,14,31,14,30,14,29,239,31,92,31,232,31,229,31,248,31,248,30,122,31,122,30,53,31,142,31,142,30,168,31,186,31,226,31,59,31,210,31,210,30,227,31,209,31,43,31,229,31,49,31,239,31,24,31,188,31,211,31,58,31,210,31,192,31,9,31,159,31,63,31,146,31,114,31,43,31,150,31,133,31,128,31,53,31,128,31,128,30,98,31,130,31,130,30,130,29,225,31,107,31,139,31,77,31,135,31,236,31,43,31,106,31,210,31,55,31,54,31,117,31,216,31,216,30,216,29,96,31,184,31,233,31,39,31,51,31,108,31,229,31,107,31,161,31,161,30,161,29,24,31,62,31,220,31,197,31,197,30,248,31,48,31,143,31,17,31,116,31,116,30,113,31,134,31,194,31,156,31,156,30,103,31,244,31,70,31,35,31,130,31,104,31,28,31,168,31,74,31,248,31,34,31,34,30,223,31,180,31,134,31,126,31,171,31,171,30,101,31,174,31,174,30,108,31,67,31,255,31,19,31,19,30,68,31,137,31,137,30,49,31,36,31,185,31,72,31,71,31,188,31,225,31,254,31,169,31,169,30,169,29,37,31,159,31,172,31,46,31,46,30,46,29,46,28,39,31,23,31,186,31,186,30,84,31,106,31,65,31,29,31,29,30,29,29,205,31,246,31,227,31,243,31,199,31,174,31,174,30,156,31,156,30,236,31,63,31,227,31,70,31,84,31,98,31,9,31,53,31,38,31,255,31,83,31,83,30,217,31,221,31,83,31,75,31,149,31,160,31,160,30,80,31,46,31,180,31,180,30,181,31,181,30,157,31,141,31,84,31,168,31,168,30,157,31,109,31,241,31,86,31,79,31,167,31,177,31,7,31,95,31,224,31,224,30,233,31,203,31,203,30,195,31,81,31,45,31,168,31,64,31,91,31,169,31,19,31,122,31,10,31,10,30,186,31,28,31,72,31,231,31,120,31,120,30,120,29,90,31,123,31,26,31,195,31,30,31,237,31,67,31,169,31,62,31,62,30,245,31,167,31,130,31,50,31,112,31,45,31,113,31,84,31,112,31,112,30,196,31,150,31,89,31,255,31,106,31,130,31,44,31,10,31,179,31,179,30,88,31,182,31,71,31,215,31,62,31,62,30,73,31,118,31,143,31,228,31,198,31,98,31,36,31,70,31,230,31,214,31,214,30,239,31,100,31,100,30,184,31,53,31,53,30,179,31,195,31,244,31,252,31,21,31,121,31,157,31,157,30,157,29,96,31,136,31,232,31,33,31,78,31,70,31,171,31,62,31,206,31,251,31,3,31,189,31,252,31,120,31,120,30,120,29,195,31,1,31,132,31,129,31,19,31,72,31,127,31,127,30,15,31,161,31,161,30,161,29,109,31,192,31,180,31,196,31,16,31,16,30,204,31,242,31,211,31,211,30,170,31,107,31,43,31,42,31,61,31,93,31,44,31,144,31,229,31,52,31,75,31,111,31,184,31,124,31,235,31,235,30,245,31,38,31,195,31,180,31,233,31,255,31,250,31,192,31,31,31,31,30,48,31,243,31,94,31,172,31,201,31,94,31,55,31,156,31,33,31,92,31,39,31,133,31,200,31,121,31,78,31,16,31,231,31,231,30,169,31,150,31,143,31,240,31,240,30,59,31,93,31,197,31,197,30,194,31,115,31,71,31,71,30,71,29,220,31,7,31,226,31,47,31,47,30,201,31,201,30,184,31,184,30,249,31,249,30,158,31,254,31,50,31,150,31,88,31,34,31,34,30,34,29,3,31,238,31,238,30,123,31,68,31,4,31,4,30,54,31,30,31,30,30,67,31,227,31,157,31,168,31,193,31,246,31,19,31,19,30,19,29,147,31,249,31,249,30,64,31,64,30,116,31,116,30,116,29,217,31,27,31,97,31,192,31,254,31,255,31,255,30,255,29,74,31,221,31,91,31,91,30,91,29,19,31,231,31,12,31,54,31,240,31,120,31,225,31,91,31,252,31,59,31,59,30,59,29,251,31,77,31,77,30,55,31,131,31,226,31,68,31,74,31,198,31,26,31,39,31,19,31,132,31,168,31,190,31,186,31,198,31,45,31,125,31,37,31,35,31,27,31,27,30,7,31,185,31,141,31,40,31,40,30,172,31,146,31,74,31,140,31,140,30,243,31,229,31,229,30,250,31,250,30,40,31,226,31,223,31,223,30,223,29,223,28,120,31,120,30,47,31,47,30,47,29,15,31,156,31,198,31,40,31,231,31,124,31,250,31,106,31,170,31,218,31,237,31,83,31,83,30,174,31,148,31,64,31,145,31,145,30,183,31,217,31,217,30,164,31,164,30,9,31,168,31,54,31,40,31,68,31,127,31,184,31,24,31,209,31,209,30,27,31,25,31,28,31,28,30,190,31,178,31,46,31,28,31,111,31,129,31,129,30,21,31,131,31,102,31,198,31,212,31,212,31,139,31,161,31,161,30,104,31,28,31,28,30,245,31,178,31,204,31,82,31,207,31,185,31,125,31,167,31,33,31,33,30,197,31,124,31,200,31,106,31,17,31,169,31,169,30,195,31,125,31,237,31,237,30,224,31,229,31,140,31,140,31,140,30,140,29,236,31,64,31,64,31,64,30,31,31,174,31,204,31,204,30,7,31,68,31,68,30,70,31,75,31,223,31,80,31,247,31,11,31,10,31,10,30,158,31,97,31,210,31,50,31,30,31,201,31,113,31,198,31,196,31,177,31,78,31,78,30,81,31,213,31,47,31,11,31,112,31,163,31,180,31,136,31,42,31,242,31,242,30,253,31,192,31,192,30,37,31,28,31,210,31,231,31,53,31,53,30,183,31,145,31,116,31,116,30,116,29,148,31,170,31,5,31,230,31,221,31,53,31,74,31,27,31,144,31,209,31,90,31,175,31,73,31,143,31,147,31,54,31,163,31,186,31,194,31,194,30,194,29,66,31,227,31,71,31,71,30,83,31,79,31,229,31,229,30,6,31,17,31,17,30,121,31,137,31,150,31,150,30,56,31,93,31,93,30,64,31,205,31,205,30,237,31,237,30,15,31,89,31,157,31,157,30,123,31,123,30,38,31,15,31,15,30,13,31,15,31,181,31,124,31,124,30,53,31,228,31,228,30,215,31,16,31,169,31,39,31,246,31,20,31,20,30,25,31,230,31,63,31,63,30,13,31,241,31,13,31,132,31,3,31,3,30,123,31,130,31,223,31,3,31,11,31,167,31,199,31,199,30,88,31,180,31,180,30,235,31,243,31,243,30,23,31,124,31,35,31,35,30,35,29,162,31,148,31,175,31,175,30,160,31,167,31,238,31,225,31,21,31,157,31,217,31,184,31,126,31,252,31,174,31,179,31,39,31,48,31,48,30,215,31,22,31,118,31,118,30,245,31,162,31,195,31,184,31,63,31,175,31,4,31,4,30,4,29,183,31,183,30,24,31,56,31,182,31,182,30,168,31,168,30,185,31,243,31,243,30,54,31,236,31,236,30,68,31,253,31,253,30,66,31,66,30,132,31,132,30,165,31,34,31,34,30,118,31,7,31,7,30,192,31,171,31,172,31,172,30,124,31,156,31,55,31,134,31,134,30,7,31,230,31,230,30,147,31,166,31,190,31,190,30,197,31,227,31,125,31,229,31,223,31,64,31,10,31,79,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
