-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 261;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,208,0,134,0,0,0,159,0,0,0,249,0,0,0,91,0,229,0,214,0,130,0,148,0,189,0,229,0,0,0,85,0,69,0,219,0,0,0,217,0,221,0,142,0,230,0,45,0,47,0,0,0,0,0,26,0,226,0,30,0,175,0,94,0,172,0,5,0,0,0,124,0,7,0,237,0,41,0,26,0,252,0,235,0,0,0,0,0,114,0,145,0,229,0,242,0,0,0,224,0,0,0,48,0,3,0,173,0,190,0,0,0,244,0,184,0,91,0,130,0,195,0,136,0,0,0,242,0,0,0,0,0,39,0,191,0,160,0,0,0,0,0,64,0,250,0,195,0,27,0,110,0,0,0,218,0,169,0,15,0,139,0,142,0,0,0,0,0,192,0,114,0,179,0,176,0,94,0,163,0,222,0,0,0,157,0,11,0,208,0,189,0,158,0,0,0,222,0,212,0,156,0,237,0,184,0,222,0,242,0,0,0,77,0,154,0,0,0,37,0,0,0,255,0,12,0,244,0,184,0,156,0,77,0,27,0,14,0,234,0,0,0,1,0,123,0,158,0,177,0,15,0,213,0,252,0,0,0,65,0,82,0,0,0,86,0,174,0,111,0,51,0,83,0,55,0,218,0,0,0,177,0,94,0,107,0,246,0,0,0,17,0,190,0,139,0,27,0,0,0,14,0,0,0,151,0,82,0,125,0,124,0,147,0,31,0,0,0,250,0,60,0,115,0,232,0,126,0,122,0,201,0,0,0,0,0,184,0,90,0,108,0,0,0,117,0,61,0,151,0,43,0,0,0,136,0,149,0,0,0,0,0,199,0,110,0,221,0,100,0,43,0,225,0,222,0,109,0,147,0,182,0,197,0,207,0,1,0,0,0,36,0,102,0,248,0,108,0,13,0,0,0,0,0,151,0,145,0,126,0,105,0,234,0,0,0,197,0,0,0,87,0,91,0,133,0,0,0,0,0,7,0,0,0,18,0,114,0,192,0,75,0,229,0,76,0,21,0,0,0,120,0,58,0,124,0,29,0,173,0,0,0,191,0,204,0,175,0,111,0,24,0,243,0,81,0,94,0,190,0,33,0,104,0,95,0,123,0,238,0,0,0,0,0,137,0,167,0,213,0,77,0,0,0,157,0,33,0,0,0,214,0,199,0,73,0,241,0,156,0);
signal scenario_full  : scenario_type := (0,0,208,31,134,31,134,30,159,31,159,30,249,31,249,30,91,31,229,31,214,31,130,31,148,31,189,31,229,31,229,30,85,31,69,31,219,31,219,30,217,31,221,31,142,31,230,31,45,31,47,31,47,30,47,29,26,31,226,31,30,31,175,31,94,31,172,31,5,31,5,30,124,31,7,31,237,31,41,31,26,31,252,31,235,31,235,30,235,29,114,31,145,31,229,31,242,31,242,30,224,31,224,30,48,31,3,31,173,31,190,31,190,30,244,31,184,31,91,31,130,31,195,31,136,31,136,30,242,31,242,30,242,29,39,31,191,31,160,31,160,30,160,29,64,31,250,31,195,31,27,31,110,31,110,30,218,31,169,31,15,31,139,31,142,31,142,30,142,29,192,31,114,31,179,31,176,31,94,31,163,31,222,31,222,30,157,31,11,31,208,31,189,31,158,31,158,30,222,31,212,31,156,31,237,31,184,31,222,31,242,31,242,30,77,31,154,31,154,30,37,31,37,30,255,31,12,31,244,31,184,31,156,31,77,31,27,31,14,31,234,31,234,30,1,31,123,31,158,31,177,31,15,31,213,31,252,31,252,30,65,31,82,31,82,30,86,31,174,31,111,31,51,31,83,31,55,31,218,31,218,30,177,31,94,31,107,31,246,31,246,30,17,31,190,31,139,31,27,31,27,30,14,31,14,30,151,31,82,31,125,31,124,31,147,31,31,31,31,30,250,31,60,31,115,31,232,31,126,31,122,31,201,31,201,30,201,29,184,31,90,31,108,31,108,30,117,31,61,31,151,31,43,31,43,30,136,31,149,31,149,30,149,29,199,31,110,31,221,31,100,31,43,31,225,31,222,31,109,31,147,31,182,31,197,31,207,31,1,31,1,30,36,31,102,31,248,31,108,31,13,31,13,30,13,29,151,31,145,31,126,31,105,31,234,31,234,30,197,31,197,30,87,31,91,31,133,31,133,30,133,29,7,31,7,30,18,31,114,31,192,31,75,31,229,31,76,31,21,31,21,30,120,31,58,31,124,31,29,31,173,31,173,30,191,31,204,31,175,31,111,31,24,31,243,31,81,31,94,31,190,31,33,31,104,31,95,31,123,31,238,31,238,30,238,29,137,31,167,31,213,31,77,31,77,30,157,31,33,31,33,30,214,31,199,31,73,31,241,31,156,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
