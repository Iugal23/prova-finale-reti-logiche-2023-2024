-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 492;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (216,0,151,0,36,0,121,0,11,0,91,0,213,0,246,0,0,0,161,0,5,0,87,0,173,0,177,0,9,0,0,0,43,0,24,0,0,0,84,0,72,0,154,0,72,0,194,0,152,0,128,0,53,0,132,0,0,0,84,0,100,0,78,0,85,0,180,0,105,0,19,0,227,0,237,0,149,0,245,0,0,0,0,0,54,0,239,0,187,0,226,0,192,0,155,0,0,0,65,0,181,0,28,0,89,0,93,0,138,0,176,0,58,0,182,0,39,0,0,0,168,0,126,0,51,0,185,0,0,0,207,0,128,0,0,0,246,0,146,0,189,0,0,0,8,0,163,0,0,0,54,0,134,0,178,0,114,0,169,0,110,0,239,0,187,0,136,0,232,0,249,0,144,0,0,0,0,0,101,0,225,0,0,0,0,0,202,0,16,0,207,0,17,0,0,0,141,0,0,0,240,0,87,0,85,0,0,0,0,0,121,0,248,0,160,0,0,0,0,0,195,0,22,0,105,0,49,0,71,0,0,0,74,0,130,0,131,0,0,0,192,0,118,0,112,0,165,0,98,0,40,0,1,0,0,0,145,0,0,0,87,0,98,0,234,0,245,0,0,0,235,0,210,0,211,0,199,0,175,0,88,0,230,0,65,0,99,0,61,0,48,0,0,0,121,0,15,0,128,0,185,0,70,0,122,0,60,0,229,0,150,0,0,0,200,0,0,0,189,0,220,0,146,0,0,0,62,0,179,0,138,0,75,0,126,0,47,0,50,0,113,0,168,0,95,0,3,0,0,0,128,0,0,0,209,0,96,0,1,0,25,0,4,0,237,0,27,0,227,0,0,0,245,0,242,0,151,0,141,0,134,0,231,0,24,0,105,0,0,0,22,0,142,0,212,0,23,0,2,0,0,0,249,0,53,0,213,0,59,0,237,0,18,0,135,0,37,0,0,0,50,0,218,0,196,0,85,0,86,0,47,0,113,0,189,0,0,0,251,0,56,0,55,0,0,0,185,0,223,0,207,0,117,0,0,0,202,0,234,0,209,0,252,0,0,0,19,0,188,0,4,0,147,0,0,0,102,0,53,0,19,0,2,0,248,0,232,0,0,0,0,0,162,0,17,0,148,0,69,0,59,0,165,0,0,0,0,0,104,0,70,0,0,0,220,0,72,0,251,0,0,0,209,0,0,0,100,0,178,0,0,0,84,0,161,0,238,0,94,0,202,0,218,0,0,0,98,0,249,0,49,0,102,0,216,0,157,0,76,0,65,0,54,0,12,0,122,0,85,0,225,0,27,0,44,0,167,0,200,0,143,0,63,0,145,0,85,0,161,0,89,0,0,0,197,0,0,0,41,0,0,0,239,0,32,0,226,0,222,0,126,0,220,0,5,0,247,0,108,0,68,0,48,0,174,0,0,0,138,0,0,0,114,0,0,0,178,0,0,0,140,0,0,0,119,0,5,0,189,0,214,0,63,0,78,0,227,0,186,0,104,0,231,0,0,0,5,0,23,0,66,0,216,0,49,0,150,0,196,0,15,0,19,0,60,0,150,0,0,0,0,0,253,0,78,0,135,0,0,0,238,0,0,0,186,0,252,0,14,0,121,0,0,0,147,0,246,0,45,0,0,0,152,0,252,0,1,0,0,0,122,0,22,0,232,0,0,0,124,0,136,0,0,0,0,0,35,0,123,0,150,0,0,0,241,0,196,0,245,0,76,0,242,0,174,0,0,0,69,0,183,0,143,0,124,0,52,0,0,0,44,0,227,0,67,0,243,0,171,0,240,0,40,0,110,0,96,0,0,0,216,0,90,0,53,0,197,0,111,0,0,0,0,0,39,0,116,0,31,0,177,0,236,0,0,0,210,0,165,0,217,0,126,0,16,0,156,0,88,0,0,0,178,0,124,0,92,0,148,0,46,0,141,0,0,0,83,0,209,0,146,0,0,0,77,0,2,0,178,0,184,0,176,0,182,0,197,0,59,0,9,0,191,0,142,0,63,0,172,0,247,0,232,0,159,0,80,0,72,0,3,0,130,0,102,0,1,0,237,0,0,0,39,0,100,0,73,0,0,0,148,0,245,0,171,0,164,0,170,0,219,0,0,0,123,0,252,0,99,0,244,0,22,0,248,0,0,0,242,0,130,0,27,0,200,0,149,0,217,0,0,0,50,0,211,0,46,0,222,0,0,0,117,0,123,0,67,0,4,0,37,0,183,0);
signal scenario_full  : scenario_type := (216,31,151,31,36,31,121,31,11,31,91,31,213,31,246,31,246,30,161,31,5,31,87,31,173,31,177,31,9,31,9,30,43,31,24,31,24,30,84,31,72,31,154,31,72,31,194,31,152,31,128,31,53,31,132,31,132,30,84,31,100,31,78,31,85,31,180,31,105,31,19,31,227,31,237,31,149,31,245,31,245,30,245,29,54,31,239,31,187,31,226,31,192,31,155,31,155,30,65,31,181,31,28,31,89,31,93,31,138,31,176,31,58,31,182,31,39,31,39,30,168,31,126,31,51,31,185,31,185,30,207,31,128,31,128,30,246,31,146,31,189,31,189,30,8,31,163,31,163,30,54,31,134,31,178,31,114,31,169,31,110,31,239,31,187,31,136,31,232,31,249,31,144,31,144,30,144,29,101,31,225,31,225,30,225,29,202,31,16,31,207,31,17,31,17,30,141,31,141,30,240,31,87,31,85,31,85,30,85,29,121,31,248,31,160,31,160,30,160,29,195,31,22,31,105,31,49,31,71,31,71,30,74,31,130,31,131,31,131,30,192,31,118,31,112,31,165,31,98,31,40,31,1,31,1,30,145,31,145,30,87,31,98,31,234,31,245,31,245,30,235,31,210,31,211,31,199,31,175,31,88,31,230,31,65,31,99,31,61,31,48,31,48,30,121,31,15,31,128,31,185,31,70,31,122,31,60,31,229,31,150,31,150,30,200,31,200,30,189,31,220,31,146,31,146,30,62,31,179,31,138,31,75,31,126,31,47,31,50,31,113,31,168,31,95,31,3,31,3,30,128,31,128,30,209,31,96,31,1,31,25,31,4,31,237,31,27,31,227,31,227,30,245,31,242,31,151,31,141,31,134,31,231,31,24,31,105,31,105,30,22,31,142,31,212,31,23,31,2,31,2,30,249,31,53,31,213,31,59,31,237,31,18,31,135,31,37,31,37,30,50,31,218,31,196,31,85,31,86,31,47,31,113,31,189,31,189,30,251,31,56,31,55,31,55,30,185,31,223,31,207,31,117,31,117,30,202,31,234,31,209,31,252,31,252,30,19,31,188,31,4,31,147,31,147,30,102,31,53,31,19,31,2,31,248,31,232,31,232,30,232,29,162,31,17,31,148,31,69,31,59,31,165,31,165,30,165,29,104,31,70,31,70,30,220,31,72,31,251,31,251,30,209,31,209,30,100,31,178,31,178,30,84,31,161,31,238,31,94,31,202,31,218,31,218,30,98,31,249,31,49,31,102,31,216,31,157,31,76,31,65,31,54,31,12,31,122,31,85,31,225,31,27,31,44,31,167,31,200,31,143,31,63,31,145,31,85,31,161,31,89,31,89,30,197,31,197,30,41,31,41,30,239,31,32,31,226,31,222,31,126,31,220,31,5,31,247,31,108,31,68,31,48,31,174,31,174,30,138,31,138,30,114,31,114,30,178,31,178,30,140,31,140,30,119,31,5,31,189,31,214,31,63,31,78,31,227,31,186,31,104,31,231,31,231,30,5,31,23,31,66,31,216,31,49,31,150,31,196,31,15,31,19,31,60,31,150,31,150,30,150,29,253,31,78,31,135,31,135,30,238,31,238,30,186,31,252,31,14,31,121,31,121,30,147,31,246,31,45,31,45,30,152,31,252,31,1,31,1,30,122,31,22,31,232,31,232,30,124,31,136,31,136,30,136,29,35,31,123,31,150,31,150,30,241,31,196,31,245,31,76,31,242,31,174,31,174,30,69,31,183,31,143,31,124,31,52,31,52,30,44,31,227,31,67,31,243,31,171,31,240,31,40,31,110,31,96,31,96,30,216,31,90,31,53,31,197,31,111,31,111,30,111,29,39,31,116,31,31,31,177,31,236,31,236,30,210,31,165,31,217,31,126,31,16,31,156,31,88,31,88,30,178,31,124,31,92,31,148,31,46,31,141,31,141,30,83,31,209,31,146,31,146,30,77,31,2,31,178,31,184,31,176,31,182,31,197,31,59,31,9,31,191,31,142,31,63,31,172,31,247,31,232,31,159,31,80,31,72,31,3,31,130,31,102,31,1,31,237,31,237,30,39,31,100,31,73,31,73,30,148,31,245,31,171,31,164,31,170,31,219,31,219,30,123,31,252,31,99,31,244,31,22,31,248,31,248,30,242,31,130,31,27,31,200,31,149,31,217,31,217,30,50,31,211,31,46,31,222,31,222,30,117,31,123,31,67,31,4,31,37,31,183,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
