-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_552 is
end project_tb_552;

architecture project_tb_arch_552 of project_tb_552 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 714;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,21,0,202,0,0,0,163,0,0,0,193,0,147,0,47,0,106,0,22,0,12,0,118,0,152,0,197,0,151,0,200,0,0,0,178,0,123,0,226,0,28,0,166,0,124,0,199,0,0,0,0,0,0,0,165,0,194,0,171,0,19,0,90,0,253,0,253,0,61,0,254,0,33,0,106,0,0,0,54,0,0,0,0,0,43,0,52,0,160,0,20,0,251,0,167,0,134,0,41,0,243,0,0,0,217,0,102,0,10,0,69,0,0,0,0,0,137,0,179,0,88,0,98,0,220,0,43,0,175,0,115,0,83,0,173,0,0,0,97,0,0,0,215,0,0,0,103,0,0,0,114,0,46,0,230,0,193,0,78,0,173,0,0,0,102,0,0,0,182,0,229,0,0,0,140,0,131,0,0,0,71,0,240,0,0,0,32,0,163,0,0,0,163,0,138,0,161,0,128,0,183,0,0,0,0,0,99,0,82,0,0,0,17,0,87,0,217,0,114,0,95,0,166,0,30,0,191,0,62,0,205,0,133,0,0,0,32,0,141,0,106,0,45,0,0,0,171,0,72,0,65,0,201,0,105,0,213,0,239,0,72,0,236,0,233,0,57,0,188,0,161,0,31,0,0,0,48,0,0,0,0,0,232,0,227,0,96,0,187,0,155,0,138,0,77,0,253,0,0,0,250,0,27,0,166,0,181,0,239,0,124,0,97,0,116,0,12,0,123,0,0,0,0,0,12,0,0,0,79,0,42,0,143,0,0,0,0,0,226,0,0,0,157,0,0,0,13,0,0,0,77,0,0,0,186,0,143,0,92,0,249,0,218,0,240,0,39,0,90,0,0,0,0,0,43,0,98,0,0,0,212,0,166,0,179,0,45,0,82,0,254,0,186,0,214,0,245,0,179,0,96,0,224,0,239,0,111,0,3,0,248,0,0,0,0,0,136,0,119,0,168,0,147,0,51,0,0,0,162,0,55,0,28,0,19,0,251,0,103,0,0,0,143,0,98,0,201,0,0,0,245,0,79,0,0,0,103,0,35,0,104,0,8,0,0,0,24,0,80,0,125,0,0,0,89,0,0,0,150,0,186,0,45,0,161,0,0,0,3,0,97,0,92,0,0,0,90,0,192,0,188,0,39,0,0,0,89,0,181,0,172,0,232,0,31,0,72,0,6,0,151,0,0,0,0,0,236,0,35,0,81,0,0,0,4,0,172,0,55,0,181,0,243,0,100,0,54,0,225,0,249,0,253,0,119,0,174,0,206,0,230,0,6,0,184,0,15,0,0,0,177,0,66,0,134,0,74,0,0,0,40,0,128,0,158,0,0,0,193,0,46,0,220,0,35,0,52,0,0,0,113,0,36,0,109,0,204,0,89,0,223,0,0,0,71,0,59,0,243,0,74,0,98,0,21,0,124,0,168,0,0,0,5,0,49,0,6,0,3,0,247,0,210,0,229,0,0,0,203,0,0,0,247,0,215,0,0,0,27,0,135,0,82,0,84,0,175,0,0,0,114,0,144,0,0,0,0,0,43,0,18,0,0,0,81,0,249,0,101,0,82,0,8,0,22,0,215,0,83,0,180,0,1,0,88,0,48,0,183,0,180,0,66,0,242,0,86,0,56,0,48,0,0,0,0,0,67,0,155,0,153,0,60,0,124,0,26,0,173,0,137,0,174,0,122,0,153,0,171,0,0,0,96,0,28,0,63,0,241,0,228,0,195,0,25,0,0,0,154,0,245,0,43,0,180,0,160,0,38,0,224,0,71,0,134,0,172,0,143,0,6,0,187,0,127,0,191,0,58,0,0,0,0,0,221,0,0,0,59,0,134,0,37,0,0,0,0,0,153,0,96,0,168,0,238,0,27,0,0,0,36,0,131,0,36,0,5,0,0,0,152,0,104,0,0,0,0,0,35,0,218,0,28,0,43,0,203,0,98,0,0,0,0,0,0,0,21,0,126,0,77,0,167,0,207,0,80,0,124,0,235,0,67,0,196,0,0,0,0,0,22,0,50,0,56,0,0,0,127,0,247,0,0,0,0,0,0,0,183,0,0,0,76,0,0,0,0,0,24,0,143,0,43,0,199,0,232,0,241,0,0,0,0,0,206,0,137,0,152,0,229,0,225,0,0,0,59,0,220,0,0,0,139,0,0,0,177,0,23,0,29,0,125,0,172,0,7,0,25,0,97,0,187,0,128,0,14,0,50,0,6,0,146,0,78,0,43,0,37,0,239,0,117,0,171,0,110,0,0,0,145,0,47,0,0,0,116,0,53,0,99,0,0,0,67,0,13,0,0,0,78,0,111,0,0,0,2,0,65,0,0,0,62,0,160,0,50,0,70,0,10,0,41,0,65,0,48,0,132,0,208,0,207,0,233,0,125,0,0,0,119,0,16,0,155,0,231,0,239,0,38,0,24,0,108,0,52,0,55,0,29,0,46,0,215,0,122,0,199,0,81,0,166,0,89,0,204,0,207,0,27,0,156,0,0,0,90,0,97,0,47,0,177,0,31,0,215,0,22,0,44,0,3,0,223,0,106,0,21,0,120,0,197,0,110,0,147,0,207,0,81,0,90,0,26,0,47,0,52,0,38,0,0,0,73,0,62,0,108,0,179,0,0,0,120,0,0,0,204,0,0,0,160,0,0,0,0,0,173,0,0,0,240,0,216,0,0,0,178,0,55,0,174,0,118,0,121,0,34,0,128,0,170,0,0,0,0,0,141,0,149,0,0,0,0,0,227,0,201,0,0,0,20,0,0,0,197,0,145,0,117,0,139,0,95,0,215,0,6,0,251,0,62,0,0,0,0,0,240,0,0,0,105,0,64,0,0,0,134,0,162,0,71,0,0,0,0,0,11,0,12,0,251,0,207,0,204,0,102,0,7,0,41,0,23,0,110,0,133,0,67,0,144,0,249,0,184,0,0,0,177,0,0,0,21,0,0,0,11,0,71,0,138,0,58,0,0,0,0,0,248,0,29,0,0,0,0,0,0,0,142,0,40,0,0,0,82,0,127,0,0,0,173,0,148,0,187,0,16,0,204,0,167,0,12,0,223,0,0,0,198,0,2,0,41,0,57,0,112,0,130,0,180,0,0,0,230,0,114,0,59,0,65,0,57,0,119,0,56,0,0,0,107,0,134,0,134,0,65,0,0,0,166,0,0,0,170,0,218,0,208,0,120,0,169,0,13,0,0,0,129,0,0,0,114,0);
signal scenario_full  : scenario_type := (0,0,21,31,202,31,202,30,163,31,163,30,193,31,147,31,47,31,106,31,22,31,12,31,118,31,152,31,197,31,151,31,200,31,200,30,178,31,123,31,226,31,28,31,166,31,124,31,199,31,199,30,199,29,199,28,165,31,194,31,171,31,19,31,90,31,253,31,253,31,61,31,254,31,33,31,106,31,106,30,54,31,54,30,54,29,43,31,52,31,160,31,20,31,251,31,167,31,134,31,41,31,243,31,243,30,217,31,102,31,10,31,69,31,69,30,69,29,137,31,179,31,88,31,98,31,220,31,43,31,175,31,115,31,83,31,173,31,173,30,97,31,97,30,215,31,215,30,103,31,103,30,114,31,46,31,230,31,193,31,78,31,173,31,173,30,102,31,102,30,182,31,229,31,229,30,140,31,131,31,131,30,71,31,240,31,240,30,32,31,163,31,163,30,163,31,138,31,161,31,128,31,183,31,183,30,183,29,99,31,82,31,82,30,17,31,87,31,217,31,114,31,95,31,166,31,30,31,191,31,62,31,205,31,133,31,133,30,32,31,141,31,106,31,45,31,45,30,171,31,72,31,65,31,201,31,105,31,213,31,239,31,72,31,236,31,233,31,57,31,188,31,161,31,31,31,31,30,48,31,48,30,48,29,232,31,227,31,96,31,187,31,155,31,138,31,77,31,253,31,253,30,250,31,27,31,166,31,181,31,239,31,124,31,97,31,116,31,12,31,123,31,123,30,123,29,12,31,12,30,79,31,42,31,143,31,143,30,143,29,226,31,226,30,157,31,157,30,13,31,13,30,77,31,77,30,186,31,143,31,92,31,249,31,218,31,240,31,39,31,90,31,90,30,90,29,43,31,98,31,98,30,212,31,166,31,179,31,45,31,82,31,254,31,186,31,214,31,245,31,179,31,96,31,224,31,239,31,111,31,3,31,248,31,248,30,248,29,136,31,119,31,168,31,147,31,51,31,51,30,162,31,55,31,28,31,19,31,251,31,103,31,103,30,143,31,98,31,201,31,201,30,245,31,79,31,79,30,103,31,35,31,104,31,8,31,8,30,24,31,80,31,125,31,125,30,89,31,89,30,150,31,186,31,45,31,161,31,161,30,3,31,97,31,92,31,92,30,90,31,192,31,188,31,39,31,39,30,89,31,181,31,172,31,232,31,31,31,72,31,6,31,151,31,151,30,151,29,236,31,35,31,81,31,81,30,4,31,172,31,55,31,181,31,243,31,100,31,54,31,225,31,249,31,253,31,119,31,174,31,206,31,230,31,6,31,184,31,15,31,15,30,177,31,66,31,134,31,74,31,74,30,40,31,128,31,158,31,158,30,193,31,46,31,220,31,35,31,52,31,52,30,113,31,36,31,109,31,204,31,89,31,223,31,223,30,71,31,59,31,243,31,74,31,98,31,21,31,124,31,168,31,168,30,5,31,49,31,6,31,3,31,247,31,210,31,229,31,229,30,203,31,203,30,247,31,215,31,215,30,27,31,135,31,82,31,84,31,175,31,175,30,114,31,144,31,144,30,144,29,43,31,18,31,18,30,81,31,249,31,101,31,82,31,8,31,22,31,215,31,83,31,180,31,1,31,88,31,48,31,183,31,180,31,66,31,242,31,86,31,56,31,48,31,48,30,48,29,67,31,155,31,153,31,60,31,124,31,26,31,173,31,137,31,174,31,122,31,153,31,171,31,171,30,96,31,28,31,63,31,241,31,228,31,195,31,25,31,25,30,154,31,245,31,43,31,180,31,160,31,38,31,224,31,71,31,134,31,172,31,143,31,6,31,187,31,127,31,191,31,58,31,58,30,58,29,221,31,221,30,59,31,134,31,37,31,37,30,37,29,153,31,96,31,168,31,238,31,27,31,27,30,36,31,131,31,36,31,5,31,5,30,152,31,104,31,104,30,104,29,35,31,218,31,28,31,43,31,203,31,98,31,98,30,98,29,98,28,21,31,126,31,77,31,167,31,207,31,80,31,124,31,235,31,67,31,196,31,196,30,196,29,22,31,50,31,56,31,56,30,127,31,247,31,247,30,247,29,247,28,183,31,183,30,76,31,76,30,76,29,24,31,143,31,43,31,199,31,232,31,241,31,241,30,241,29,206,31,137,31,152,31,229,31,225,31,225,30,59,31,220,31,220,30,139,31,139,30,177,31,23,31,29,31,125,31,172,31,7,31,25,31,97,31,187,31,128,31,14,31,50,31,6,31,146,31,78,31,43,31,37,31,239,31,117,31,171,31,110,31,110,30,145,31,47,31,47,30,116,31,53,31,99,31,99,30,67,31,13,31,13,30,78,31,111,31,111,30,2,31,65,31,65,30,62,31,160,31,50,31,70,31,10,31,41,31,65,31,48,31,132,31,208,31,207,31,233,31,125,31,125,30,119,31,16,31,155,31,231,31,239,31,38,31,24,31,108,31,52,31,55,31,29,31,46,31,215,31,122,31,199,31,81,31,166,31,89,31,204,31,207,31,27,31,156,31,156,30,90,31,97,31,47,31,177,31,31,31,215,31,22,31,44,31,3,31,223,31,106,31,21,31,120,31,197,31,110,31,147,31,207,31,81,31,90,31,26,31,47,31,52,31,38,31,38,30,73,31,62,31,108,31,179,31,179,30,120,31,120,30,204,31,204,30,160,31,160,30,160,29,173,31,173,30,240,31,216,31,216,30,178,31,55,31,174,31,118,31,121,31,34,31,128,31,170,31,170,30,170,29,141,31,149,31,149,30,149,29,227,31,201,31,201,30,20,31,20,30,197,31,145,31,117,31,139,31,95,31,215,31,6,31,251,31,62,31,62,30,62,29,240,31,240,30,105,31,64,31,64,30,134,31,162,31,71,31,71,30,71,29,11,31,12,31,251,31,207,31,204,31,102,31,7,31,41,31,23,31,110,31,133,31,67,31,144,31,249,31,184,31,184,30,177,31,177,30,21,31,21,30,11,31,71,31,138,31,58,31,58,30,58,29,248,31,29,31,29,30,29,29,29,28,142,31,40,31,40,30,82,31,127,31,127,30,173,31,148,31,187,31,16,31,204,31,167,31,12,31,223,31,223,30,198,31,2,31,41,31,57,31,112,31,130,31,180,31,180,30,230,31,114,31,59,31,65,31,57,31,119,31,56,31,56,30,107,31,134,31,134,31,65,31,65,30,166,31,166,30,170,31,218,31,208,31,120,31,169,31,13,31,13,30,129,31,129,30,114,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
