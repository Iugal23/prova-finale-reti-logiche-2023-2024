-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_181 is
end project_tb_181;

architecture project_tb_arch_181 of project_tb_181 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 215;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (162,0,254,0,54,0,183,0,231,0,62,0,247,0,183,0,43,0,151,0,0,0,252,0,120,0,58,0,214,0,192,0,0,0,0,0,0,0,0,0,39,0,70,0,0,0,28,0,62,0,123,0,254,0,10,0,0,0,66,0,0,0,17,0,0,0,86,0,53,0,0,0,68,0,25,0,0,0,209,0,153,0,212,0,125,0,187,0,1,0,9,0,215,0,118,0,130,0,226,0,112,0,0,0,38,0,16,0,0,0,25,0,0,0,38,0,0,0,248,0,100,0,40,0,0,0,0,0,153,0,0,0,11,0,0,0,234,0,0,0,12,0,0,0,196,0,0,0,208,0,228,0,53,0,177,0,205,0,150,0,166,0,208,0,0,0,224,0,233,0,103,0,42,0,99,0,0,0,107,0,0,0,77,0,27,0,22,0,34,0,3,0,69,0,126,0,0,0,13,0,179,0,68,0,0,0,134,0,149,0,121,0,0,0,0,0,221,0,42,0,0,0,27,0,211,0,174,0,26,0,0,0,70,0,0,0,0,0,34,0,39,0,224,0,142,0,173,0,144,0,25,0,252,0,27,0,253,0,4,0,54,0,0,0,248,0,180,0,209,0,188,0,189,0,46,0,121,0,13,0,233,0,124,0,85,0,206,0,89,0,153,0,135,0,136,0,183,0,71,0,63,0,189,0,121,0,178,0,11,0,126,0,2,0,25,0,147,0,0,0,30,0,180,0,160,0,26,0,159,0,0,0,50,0,217,0,0,0,0,0,0,0,255,0,0,0,170,0,226,0,204,0,0,0,111,0,160,0,143,0,211,0,172,0,121,0,174,0,212,0,184,0,238,0,0,0,98,0,236,0,255,0,230,0,144,0,96,0,102,0,3,0,154,0,0,0,208,0,215,0,240,0,144,0,120,0,0,0,39,0,89,0,173,0,0,0,0,0,225,0,0,0,0,0,43,0,60,0,35,0);
signal scenario_full  : scenario_type := (162,31,254,31,54,31,183,31,231,31,62,31,247,31,183,31,43,31,151,31,151,30,252,31,120,31,58,31,214,31,192,31,192,30,192,29,192,28,192,27,39,31,70,31,70,30,28,31,62,31,123,31,254,31,10,31,10,30,66,31,66,30,17,31,17,30,86,31,53,31,53,30,68,31,25,31,25,30,209,31,153,31,212,31,125,31,187,31,1,31,9,31,215,31,118,31,130,31,226,31,112,31,112,30,38,31,16,31,16,30,25,31,25,30,38,31,38,30,248,31,100,31,40,31,40,30,40,29,153,31,153,30,11,31,11,30,234,31,234,30,12,31,12,30,196,31,196,30,208,31,228,31,53,31,177,31,205,31,150,31,166,31,208,31,208,30,224,31,233,31,103,31,42,31,99,31,99,30,107,31,107,30,77,31,27,31,22,31,34,31,3,31,69,31,126,31,126,30,13,31,179,31,68,31,68,30,134,31,149,31,121,31,121,30,121,29,221,31,42,31,42,30,27,31,211,31,174,31,26,31,26,30,70,31,70,30,70,29,34,31,39,31,224,31,142,31,173,31,144,31,25,31,252,31,27,31,253,31,4,31,54,31,54,30,248,31,180,31,209,31,188,31,189,31,46,31,121,31,13,31,233,31,124,31,85,31,206,31,89,31,153,31,135,31,136,31,183,31,71,31,63,31,189,31,121,31,178,31,11,31,126,31,2,31,25,31,147,31,147,30,30,31,180,31,160,31,26,31,159,31,159,30,50,31,217,31,217,30,217,29,217,28,255,31,255,30,170,31,226,31,204,31,204,30,111,31,160,31,143,31,211,31,172,31,121,31,174,31,212,31,184,31,238,31,238,30,98,31,236,31,255,31,230,31,144,31,96,31,102,31,3,31,154,31,154,30,208,31,215,31,240,31,144,31,120,31,120,30,39,31,89,31,173,31,173,30,173,29,225,31,225,30,225,29,43,31,60,31,35,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
