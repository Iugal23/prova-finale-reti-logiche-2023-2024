-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 758;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (122,0,0,0,191,0,0,0,0,0,0,0,202,0,197,0,110,0,0,0,245,0,95,0,0,0,38,0,120,0,117,0,222,0,157,0,141,0,24,0,68,0,15,0,78,0,168,0,214,0,58,0,188,0,240,0,135,0,162,0,0,0,55,0,76,0,0,0,35,0,0,0,86,0,27,0,124,0,104,0,223,0,112,0,0,0,181,0,80,0,245,0,74,0,74,0,47,0,31,0,0,0,180,0,61,0,55,0,32,0,10,0,101,0,234,0,230,0,141,0,0,0,164,0,254,0,255,0,89,0,0,0,107,0,18,0,160,0,49,0,197,0,117,0,51,0,16,0,179,0,38,0,9,0,171,0,7,0,228,0,102,0,12,0,0,0,0,0,16,0,219,0,89,0,131,0,30,0,38,0,19,0,37,0,201,0,103,0,31,0,232,0,217,0,16,0,137,0,175,0,0,0,5,0,179,0,1,0,80,0,228,0,117,0,239,0,239,0,87,0,226,0,85,0,82,0,157,0,16,0,47,0,100,0,26,0,130,0,221,0,242,0,88,0,40,0,155,0,6,0,216,0,0,0,0,0,43,0,102,0,0,0,147,0,120,0,2,0,238,0,0,0,247,0,218,0,225,0,72,0,240,0,171,0,66,0,11,0,231,0,0,0,0,0,254,0,116,0,0,0,36,0,59,0,72,0,11,0,0,0,202,0,66,0,189,0,0,0,0,0,0,0,81,0,140,0,0,0,0,0,110,0,114,0,214,0,241,0,54,0,115,0,176,0,59,0,0,0,102,0,44,0,229,0,182,0,128,0,246,0,0,0,234,0,139,0,144,0,0,0,155,0,5,0,196,0,81,0,183,0,176,0,58,0,20,0,189,0,151,0,154,0,233,0,85,0,236,0,170,0,132,0,75,0,0,0,0,0,245,0,201,0,0,0,165,0,25,0,0,0,2,0,0,0,96,0,3,0,105,0,48,0,175,0,33,0,82,0,0,0,63,0,0,0,189,0,87,0,118,0,20,0,170,0,4,0,197,0,2,0,5,0,251,0,117,0,0,0,137,0,0,0,0,0,18,0,131,0,74,0,41,0,57,0,0,0,123,0,0,0,248,0,0,0,11,0,0,0,146,0,92,0,208,0,152,0,0,0,154,0,181,0,11,0,214,0,25,0,0,0,0,0,85,0,143,0,241,0,0,0,99,0,1,0,218,0,118,0,43,0,48,0,0,0,244,0,172,0,0,0,210,0,128,0,244,0,158,0,20,0,0,0,19,0,0,0,144,0,0,0,216,0,174,0,78,0,56,0,59,0,178,0,118,0,124,0,40,0,2,0,0,0,197,0,187,0,0,0,124,0,158,0,139,0,254,0,252,0,30,0,132,0,169,0,24,0,75,0,178,0,252,0,100,0,146,0,130,0,0,0,107,0,238,0,238,0,93,0,160,0,146,0,91,0,63,0,71,0,105,0,0,0,34,0,200,0,229,0,53,0,237,0,0,0,104,0,27,0,167,0,48,0,63,0,6,0,184,0,111,0,63,0,220,0,0,0,92,0,164,0,26,0,1,0,0,0,204,0,205,0,187,0,23,0,134,0,157,0,69,0,140,0,89,0,72,0,46,0,253,0,223,0,172,0,56,0,202,0,0,0,111,0,240,0,69,0,118,0,17,0,12,0,65,0,213,0,253,0,0,0,77,0,11,0,128,0,0,0,204,0,193,0,16,0,114,0,44,0,159,0,50,0,217,0,0,0,92,0,199,0,104,0,0,0,70,0,237,0,196,0,224,0,242,0,22,0,0,0,221,0,222,0,88,0,180,0,236,0,102,0,206,0,184,0,100,0,0,0,0,0,10,0,0,0,0,0,222,0,157,0,48,0,40,0,0,0,0,0,50,0,0,0,19,0,85,0,0,0,15,0,224,0,0,0,192,0,170,0,0,0,0,0,0,0,69,0,0,0,25,0,232,0,83,0,124,0,0,0,0,0,130,0,0,0,230,0,206,0,0,0,139,0,0,0,0,0,0,0,0,0,95,0,71,0,0,0,192,0,16,0,3,0,191,0,17,0,117,0,135,0,76,0,179,0,154,0,23,0,10,0,38,0,214,0,190,0,70,0,58,0,0,0,90,0,0,0,158,0,214,0,190,0,0,0,20,0,221,0,0,0,12,0,216,0,199,0,231,0,146,0,143,0,224,0,233,0,0,0,216,0,212,0,149,0,107,0,140,0,23,0,72,0,144,0,45,0,232,0,0,0,0,0,103,0,75,0,39,0,151,0,126,0,0,0,125,0,85,0,0,0,159,0,81,0,177,0,112,0,117,0,2,0,0,0,0,0,49,0,0,0,137,0,153,0,0,0,158,0,78,0,53,0,210,0,26,0,35,0,151,0,135,0,0,0,0,0,41,0,199,0,0,0,0,0,68,0,231,0,73,0,186,0,172,0,0,0,178,0,165,0,0,0,0,0,45,0,0,0,145,0,88,0,144,0,226,0,28,0,0,0,192,0,0,0,6,0,45,0,83,0,6,0,62,0,95,0,172,0,136,0,169,0,100,0,166,0,0,0,96,0,18,0,0,0,0,0,134,0,132,0,147,0,0,0,201,0,216,0,127,0,0,0,171,0,106,0,0,0,203,0,31,0,230,0,209,0,185,0,26,0,28,0,13,0,22,0,23,0,0,0,14,0,57,0,123,0,0,0,254,0,11,0,12,0,230,0,129,0,186,0,0,0,64,0,0,0,0,0,0,0,110,0,0,0,82,0,35,0,155,0,0,0,94,0,211,0,0,0,0,0,202,0,132,0,47,0,83,0,215,0,253,0,132,0,31,0,125,0,113,0,55,0,11,0,0,0,128,0,70,0,34,0,0,0,0,0,200,0,174,0,0,0,0,0,248,0,105,0,0,0,176,0,0,0,231,0,210,0,31,0,0,0,159,0,0,0,0,0,175,0,230,0,152,0,0,0,33,0,97,0,181,0,228,0,151,0,0,0,232,0,152,0,0,0,116,0,57,0,199,0,69,0,136,0,22,0,55,0,27,0,254,0,206,0,6,0,105,0,165,0,120,0,69,0,170,0,218,0,28,0,219,0,27,0,187,0,119,0,0,0,44,0,0,0,44,0,95,0,68,0,41,0,0,0,153,0,14,0,0,0,150,0,0,0,196,0,132,0,59,0,141,0,54,0,63,0,111,0,205,0,75,0,219,0,0,0,117,0,0,0,46,0,164,0,231,0,172,0,19,0,141,0,73,0,183,0,138,0,167,0,227,0,0,0,241,0,96,0,0,0,21,0,0,0,0,0,190,0,127,0,95,0,156,0,77,0,20,0,8,0,126,0,17,0,153,0,0,0,106,0,247,0,119,0,0,0,113,0,54,0,214,0,213,0,188,0,170,0,104,0,123,0,0,0,146,0);
signal scenario_full  : scenario_type := (122,31,122,30,191,31,191,30,191,29,191,28,202,31,197,31,110,31,110,30,245,31,95,31,95,30,38,31,120,31,117,31,222,31,157,31,141,31,24,31,68,31,15,31,78,31,168,31,214,31,58,31,188,31,240,31,135,31,162,31,162,30,55,31,76,31,76,30,35,31,35,30,86,31,27,31,124,31,104,31,223,31,112,31,112,30,181,31,80,31,245,31,74,31,74,31,47,31,31,31,31,30,180,31,61,31,55,31,32,31,10,31,101,31,234,31,230,31,141,31,141,30,164,31,254,31,255,31,89,31,89,30,107,31,18,31,160,31,49,31,197,31,117,31,51,31,16,31,179,31,38,31,9,31,171,31,7,31,228,31,102,31,12,31,12,30,12,29,16,31,219,31,89,31,131,31,30,31,38,31,19,31,37,31,201,31,103,31,31,31,232,31,217,31,16,31,137,31,175,31,175,30,5,31,179,31,1,31,80,31,228,31,117,31,239,31,239,31,87,31,226,31,85,31,82,31,157,31,16,31,47,31,100,31,26,31,130,31,221,31,242,31,88,31,40,31,155,31,6,31,216,31,216,30,216,29,43,31,102,31,102,30,147,31,120,31,2,31,238,31,238,30,247,31,218,31,225,31,72,31,240,31,171,31,66,31,11,31,231,31,231,30,231,29,254,31,116,31,116,30,36,31,59,31,72,31,11,31,11,30,202,31,66,31,189,31,189,30,189,29,189,28,81,31,140,31,140,30,140,29,110,31,114,31,214,31,241,31,54,31,115,31,176,31,59,31,59,30,102,31,44,31,229,31,182,31,128,31,246,31,246,30,234,31,139,31,144,31,144,30,155,31,5,31,196,31,81,31,183,31,176,31,58,31,20,31,189,31,151,31,154,31,233,31,85,31,236,31,170,31,132,31,75,31,75,30,75,29,245,31,201,31,201,30,165,31,25,31,25,30,2,31,2,30,96,31,3,31,105,31,48,31,175,31,33,31,82,31,82,30,63,31,63,30,189,31,87,31,118,31,20,31,170,31,4,31,197,31,2,31,5,31,251,31,117,31,117,30,137,31,137,30,137,29,18,31,131,31,74,31,41,31,57,31,57,30,123,31,123,30,248,31,248,30,11,31,11,30,146,31,92,31,208,31,152,31,152,30,154,31,181,31,11,31,214,31,25,31,25,30,25,29,85,31,143,31,241,31,241,30,99,31,1,31,218,31,118,31,43,31,48,31,48,30,244,31,172,31,172,30,210,31,128,31,244,31,158,31,20,31,20,30,19,31,19,30,144,31,144,30,216,31,174,31,78,31,56,31,59,31,178,31,118,31,124,31,40,31,2,31,2,30,197,31,187,31,187,30,124,31,158,31,139,31,254,31,252,31,30,31,132,31,169,31,24,31,75,31,178,31,252,31,100,31,146,31,130,31,130,30,107,31,238,31,238,31,93,31,160,31,146,31,91,31,63,31,71,31,105,31,105,30,34,31,200,31,229,31,53,31,237,31,237,30,104,31,27,31,167,31,48,31,63,31,6,31,184,31,111,31,63,31,220,31,220,30,92,31,164,31,26,31,1,31,1,30,204,31,205,31,187,31,23,31,134,31,157,31,69,31,140,31,89,31,72,31,46,31,253,31,223,31,172,31,56,31,202,31,202,30,111,31,240,31,69,31,118,31,17,31,12,31,65,31,213,31,253,31,253,30,77,31,11,31,128,31,128,30,204,31,193,31,16,31,114,31,44,31,159,31,50,31,217,31,217,30,92,31,199,31,104,31,104,30,70,31,237,31,196,31,224,31,242,31,22,31,22,30,221,31,222,31,88,31,180,31,236,31,102,31,206,31,184,31,100,31,100,30,100,29,10,31,10,30,10,29,222,31,157,31,48,31,40,31,40,30,40,29,50,31,50,30,19,31,85,31,85,30,15,31,224,31,224,30,192,31,170,31,170,30,170,29,170,28,69,31,69,30,25,31,232,31,83,31,124,31,124,30,124,29,130,31,130,30,230,31,206,31,206,30,139,31,139,30,139,29,139,28,139,27,95,31,71,31,71,30,192,31,16,31,3,31,191,31,17,31,117,31,135,31,76,31,179,31,154,31,23,31,10,31,38,31,214,31,190,31,70,31,58,31,58,30,90,31,90,30,158,31,214,31,190,31,190,30,20,31,221,31,221,30,12,31,216,31,199,31,231,31,146,31,143,31,224,31,233,31,233,30,216,31,212,31,149,31,107,31,140,31,23,31,72,31,144,31,45,31,232,31,232,30,232,29,103,31,75,31,39,31,151,31,126,31,126,30,125,31,85,31,85,30,159,31,81,31,177,31,112,31,117,31,2,31,2,30,2,29,49,31,49,30,137,31,153,31,153,30,158,31,78,31,53,31,210,31,26,31,35,31,151,31,135,31,135,30,135,29,41,31,199,31,199,30,199,29,68,31,231,31,73,31,186,31,172,31,172,30,178,31,165,31,165,30,165,29,45,31,45,30,145,31,88,31,144,31,226,31,28,31,28,30,192,31,192,30,6,31,45,31,83,31,6,31,62,31,95,31,172,31,136,31,169,31,100,31,166,31,166,30,96,31,18,31,18,30,18,29,134,31,132,31,147,31,147,30,201,31,216,31,127,31,127,30,171,31,106,31,106,30,203,31,31,31,230,31,209,31,185,31,26,31,28,31,13,31,22,31,23,31,23,30,14,31,57,31,123,31,123,30,254,31,11,31,12,31,230,31,129,31,186,31,186,30,64,31,64,30,64,29,64,28,110,31,110,30,82,31,35,31,155,31,155,30,94,31,211,31,211,30,211,29,202,31,132,31,47,31,83,31,215,31,253,31,132,31,31,31,125,31,113,31,55,31,11,31,11,30,128,31,70,31,34,31,34,30,34,29,200,31,174,31,174,30,174,29,248,31,105,31,105,30,176,31,176,30,231,31,210,31,31,31,31,30,159,31,159,30,159,29,175,31,230,31,152,31,152,30,33,31,97,31,181,31,228,31,151,31,151,30,232,31,152,31,152,30,116,31,57,31,199,31,69,31,136,31,22,31,55,31,27,31,254,31,206,31,6,31,105,31,165,31,120,31,69,31,170,31,218,31,28,31,219,31,27,31,187,31,119,31,119,30,44,31,44,30,44,31,95,31,68,31,41,31,41,30,153,31,14,31,14,30,150,31,150,30,196,31,132,31,59,31,141,31,54,31,63,31,111,31,205,31,75,31,219,31,219,30,117,31,117,30,46,31,164,31,231,31,172,31,19,31,141,31,73,31,183,31,138,31,167,31,227,31,227,30,241,31,96,31,96,30,21,31,21,30,21,29,190,31,127,31,95,31,156,31,77,31,20,31,8,31,126,31,17,31,153,31,153,30,106,31,247,31,119,31,119,30,113,31,54,31,214,31,213,31,188,31,170,31,104,31,123,31,123,30,146,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
