-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_520 is
end project_tb_520;

architecture project_tb_arch_520 of project_tb_520 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 667;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,136,0,130,0,28,0,202,0,0,0,243,0,126,0,194,0,0,0,239,0,74,0,130,0,161,0,0,0,0,0,61,0,107,0,0,0,90,0,0,0,64,0,212,0,0,0,116,0,154,0,0,0,34,0,0,0,123,0,164,0,0,0,0,0,180,0,62,0,249,0,0,0,163,0,232,0,255,0,209,0,0,0,0,0,0,0,87,0,0,0,34,0,195,0,78,0,41,0,0,0,95,0,174,0,138,0,144,0,220,0,0,0,209,0,0,0,44,0,171,0,154,0,204,0,26,0,74,0,138,0,173,0,181,0,73,0,0,0,121,0,0,0,0,0,252,0,15,0,176,0,213,0,0,0,147,0,53,0,58,0,0,0,30,0,95,0,111,0,222,0,218,0,121,0,132,0,0,0,77,0,184,0,117,0,166,0,0,0,222,0,59,0,0,0,223,0,91,0,141,0,204,0,85,0,168,0,0,0,0,0,162,0,238,0,73,0,73,0,47,0,228,0,127,0,118,0,48,0,56,0,90,0,74,0,215,0,0,0,0,0,106,0,68,0,41,0,0,0,42,0,0,0,0,0,1,0,5,0,0,0,60,0,226,0,25,0,157,0,149,0,192,0,241,0,234,0,199,0,0,0,0,0,209,0,226,0,86,0,236,0,0,0,187,0,0,0,0,0,1,0,245,0,0,0,0,0,99,0,14,0,29,0,0,0,76,0,158,0,0,0,0,0,178,0,83,0,135,0,50,0,105,0,192,0,94,0,55,0,185,0,71,0,0,0,12,0,143,0,243,0,201,0,22,0,150,0,135,0,0,0,0,0,0,0,79,0,192,0,0,0,238,0,237,0,0,0,105,0,40,0,174,0,172,0,60,0,0,0,0,0,64,0,248,0,22,0,232,0,195,0,131,0,132,0,217,0,142,0,0,0,248,0,42,0,0,0,38,0,29,0,90,0,94,0,0,0,98,0,0,0,136,0,0,0,14,0,216,0,21,0,217,0,131,0,0,0,125,0,0,0,181,0,53,0,100,0,57,0,51,0,214,0,136,0,173,0,0,0,252,0,254,0,133,0,57,0,0,0,230,0,180,0,1,0,0,0,10,0,59,0,86,0,0,0,0,0,0,0,8,0,186,0,210,0,30,0,139,0,17,0,94,0,138,0,7,0,179,0,0,0,76,0,152,0,111,0,20,0,35,0,37,0,200,0,63,0,0,0,26,0,75,0,49,0,0,0,179,0,213,0,205,0,0,0,81,0,105,0,228,0,29,0,244,0,0,0,151,0,0,0,189,0,201,0,0,0,177,0,218,0,6,0,114,0,4,0,154,0,213,0,82,0,193,0,0,0,49,0,198,0,0,0,146,0,180,0,0,0,63,0,228,0,68,0,0,0,78,0,27,0,0,0,77,0,44,0,0,0,247,0,190,0,95,0,84,0,58,0,191,0,199,0,0,0,0,0,17,0,185,0,54,0,0,0,98,0,0,0,0,0,140,0,86,0,179,0,4,0,0,0,139,0,158,0,0,0,83,0,0,0,212,0,234,0,0,0,0,0,51,0,0,0,0,0,0,0,192,0,104,0,67,0,24,0,253,0,118,0,154,0,0,0,245,0,150,0,0,0,0,0,119,0,6,0,145,0,0,0,1,0,101,0,218,0,75,0,100,0,148,0,53,0,160,0,31,0,2,0,46,0,51,0,158,0,249,0,243,0,7,0,117,0,238,0,212,0,176,0,0,0,50,0,123,0,34,0,153,0,0,0,115,0,111,0,61,0,228,0,0,0,205,0,226,0,65,0,84,0,74,0,74,0,159,0,0,0,0,0,122,0,0,0,175,0,251,0,78,0,0,0,217,0,72,0,232,0,0,0,154,0,178,0,206,0,0,0,166,0,0,0,148,0,21,0,102,0,224,0,193,0,185,0,61,0,129,0,56,0,149,0,92,0,103,0,0,0,246,0,135,0,231,0,143,0,3,0,0,0,236,0,45,0,9,0,0,0,134,0,168,0,187,0,135,0,4,0,114,0,252,0,236,0,203,0,217,0,123,0,181,0,106,0,122,0,229,0,167,0,178,0,0,0,251,0,17,0,251,0,183,0,22,0,34,0,0,0,189,0,194,0,0,0,13,0,0,0,89,0,134,0,197,0,206,0,132,0,84,0,143,0,79,0,164,0,42,0,110,0,0,0,0,0,86,0,227,0,122,0,0,0,234,0,0,0,151,0,198,0,6,0,179,0,155,0,0,0,178,0,97,0,0,0,119,0,143,0,250,0,0,0,118,0,180,0,121,0,0,0,0,0,105,0,71,0,127,0,16,0,247,0,97,0,117,0,36,0,68,0,22,0,0,0,107,0,127,0,123,0,136,0,91,0,0,0,141,0,9,0,0,0,26,0,0,0,0,0,89,0,106,0,124,0,186,0,60,0,9,0,121,0,84,0,159,0,63,0,53,0,218,0,124,0,103,0,108,0,0,0,172,0,155,0,49,0,21,0,0,0,195,0,57,0,229,0,0,0,0,0,87,0,249,0,122,0,1,0,164,0,147,0,154,0,57,0,0,0,194,0,33,0,193,0,62,0,105,0,110,0,159,0,0,0,149,0,177,0,249,0,0,0,133,0,200,0,53,0,189,0,0,0,0,0,51,0,46,0,0,0,23,0,190,0,0,0,0,0,82,0,152,0,0,0,170,0,20,0,144,0,76,0,65,0,48,0,249,0,47,0,204,0,196,0,217,0,97,0,85,0,251,0,103,0,222,0,230,0,211,0,200,0,195,0,0,0,172,0,94,0,0,0,146,0,143,0,96,0,52,0,47,0,178,0,148,0,214,0,247,0,0,0,222,0,235,0,73,0,54,0,9,0,50,0,247,0,140,0,49,0,175,0,122,0,0,0,216,0,254,0,80,0,252,0,24,0,209,0,113,0,253,0,94,0,218,0,121,0,0,0,5,0,235,0,134,0,0,0,0,0,49,0,59,0,185,0,243,0,156,0,34,0);
signal scenario_full  : scenario_type := (0,0,0,0,136,31,130,31,28,31,202,31,202,30,243,31,126,31,194,31,194,30,239,31,74,31,130,31,161,31,161,30,161,29,61,31,107,31,107,30,90,31,90,30,64,31,212,31,212,30,116,31,154,31,154,30,34,31,34,30,123,31,164,31,164,30,164,29,180,31,62,31,249,31,249,30,163,31,232,31,255,31,209,31,209,30,209,29,209,28,87,31,87,30,34,31,195,31,78,31,41,31,41,30,95,31,174,31,138,31,144,31,220,31,220,30,209,31,209,30,44,31,171,31,154,31,204,31,26,31,74,31,138,31,173,31,181,31,73,31,73,30,121,31,121,30,121,29,252,31,15,31,176,31,213,31,213,30,147,31,53,31,58,31,58,30,30,31,95,31,111,31,222,31,218,31,121,31,132,31,132,30,77,31,184,31,117,31,166,31,166,30,222,31,59,31,59,30,223,31,91,31,141,31,204,31,85,31,168,31,168,30,168,29,162,31,238,31,73,31,73,31,47,31,228,31,127,31,118,31,48,31,56,31,90,31,74,31,215,31,215,30,215,29,106,31,68,31,41,31,41,30,42,31,42,30,42,29,1,31,5,31,5,30,60,31,226,31,25,31,157,31,149,31,192,31,241,31,234,31,199,31,199,30,199,29,209,31,226,31,86,31,236,31,236,30,187,31,187,30,187,29,1,31,245,31,245,30,245,29,99,31,14,31,29,31,29,30,76,31,158,31,158,30,158,29,178,31,83,31,135,31,50,31,105,31,192,31,94,31,55,31,185,31,71,31,71,30,12,31,143,31,243,31,201,31,22,31,150,31,135,31,135,30,135,29,135,28,79,31,192,31,192,30,238,31,237,31,237,30,105,31,40,31,174,31,172,31,60,31,60,30,60,29,64,31,248,31,22,31,232,31,195,31,131,31,132,31,217,31,142,31,142,30,248,31,42,31,42,30,38,31,29,31,90,31,94,31,94,30,98,31,98,30,136,31,136,30,14,31,216,31,21,31,217,31,131,31,131,30,125,31,125,30,181,31,53,31,100,31,57,31,51,31,214,31,136,31,173,31,173,30,252,31,254,31,133,31,57,31,57,30,230,31,180,31,1,31,1,30,10,31,59,31,86,31,86,30,86,29,86,28,8,31,186,31,210,31,30,31,139,31,17,31,94,31,138,31,7,31,179,31,179,30,76,31,152,31,111,31,20,31,35,31,37,31,200,31,63,31,63,30,26,31,75,31,49,31,49,30,179,31,213,31,205,31,205,30,81,31,105,31,228,31,29,31,244,31,244,30,151,31,151,30,189,31,201,31,201,30,177,31,218,31,6,31,114,31,4,31,154,31,213,31,82,31,193,31,193,30,49,31,198,31,198,30,146,31,180,31,180,30,63,31,228,31,68,31,68,30,78,31,27,31,27,30,77,31,44,31,44,30,247,31,190,31,95,31,84,31,58,31,191,31,199,31,199,30,199,29,17,31,185,31,54,31,54,30,98,31,98,30,98,29,140,31,86,31,179,31,4,31,4,30,139,31,158,31,158,30,83,31,83,30,212,31,234,31,234,30,234,29,51,31,51,30,51,29,51,28,192,31,104,31,67,31,24,31,253,31,118,31,154,31,154,30,245,31,150,31,150,30,150,29,119,31,6,31,145,31,145,30,1,31,101,31,218,31,75,31,100,31,148,31,53,31,160,31,31,31,2,31,46,31,51,31,158,31,249,31,243,31,7,31,117,31,238,31,212,31,176,31,176,30,50,31,123,31,34,31,153,31,153,30,115,31,111,31,61,31,228,31,228,30,205,31,226,31,65,31,84,31,74,31,74,31,159,31,159,30,159,29,122,31,122,30,175,31,251,31,78,31,78,30,217,31,72,31,232,31,232,30,154,31,178,31,206,31,206,30,166,31,166,30,148,31,21,31,102,31,224,31,193,31,185,31,61,31,129,31,56,31,149,31,92,31,103,31,103,30,246,31,135,31,231,31,143,31,3,31,3,30,236,31,45,31,9,31,9,30,134,31,168,31,187,31,135,31,4,31,114,31,252,31,236,31,203,31,217,31,123,31,181,31,106,31,122,31,229,31,167,31,178,31,178,30,251,31,17,31,251,31,183,31,22,31,34,31,34,30,189,31,194,31,194,30,13,31,13,30,89,31,134,31,197,31,206,31,132,31,84,31,143,31,79,31,164,31,42,31,110,31,110,30,110,29,86,31,227,31,122,31,122,30,234,31,234,30,151,31,198,31,6,31,179,31,155,31,155,30,178,31,97,31,97,30,119,31,143,31,250,31,250,30,118,31,180,31,121,31,121,30,121,29,105,31,71,31,127,31,16,31,247,31,97,31,117,31,36,31,68,31,22,31,22,30,107,31,127,31,123,31,136,31,91,31,91,30,141,31,9,31,9,30,26,31,26,30,26,29,89,31,106,31,124,31,186,31,60,31,9,31,121,31,84,31,159,31,63,31,53,31,218,31,124,31,103,31,108,31,108,30,172,31,155,31,49,31,21,31,21,30,195,31,57,31,229,31,229,30,229,29,87,31,249,31,122,31,1,31,164,31,147,31,154,31,57,31,57,30,194,31,33,31,193,31,62,31,105,31,110,31,159,31,159,30,149,31,177,31,249,31,249,30,133,31,200,31,53,31,189,31,189,30,189,29,51,31,46,31,46,30,23,31,190,31,190,30,190,29,82,31,152,31,152,30,170,31,20,31,144,31,76,31,65,31,48,31,249,31,47,31,204,31,196,31,217,31,97,31,85,31,251,31,103,31,222,31,230,31,211,31,200,31,195,31,195,30,172,31,94,31,94,30,146,31,143,31,96,31,52,31,47,31,178,31,148,31,214,31,247,31,247,30,222,31,235,31,73,31,54,31,9,31,50,31,247,31,140,31,49,31,175,31,122,31,122,30,216,31,254,31,80,31,252,31,24,31,209,31,113,31,253,31,94,31,218,31,121,31,121,30,5,31,235,31,134,31,134,30,134,29,49,31,59,31,185,31,243,31,156,31,34,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
