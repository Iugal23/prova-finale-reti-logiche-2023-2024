-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 631;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (235,0,68,0,82,0,112,0,217,0,100,0,118,0,174,0,78,0,0,0,197,0,66,0,0,0,143,0,13,0,128,0,100,0,60,0,24,0,0,0,58,0,147,0,199,0,157,0,56,0,0,0,194,0,234,0,0,0,156,0,120,0,95,0,250,0,225,0,134,0,118,0,141,0,0,0,183,0,145,0,150,0,0,0,149,0,0,0,102,0,201,0,56,0,0,0,0,0,59,0,0,0,200,0,106,0,242,0,139,0,10,0,199,0,27,0,148,0,226,0,135,0,0,0,47,0,204,0,104,0,2,0,80,0,207,0,114,0,194,0,0,0,209,0,229,0,145,0,80,0,0,0,50,0,224,0,239,0,65,0,98,0,0,0,194,0,174,0,139,0,59,0,84,0,84,0,84,0,104,0,51,0,156,0,0,0,127,0,0,0,0,0,192,0,191,0,237,0,0,0,206,0,78,0,78,0,172,0,117,0,96,0,126,0,29,0,38,0,128,0,171,0,132,0,120,0,83,0,232,0,0,0,0,0,0,0,18,0,242,0,82,0,41,0,149,0,93,0,215,0,224,0,43,0,163,0,98,0,247,0,221,0,168,0,0,0,180,0,47,0,52,0,222,0,46,0,34,0,38,0,0,0,162,0,0,0,230,0,85,0,180,0,178,0,0,0,148,0,193,0,0,0,112,0,0,0,138,0,200,0,152,0,214,0,241,0,170,0,179,0,43,0,33,0,0,0,13,0,39,0,11,0,51,0,66,0,183,0,192,0,45,0,0,0,184,0,231,0,59,0,236,0,195,0,205,0,116,0,162,0,0,0,212,0,196,0,91,0,161,0,157,0,176,0,225,0,139,0,5,0,228,0,0,0,0,0,55,0,54,0,27,0,2,0,212,0,111,0,70,0,39,0,43,0,0,0,167,0,147,0,0,0,119,0,46,0,35,0,16,0,0,0,82,0,225,0,0,0,60,0,111,0,72,0,38,0,177,0,163,0,0,0,234,0,0,0,0,0,50,0,160,0,133,0,123,0,59,0,87,0,96,0,153,0,101,0,13,0,0,0,0,0,251,0,238,0,16,0,176,0,71,0,123,0,159,0,161,0,0,0,158,0,255,0,140,0,75,0,141,0,19,0,9,0,199,0,183,0,224,0,0,0,173,0,0,0,68,0,98,0,227,0,169,0,155,0,235,0,43,0,85,0,2,0,173,0,79,0,125,0,208,0,77,0,241,0,218,0,164,0,0,0,111,0,47,0,134,0,137,0,207,0,189,0,231,0,59,0,204,0,237,0,92,0,119,0,38,0,211,0,160,0,205,0,81,0,211,0,121,0,64,0,185,0,199,0,111,0,0,0,152,0,0,0,43,0,0,0,90,0,116,0,135,0,126,0,164,0,0,0,64,0,0,0,8,0,0,0,180,0,30,0,45,0,0,0,143,0,130,0,189,0,18,0,110,0,210,0,143,0,184,0,241,0,106,0,199,0,205,0,61,0,139,0,5,0,99,0,53,0,0,0,116,0,182,0,173,0,67,0,145,0,162,0,26,0,48,0,37,0,216,0,153,0,131,0,0,0,40,0,25,0,0,0,48,0,7,0,222,0,193,0,51,0,114,0,112,0,0,0,41,0,250,0,119,0,0,0,174,0,48,0,55,0,37,0,28,0,199,0,106,0,0,0,31,0,14,0,21,0,0,0,0,0,234,0,100,0,99,0,10,0,242,0,43,0,44,0,159,0,224,0,208,0,240,0,96,0,53,0,129,0,0,0,0,0,59,0,70,0,107,0,24,0,0,0,157,0,0,0,0,0,0,0,74,0,31,0,24,0,120,0,45,0,20,0,0,0,106,0,26,0,215,0,39,0,46,0,206,0,7,0,58,0,248,0,49,0,130,0,250,0,0,0,147,0,0,0,177,0,12,0,229,0,195,0,176,0,124,0,141,0,245,0,99,0,0,0,51,0,191,0,215,0,255,0,176,0,183,0,243,0,94,0,37,0,224,0,144,0,109,0,213,0,19,0,66,0,188,0,10,0,0,0,0,0,255,0,0,0,11,0,239,0,226,0,220,0,69,0,117,0,0,0,158,0,199,0,0,0,0,0,12,0,110,0,45,0,105,0,0,0,93,0,11,0,125,0,60,0,47,0,237,0,165,0,107,0,100,0,206,0,51,0,170,0,5,0,140,0,145,0,47,0,190,0,10,0,135,0,18,0,0,0,148,0,99,0,88,0,0,0,174,0,0,0,253,0,0,0,235,0,204,0,76,0,249,0,0,0,246,0,87,0,200,0,181,0,101,0,20,0,131,0,46,0,0,0,123,0,0,0,137,0,192,0,69,0,0,0,200,0,243,0,0,0,54,0,142,0,203,0,155,0,32,0,222,0,6,0,42,0,133,0,115,0,236,0,0,0,0,0,131,0,95,0,196,0,185,0,145,0,0,0,8,0,232,0,0,0,17,0,144,0,15,0,167,0,195,0,66,0,223,0,54,0,0,0,176,0,75,0,160,0,192,0,2,0,50,0,59,0,2,0,244,0,253,0,123,0,138,0,75,0,242,0,41,0,158,0,162,0,246,0,0,0,70,0,0,0,127,0,0,0,0,0,0,0,139,0,43,0,0,0,242,0,86,0,153,0,0,0,191,0,0,0,76,0,238,0,130,0,142,0,34,0,197,0,128,0,131,0,132,0,21,0,30,0,0,0,177,0,5,0,0,0,219,0,238,0,155,0,220,0,103,0,198,0,69,0,167,0,231,0,0,0,111,0,0,0,0,0,0,0,63,0,45,0,251,0,101,0,0,0,134,0,220,0,199,0,227,0,64,0,183,0,0,0,142,0,0,0);
signal scenario_full  : scenario_type := (235,31,68,31,82,31,112,31,217,31,100,31,118,31,174,31,78,31,78,30,197,31,66,31,66,30,143,31,13,31,128,31,100,31,60,31,24,31,24,30,58,31,147,31,199,31,157,31,56,31,56,30,194,31,234,31,234,30,156,31,120,31,95,31,250,31,225,31,134,31,118,31,141,31,141,30,183,31,145,31,150,31,150,30,149,31,149,30,102,31,201,31,56,31,56,30,56,29,59,31,59,30,200,31,106,31,242,31,139,31,10,31,199,31,27,31,148,31,226,31,135,31,135,30,47,31,204,31,104,31,2,31,80,31,207,31,114,31,194,31,194,30,209,31,229,31,145,31,80,31,80,30,50,31,224,31,239,31,65,31,98,31,98,30,194,31,174,31,139,31,59,31,84,31,84,31,84,31,104,31,51,31,156,31,156,30,127,31,127,30,127,29,192,31,191,31,237,31,237,30,206,31,78,31,78,31,172,31,117,31,96,31,126,31,29,31,38,31,128,31,171,31,132,31,120,31,83,31,232,31,232,30,232,29,232,28,18,31,242,31,82,31,41,31,149,31,93,31,215,31,224,31,43,31,163,31,98,31,247,31,221,31,168,31,168,30,180,31,47,31,52,31,222,31,46,31,34,31,38,31,38,30,162,31,162,30,230,31,85,31,180,31,178,31,178,30,148,31,193,31,193,30,112,31,112,30,138,31,200,31,152,31,214,31,241,31,170,31,179,31,43,31,33,31,33,30,13,31,39,31,11,31,51,31,66,31,183,31,192,31,45,31,45,30,184,31,231,31,59,31,236,31,195,31,205,31,116,31,162,31,162,30,212,31,196,31,91,31,161,31,157,31,176,31,225,31,139,31,5,31,228,31,228,30,228,29,55,31,54,31,27,31,2,31,212,31,111,31,70,31,39,31,43,31,43,30,167,31,147,31,147,30,119,31,46,31,35,31,16,31,16,30,82,31,225,31,225,30,60,31,111,31,72,31,38,31,177,31,163,31,163,30,234,31,234,30,234,29,50,31,160,31,133,31,123,31,59,31,87,31,96,31,153,31,101,31,13,31,13,30,13,29,251,31,238,31,16,31,176,31,71,31,123,31,159,31,161,31,161,30,158,31,255,31,140,31,75,31,141,31,19,31,9,31,199,31,183,31,224,31,224,30,173,31,173,30,68,31,98,31,227,31,169,31,155,31,235,31,43,31,85,31,2,31,173,31,79,31,125,31,208,31,77,31,241,31,218,31,164,31,164,30,111,31,47,31,134,31,137,31,207,31,189,31,231,31,59,31,204,31,237,31,92,31,119,31,38,31,211,31,160,31,205,31,81,31,211,31,121,31,64,31,185,31,199,31,111,31,111,30,152,31,152,30,43,31,43,30,90,31,116,31,135,31,126,31,164,31,164,30,64,31,64,30,8,31,8,30,180,31,30,31,45,31,45,30,143,31,130,31,189,31,18,31,110,31,210,31,143,31,184,31,241,31,106,31,199,31,205,31,61,31,139,31,5,31,99,31,53,31,53,30,116,31,182,31,173,31,67,31,145,31,162,31,26,31,48,31,37,31,216,31,153,31,131,31,131,30,40,31,25,31,25,30,48,31,7,31,222,31,193,31,51,31,114,31,112,31,112,30,41,31,250,31,119,31,119,30,174,31,48,31,55,31,37,31,28,31,199,31,106,31,106,30,31,31,14,31,21,31,21,30,21,29,234,31,100,31,99,31,10,31,242,31,43,31,44,31,159,31,224,31,208,31,240,31,96,31,53,31,129,31,129,30,129,29,59,31,70,31,107,31,24,31,24,30,157,31,157,30,157,29,157,28,74,31,31,31,24,31,120,31,45,31,20,31,20,30,106,31,26,31,215,31,39,31,46,31,206,31,7,31,58,31,248,31,49,31,130,31,250,31,250,30,147,31,147,30,177,31,12,31,229,31,195,31,176,31,124,31,141,31,245,31,99,31,99,30,51,31,191,31,215,31,255,31,176,31,183,31,243,31,94,31,37,31,224,31,144,31,109,31,213,31,19,31,66,31,188,31,10,31,10,30,10,29,255,31,255,30,11,31,239,31,226,31,220,31,69,31,117,31,117,30,158,31,199,31,199,30,199,29,12,31,110,31,45,31,105,31,105,30,93,31,11,31,125,31,60,31,47,31,237,31,165,31,107,31,100,31,206,31,51,31,170,31,5,31,140,31,145,31,47,31,190,31,10,31,135,31,18,31,18,30,148,31,99,31,88,31,88,30,174,31,174,30,253,31,253,30,235,31,204,31,76,31,249,31,249,30,246,31,87,31,200,31,181,31,101,31,20,31,131,31,46,31,46,30,123,31,123,30,137,31,192,31,69,31,69,30,200,31,243,31,243,30,54,31,142,31,203,31,155,31,32,31,222,31,6,31,42,31,133,31,115,31,236,31,236,30,236,29,131,31,95,31,196,31,185,31,145,31,145,30,8,31,232,31,232,30,17,31,144,31,15,31,167,31,195,31,66,31,223,31,54,31,54,30,176,31,75,31,160,31,192,31,2,31,50,31,59,31,2,31,244,31,253,31,123,31,138,31,75,31,242,31,41,31,158,31,162,31,246,31,246,30,70,31,70,30,127,31,127,30,127,29,127,28,139,31,43,31,43,30,242,31,86,31,153,31,153,30,191,31,191,30,76,31,238,31,130,31,142,31,34,31,197,31,128,31,131,31,132,31,21,31,30,31,30,30,177,31,5,31,5,30,219,31,238,31,155,31,220,31,103,31,198,31,69,31,167,31,231,31,231,30,111,31,111,30,111,29,111,28,63,31,45,31,251,31,101,31,101,30,134,31,220,31,199,31,227,31,64,31,183,31,183,30,142,31,142,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
