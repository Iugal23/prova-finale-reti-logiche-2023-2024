-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_168 is
end project_tb_168;

architecture project_tb_arch_168 of project_tb_168 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 650;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (140,0,127,0,0,0,0,0,167,0,149,0,196,0,54,0,0,0,77,0,216,0,94,0,85,0,210,0,171,0,2,0,0,0,41,0,164,0,133,0,198,0,78,0,112,0,255,0,0,0,151,0,0,0,74,0,143,0,50,0,247,0,0,0,202,0,212,0,167,0,122,0,19,0,132,0,106,0,59,0,0,0,33,0,225,0,79,0,0,0,134,0,0,0,55,0,196,0,185,0,0,0,0,0,72,0,0,0,78,0,112,0,107,0,18,0,0,0,0,0,0,0,71,0,0,0,25,0,0,0,198,0,3,0,76,0,168,0,6,0,244,0,160,0,54,0,60,0,182,0,114,0,127,0,0,0,32,0,161,0,254,0,0,0,253,0,182,0,169,0,161,0,119,0,235,0,0,0,221,0,0,0,194,0,141,0,255,0,0,0,0,0,98,0,165,0,217,0,62,0,118,0,111,0,78,0,16,0,96,0,171,0,0,0,15,0,16,0,19,0,5,0,84,0,239,0,141,0,196,0,28,0,70,0,0,0,54,0,228,0,139,0,94,0,254,0,0,0,129,0,0,0,116,0,74,0,248,0,139,0,247,0,171,0,27,0,244,0,123,0,0,0,84,0,143,0,253,0,88,0,74,0,192,0,0,0,238,0,241,0,59,0,120,0,120,0,131,0,177,0,8,0,103,0,157,0,29,0,38,0,214,0,122,0,56,0,226,0,225,0,188,0,193,0,251,0,54,0,10,0,191,0,204,0,0,0,69,0,248,0,202,0,49,0,22,0,237,0,0,0,0,0,0,0,216,0,0,0,0,0,161,0,200,0,91,0,241,0,35,0,78,0,10,0,0,0,73,0,183,0,153,0,105,0,171,0,146,0,16,0,230,0,82,0,198,0,157,0,77,0,185,0,10,0,41,0,0,0,202,0,180,0,86,0,0,0,110,0,251,0,25,0,99,0,181,0,3,0,58,0,245,0,187,0,191,0,236,0,57,0,155,0,0,0,248,0,11,0,0,0,47,0,129,0,68,0,127,0,207,0,0,0,231,0,36,0,255,0,157,0,197,0,116,0,188,0,224,0,0,0,65,0,0,0,28,0,164,0,107,0,34,0,45,0,161,0,74,0,0,0,183,0,116,0,248,0,0,0,23,0,208,0,177,0,105,0,17,0,95,0,95,0,165,0,239,0,144,0,201,0,0,0,0,0,86,0,0,0,199,0,0,0,0,0,135,0,24,0,177,0,31,0,13,0,57,0,0,0,56,0,245,0,228,0,48,0,0,0,61,0,174,0,97,0,162,0,236,0,90,0,207,0,223,0,192,0,255,0,152,0,0,0,0,0,178,0,215,0,0,0,247,0,250,0,0,0,168,0,7,0,133,0,76,0,181,0,80,0,36,0,198,0,0,0,0,0,20,0,0,0,200,0,130,0,64,0,75,0,5,0,116,0,13,0,0,0,0,0,221,0,250,0,0,0,148,0,36,0,154,0,217,0,181,0,245,0,118,0,55,0,218,0,107,0,0,0,0,0,249,0,0,0,217,0,60,0,0,0,126,0,22,0,27,0,108,0,99,0,151,0,249,0,53,0,112,0,132,0,166,0,70,0,180,0,84,0,112,0,213,0,220,0,0,0,118,0,0,0,188,0,82,0,65,0,0,0,174,0,29,0,33,0,177,0,0,0,0,0,0,0,255,0,214,0,121,0,249,0,8,0,127,0,0,0,143,0,170,0,0,0,211,0,179,0,0,0,18,0,90,0,79,0,109,0,36,0,88,0,63,0,157,0,91,0,78,0,197,0,160,0,241,0,253,0,248,0,197,0,0,0,0,0,0,0,26,0,12,0,0,0,239,0,0,0,0,0,0,0,183,0,151,0,76,0,47,0,181,0,248,0,103,0,0,0,155,0,0,0,240,0,213,0,155,0,75,0,69,0,124,0,227,0,197,0,134,0,219,0,251,0,249,0,224,0,150,0,69,0,240,0,210,0,118,0,175,0,27,0,41,0,246,0,68,0,111,0,0,0,202,0,124,0,2,0,58,0,32,0,122,0,143,0,216,0,127,0,24,0,251,0,0,0,0,0,6,0,31,0,241,0,242,0,216,0,217,0,0,0,105,0,0,0,0,0,116,0,182,0,217,0,54,0,173,0,0,0,31,0,156,0,238,0,250,0,208,0,12,0,0,0,34,0,142,0,133,0,0,0,9,0,239,0,248,0,116,0,2,0,111,0,180,0,0,0,48,0,115,0,112,0,125,0,93,0,113,0,206,0,152,0,65,0,55,0,171,0,71,0,125,0,244,0,240,0,244,0,245,0,64,0,0,0,26,0,0,0,205,0,133,0,0,0,0,0,165,0,5,0,116,0,80,0,152,0,211,0,0,0,134,0,0,0,172,0,0,0,0,0,208,0,147,0,5,0,0,0,148,0,0,0,36,0,176,0,24,0,195,0,197,0,0,0,87,0,19,0,8,0,213,0,0,0,54,0,0,0,8,0,190,0,62,0,116,0,223,0,89,0,0,0,17,0,205,0,87,0,162,0,196,0,151,0,41,0,244,0,145,0,170,0,133,0,0,0,251,0,186,0,94,0,137,0,20,0,187,0,249,0,80,0,0,0,90,0,0,0,188,0,107,0,254,0,255,0,87,0,43,0,147,0,111,0,148,0,235,0,131,0,38,0,219,0,0,0,131,0,0,0,75,0,220,0,0,0,100,0,0,0,10,0,128,0,0,0,212,0,68,0,10,0,131,0,240,0,151,0,73,0,204,0,0,0,2,0,0,0,45,0,74,0,119,0,66,0,0,0,109,0,0,0,142,0,57,0,0,0,250,0,127,0,70,0,128,0,108,0,143,0,147,0,0,0,0,0,0,0,211,0,37,0,202,0,3,0,0,0,17,0,50,0,70,0,0,0,230,0,17,0,211,0);
signal scenario_full  : scenario_type := (140,31,127,31,127,30,127,29,167,31,149,31,196,31,54,31,54,30,77,31,216,31,94,31,85,31,210,31,171,31,2,31,2,30,41,31,164,31,133,31,198,31,78,31,112,31,255,31,255,30,151,31,151,30,74,31,143,31,50,31,247,31,247,30,202,31,212,31,167,31,122,31,19,31,132,31,106,31,59,31,59,30,33,31,225,31,79,31,79,30,134,31,134,30,55,31,196,31,185,31,185,30,185,29,72,31,72,30,78,31,112,31,107,31,18,31,18,30,18,29,18,28,71,31,71,30,25,31,25,30,198,31,3,31,76,31,168,31,6,31,244,31,160,31,54,31,60,31,182,31,114,31,127,31,127,30,32,31,161,31,254,31,254,30,253,31,182,31,169,31,161,31,119,31,235,31,235,30,221,31,221,30,194,31,141,31,255,31,255,30,255,29,98,31,165,31,217,31,62,31,118,31,111,31,78,31,16,31,96,31,171,31,171,30,15,31,16,31,19,31,5,31,84,31,239,31,141,31,196,31,28,31,70,31,70,30,54,31,228,31,139,31,94,31,254,31,254,30,129,31,129,30,116,31,74,31,248,31,139,31,247,31,171,31,27,31,244,31,123,31,123,30,84,31,143,31,253,31,88,31,74,31,192,31,192,30,238,31,241,31,59,31,120,31,120,31,131,31,177,31,8,31,103,31,157,31,29,31,38,31,214,31,122,31,56,31,226,31,225,31,188,31,193,31,251,31,54,31,10,31,191,31,204,31,204,30,69,31,248,31,202,31,49,31,22,31,237,31,237,30,237,29,237,28,216,31,216,30,216,29,161,31,200,31,91,31,241,31,35,31,78,31,10,31,10,30,73,31,183,31,153,31,105,31,171,31,146,31,16,31,230,31,82,31,198,31,157,31,77,31,185,31,10,31,41,31,41,30,202,31,180,31,86,31,86,30,110,31,251,31,25,31,99,31,181,31,3,31,58,31,245,31,187,31,191,31,236,31,57,31,155,31,155,30,248,31,11,31,11,30,47,31,129,31,68,31,127,31,207,31,207,30,231,31,36,31,255,31,157,31,197,31,116,31,188,31,224,31,224,30,65,31,65,30,28,31,164,31,107,31,34,31,45,31,161,31,74,31,74,30,183,31,116,31,248,31,248,30,23,31,208,31,177,31,105,31,17,31,95,31,95,31,165,31,239,31,144,31,201,31,201,30,201,29,86,31,86,30,199,31,199,30,199,29,135,31,24,31,177,31,31,31,13,31,57,31,57,30,56,31,245,31,228,31,48,31,48,30,61,31,174,31,97,31,162,31,236,31,90,31,207,31,223,31,192,31,255,31,152,31,152,30,152,29,178,31,215,31,215,30,247,31,250,31,250,30,168,31,7,31,133,31,76,31,181,31,80,31,36,31,198,31,198,30,198,29,20,31,20,30,200,31,130,31,64,31,75,31,5,31,116,31,13,31,13,30,13,29,221,31,250,31,250,30,148,31,36,31,154,31,217,31,181,31,245,31,118,31,55,31,218,31,107,31,107,30,107,29,249,31,249,30,217,31,60,31,60,30,126,31,22,31,27,31,108,31,99,31,151,31,249,31,53,31,112,31,132,31,166,31,70,31,180,31,84,31,112,31,213,31,220,31,220,30,118,31,118,30,188,31,82,31,65,31,65,30,174,31,29,31,33,31,177,31,177,30,177,29,177,28,255,31,214,31,121,31,249,31,8,31,127,31,127,30,143,31,170,31,170,30,211,31,179,31,179,30,18,31,90,31,79,31,109,31,36,31,88,31,63,31,157,31,91,31,78,31,197,31,160,31,241,31,253,31,248,31,197,31,197,30,197,29,197,28,26,31,12,31,12,30,239,31,239,30,239,29,239,28,183,31,151,31,76,31,47,31,181,31,248,31,103,31,103,30,155,31,155,30,240,31,213,31,155,31,75,31,69,31,124,31,227,31,197,31,134,31,219,31,251,31,249,31,224,31,150,31,69,31,240,31,210,31,118,31,175,31,27,31,41,31,246,31,68,31,111,31,111,30,202,31,124,31,2,31,58,31,32,31,122,31,143,31,216,31,127,31,24,31,251,31,251,30,251,29,6,31,31,31,241,31,242,31,216,31,217,31,217,30,105,31,105,30,105,29,116,31,182,31,217,31,54,31,173,31,173,30,31,31,156,31,238,31,250,31,208,31,12,31,12,30,34,31,142,31,133,31,133,30,9,31,239,31,248,31,116,31,2,31,111,31,180,31,180,30,48,31,115,31,112,31,125,31,93,31,113,31,206,31,152,31,65,31,55,31,171,31,71,31,125,31,244,31,240,31,244,31,245,31,64,31,64,30,26,31,26,30,205,31,133,31,133,30,133,29,165,31,5,31,116,31,80,31,152,31,211,31,211,30,134,31,134,30,172,31,172,30,172,29,208,31,147,31,5,31,5,30,148,31,148,30,36,31,176,31,24,31,195,31,197,31,197,30,87,31,19,31,8,31,213,31,213,30,54,31,54,30,8,31,190,31,62,31,116,31,223,31,89,31,89,30,17,31,205,31,87,31,162,31,196,31,151,31,41,31,244,31,145,31,170,31,133,31,133,30,251,31,186,31,94,31,137,31,20,31,187,31,249,31,80,31,80,30,90,31,90,30,188,31,107,31,254,31,255,31,87,31,43,31,147,31,111,31,148,31,235,31,131,31,38,31,219,31,219,30,131,31,131,30,75,31,220,31,220,30,100,31,100,30,10,31,128,31,128,30,212,31,68,31,10,31,131,31,240,31,151,31,73,31,204,31,204,30,2,31,2,30,45,31,74,31,119,31,66,31,66,30,109,31,109,30,142,31,57,31,57,30,250,31,127,31,70,31,128,31,108,31,143,31,147,31,147,30,147,29,147,28,211,31,37,31,202,31,3,31,3,30,17,31,50,31,70,31,70,30,230,31,17,31,211,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
