-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_221 is
end project_tb_221;

architecture project_tb_arch_221 of project_tb_221 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (17,0,173,0,24,0,233,0,0,0,172,0,61,0,0,0,169,0,200,0,2,0,201,0,105,0,0,0,137,0,196,0,181,0,0,0,0,0,19,0,0,0,153,0,137,0,244,0,0,0,170,0,38,0,51,0,0,0,170,0,71,0,57,0,0,0,239,0,29,0,132,0,206,0,110,0,115,0,245,0,0,0,153,0,81,0,182,0,0,0,42,0,253,0,37,0,11,0,239,0,29,0,219,0,117,0,214,0,205,0,0,0,169,0,82,0,40,0,157,0,213,0,73,0,0,0,154,0,35,0,171,0,39,0,125,0,252,0,245,0,0,0,0,0,49,0,254,0,0,0,254,0,72,0,113,0,125,0,62,0,0,0,185,0,140,0,22,0,161,0,0,0,70,0,121,0,0,0,0,0,215,0,31,0,0,0,52,0,106,0,58,0,255,0,0,0,169,0,192,0,232,0,87,0,127,0,122,0,45,0,0,0,235,0,196,0,23,0,0,0,0,0,97,0,188,0,0,0,254,0,0,0,0,0,50,0,128,0,178,0,162,0,0,0,66,0,164,0,0,0,0,0,0,0,138,0,0,0,14,0,14,0,220,0,74,0,92,0,162,0,236,0,61,0,95,0,0,0,35,0,148,0,25,0,18,0,233,0,0,0,224,0,31,0,109,0,126,0,218,0,131,0,253,0,199,0,50,0,36,0,206,0,255,0,181,0,0,0,0,0,0,0,8,0,225,0,22,0,0,0,18,0,156,0,149,0,98,0,207,0,30,0,145,0,231,0,202,0,30,0,13,0,0,0,0,0,0,0,133,0,228,0,122,0,173,0,9,0,203,0,39,0,74,0,176,0,102,0,44,0,0,0,196,0,150,0,129,0,153,0,173,0,0,0,99,0,199,0,187,0,49,0,183,0,171,0,112,0,0,0,0,0,157,0,221,0,100,0,110,0,241,0,55,0,62,0,0,0,195,0,47,0,141,0,0,0,149,0,53,0,252,0,20,0,28,0,31,0,190,0,215,0,25,0,0,0,7,0,154,0,153,0,68,0,17,0,118,0,234,0,106,0,218,0,0,0,199,0,5,0,0,0,0,0,115,0,122,0,0,0,147,0,30,0,250,0,148,0,193,0,66,0,0,0,0,0,248,0,0,0,0,0,159,0,1,0,89,0,56,0,15,0,6,0,70,0,168,0,15,0,0,0,37,0,178,0,14,0,73,0,182,0,104,0,116,0,0,0,106,0,2,0,14,0,246,0,179,0,132,0,162,0,165,0,82,0,0,0,97,0,0,0,252,0,123,0,103,0,1,0,114,0,231,0,85,0,87,0,215,0,56,0,243,0,77,0,30,0,17,0,117,0,58,0,222,0,21,0,93,0,52,0,0,0,69,0,83,0,59,0,248,0,74,0,73,0,24,0,215,0,6,0,0,0,0,0,180,0,92,0,0,0,0,0,0,0,0,0,48,0,0,0,63,0,51,0,0,0,81,0,174,0,16,0,38,0,138,0,58,0,72,0,197,0,0,0,15,0,0,0,139,0,16,0,0,0,14,0,83,0,185,0,121,0,94,0,0,0,0,0,170,0,196,0,14,0,7,0,14,0,35,0,86,0,162,0,0,0,123,0,0,0,54,0,0,0,45,0,225,0,198,0,79,0,133,0,24,0,0,0,76,0,128,0,0,0,137,0,238,0,0,0,24,0,0,0,6,0,177,0,0,0,230,0,46,0,113,0,42,0,0,0,9,0,100,0,240,0,26,0,100,0,0,0,0,0,212,0,0,0,210,0,161,0,192,0,126,0,106,0,100,0,82,0,253,0,91,0,20,0,229,0,0,0,88,0,218,0,244,0,108,0,141,0,173,0,0,0,28,0,4,0,83,0,173,0,167,0,197,0,0,0,159,0,0,0,194,0,24,0,197,0,237,0,83,0,191,0,189,0,225,0,141,0,169,0,75,0,0,0,17,0,31,0,146,0,145,0,40,0,174,0,50,0,139,0,14,0,16,0,244,0,54,0,28,0,215,0,14,0,190,0,122,0,73,0,0,0,0,0,38,0,188,0,165,0,144,0,53,0,32,0,252,0,236,0,0,0,108,0,173,0,24,0,93,0,216,0,0,0,0,0,118,0,57,0,47,0,0,0,175,0,193,0,162,0,0,0,232,0,0,0,0,0,193,0,72,0,0,0,117,0,254,0,0,0,215,0,67,0,130,0,0,0,147,0,1,0,5,0,230,0,64,0,123,0,202,0,131,0,71,0,0,0,124,0,70,0,205,0,0,0,173,0,0,0,235,0,21,0,251,0,183,0,0,0,0,0,39,0,245,0,213,0,0,0,0,0,227,0,143,0,0,0,37,0,175,0,18,0,13,0,38,0,114,0,38,0,35,0,0,0,0,0,0,0,13,0,0,0,178,0,223,0,69,0,55,0,175,0,0,0,219,0,43,0,83,0,0,0,187,0,56,0,77,0,0,0,110,0,128,0,210,0,51,0,192,0,78,0,91,0,227,0,248,0,102,0,1,0,97,0,62,0,0,0,180,0,0,0,204,0,42,0,0,0,38,0,243,0,192,0,209,0,255,0,222,0,132,0,127,0,0,0,161,0,51,0,108,0,179,0,5,0,215,0,198,0,205,0,112,0,192,0,0,0,254,0,111,0,0,0,140,0,87,0,88,0,119,0,162,0,0,0,96,0,121,0,160,0,0,0,94,0,188,0,84,0,180,0,97,0,100,0,0,0,15,0,0,0,212,0,125,0,229,0,154,0,57,0,59,0,173,0,19,0,114,0,107,0,190,0,176,0,0,0,117,0,72,0,95,0,147,0,155,0,0,0,58,0,0,0,14,0,131,0,4,0,47,0,23,0,0,0,195,0,0,0,0,0,239,0,0,0,178,0,47,0,143,0,150,0,176,0,0,0,0,0,168,0,220,0,162,0,113,0,0,0,95,0,0,0,0,0,226,0,219,0,186,0,33,0,0,0,67,0,0,0,123,0,29,0,129,0,73,0,0,0,134,0,217,0,130,0,193,0,126,0,209,0,0,0,101,0,232,0,117,0,0,0,40,0,151,0,245,0,144,0,44,0,111,0,130,0,158,0,0,0,216,0,254,0,114,0,18,0,175,0,33,0,190,0,243,0,138,0,56,0,121,0,121,0,153,0,11,0,244,0,0,0,212,0,240,0,0,0,1,0,193,0,2,0,135,0,0,0,145,0,22,0,204,0,85,0,115,0,184,0,152,0,100,0,0,0,21,0,63,0,151,0,138,0,206,0,0,0,231,0,32,0,59,0,135,0,0,0,163,0,231,0,145,0,127,0,0,0,14,0,132,0,0,0,58,0,0,0,196,0,186,0,0,0,79,0,0,0,225,0,0,0,0,0,0,0,40,0,242,0,166,0,0,0,162,0,22,0,107,0,79,0,0,0,98,0,0,0,0,0,126,0,234,0,130,0,42,0,238,0,177,0,110,0,194,0,191,0,103,0,193,0,33,0,0,0,132,0,230,0,68,0,239,0,51,0,93,0,160,0,111,0,71,0,167,0,0,0,220,0,0,0,24,0,243,0,0,0,110,0,0,0,99,0,177,0,46,0,240,0,54,0,123,0,230,0,183,0,84,0,116,0,27,0,112,0,111,0,233,0,0,0,142,0,0,0,57,0,0,0,223,0,45,0,198,0,99,0,48,0,110,0,201,0,29,0,0,0,240,0,50,0,83,0,102,0,208,0,0,0,0,0,53,0,0,0,133,0,226,0,0,0,0,0,74,0,115,0,61,0,60,0,134,0,38,0,175,0,0,0,145,0,8,0,7,0,242,0,158,0,158,0,220,0,175,0,118,0,202,0,0,0,6,0,98,0);
signal scenario_full  : scenario_type := (17,31,173,31,24,31,233,31,233,30,172,31,61,31,61,30,169,31,200,31,2,31,201,31,105,31,105,30,137,31,196,31,181,31,181,30,181,29,19,31,19,30,153,31,137,31,244,31,244,30,170,31,38,31,51,31,51,30,170,31,71,31,57,31,57,30,239,31,29,31,132,31,206,31,110,31,115,31,245,31,245,30,153,31,81,31,182,31,182,30,42,31,253,31,37,31,11,31,239,31,29,31,219,31,117,31,214,31,205,31,205,30,169,31,82,31,40,31,157,31,213,31,73,31,73,30,154,31,35,31,171,31,39,31,125,31,252,31,245,31,245,30,245,29,49,31,254,31,254,30,254,31,72,31,113,31,125,31,62,31,62,30,185,31,140,31,22,31,161,31,161,30,70,31,121,31,121,30,121,29,215,31,31,31,31,30,52,31,106,31,58,31,255,31,255,30,169,31,192,31,232,31,87,31,127,31,122,31,45,31,45,30,235,31,196,31,23,31,23,30,23,29,97,31,188,31,188,30,254,31,254,30,254,29,50,31,128,31,178,31,162,31,162,30,66,31,164,31,164,30,164,29,164,28,138,31,138,30,14,31,14,31,220,31,74,31,92,31,162,31,236,31,61,31,95,31,95,30,35,31,148,31,25,31,18,31,233,31,233,30,224,31,31,31,109,31,126,31,218,31,131,31,253,31,199,31,50,31,36,31,206,31,255,31,181,31,181,30,181,29,181,28,8,31,225,31,22,31,22,30,18,31,156,31,149,31,98,31,207,31,30,31,145,31,231,31,202,31,30,31,13,31,13,30,13,29,13,28,133,31,228,31,122,31,173,31,9,31,203,31,39,31,74,31,176,31,102,31,44,31,44,30,196,31,150,31,129,31,153,31,173,31,173,30,99,31,199,31,187,31,49,31,183,31,171,31,112,31,112,30,112,29,157,31,221,31,100,31,110,31,241,31,55,31,62,31,62,30,195,31,47,31,141,31,141,30,149,31,53,31,252,31,20,31,28,31,31,31,190,31,215,31,25,31,25,30,7,31,154,31,153,31,68,31,17,31,118,31,234,31,106,31,218,31,218,30,199,31,5,31,5,30,5,29,115,31,122,31,122,30,147,31,30,31,250,31,148,31,193,31,66,31,66,30,66,29,248,31,248,30,248,29,159,31,1,31,89,31,56,31,15,31,6,31,70,31,168,31,15,31,15,30,37,31,178,31,14,31,73,31,182,31,104,31,116,31,116,30,106,31,2,31,14,31,246,31,179,31,132,31,162,31,165,31,82,31,82,30,97,31,97,30,252,31,123,31,103,31,1,31,114,31,231,31,85,31,87,31,215,31,56,31,243,31,77,31,30,31,17,31,117,31,58,31,222,31,21,31,93,31,52,31,52,30,69,31,83,31,59,31,248,31,74,31,73,31,24,31,215,31,6,31,6,30,6,29,180,31,92,31,92,30,92,29,92,28,92,27,48,31,48,30,63,31,51,31,51,30,81,31,174,31,16,31,38,31,138,31,58,31,72,31,197,31,197,30,15,31,15,30,139,31,16,31,16,30,14,31,83,31,185,31,121,31,94,31,94,30,94,29,170,31,196,31,14,31,7,31,14,31,35,31,86,31,162,31,162,30,123,31,123,30,54,31,54,30,45,31,225,31,198,31,79,31,133,31,24,31,24,30,76,31,128,31,128,30,137,31,238,31,238,30,24,31,24,30,6,31,177,31,177,30,230,31,46,31,113,31,42,31,42,30,9,31,100,31,240,31,26,31,100,31,100,30,100,29,212,31,212,30,210,31,161,31,192,31,126,31,106,31,100,31,82,31,253,31,91,31,20,31,229,31,229,30,88,31,218,31,244,31,108,31,141,31,173,31,173,30,28,31,4,31,83,31,173,31,167,31,197,31,197,30,159,31,159,30,194,31,24,31,197,31,237,31,83,31,191,31,189,31,225,31,141,31,169,31,75,31,75,30,17,31,31,31,146,31,145,31,40,31,174,31,50,31,139,31,14,31,16,31,244,31,54,31,28,31,215,31,14,31,190,31,122,31,73,31,73,30,73,29,38,31,188,31,165,31,144,31,53,31,32,31,252,31,236,31,236,30,108,31,173,31,24,31,93,31,216,31,216,30,216,29,118,31,57,31,47,31,47,30,175,31,193,31,162,31,162,30,232,31,232,30,232,29,193,31,72,31,72,30,117,31,254,31,254,30,215,31,67,31,130,31,130,30,147,31,1,31,5,31,230,31,64,31,123,31,202,31,131,31,71,31,71,30,124,31,70,31,205,31,205,30,173,31,173,30,235,31,21,31,251,31,183,31,183,30,183,29,39,31,245,31,213,31,213,30,213,29,227,31,143,31,143,30,37,31,175,31,18,31,13,31,38,31,114,31,38,31,35,31,35,30,35,29,35,28,13,31,13,30,178,31,223,31,69,31,55,31,175,31,175,30,219,31,43,31,83,31,83,30,187,31,56,31,77,31,77,30,110,31,128,31,210,31,51,31,192,31,78,31,91,31,227,31,248,31,102,31,1,31,97,31,62,31,62,30,180,31,180,30,204,31,42,31,42,30,38,31,243,31,192,31,209,31,255,31,222,31,132,31,127,31,127,30,161,31,51,31,108,31,179,31,5,31,215,31,198,31,205,31,112,31,192,31,192,30,254,31,111,31,111,30,140,31,87,31,88,31,119,31,162,31,162,30,96,31,121,31,160,31,160,30,94,31,188,31,84,31,180,31,97,31,100,31,100,30,15,31,15,30,212,31,125,31,229,31,154,31,57,31,59,31,173,31,19,31,114,31,107,31,190,31,176,31,176,30,117,31,72,31,95,31,147,31,155,31,155,30,58,31,58,30,14,31,131,31,4,31,47,31,23,31,23,30,195,31,195,30,195,29,239,31,239,30,178,31,47,31,143,31,150,31,176,31,176,30,176,29,168,31,220,31,162,31,113,31,113,30,95,31,95,30,95,29,226,31,219,31,186,31,33,31,33,30,67,31,67,30,123,31,29,31,129,31,73,31,73,30,134,31,217,31,130,31,193,31,126,31,209,31,209,30,101,31,232,31,117,31,117,30,40,31,151,31,245,31,144,31,44,31,111,31,130,31,158,31,158,30,216,31,254,31,114,31,18,31,175,31,33,31,190,31,243,31,138,31,56,31,121,31,121,31,153,31,11,31,244,31,244,30,212,31,240,31,240,30,1,31,193,31,2,31,135,31,135,30,145,31,22,31,204,31,85,31,115,31,184,31,152,31,100,31,100,30,21,31,63,31,151,31,138,31,206,31,206,30,231,31,32,31,59,31,135,31,135,30,163,31,231,31,145,31,127,31,127,30,14,31,132,31,132,30,58,31,58,30,196,31,186,31,186,30,79,31,79,30,225,31,225,30,225,29,225,28,40,31,242,31,166,31,166,30,162,31,22,31,107,31,79,31,79,30,98,31,98,30,98,29,126,31,234,31,130,31,42,31,238,31,177,31,110,31,194,31,191,31,103,31,193,31,33,31,33,30,132,31,230,31,68,31,239,31,51,31,93,31,160,31,111,31,71,31,167,31,167,30,220,31,220,30,24,31,243,31,243,30,110,31,110,30,99,31,177,31,46,31,240,31,54,31,123,31,230,31,183,31,84,31,116,31,27,31,112,31,111,31,233,31,233,30,142,31,142,30,57,31,57,30,223,31,45,31,198,31,99,31,48,31,110,31,201,31,29,31,29,30,240,31,50,31,83,31,102,31,208,31,208,30,208,29,53,31,53,30,133,31,226,31,226,30,226,29,74,31,115,31,61,31,60,31,134,31,38,31,175,31,175,30,145,31,8,31,7,31,242,31,158,31,158,31,220,31,175,31,118,31,202,31,202,30,6,31,98,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
