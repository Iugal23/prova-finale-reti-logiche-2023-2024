-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 610;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (124,0,61,0,173,0,155,0,91,0,213,0,50,0,181,0,33,0,211,0,178,0,0,0,142,0,121,0,0,0,97,0,217,0,0,0,102,0,192,0,0,0,151,0,226,0,239,0,8,0,249,0,0,0,196,0,240,0,53,0,0,0,89,0,231,0,252,0,33,0,0,0,0,0,131,0,93,0,169,0,0,0,244,0,0,0,251,0,9,0,128,0,92,0,59,0,155,0,234,0,213,0,56,0,8,0,123,0,146,0,220,0,55,0,211,0,230,0,3,0,134,0,0,0,199,0,21,0,4,0,0,0,0,0,149,0,63,0,0,0,238,0,63,0,107,0,183,0,79,0,25,0,221,0,23,0,0,0,55,0,192,0,178,0,0,0,216,0,90,0,166,0,0,0,155,0,134,0,15,0,119,0,76,0,121,0,132,0,114,0,244,0,180,0,229,0,177,0,37,0,230,0,73,0,75,0,173,0,123,0,243,0,166,0,245,0,0,0,13,0,231,0,106,0,67,0,141,0,142,0,62,0,193,0,36,0,192,0,170,0,240,0,25,0,203,0,40,0,74,0,59,0,14,0,173,0,134,0,38,0,179,0,246,0,164,0,0,0,177,0,70,0,38,0,96,0,87,0,148,0,13,0,231,0,137,0,0,0,17,0,0,0,214,0,113,0,0,0,197,0,236,0,117,0,107,0,226,0,78,0,232,0,39,0,126,0,72,0,158,0,240,0,184,0,0,0,186,0,0,0,191,0,160,0,203,0,11,0,190,0,237,0,208,0,0,0,125,0,254,0,221,0,73,0,118,0,194,0,155,0,248,0,130,0,36,0,150,0,129,0,152,0,73,0,85,0,62,0,0,0,14,0,23,0,0,0,0,0,0,0,173,0,97,0,0,0,67,0,181,0,59,0,23,0,34,0,72,0,114,0,88,0,2,0,11,0,68,0,33,0,16,0,153,0,77,0,115,0,0,0,211,0,82,0,189,0,186,0,205,0,0,0,248,0,161,0,38,0,41,0,156,0,48,0,25,0,251,0,70,0,124,0,236,0,17,0,254,0,125,0,111,0,0,0,144,0,112,0,242,0,228,0,120,0,122,0,230,0,23,0,119,0,196,0,163,0,250,0,89,0,0,0,102,0,32,0,161,0,0,0,7,0,11,0,100,0,91,0,148,0,224,0,0,0,163,0,25,0,0,0,0,0,216,0,179,0,247,0,0,0,136,0,0,0,0,0,231,0,125,0,0,0,175,0,0,0,212,0,91,0,67,0,115,0,211,0,197,0,128,0,156,0,0,0,247,0,45,0,156,0,0,0,24,0,155,0,90,0,33,0,247,0,0,0,0,0,229,0,0,0,0,0,181,0,145,0,154,0,61,0,0,0,228,0,103,0,165,0,223,0,1,0,62,0,246,0,52,0,252,0,245,0,175,0,104,0,67,0,215,0,183,0,132,0,16,0,0,0,219,0,68,0,122,0,0,0,0,0,0,0,34,0,0,0,0,0,119,0,68,0,122,0,223,0,198,0,0,0,29,0,0,0,46,0,54,0,149,0,0,0,43,0,0,0,80,0,113,0,149,0,221,0,218,0,0,0,238,0,240,0,160,0,89,0,118,0,0,0,118,0,40,0,109,0,32,0,0,0,9,0,107,0,97,0,111,0,244,0,224,0,200,0,193,0,250,0,59,0,22,0,5,0,37,0,0,0,37,0,114,0,123,0,131,0,65,0,216,0,126,0,89,0,126,0,232,0,86,0,212,0,69,0,131,0,148,0,135,0,194,0,0,0,28,0,0,0,146,0,93,0,172,0,197,0,115,0,0,0,194,0,216,0,71,0,248,0,98,0,65,0,0,0,189,0,237,0,0,0,117,0,117,0,0,0,235,0,194,0,0,0,152,0,44,0,65,0,106,0,243,0,247,0,10,0,85,0,238,0,205,0,87,0,155,0,204,0,216,0,102,0,203,0,215,0,110,0,0,0,161,0,41,0,83,0,42,0,0,0,105,0,35,0,204,0,34,0,104,0,10,0,65,0,166,0,200,0,49,0,0,0,200,0,0,0,113,0,193,0,224,0,223,0,127,0,145,0,16,0,240,0,244,0,118,0,183,0,82,0,0,0,6,0,225,0,214,0,28,0,0,0,134,0,0,0,178,0,214,0,9,0,233,0,117,0,215,0,114,0,97,0,7,0,210,0,54,0,157,0,153,0,252,0,0,0,128,0,205,0,0,0,242,0,92,0,103,0,0,0,182,0,121,0,137,0,0,0,0,0,8,0,57,0,86,0,0,0,13,0,193,0,59,0,227,0,222,0,3,0,132,0,0,0,44,0,18,0,0,0,0,0,65,0,193,0,32,0,125,0,173,0,0,0,62,0,158,0,107,0,77,0,0,0,239,0,120,0,223,0,184,0,222,0,45,0,18,0,109,0,77,0,79,0,220,0,228,0,98,0,0,0,57,0,220,0,99,0,187,0,5,0,0,0,23,0,0,0,185,0,0,0,0,0,94,0,222,0,110,0,0,0,164,0,11,0,206,0,0,0,31,0,42,0,160,0,91,0,0,0,128,0,161,0,148,0,121,0,59,0,42,0,163,0,0,0,254,0,0,0,20,0,97,0,242,0,205,0,49,0,0,0,228,0,120,0,90,0,0,0,17,0,97,0,111,0,245,0,198,0,71,0,132,0,117,0,245,0,206,0,0,0,0,0,0,0,206,0,0,0,0,0,96,0,178,0,0,0,70,0,136,0);
signal scenario_full  : scenario_type := (124,31,61,31,173,31,155,31,91,31,213,31,50,31,181,31,33,31,211,31,178,31,178,30,142,31,121,31,121,30,97,31,217,31,217,30,102,31,192,31,192,30,151,31,226,31,239,31,8,31,249,31,249,30,196,31,240,31,53,31,53,30,89,31,231,31,252,31,33,31,33,30,33,29,131,31,93,31,169,31,169,30,244,31,244,30,251,31,9,31,128,31,92,31,59,31,155,31,234,31,213,31,56,31,8,31,123,31,146,31,220,31,55,31,211,31,230,31,3,31,134,31,134,30,199,31,21,31,4,31,4,30,4,29,149,31,63,31,63,30,238,31,63,31,107,31,183,31,79,31,25,31,221,31,23,31,23,30,55,31,192,31,178,31,178,30,216,31,90,31,166,31,166,30,155,31,134,31,15,31,119,31,76,31,121,31,132,31,114,31,244,31,180,31,229,31,177,31,37,31,230,31,73,31,75,31,173,31,123,31,243,31,166,31,245,31,245,30,13,31,231,31,106,31,67,31,141,31,142,31,62,31,193,31,36,31,192,31,170,31,240,31,25,31,203,31,40,31,74,31,59,31,14,31,173,31,134,31,38,31,179,31,246,31,164,31,164,30,177,31,70,31,38,31,96,31,87,31,148,31,13,31,231,31,137,31,137,30,17,31,17,30,214,31,113,31,113,30,197,31,236,31,117,31,107,31,226,31,78,31,232,31,39,31,126,31,72,31,158,31,240,31,184,31,184,30,186,31,186,30,191,31,160,31,203,31,11,31,190,31,237,31,208,31,208,30,125,31,254,31,221,31,73,31,118,31,194,31,155,31,248,31,130,31,36,31,150,31,129,31,152,31,73,31,85,31,62,31,62,30,14,31,23,31,23,30,23,29,23,28,173,31,97,31,97,30,67,31,181,31,59,31,23,31,34,31,72,31,114,31,88,31,2,31,11,31,68,31,33,31,16,31,153,31,77,31,115,31,115,30,211,31,82,31,189,31,186,31,205,31,205,30,248,31,161,31,38,31,41,31,156,31,48,31,25,31,251,31,70,31,124,31,236,31,17,31,254,31,125,31,111,31,111,30,144,31,112,31,242,31,228,31,120,31,122,31,230,31,23,31,119,31,196,31,163,31,250,31,89,31,89,30,102,31,32,31,161,31,161,30,7,31,11,31,100,31,91,31,148,31,224,31,224,30,163,31,25,31,25,30,25,29,216,31,179,31,247,31,247,30,136,31,136,30,136,29,231,31,125,31,125,30,175,31,175,30,212,31,91,31,67,31,115,31,211,31,197,31,128,31,156,31,156,30,247,31,45,31,156,31,156,30,24,31,155,31,90,31,33,31,247,31,247,30,247,29,229,31,229,30,229,29,181,31,145,31,154,31,61,31,61,30,228,31,103,31,165,31,223,31,1,31,62,31,246,31,52,31,252,31,245,31,175,31,104,31,67,31,215,31,183,31,132,31,16,31,16,30,219,31,68,31,122,31,122,30,122,29,122,28,34,31,34,30,34,29,119,31,68,31,122,31,223,31,198,31,198,30,29,31,29,30,46,31,54,31,149,31,149,30,43,31,43,30,80,31,113,31,149,31,221,31,218,31,218,30,238,31,240,31,160,31,89,31,118,31,118,30,118,31,40,31,109,31,32,31,32,30,9,31,107,31,97,31,111,31,244,31,224,31,200,31,193,31,250,31,59,31,22,31,5,31,37,31,37,30,37,31,114,31,123,31,131,31,65,31,216,31,126,31,89,31,126,31,232,31,86,31,212,31,69,31,131,31,148,31,135,31,194,31,194,30,28,31,28,30,146,31,93,31,172,31,197,31,115,31,115,30,194,31,216,31,71,31,248,31,98,31,65,31,65,30,189,31,237,31,237,30,117,31,117,31,117,30,235,31,194,31,194,30,152,31,44,31,65,31,106,31,243,31,247,31,10,31,85,31,238,31,205,31,87,31,155,31,204,31,216,31,102,31,203,31,215,31,110,31,110,30,161,31,41,31,83,31,42,31,42,30,105,31,35,31,204,31,34,31,104,31,10,31,65,31,166,31,200,31,49,31,49,30,200,31,200,30,113,31,193,31,224,31,223,31,127,31,145,31,16,31,240,31,244,31,118,31,183,31,82,31,82,30,6,31,225,31,214,31,28,31,28,30,134,31,134,30,178,31,214,31,9,31,233,31,117,31,215,31,114,31,97,31,7,31,210,31,54,31,157,31,153,31,252,31,252,30,128,31,205,31,205,30,242,31,92,31,103,31,103,30,182,31,121,31,137,31,137,30,137,29,8,31,57,31,86,31,86,30,13,31,193,31,59,31,227,31,222,31,3,31,132,31,132,30,44,31,18,31,18,30,18,29,65,31,193,31,32,31,125,31,173,31,173,30,62,31,158,31,107,31,77,31,77,30,239,31,120,31,223,31,184,31,222,31,45,31,18,31,109,31,77,31,79,31,220,31,228,31,98,31,98,30,57,31,220,31,99,31,187,31,5,31,5,30,23,31,23,30,185,31,185,30,185,29,94,31,222,31,110,31,110,30,164,31,11,31,206,31,206,30,31,31,42,31,160,31,91,31,91,30,128,31,161,31,148,31,121,31,59,31,42,31,163,31,163,30,254,31,254,30,20,31,97,31,242,31,205,31,49,31,49,30,228,31,120,31,90,31,90,30,17,31,97,31,111,31,245,31,198,31,71,31,132,31,117,31,245,31,206,31,206,30,206,29,206,28,206,31,206,30,206,29,96,31,178,31,178,30,70,31,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
