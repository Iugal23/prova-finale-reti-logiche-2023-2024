-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 877;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (19,0,0,0,3,0,53,0,65,0,74,0,251,0,61,0,7,0,176,0,0,0,255,0,0,0,65,0,0,0,234,0,107,0,59,0,158,0,88,0,0,0,47,0,0,0,145,0,6,0,0,0,44,0,135,0,211,0,116,0,61,0,148,0,209,0,183,0,71,0,9,0,0,0,176,0,7,0,0,0,47,0,2,0,153,0,215,0,0,0,179,0,194,0,226,0,121,0,147,0,0,0,229,0,245,0,195,0,7,0,6,0,198,0,0,0,212,0,121,0,0,0,0,0,138,0,97,0,0,0,0,0,0,0,23,0,198,0,0,0,0,0,0,0,93,0,0,0,157,0,0,0,140,0,166,0,234,0,0,0,66,0,90,0,195,0,103,0,1,0,216,0,23,0,249,0,43,0,128,0,68,0,37,0,58,0,157,0,98,0,71,0,0,0,3,0,125,0,223,0,186,0,188,0,0,0,135,0,124,0,225,0,0,0,143,0,227,0,179,0,252,0,218,0,39,0,0,0,41,0,141,0,0,0,179,0,241,0,0,0,143,0,0,0,107,0,37,0,0,0,0,0,142,0,0,0,23,0,0,0,112,0,0,0,0,0,0,0,0,0,210,0,64,0,8,0,249,0,41,0,27,0,76,0,111,0,56,0,208,0,18,0,110,0,69,0,27,0,228,0,22,0,3,0,237,0,0,0,0,0,221,0,44,0,0,0,90,0,147,0,94,0,4,0,0,0,0,0,0,0,149,0,32,0,255,0,110,0,88,0,246,0,128,0,3,0,193,0,249,0,18,0,106,0,0,0,36,0,243,0,13,0,140,0,0,0,61,0,238,0,77,0,18,0,0,0,43,0,0,0,158,0,107,0,198,0,73,0,218,0,0,0,138,0,161,0,57,0,82,0,0,0,93,0,123,0,117,0,183,0,249,0,80,0,3,0,0,0,175,0,103,0,13,0,134,0,0,0,0,0,61,0,0,0,0,0,194,0,149,0,252,0,32,0,0,0,0,0,7,0,76,0,102,0,202,0,0,0,116,0,140,0,0,0,246,0,56,0,27,0,0,0,32,0,47,0,218,0,143,0,160,0,0,0,1,0,27,0,66,0,182,0,47,0,53,0,92,0,0,0,0,0,0,0,102,0,220,0,191,0,248,0,240,0,225,0,31,0,238,0,251,0,0,0,21,0,222,0,225,0,153,0,49,0,155,0,0,0,23,0,165,0,20,0,209,0,74,0,0,0,104,0,0,0,112,0,214,0,0,0,191,0,0,0,66,0,60,0,172,0,199,0,80,0,119,0,92,0,202,0,3,0,47,0,192,0,172,0,146,0,212,0,128,0,65,0,209,0,159,0,174,0,202,0,20,0,165,0,104,0,19,0,95,0,132,0,163,0,163,0,0,0,226,0,86,0,29,0,114,0,139,0,202,0,0,0,178,0,56,0,197,0,0,0,15,0,141,0,96,0,160,0,29,0,0,0,227,0,0,0,0,0,125,0,175,0,69,0,0,0,0,0,81,0,0,0,206,0,122,0,0,0,211,0,155,0,6,0,50,0,237,0,47,0,0,0,112,0,173,0,88,0,106,0,73,0,0,0,19,0,234,0,0,0,235,0,8,0,59,0,0,0,254,0,176,0,110,0,0,0,187,0,208,0,233,0,0,0,111,0,38,0,126,0,229,0,148,0,0,0,154,0,0,0,52,0,82,0,0,0,46,0,118,0,166,0,84,0,214,0,70,0,167,0,156,0,0,0,131,0,107,0,144,0,19,0,131,0,174,0,0,0,15,0,0,0,33,0,217,0,0,0,53,0,65,0,66,0,50,0,0,0,177,0,120,0,77,0,152,0,0,0,112,0,167,0,185,0,84,0,98,0,242,0,85,0,149,0,246,0,55,0,217,0,173,0,1,0,202,0,0,0,102,0,9,0,209,0,150,0,25,0,14,0,135,0,0,0,51,0,18,0,239,0,130,0,13,0,24,0,28,0,76,0,0,0,168,0,249,0,143,0,218,0,215,0,124,0,0,0,82,0,4,0,0,0,0,0,78,0,20,0,201,0,54,0,56,0,14,0,166,0,164,0,138,0,17,0,13,0,103,0,249,0,239,0,0,0,16,0,0,0,63,0,227,0,121,0,26,0,77,0,150,0,248,0,200,0,195,0,0,0,0,0,243,0,160,0,154,0,151,0,152,0,18,0,101,0,79,0,0,0,60,0,230,0,104,0,124,0,0,0,109,0,220,0,49,0,251,0,42,0,160,0,32,0,221,0,91,0,135,0,40,0,117,0,50,0,40,0,58,0,154,0,66,0,101,0,0,0,108,0,60,0,0,0,211,0,13,0,2,0,14,0,61,0,175,0,8,0,0,0,0,0,147,0,90,0,207,0,100,0,78,0,251,0,184,0,146,0,63,0,33,0,15,0,0,0,119,0,132,0,0,0,9,0,211,0,179,0,0,0,223,0,175,0,0,0,208,0,15,0,120,0,49,0,48,0,0,0,82,0,232,0,0,0,0,0,51,0,162,0,231,0,39,0,1,0,126,0,0,0,0,0,42,0,0,0,35,0,31,0,51,0,120,0,147,0,90,0,57,0,146,0,31,0,152,0,0,0,0,0,99,0,125,0,116,0,188,0,0,0,143,0,244,0,0,0,150,0,186,0,0,0,134,0,246,0,181,0,0,0,141,0,0,0,172,0,148,0,78,0,54,0,223,0,41,0,160,0,24,0,135,0,0,0,26,0,48,0,240,0,42,0,142,0,40,0,129,0,235,0,52,0,158,0,181,0,134,0,0,0,18,0,0,0,81,0,181,0,74,0,151,0,0,0,113,0,148,0,245,0,111,0,145,0,0,0,131,0,2,0,116,0,179,0,140,0,0,0,242,0,0,0,0,0,10,0,98,0,149,0,0,0,245,0,169,0,173,0,18,0,225,0,5,0,208,0,0,0,6,0,0,0,0,0,50,0,0,0,0,0,156,0,70,0,120,0,0,0,163,0,162,0,0,0,0,0,41,0,113,0,156,0,160,0,85,0,253,0,235,0,75,0,116,0,51,0,38,0,191,0,109,0,116,0,5,0,95,0,100,0,244,0,130,0,236,0,128,0,182,0,33,0,161,0,0,0,76,0,0,0,137,0,73,0,174,0,105,0,0,0,116,0,83,0,157,0,50,0,120,0,74,0,165,0,20,0,151,0,29,0,180,0,110,0,88,0,208,0,193,0,0,0,0,0,114,0,159,0,53,0,61,0,0,0,58,0,0,0,205,0,21,0,139,0,39,0,64,0,41,0,93,0,206,0,247,0,101,0,32,0,236,0,223,0,157,0,0,0,0,0,0,0,0,0,175,0,0,0,121,0,17,0,47,0,232,0,63,0,20,0,0,0,0,0,0,0,98,0,100,0,28,0,0,0,58,0,0,0,229,0,117,0,0,0,130,0,0,0,0,0,76,0,70,0,74,0,95,0,244,0,80,0,203,0,183,0,0,0,153,0,25,0,190,0,51,0,0,0,232,0,217,0,239,0,183,0,123,0,0,0,234,0,225,0,188,0,0,0,186,0,93,0,0,0,122,0,5,0,74,0,94,0,244,0,136,0,62,0,0,0,202,0,239,0,134,0,142,0,0,0,92,0,20,0,229,0,51,0,102,0,245,0,0,0,122,0,0,0,210,0,210,0,228,0,209,0,28,0,18,0,135,0,214,0,0,0,173,0,108,0,31,0,205,0,94,0,113,0,2,0,0,0,19,0,79,0,112,0,0,0,72,0,229,0,191,0,0,0,0,0,93,0,247,0,0,0,0,0,251,0,0,0,0,0,246,0,227,0,141,0,252,0,69,0,198,0,231,0,96,0,215,0,51,0,83,0,124,0,13,0,104,0,251,0,0,0,0,0,0,0,248,0,53,0,43,0,3,0,92,0,25,0,95,0,70,0,86,0,0,0,0,0);
signal scenario_full  : scenario_type := (19,31,19,30,3,31,53,31,65,31,74,31,251,31,61,31,7,31,176,31,176,30,255,31,255,30,65,31,65,30,234,31,107,31,59,31,158,31,88,31,88,30,47,31,47,30,145,31,6,31,6,30,44,31,135,31,211,31,116,31,61,31,148,31,209,31,183,31,71,31,9,31,9,30,176,31,7,31,7,30,47,31,2,31,153,31,215,31,215,30,179,31,194,31,226,31,121,31,147,31,147,30,229,31,245,31,195,31,7,31,6,31,198,31,198,30,212,31,121,31,121,30,121,29,138,31,97,31,97,30,97,29,97,28,23,31,198,31,198,30,198,29,198,28,93,31,93,30,157,31,157,30,140,31,166,31,234,31,234,30,66,31,90,31,195,31,103,31,1,31,216,31,23,31,249,31,43,31,128,31,68,31,37,31,58,31,157,31,98,31,71,31,71,30,3,31,125,31,223,31,186,31,188,31,188,30,135,31,124,31,225,31,225,30,143,31,227,31,179,31,252,31,218,31,39,31,39,30,41,31,141,31,141,30,179,31,241,31,241,30,143,31,143,30,107,31,37,31,37,30,37,29,142,31,142,30,23,31,23,30,112,31,112,30,112,29,112,28,112,27,210,31,64,31,8,31,249,31,41,31,27,31,76,31,111,31,56,31,208,31,18,31,110,31,69,31,27,31,228,31,22,31,3,31,237,31,237,30,237,29,221,31,44,31,44,30,90,31,147,31,94,31,4,31,4,30,4,29,4,28,149,31,32,31,255,31,110,31,88,31,246,31,128,31,3,31,193,31,249,31,18,31,106,31,106,30,36,31,243,31,13,31,140,31,140,30,61,31,238,31,77,31,18,31,18,30,43,31,43,30,158,31,107,31,198,31,73,31,218,31,218,30,138,31,161,31,57,31,82,31,82,30,93,31,123,31,117,31,183,31,249,31,80,31,3,31,3,30,175,31,103,31,13,31,134,31,134,30,134,29,61,31,61,30,61,29,194,31,149,31,252,31,32,31,32,30,32,29,7,31,76,31,102,31,202,31,202,30,116,31,140,31,140,30,246,31,56,31,27,31,27,30,32,31,47,31,218,31,143,31,160,31,160,30,1,31,27,31,66,31,182,31,47,31,53,31,92,31,92,30,92,29,92,28,102,31,220,31,191,31,248,31,240,31,225,31,31,31,238,31,251,31,251,30,21,31,222,31,225,31,153,31,49,31,155,31,155,30,23,31,165,31,20,31,209,31,74,31,74,30,104,31,104,30,112,31,214,31,214,30,191,31,191,30,66,31,60,31,172,31,199,31,80,31,119,31,92,31,202,31,3,31,47,31,192,31,172,31,146,31,212,31,128,31,65,31,209,31,159,31,174,31,202,31,20,31,165,31,104,31,19,31,95,31,132,31,163,31,163,31,163,30,226,31,86,31,29,31,114,31,139,31,202,31,202,30,178,31,56,31,197,31,197,30,15,31,141,31,96,31,160,31,29,31,29,30,227,31,227,30,227,29,125,31,175,31,69,31,69,30,69,29,81,31,81,30,206,31,122,31,122,30,211,31,155,31,6,31,50,31,237,31,47,31,47,30,112,31,173,31,88,31,106,31,73,31,73,30,19,31,234,31,234,30,235,31,8,31,59,31,59,30,254,31,176,31,110,31,110,30,187,31,208,31,233,31,233,30,111,31,38,31,126,31,229,31,148,31,148,30,154,31,154,30,52,31,82,31,82,30,46,31,118,31,166,31,84,31,214,31,70,31,167,31,156,31,156,30,131,31,107,31,144,31,19,31,131,31,174,31,174,30,15,31,15,30,33,31,217,31,217,30,53,31,65,31,66,31,50,31,50,30,177,31,120,31,77,31,152,31,152,30,112,31,167,31,185,31,84,31,98,31,242,31,85,31,149,31,246,31,55,31,217,31,173,31,1,31,202,31,202,30,102,31,9,31,209,31,150,31,25,31,14,31,135,31,135,30,51,31,18,31,239,31,130,31,13,31,24,31,28,31,76,31,76,30,168,31,249,31,143,31,218,31,215,31,124,31,124,30,82,31,4,31,4,30,4,29,78,31,20,31,201,31,54,31,56,31,14,31,166,31,164,31,138,31,17,31,13,31,103,31,249,31,239,31,239,30,16,31,16,30,63,31,227,31,121,31,26,31,77,31,150,31,248,31,200,31,195,31,195,30,195,29,243,31,160,31,154,31,151,31,152,31,18,31,101,31,79,31,79,30,60,31,230,31,104,31,124,31,124,30,109,31,220,31,49,31,251,31,42,31,160,31,32,31,221,31,91,31,135,31,40,31,117,31,50,31,40,31,58,31,154,31,66,31,101,31,101,30,108,31,60,31,60,30,211,31,13,31,2,31,14,31,61,31,175,31,8,31,8,30,8,29,147,31,90,31,207,31,100,31,78,31,251,31,184,31,146,31,63,31,33,31,15,31,15,30,119,31,132,31,132,30,9,31,211,31,179,31,179,30,223,31,175,31,175,30,208,31,15,31,120,31,49,31,48,31,48,30,82,31,232,31,232,30,232,29,51,31,162,31,231,31,39,31,1,31,126,31,126,30,126,29,42,31,42,30,35,31,31,31,51,31,120,31,147,31,90,31,57,31,146,31,31,31,152,31,152,30,152,29,99,31,125,31,116,31,188,31,188,30,143,31,244,31,244,30,150,31,186,31,186,30,134,31,246,31,181,31,181,30,141,31,141,30,172,31,148,31,78,31,54,31,223,31,41,31,160,31,24,31,135,31,135,30,26,31,48,31,240,31,42,31,142,31,40,31,129,31,235,31,52,31,158,31,181,31,134,31,134,30,18,31,18,30,81,31,181,31,74,31,151,31,151,30,113,31,148,31,245,31,111,31,145,31,145,30,131,31,2,31,116,31,179,31,140,31,140,30,242,31,242,30,242,29,10,31,98,31,149,31,149,30,245,31,169,31,173,31,18,31,225,31,5,31,208,31,208,30,6,31,6,30,6,29,50,31,50,30,50,29,156,31,70,31,120,31,120,30,163,31,162,31,162,30,162,29,41,31,113,31,156,31,160,31,85,31,253,31,235,31,75,31,116,31,51,31,38,31,191,31,109,31,116,31,5,31,95,31,100,31,244,31,130,31,236,31,128,31,182,31,33,31,161,31,161,30,76,31,76,30,137,31,73,31,174,31,105,31,105,30,116,31,83,31,157,31,50,31,120,31,74,31,165,31,20,31,151,31,29,31,180,31,110,31,88,31,208,31,193,31,193,30,193,29,114,31,159,31,53,31,61,31,61,30,58,31,58,30,205,31,21,31,139,31,39,31,64,31,41,31,93,31,206,31,247,31,101,31,32,31,236,31,223,31,157,31,157,30,157,29,157,28,157,27,175,31,175,30,121,31,17,31,47,31,232,31,63,31,20,31,20,30,20,29,20,28,98,31,100,31,28,31,28,30,58,31,58,30,229,31,117,31,117,30,130,31,130,30,130,29,76,31,70,31,74,31,95,31,244,31,80,31,203,31,183,31,183,30,153,31,25,31,190,31,51,31,51,30,232,31,217,31,239,31,183,31,123,31,123,30,234,31,225,31,188,31,188,30,186,31,93,31,93,30,122,31,5,31,74,31,94,31,244,31,136,31,62,31,62,30,202,31,239,31,134,31,142,31,142,30,92,31,20,31,229,31,51,31,102,31,245,31,245,30,122,31,122,30,210,31,210,31,228,31,209,31,28,31,18,31,135,31,214,31,214,30,173,31,108,31,31,31,205,31,94,31,113,31,2,31,2,30,19,31,79,31,112,31,112,30,72,31,229,31,191,31,191,30,191,29,93,31,247,31,247,30,247,29,251,31,251,30,251,29,246,31,227,31,141,31,252,31,69,31,198,31,231,31,96,31,215,31,51,31,83,31,124,31,13,31,104,31,251,31,251,30,251,29,251,28,248,31,53,31,43,31,3,31,92,31,25,31,95,31,70,31,86,31,86,30,86,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
