-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 883;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,24,0,0,0,69,0,139,0,133,0,133,0,70,0,226,0,224,0,55,0,0,0,243,0,189,0,16,0,0,0,182,0,0,0,139,0,2,0,0,0,180,0,1,0,200,0,146,0,131,0,0,0,14,0,0,0,0,0,0,0,0,0,78,0,165,0,22,0,0,0,3,0,34,0,87,0,98,0,248,0,245,0,143,0,223,0,183,0,176,0,93,0,193,0,105,0,180,0,105,0,209,0,0,0,216,0,111,0,138,0,79,0,205,0,12,0,0,0,95,0,0,0,126,0,85,0,70,0,75,0,188,0,14,0,213,0,0,0,0,0,123,0,93,0,241,0,0,0,192,0,125,0,0,0,100,0,99,0,3,0,240,0,0,0,182,0,208,0,213,0,218,0,0,0,235,0,252,0,72,0,175,0,71,0,27,0,12,0,198,0,0,0,135,0,193,0,213,0,15,0,8,0,190,0,17,0,90,0,0,0,55,0,162,0,0,0,117,0,242,0,130,0,129,0,215,0,230,0,240,0,17,0,195,0,43,0,137,0,254,0,81,0,112,0,198,0,84,0,0,0,79,0,246,0,201,0,0,0,29,0,47,0,249,0,46,0,68,0,6,0,53,0,221,0,121,0,207,0,122,0,156,0,23,0,56,0,40,0,224,0,67,0,7,0,195,0,243,0,6,0,0,0,8,0,45,0,203,0,210,0,252,0,95,0,0,0,0,0,0,0,47,0,242,0,123,0,9,0,26,0,163,0,254,0,0,0,81,0,113,0,209,0,243,0,42,0,176,0,134,0,242,0,241,0,0,0,71,0,111,0,96,0,9,0,0,0,214,0,249,0,200,0,104,0,86,0,121,0,106,0,220,0,122,0,76,0,162,0,211,0,241,0,136,0,0,0,163,0,140,0,227,0,222,0,0,0,23,0,86,0,74,0,249,0,40,0,148,0,38,0,210,0,188,0,26,0,109,0,0,0,83,0,42,0,146,0,133,0,48,0,0,0,239,0,0,0,119,0,6,0,126,0,208,0,3,0,0,0,205,0,194,0,0,0,45,0,119,0,107,0,201,0,79,0,39,0,0,0,185,0,61,0,93,0,0,0,133,0,254,0,80,0,12,0,243,0,18,0,38,0,214,0,172,0,0,0,32,0,0,0,233,0,0,0,133,0,103,0,0,0,134,0,0,0,110,0,53,0,92,0,20,0,0,0,0,0,22,0,89,0,20,0,0,0,228,0,122,0,238,0,212,0,23,0,184,0,214,0,136,0,99,0,80,0,238,0,209,0,160,0,238,0,45,0,169,0,0,0,210,0,123,0,0,0,219,0,64,0,23,0,101,0,237,0,240,0,213,0,55,0,117,0,181,0,0,0,240,0,33,0,0,0,45,0,49,0,46,0,0,0,80,0,115,0,78,0,159,0,94,0,49,0,243,0,191,0,202,0,0,0,33,0,0,0,64,0,227,0,0,0,135,0,211,0,125,0,41,0,173,0,53,0,241,0,0,0,0,0,11,0,0,0,0,0,14,0,84,0,0,0,0,0,109,0,0,0,37,0,204,0,130,0,120,0,0,0,126,0,0,0,232,0,158,0,140,0,202,0,184,0,51,0,174,0,0,0,134,0,162,0,0,0,0,0,191,0,196,0,216,0,223,0,100,0,168,0,62,0,123,0,162,0,156,0,155,0,107,0,142,0,89,0,0,0,120,0,42,0,44,0,239,0,201,0,0,0,0,0,0,0,141,0,0,0,217,0,83,0,50,0,0,0,0,0,182,0,207,0,50,0,0,0,214,0,246,0,0,0,174,0,125,0,87,0,122,0,11,0,226,0,147,0,10,0,91,0,106,0,169,0,0,0,21,0,30,0,85,0,43,0,5,0,52,0,173,0,49,0,59,0,106,0,0,0,40,0,212,0,255,0,13,0,0,0,245,0,0,0,176,0,143,0,219,0,91,0,165,0,121,0,70,0,0,0,70,0,0,0,242,0,160,0,135,0,236,0,239,0,140,0,155,0,0,0,130,0,76,0,176,0,0,0,254,0,0,0,118,0,0,0,0,0,246,0,156,0,212,0,2,0,171,0,103,0,123,0,251,0,61,0,203,0,146,0,0,0,14,0,0,0,204,0,115,0,129,0,58,0,0,0,34,0,55,0,114,0,0,0,83,0,0,0,0,0,194,0,248,0,60,0,54,0,227,0,253,0,0,0,64,0,114,0,6,0,0,0,37,0,0,0,240,0,13,0,119,0,70,0,99,0,76,0,38,0,103,0,237,0,177,0,46,0,133,0,242,0,0,0,135,0,157,0,155,0,29,0,107,0,160,0,201,0,136,0,190,0,25,0,0,0,130,0,0,0,223,0,132,0,147,0,212,0,11,0,240,0,31,0,174,0,73,0,182,0,114,0,214,0,189,0,222,0,0,0,147,0,95,0,214,0,8,0,151,0,163,0,19,0,69,0,179,0,0,0,131,0,0,0,58,0,156,0,68,0,0,0,165,0,54,0,161,0,216,0,182,0,105,0,84,0,38,0,149,0,245,0,23,0,98,0,56,0,240,0,245,0,232,0,0,0,0,0,0,0,0,0,242,0,0,0,125,0,28,0,123,0,98,0,215,0,0,0,0,0,0,0,117,0,0,0,172,0,127,0,1,0,0,0,189,0,50,0,85,0,134,0,251,0,234,0,0,0,53,0,78,0,72,0,207,0,61,0,5,0,134,0,14,0,0,0,0,0,0,0,61,0,196,0,120,0,15,0,49,0,192,0,57,0,249,0,46,0,25,0,214,0,183,0,0,0,0,0,0,0,150,0,0,0,62,0,128,0,199,0,51,0,205,0,0,0,61,0,0,0,153,0,0,0,113,0,63,0,0,0,135,0,194,0,86,0,44,0,147,0,79,0,232,0,179,0,49,0,96,0,133,0,56,0,110,0,178,0,170,0,130,0,250,0,18,0,0,0,54,0,140,0,126,0,130,0,176,0,241,0,41,0,178,0,29,0,167,0,122,0,37,0,150,0,113,0,1,0,44,0,117,0,88,0,0,0,221,0,200,0,0,0,80,0,196,0,134,0,119,0,33,0,32,0,5,0,72,0,140,0,119,0,209,0,104,0,223,0,134,0,152,0,3,0,253,0,0,0,133,0,20,0,227,0,0,0,241,0,0,0,0,0,0,0,21,0,137,0,147,0,151,0,75,0,26,0,55,0,168,0,198,0,184,0,0,0,97,0,126,0,106,0,53,0,0,0,0,0,131,0,238,0,12,0,172,0,95,0,31,0,25,0,112,0,0,0,0,0,15,0,33,0,135,0,227,0,135,0,117,0,163,0,129,0,0,0,232,0,0,0,16,0,94,0,78,0,153,0,174,0,60,0,0,0,143,0,98,0,10,0,35,0,0,0,245,0,0,0,148,0,59,0,216,0,0,0,155,0,10,0,46,0,76,0,158,0,0,0,135,0,0,0,184,0,0,0,231,0,218,0,0,0,24,0,182,0,41,0,161,0,174,0,180,0,73,0,156,0,19,0,210,0,190,0,40,0,146,0,158,0,66,0,0,0,0,0,6,0,42,0,203,0,0,0,56,0,154,0,23,0,154,0,98,0,29,0,231,0,0,0,167,0,172,0,36,0,200,0,237,0,156,0,216,0,0,0,0,0,185,0,88,0,0,0,142,0,243,0,36,0,138,0,229,0,42,0,0,0,2,0,11,0,231,0,251,0,67,0,220,0,39,0,132,0,87,0,0,0,135,0,30,0,22,0,80,0,55,0,149,0,143,0,0,0,0,0,141,0,197,0,251,0,186,0,150,0,113,0,88,0,229,0,117,0,0,0,174,0,0,0,0,0,0,0,0,0,33,0,61,0,0,0,113,0,225,0,214,0,247,0,104,0,0,0,198,0,0,0,84,0,199,0,129,0,9,0,76,0,142,0,0,0,135,0,0,0,0,0,42,0,0,0,51,0,139,0,0,0,213,0);
signal scenario_full  : scenario_type := (0,0,24,31,24,30,69,31,139,31,133,31,133,31,70,31,226,31,224,31,55,31,55,30,243,31,189,31,16,31,16,30,182,31,182,30,139,31,2,31,2,30,180,31,1,31,200,31,146,31,131,31,131,30,14,31,14,30,14,29,14,28,14,27,78,31,165,31,22,31,22,30,3,31,34,31,87,31,98,31,248,31,245,31,143,31,223,31,183,31,176,31,93,31,193,31,105,31,180,31,105,31,209,31,209,30,216,31,111,31,138,31,79,31,205,31,12,31,12,30,95,31,95,30,126,31,85,31,70,31,75,31,188,31,14,31,213,31,213,30,213,29,123,31,93,31,241,31,241,30,192,31,125,31,125,30,100,31,99,31,3,31,240,31,240,30,182,31,208,31,213,31,218,31,218,30,235,31,252,31,72,31,175,31,71,31,27,31,12,31,198,31,198,30,135,31,193,31,213,31,15,31,8,31,190,31,17,31,90,31,90,30,55,31,162,31,162,30,117,31,242,31,130,31,129,31,215,31,230,31,240,31,17,31,195,31,43,31,137,31,254,31,81,31,112,31,198,31,84,31,84,30,79,31,246,31,201,31,201,30,29,31,47,31,249,31,46,31,68,31,6,31,53,31,221,31,121,31,207,31,122,31,156,31,23,31,56,31,40,31,224,31,67,31,7,31,195,31,243,31,6,31,6,30,8,31,45,31,203,31,210,31,252,31,95,31,95,30,95,29,95,28,47,31,242,31,123,31,9,31,26,31,163,31,254,31,254,30,81,31,113,31,209,31,243,31,42,31,176,31,134,31,242,31,241,31,241,30,71,31,111,31,96,31,9,31,9,30,214,31,249,31,200,31,104,31,86,31,121,31,106,31,220,31,122,31,76,31,162,31,211,31,241,31,136,31,136,30,163,31,140,31,227,31,222,31,222,30,23,31,86,31,74,31,249,31,40,31,148,31,38,31,210,31,188,31,26,31,109,31,109,30,83,31,42,31,146,31,133,31,48,31,48,30,239,31,239,30,119,31,6,31,126,31,208,31,3,31,3,30,205,31,194,31,194,30,45,31,119,31,107,31,201,31,79,31,39,31,39,30,185,31,61,31,93,31,93,30,133,31,254,31,80,31,12,31,243,31,18,31,38,31,214,31,172,31,172,30,32,31,32,30,233,31,233,30,133,31,103,31,103,30,134,31,134,30,110,31,53,31,92,31,20,31,20,30,20,29,22,31,89,31,20,31,20,30,228,31,122,31,238,31,212,31,23,31,184,31,214,31,136,31,99,31,80,31,238,31,209,31,160,31,238,31,45,31,169,31,169,30,210,31,123,31,123,30,219,31,64,31,23,31,101,31,237,31,240,31,213,31,55,31,117,31,181,31,181,30,240,31,33,31,33,30,45,31,49,31,46,31,46,30,80,31,115,31,78,31,159,31,94,31,49,31,243,31,191,31,202,31,202,30,33,31,33,30,64,31,227,31,227,30,135,31,211,31,125,31,41,31,173,31,53,31,241,31,241,30,241,29,11,31,11,30,11,29,14,31,84,31,84,30,84,29,109,31,109,30,37,31,204,31,130,31,120,31,120,30,126,31,126,30,232,31,158,31,140,31,202,31,184,31,51,31,174,31,174,30,134,31,162,31,162,30,162,29,191,31,196,31,216,31,223,31,100,31,168,31,62,31,123,31,162,31,156,31,155,31,107,31,142,31,89,31,89,30,120,31,42,31,44,31,239,31,201,31,201,30,201,29,201,28,141,31,141,30,217,31,83,31,50,31,50,30,50,29,182,31,207,31,50,31,50,30,214,31,246,31,246,30,174,31,125,31,87,31,122,31,11,31,226,31,147,31,10,31,91,31,106,31,169,31,169,30,21,31,30,31,85,31,43,31,5,31,52,31,173,31,49,31,59,31,106,31,106,30,40,31,212,31,255,31,13,31,13,30,245,31,245,30,176,31,143,31,219,31,91,31,165,31,121,31,70,31,70,30,70,31,70,30,242,31,160,31,135,31,236,31,239,31,140,31,155,31,155,30,130,31,76,31,176,31,176,30,254,31,254,30,118,31,118,30,118,29,246,31,156,31,212,31,2,31,171,31,103,31,123,31,251,31,61,31,203,31,146,31,146,30,14,31,14,30,204,31,115,31,129,31,58,31,58,30,34,31,55,31,114,31,114,30,83,31,83,30,83,29,194,31,248,31,60,31,54,31,227,31,253,31,253,30,64,31,114,31,6,31,6,30,37,31,37,30,240,31,13,31,119,31,70,31,99,31,76,31,38,31,103,31,237,31,177,31,46,31,133,31,242,31,242,30,135,31,157,31,155,31,29,31,107,31,160,31,201,31,136,31,190,31,25,31,25,30,130,31,130,30,223,31,132,31,147,31,212,31,11,31,240,31,31,31,174,31,73,31,182,31,114,31,214,31,189,31,222,31,222,30,147,31,95,31,214,31,8,31,151,31,163,31,19,31,69,31,179,31,179,30,131,31,131,30,58,31,156,31,68,31,68,30,165,31,54,31,161,31,216,31,182,31,105,31,84,31,38,31,149,31,245,31,23,31,98,31,56,31,240,31,245,31,232,31,232,30,232,29,232,28,232,27,242,31,242,30,125,31,28,31,123,31,98,31,215,31,215,30,215,29,215,28,117,31,117,30,172,31,127,31,1,31,1,30,189,31,50,31,85,31,134,31,251,31,234,31,234,30,53,31,78,31,72,31,207,31,61,31,5,31,134,31,14,31,14,30,14,29,14,28,61,31,196,31,120,31,15,31,49,31,192,31,57,31,249,31,46,31,25,31,214,31,183,31,183,30,183,29,183,28,150,31,150,30,62,31,128,31,199,31,51,31,205,31,205,30,61,31,61,30,153,31,153,30,113,31,63,31,63,30,135,31,194,31,86,31,44,31,147,31,79,31,232,31,179,31,49,31,96,31,133,31,56,31,110,31,178,31,170,31,130,31,250,31,18,31,18,30,54,31,140,31,126,31,130,31,176,31,241,31,41,31,178,31,29,31,167,31,122,31,37,31,150,31,113,31,1,31,44,31,117,31,88,31,88,30,221,31,200,31,200,30,80,31,196,31,134,31,119,31,33,31,32,31,5,31,72,31,140,31,119,31,209,31,104,31,223,31,134,31,152,31,3,31,253,31,253,30,133,31,20,31,227,31,227,30,241,31,241,30,241,29,241,28,21,31,137,31,147,31,151,31,75,31,26,31,55,31,168,31,198,31,184,31,184,30,97,31,126,31,106,31,53,31,53,30,53,29,131,31,238,31,12,31,172,31,95,31,31,31,25,31,112,31,112,30,112,29,15,31,33,31,135,31,227,31,135,31,117,31,163,31,129,31,129,30,232,31,232,30,16,31,94,31,78,31,153,31,174,31,60,31,60,30,143,31,98,31,10,31,35,31,35,30,245,31,245,30,148,31,59,31,216,31,216,30,155,31,10,31,46,31,76,31,158,31,158,30,135,31,135,30,184,31,184,30,231,31,218,31,218,30,24,31,182,31,41,31,161,31,174,31,180,31,73,31,156,31,19,31,210,31,190,31,40,31,146,31,158,31,66,31,66,30,66,29,6,31,42,31,203,31,203,30,56,31,154,31,23,31,154,31,98,31,29,31,231,31,231,30,167,31,172,31,36,31,200,31,237,31,156,31,216,31,216,30,216,29,185,31,88,31,88,30,142,31,243,31,36,31,138,31,229,31,42,31,42,30,2,31,11,31,231,31,251,31,67,31,220,31,39,31,132,31,87,31,87,30,135,31,30,31,22,31,80,31,55,31,149,31,143,31,143,30,143,29,141,31,197,31,251,31,186,31,150,31,113,31,88,31,229,31,117,31,117,30,174,31,174,30,174,29,174,28,174,27,33,31,61,31,61,30,113,31,225,31,214,31,247,31,104,31,104,30,198,31,198,30,84,31,199,31,129,31,9,31,76,31,142,31,142,30,135,31,135,30,135,29,42,31,42,30,51,31,139,31,139,30,213,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
