-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_694 is
end project_tb_694;

architecture project_tb_arch_694 of project_tb_694 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 308;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,169,0,0,0,71,0,3,0,163,0,59,0,216,0,0,0,173,0,252,0,107,0,136,0,108,0,150,0,155,0,188,0,68,0,223,0,239,0,44,0,194,0,26,0,171,0,72,0,222,0,165,0,88,0,6,0,162,0,177,0,54,0,28,0,250,0,167,0,72,0,91,0,169,0,138,0,32,0,0,0,168,0,31,0,83,0,169,0,158,0,90,0,118,0,42,0,150,0,22,0,119,0,213,0,76,0,46,0,190,0,79,0,95,0,67,0,142,0,143,0,0,0,111,0,246,0,9,0,34,0,90,0,151,0,0,0,215,0,0,0,63,0,45,0,192,0,0,0,136,0,232,0,0,0,220,0,165,0,197,0,226,0,0,0,144,0,114,0,107,0,36,0,92,0,225,0,0,0,67,0,83,0,0,0,212,0,0,0,2,0,4,0,91,0,8,0,222,0,76,0,167,0,208,0,201,0,196,0,246,0,65,0,129,0,240,0,0,0,56,0,178,0,96,0,104,0,184,0,0,0,158,0,114,0,0,0,58,0,194,0,179,0,125,0,85,0,55,0,2,0,40,0,146,0,29,0,0,0,218,0,0,0,151,0,198,0,141,0,218,0,217,0,108,0,212,0,228,0,3,0,54,0,26,0,103,0,0,0,0,0,124,0,0,0,42,0,0,0,0,0,0,0,0,0,0,0,188,0,247,0,39,0,151,0,165,0,63,0,0,0,93,0,0,0,197,0,16,0,96,0,0,0,109,0,0,0,182,0,70,0,221,0,161,0,0,0,23,0,82,0,89,0,130,0,136,0,233,0,8,0,0,0,0,0,22,0,89,0,0,0,154,0,0,0,79,0,0,0,41,0,209,0,159,0,236,0,169,0,26,0,100,0,0,0,232,0,0,0,96,0,63,0,190,0,0,0,18,0,0,0,127,0,230,0,59,0,1,0,200,0,222,0,144,0,124,0,146,0,104,0,215,0,75,0,226,0,118,0,41,0,11,0,0,0,62,0,9,0,118,0,166,0,89,0,77,0,0,0,0,0,0,0,3,0,0,0,0,0,166,0,233,0,160,0,0,0,112,0,223,0,120,0,136,0,231,0,193,0,1,0,49,0,171,0,0,0,60,0,210,0,46,0,158,0,135,0,106,0,0,0,83,0,181,0,213,0,17,0,0,0,91,0,189,0,89,0,182,0,124,0,167,0,75,0,159,0,12,0,27,0,4,0,216,0,170,0,32,0,182,0,110,0,0,0,122,0,87,0,70,0,154,0,193,0,175,0,211,0,54,0,197,0,187,0,67,0,112,0,132,0,245,0,120,0,0,0,214,0,178,0,196,0,119,0,246,0,163,0,33,0,153,0,47,0,64,0,169,0,249,0,0,0,115,0);
signal scenario_full  : scenario_type := (0,0,169,31,169,30,71,31,3,31,163,31,59,31,216,31,216,30,173,31,252,31,107,31,136,31,108,31,150,31,155,31,188,31,68,31,223,31,239,31,44,31,194,31,26,31,171,31,72,31,222,31,165,31,88,31,6,31,162,31,177,31,54,31,28,31,250,31,167,31,72,31,91,31,169,31,138,31,32,31,32,30,168,31,31,31,83,31,169,31,158,31,90,31,118,31,42,31,150,31,22,31,119,31,213,31,76,31,46,31,190,31,79,31,95,31,67,31,142,31,143,31,143,30,111,31,246,31,9,31,34,31,90,31,151,31,151,30,215,31,215,30,63,31,45,31,192,31,192,30,136,31,232,31,232,30,220,31,165,31,197,31,226,31,226,30,144,31,114,31,107,31,36,31,92,31,225,31,225,30,67,31,83,31,83,30,212,31,212,30,2,31,4,31,91,31,8,31,222,31,76,31,167,31,208,31,201,31,196,31,246,31,65,31,129,31,240,31,240,30,56,31,178,31,96,31,104,31,184,31,184,30,158,31,114,31,114,30,58,31,194,31,179,31,125,31,85,31,55,31,2,31,40,31,146,31,29,31,29,30,218,31,218,30,151,31,198,31,141,31,218,31,217,31,108,31,212,31,228,31,3,31,54,31,26,31,103,31,103,30,103,29,124,31,124,30,42,31,42,30,42,29,42,28,42,27,42,26,188,31,247,31,39,31,151,31,165,31,63,31,63,30,93,31,93,30,197,31,16,31,96,31,96,30,109,31,109,30,182,31,70,31,221,31,161,31,161,30,23,31,82,31,89,31,130,31,136,31,233,31,8,31,8,30,8,29,22,31,89,31,89,30,154,31,154,30,79,31,79,30,41,31,209,31,159,31,236,31,169,31,26,31,100,31,100,30,232,31,232,30,96,31,63,31,190,31,190,30,18,31,18,30,127,31,230,31,59,31,1,31,200,31,222,31,144,31,124,31,146,31,104,31,215,31,75,31,226,31,118,31,41,31,11,31,11,30,62,31,9,31,118,31,166,31,89,31,77,31,77,30,77,29,77,28,3,31,3,30,3,29,166,31,233,31,160,31,160,30,112,31,223,31,120,31,136,31,231,31,193,31,1,31,49,31,171,31,171,30,60,31,210,31,46,31,158,31,135,31,106,31,106,30,83,31,181,31,213,31,17,31,17,30,91,31,189,31,89,31,182,31,124,31,167,31,75,31,159,31,12,31,27,31,4,31,216,31,170,31,32,31,182,31,110,31,110,30,122,31,87,31,70,31,154,31,193,31,175,31,211,31,54,31,197,31,187,31,67,31,112,31,132,31,245,31,120,31,120,30,214,31,178,31,196,31,119,31,246,31,163,31,33,31,153,31,47,31,64,31,169,31,249,31,249,30,115,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
