-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_452 is
end project_tb_452;

architecture project_tb_arch_452 of project_tb_452 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 637;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,0,0,10,0,202,0,41,0,137,0,0,0,31,0,165,0,0,0,73,0,172,0,1,0,64,0,77,0,65,0,243,0,102,0,75,0,3,0,31,0,248,0,97,0,183,0,88,0,236,0,169,0,149,0,0,0,87,0,204,0,0,0,70,0,10,0,0,0,133,0,150,0,161,0,233,0,155,0,0,0,222,0,217,0,155,0,250,0,176,0,84,0,23,0,250,0,166,0,209,0,108,0,18,0,70,0,38,0,81,0,242,0,21,0,0,0,62,0,79,0,169,0,56,0,0,0,51,0,214,0,173,0,126,0,144,0,142,0,14,0,0,0,150,0,0,0,193,0,242,0,177,0,180,0,83,0,0,0,100,0,17,0,0,0,94,0,109,0,1,0,0,0,218,0,228,0,38,0,40,0,18,0,171,0,16,0,47,0,215,0,68,0,35,0,82,0,53,0,31,0,57,0,111,0,131,0,112,0,204,0,0,0,214,0,97,0,130,0,193,0,191,0,0,0,82,0,0,0,86,0,0,0,156,0,0,0,0,0,0,0,195,0,0,0,65,0,0,0,100,0,29,0,0,0,107,0,71,0,0,0,0,0,242,0,202,0,32,0,0,0,148,0,0,0,0,0,0,0,0,0,4,0,167,0,0,0,0,0,190,0,187,0,0,0,95,0,95,0,0,0,0,0,0,0,0,0,170,0,31,0,197,0,6,0,0,0,182,0,0,0,176,0,0,0,27,0,132,0,248,0,27,0,91,0,214,0,0,0,86,0,113,0,60,0,144,0,0,0,204,0,216,0,100,0,0,0,158,0,1,0,179,0,181,0,0,0,250,0,122,0,73,0,216,0,0,0,6,0,0,0,12,0,47,0,213,0,60,0,84,0,182,0,0,0,183,0,217,0,147,0,172,0,0,0,92,0,141,0,121,0,152,0,211,0,227,0,234,0,234,0,0,0,160,0,0,0,112,0,182,0,89,0,165,0,95,0,44,0,187,0,3,0,133,0,91,0,99,0,172,0,97,0,92,0,45,0,73,0,0,0,250,0,0,0,165,0,154,0,120,0,0,0,205,0,48,0,62,0,56,0,112,0,151,0,21,0,0,0,107,0,249,0,119,0,87,0,168,0,0,0,4,0,25,0,137,0,59,0,0,0,6,0,167,0,249,0,0,0,173,0,154,0,202,0,0,0,160,0,210,0,255,0,0,0,210,0,233,0,0,0,3,0,0,0,123,0,126,0,165,0,0,0,202,0,220,0,0,0,0,0,41,0,0,0,140,0,87,0,167,0,120,0,0,0,52,0,43,0,203,0,22,0,36,0,6,0,86,0,88,0,186,0,0,0,112,0,0,0,0,0,158,0,108,0,194,0,104,0,79,0,220,0,83,0,193,0,0,0,192,0,5,0,0,0,0,0,0,0,179,0,0,0,0,0,0,0,0,0,208,0,0,0,11,0,162,0,230,0,107,0,2,0,222,0,41,0,205,0,116,0,64,0,231,0,88,0,35,0,247,0,134,0,0,0,44,0,128,0,116,0,0,0,23,0,128,0,210,0,0,0,0,0,222,0,216,0,88,0,49,0,201,0,208,0,70,0,61,0,230,0,245,0,83,0,0,0,0,0,64,0,54,0,101,0,226,0,100,0,148,0,0,0,0,0,0,0,95,0,100,0,0,0,152,0,15,0,145,0,178,0,4,0,184,0,249,0,0,0,166,0,64,0,8,0,208,0,98,0,0,0,154,0,0,0,0,0,99,0,133,0,0,0,0,0,0,0,188,0,228,0,0,0,0,0,214,0,236,0,140,0,6,0,185,0,173,0,16,0,0,0,0,0,4,0,242,0,139,0,0,0,158,0,170,0,246,0,180,0,119,0,155,0,0,0,230,0,0,0,4,0,64,0,0,0,0,0,184,0,54,0,181,0,233,0,22,0,0,0,175,0,191,0,49,0,0,0,0,0,105,0,208,0,215,0,78,0,160,0,231,0,88,0,174,0,229,0,0,0,147,0,161,0,14,0,8,0,232,0,11,0,132,0,12,0,0,0,167,0,213,0,205,0,140,0,129,0,202,0,247,0,0,0,208,0,34,0,0,0,249,0,17,0,243,0,209,0,57,0,60,0,86,0,0,0,0,0,13,0,228,0,44,0,239,0,2,0,100,0,173,0,0,0,134,0,211,0,0,0,253,0,16,0,164,0,0,0,0,0,59,0,0,0,60,0,0,0,0,0,0,0,28,0,210,0,177,0,159,0,125,0,0,0,0,0,0,0,0,0,150,0,74,0,0,0,0,0,67,0,255,0,88,0,0,0,168,0,0,0,176,0,0,0,123,0,179,0,147,0,222,0,208,0,127,0,0,0,0,0,100,0,0,0,231,0,165,0,70,0,167,0,41,0,0,0,180,0,216,0,59,0,214,0,140,0,16,0,193,0,80,0,38,0,238,0,200,0,190,0,126,0,0,0,172,0,0,0,177,0,199,0,138,0,248,0,0,0,46,0,0,0,6,0,0,0,0,0,116,0,0,0,0,0,127,0,0,0,154,0,0,0,0,0,228,0,179,0,224,0,34,0,36,0,0,0,115,0,0,0,101,0,20,0,123,0,51,0,215,0,119,0,37,0,146,0,116,0,224,0,158,0,0,0,0,0,0,0,159,0,46,0,28,0,29,0,0,0,122,0,34,0,100,0,156,0,12,0,73,0,81,0,0,0,0,0,153,0,43,0,51,0,243,0,131,0,144,0,138,0,0,0,18,0,0,0,56,0,226,0,131,0,0,0,196,0,160,0,209,0,201,0,158,0,219,0,154,0,200,0,249,0,41,0,77,0,82,0,98,0,242,0,0,0,110,0,0,0,107,0,0,0,24,0);
signal scenario_full  : scenario_type := (245,31,245,30,10,31,202,31,41,31,137,31,137,30,31,31,165,31,165,30,73,31,172,31,1,31,64,31,77,31,65,31,243,31,102,31,75,31,3,31,31,31,248,31,97,31,183,31,88,31,236,31,169,31,149,31,149,30,87,31,204,31,204,30,70,31,10,31,10,30,133,31,150,31,161,31,233,31,155,31,155,30,222,31,217,31,155,31,250,31,176,31,84,31,23,31,250,31,166,31,209,31,108,31,18,31,70,31,38,31,81,31,242,31,21,31,21,30,62,31,79,31,169,31,56,31,56,30,51,31,214,31,173,31,126,31,144,31,142,31,14,31,14,30,150,31,150,30,193,31,242,31,177,31,180,31,83,31,83,30,100,31,17,31,17,30,94,31,109,31,1,31,1,30,218,31,228,31,38,31,40,31,18,31,171,31,16,31,47,31,215,31,68,31,35,31,82,31,53,31,31,31,57,31,111,31,131,31,112,31,204,31,204,30,214,31,97,31,130,31,193,31,191,31,191,30,82,31,82,30,86,31,86,30,156,31,156,30,156,29,156,28,195,31,195,30,65,31,65,30,100,31,29,31,29,30,107,31,71,31,71,30,71,29,242,31,202,31,32,31,32,30,148,31,148,30,148,29,148,28,148,27,4,31,167,31,167,30,167,29,190,31,187,31,187,30,95,31,95,31,95,30,95,29,95,28,95,27,170,31,31,31,197,31,6,31,6,30,182,31,182,30,176,31,176,30,27,31,132,31,248,31,27,31,91,31,214,31,214,30,86,31,113,31,60,31,144,31,144,30,204,31,216,31,100,31,100,30,158,31,1,31,179,31,181,31,181,30,250,31,122,31,73,31,216,31,216,30,6,31,6,30,12,31,47,31,213,31,60,31,84,31,182,31,182,30,183,31,217,31,147,31,172,31,172,30,92,31,141,31,121,31,152,31,211,31,227,31,234,31,234,31,234,30,160,31,160,30,112,31,182,31,89,31,165,31,95,31,44,31,187,31,3,31,133,31,91,31,99,31,172,31,97,31,92,31,45,31,73,31,73,30,250,31,250,30,165,31,154,31,120,31,120,30,205,31,48,31,62,31,56,31,112,31,151,31,21,31,21,30,107,31,249,31,119,31,87,31,168,31,168,30,4,31,25,31,137,31,59,31,59,30,6,31,167,31,249,31,249,30,173,31,154,31,202,31,202,30,160,31,210,31,255,31,255,30,210,31,233,31,233,30,3,31,3,30,123,31,126,31,165,31,165,30,202,31,220,31,220,30,220,29,41,31,41,30,140,31,87,31,167,31,120,31,120,30,52,31,43,31,203,31,22,31,36,31,6,31,86,31,88,31,186,31,186,30,112,31,112,30,112,29,158,31,108,31,194,31,104,31,79,31,220,31,83,31,193,31,193,30,192,31,5,31,5,30,5,29,5,28,179,31,179,30,179,29,179,28,179,27,208,31,208,30,11,31,162,31,230,31,107,31,2,31,222,31,41,31,205,31,116,31,64,31,231,31,88,31,35,31,247,31,134,31,134,30,44,31,128,31,116,31,116,30,23,31,128,31,210,31,210,30,210,29,222,31,216,31,88,31,49,31,201,31,208,31,70,31,61,31,230,31,245,31,83,31,83,30,83,29,64,31,54,31,101,31,226,31,100,31,148,31,148,30,148,29,148,28,95,31,100,31,100,30,152,31,15,31,145,31,178,31,4,31,184,31,249,31,249,30,166,31,64,31,8,31,208,31,98,31,98,30,154,31,154,30,154,29,99,31,133,31,133,30,133,29,133,28,188,31,228,31,228,30,228,29,214,31,236,31,140,31,6,31,185,31,173,31,16,31,16,30,16,29,4,31,242,31,139,31,139,30,158,31,170,31,246,31,180,31,119,31,155,31,155,30,230,31,230,30,4,31,64,31,64,30,64,29,184,31,54,31,181,31,233,31,22,31,22,30,175,31,191,31,49,31,49,30,49,29,105,31,208,31,215,31,78,31,160,31,231,31,88,31,174,31,229,31,229,30,147,31,161,31,14,31,8,31,232,31,11,31,132,31,12,31,12,30,167,31,213,31,205,31,140,31,129,31,202,31,247,31,247,30,208,31,34,31,34,30,249,31,17,31,243,31,209,31,57,31,60,31,86,31,86,30,86,29,13,31,228,31,44,31,239,31,2,31,100,31,173,31,173,30,134,31,211,31,211,30,253,31,16,31,164,31,164,30,164,29,59,31,59,30,60,31,60,30,60,29,60,28,28,31,210,31,177,31,159,31,125,31,125,30,125,29,125,28,125,27,150,31,74,31,74,30,74,29,67,31,255,31,88,31,88,30,168,31,168,30,176,31,176,30,123,31,179,31,147,31,222,31,208,31,127,31,127,30,127,29,100,31,100,30,231,31,165,31,70,31,167,31,41,31,41,30,180,31,216,31,59,31,214,31,140,31,16,31,193,31,80,31,38,31,238,31,200,31,190,31,126,31,126,30,172,31,172,30,177,31,199,31,138,31,248,31,248,30,46,31,46,30,6,31,6,30,6,29,116,31,116,30,116,29,127,31,127,30,154,31,154,30,154,29,228,31,179,31,224,31,34,31,36,31,36,30,115,31,115,30,101,31,20,31,123,31,51,31,215,31,119,31,37,31,146,31,116,31,224,31,158,31,158,30,158,29,158,28,159,31,46,31,28,31,29,31,29,30,122,31,34,31,100,31,156,31,12,31,73,31,81,31,81,30,81,29,153,31,43,31,51,31,243,31,131,31,144,31,138,31,138,30,18,31,18,30,56,31,226,31,131,31,131,30,196,31,160,31,209,31,201,31,158,31,219,31,154,31,200,31,249,31,41,31,77,31,82,31,98,31,242,31,242,30,110,31,110,30,107,31,107,30,24,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
