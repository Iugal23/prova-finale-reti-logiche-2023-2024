-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 951;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (113,0,188,0,94,0,199,0,39,0,199,0,69,0,220,0,0,0,221,0,0,0,174,0,109,0,124,0,196,0,192,0,17,0,0,0,150,0,10,0,0,0,44,0,107,0,248,0,50,0,180,0,56,0,0,0,95,0,20,0,203,0,242,0,252,0,0,0,4,0,216,0,155,0,21,0,50,0,0,0,97,0,0,0,248,0,33,0,0,0,253,0,223,0,148,0,140,0,0,0,0,0,165,0,175,0,0,0,7,0,86,0,0,0,0,0,0,0,132,0,47,0,135,0,189,0,0,0,93,0,207,0,6,0,225,0,249,0,226,0,0,0,63,0,0,0,54,0,18,0,0,0,0,0,37,0,230,0,10,0,49,0,34,0,176,0,246,0,0,0,0,0,221,0,0,0,0,0,120,0,0,0,52,0,127,0,109,0,104,0,0,0,23,0,93,0,0,0,0,0,0,0,233,0,111,0,0,0,65,0,56,0,58,0,110,0,0,0,25,0,0,0,41,0,136,0,198,0,167,0,15,0,156,0,139,0,16,0,152,0,0,0,0,0,0,0,237,0,133,0,179,0,0,0,0,0,110,0,64,0,30,0,141,0,0,0,184,0,247,0,230,0,136,0,96,0,219,0,53,0,46,0,113,0,218,0,194,0,205,0,120,0,127,0,47,0,0,0,137,0,207,0,251,0,110,0,5,0,115,0,173,0,163,0,172,0,0,0,242,0,13,0,209,0,200,0,133,0,128,0,28,0,0,0,0,0,154,0,245,0,173,0,0,0,0,0,36,0,93,0,0,0,24,0,212,0,201,0,120,0,208,0,0,0,32,0,234,0,152,0,0,0,80,0,215,0,0,0,233,0,38,0,199,0,249,0,108,0,61,0,255,0,0,0,195,0,81,0,0,0,63,0,28,0,32,0,121,0,148,0,37,0,48,0,229,0,216,0,83,0,159,0,235,0,162,0,22,0,163,0,0,0,34,0,122,0,173,0,213,0,54,0,155,0,132,0,111,0,203,0,25,0,40,0,44,0,225,0,54,0,0,0,64,0,180,0,180,0,97,0,0,0,0,0,0,0,51,0,0,0,58,0,241,0,154,0,144,0,219,0,11,0,197,0,248,0,125,0,218,0,58,0,216,0,0,0,64,0,32,0,0,0,79,0,116,0,0,0,0,0,107,0,0,0,233,0,225,0,231,0,99,0,70,0,86,0,98,0,249,0,164,0,85,0,81,0,254,0,173,0,105,0,222,0,0,0,154,0,188,0,104,0,67,0,0,0,110,0,1,0,91,0,39,0,1,0,241,0,0,0,0,0,214,0,24,0,229,0,27,0,171,0,0,0,144,0,190,0,88,0,28,0,0,0,37,0,129,0,141,0,50,0,78,0,213,0,227,0,0,0,115,0,0,0,0,0,19,0,37,0,220,0,42,0,95,0,218,0,104,0,142,0,206,0,162,0,0,0,8,0,82,0,209,0,0,0,65,0,127,0,253,0,0,0,1,0,208,0,112,0,132,0,163,0,0,0,6,0,109,0,21,0,69,0,0,0,115,0,125,0,143,0,195,0,0,0,188,0,201,0,200,0,123,0,28,0,73,0,20,0,189,0,253,0,75,0,0,0,246,0,42,0,53,0,251,0,201,0,241,0,112,0,0,0,247,0,167,0,141,0,0,0,147,0,220,0,65,0,255,0,219,0,132,0,205,0,87,0,230,0,36,0,167,0,112,0,183,0,161,0,41,0,254,0,38,0,99,0,224,0,55,0,148,0,0,0,0,0,81,0,139,0,39,0,150,0,29,0,0,0,0,0,146,0,214,0,0,0,0,0,54,0,60,0,114,0,35,0,12,0,101,0,0,0,150,0,124,0,0,0,5,0,0,0,205,0,166,0,213,0,52,0,215,0,150,0,225,0,221,0,0,0,38,0,0,0,127,0,204,0,52,0,179,0,19,0,25,0,159,0,0,0,62,0,153,0,230,0,123,0,0,0,67,0,0,0,0,0,161,0,0,0,0,0,214,0,33,0,33,0,84,0,116,0,178,0,7,0,0,0,3,0,144,0,223,0,0,0,22,0,121,0,48,0,254,0,184,0,192,0,228,0,0,0,127,0,243,0,79,0,236,0,100,0,59,0,177,0,32,0,220,0,201,0,48,0,245,0,44,0,105,0,0,0,0,0,15,0,96,0,76,0,114,0,160,0,176,0,232,0,49,0,116,0,110,0,3,0,71,0,1,0,51,0,0,0,0,0,8,0,60,0,169,0,87,0,42,0,0,0,0,0,55,0,225,0,245,0,0,0,100,0,245,0,0,0,208,0,145,0,140,0,218,0,104,0,244,0,154,0,55,0,108,0,122,0,47,0,125,0,146,0,57,0,154,0,198,0,134,0,159,0,38,0,8,0,25,0,0,0,68,0,25,0,0,0,200,0,97,0,101,0,0,0,226,0,81,0,67,0,195,0,0,0,150,0,75,0,217,0,165,0,164,0,56,0,142,0,0,0,159,0,156,0,183,0,172,0,127,0,200,0,130,0,0,0,92,0,4,0,166,0,254,0,32,0,228,0,130,0,110,0,69,0,116,0,210,0,0,0,16,0,153,0,63,0,80,0,118,0,178,0,72,0,59,0,234,0,0,0,158,0,94,0,99,0,112,0,90,0,146,0,0,0,112,0,105,0,97,0,195,0,46,0,0,0,246,0,0,0,50,0,176,0,201,0,252,0,65,0,66,0,22,0,80,0,111,0,241,0,226,0,5,0,188,0,234,0,0,0,226,0,107,0,127,0,199,0,148,0,0,0,129,0,27,0,99,0,104,0,0,0,58,0,38,0,0,0,58,0,226,0,205,0,84,0,48,0,104,0,123,0,214,0,167,0,0,0,221,0,194,0,152,0,29,0,0,0,21,0,158,0,193,0,169,0,60,0,0,0,29,0,115,0,228,0,0,0,254,0,19,0,173,0,0,0,59,0,0,0,211,0,227,0,118,0,88,0,251,0,50,0,85,0,191,0,0,0,60,0,85,0,92,0,48,0,0,0,252,0,223,0,90,0,0,0,51,0,9,0,65,0,237,0,124,0,198,0,0,0,230,0,69,0,19,0,178,0,17,0,121,0,162,0,80,0,0,0,236,0,0,0,29,0,201,0,0,0,92,0,97,0,98,0,0,0,143,0,123,0,207,0,193,0,0,0,106,0,36,0,144,0,52,0,41,0,56,0,188,0,143,0,0,0,0,0,240,0,0,0,13,0,0,0,227,0,182,0,63,0,28,0,68,0,202,0,164,0,0,0,53,0,0,0,169,0,199,0,0,0,13,0,129,0,178,0,137,0,196,0,175,0,128,0,229,0,122,0,166,0,197,0,246,0,42,0,148,0,65,0,184,0,95,0,196,0,0,0,216,0,185,0,141,0,69,0,41,0,0,0,89,0,186,0,115,0,127,0,254,0,38,0,60,0,122,0,42,0,0,0,250,0,0,0,132,0,82,0,170,0,171,0,227,0,161,0,198,0,146,0,194,0,40,0,58,0,60,0,0,0,0,0,13,0,234,0,154,0,83,0,0,0,66,0,135,0,213,0,169,0,168,0,247,0,157,0,101,0,132,0,241,0,0,0,35,0,253,0,231,0,175,0,202,0,215,0,42,0,57,0,130,0,148,0,104,0,194,0,188,0,196,0,44,0,255,0,84,0,210,0,111,0,0,0,0,0,104,0,147,0,145,0,0,0,0,0,80,0,227,0,203,0,160,0,53,0,73,0,201,0,34,0,171,0,38,0,69,0,0,0,17,0,0,0,131,0,254,0,68,0,119,0,13,0,0,0,140,0,69,0,193,0,77,0,65,0,33,0,165,0,201,0,150,0,101,0,87,0,165,0,215,0,223,0,0,0,0,0,81,0,0,0,169,0,0,0,193,0,180,0,0,0,1,0,0,0,166,0,30,0,0,0,0,0,210,0,79,0,17,0,62,0,92,0,252,0,0,0,0,0,0,0,0,0,96,0,0,0,226,0,137,0,58,0,205,0,232,0,0,0,60,0,77,0,32,0,0,0,0,0,32,0,0,0,64,0,57,0,112,0,123,0,0,0,239,0,207,0,74,0,100,0,202,0,0,0,0,0,45,0,0,0,80,0,0,0,0,0,119,0,63,0,186,0,0,0,92,0,50,0,58,0,179,0,0,0,228,0,0,0,0,0,0,0,125,0,0,0,187,0,144,0,105,0,232,0,0,0,112,0,224,0,0,0,148,0,238,0,19,0,0,0,32,0,163,0,136,0,119,0,102,0);
signal scenario_full  : scenario_type := (113,31,188,31,94,31,199,31,39,31,199,31,69,31,220,31,220,30,221,31,221,30,174,31,109,31,124,31,196,31,192,31,17,31,17,30,150,31,10,31,10,30,44,31,107,31,248,31,50,31,180,31,56,31,56,30,95,31,20,31,203,31,242,31,252,31,252,30,4,31,216,31,155,31,21,31,50,31,50,30,97,31,97,30,248,31,33,31,33,30,253,31,223,31,148,31,140,31,140,30,140,29,165,31,175,31,175,30,7,31,86,31,86,30,86,29,86,28,132,31,47,31,135,31,189,31,189,30,93,31,207,31,6,31,225,31,249,31,226,31,226,30,63,31,63,30,54,31,18,31,18,30,18,29,37,31,230,31,10,31,49,31,34,31,176,31,246,31,246,30,246,29,221,31,221,30,221,29,120,31,120,30,52,31,127,31,109,31,104,31,104,30,23,31,93,31,93,30,93,29,93,28,233,31,111,31,111,30,65,31,56,31,58,31,110,31,110,30,25,31,25,30,41,31,136,31,198,31,167,31,15,31,156,31,139,31,16,31,152,31,152,30,152,29,152,28,237,31,133,31,179,31,179,30,179,29,110,31,64,31,30,31,141,31,141,30,184,31,247,31,230,31,136,31,96,31,219,31,53,31,46,31,113,31,218,31,194,31,205,31,120,31,127,31,47,31,47,30,137,31,207,31,251,31,110,31,5,31,115,31,173,31,163,31,172,31,172,30,242,31,13,31,209,31,200,31,133,31,128,31,28,31,28,30,28,29,154,31,245,31,173,31,173,30,173,29,36,31,93,31,93,30,24,31,212,31,201,31,120,31,208,31,208,30,32,31,234,31,152,31,152,30,80,31,215,31,215,30,233,31,38,31,199,31,249,31,108,31,61,31,255,31,255,30,195,31,81,31,81,30,63,31,28,31,32,31,121,31,148,31,37,31,48,31,229,31,216,31,83,31,159,31,235,31,162,31,22,31,163,31,163,30,34,31,122,31,173,31,213,31,54,31,155,31,132,31,111,31,203,31,25,31,40,31,44,31,225,31,54,31,54,30,64,31,180,31,180,31,97,31,97,30,97,29,97,28,51,31,51,30,58,31,241,31,154,31,144,31,219,31,11,31,197,31,248,31,125,31,218,31,58,31,216,31,216,30,64,31,32,31,32,30,79,31,116,31,116,30,116,29,107,31,107,30,233,31,225,31,231,31,99,31,70,31,86,31,98,31,249,31,164,31,85,31,81,31,254,31,173,31,105,31,222,31,222,30,154,31,188,31,104,31,67,31,67,30,110,31,1,31,91,31,39,31,1,31,241,31,241,30,241,29,214,31,24,31,229,31,27,31,171,31,171,30,144,31,190,31,88,31,28,31,28,30,37,31,129,31,141,31,50,31,78,31,213,31,227,31,227,30,115,31,115,30,115,29,19,31,37,31,220,31,42,31,95,31,218,31,104,31,142,31,206,31,162,31,162,30,8,31,82,31,209,31,209,30,65,31,127,31,253,31,253,30,1,31,208,31,112,31,132,31,163,31,163,30,6,31,109,31,21,31,69,31,69,30,115,31,125,31,143,31,195,31,195,30,188,31,201,31,200,31,123,31,28,31,73,31,20,31,189,31,253,31,75,31,75,30,246,31,42,31,53,31,251,31,201,31,241,31,112,31,112,30,247,31,167,31,141,31,141,30,147,31,220,31,65,31,255,31,219,31,132,31,205,31,87,31,230,31,36,31,167,31,112,31,183,31,161,31,41,31,254,31,38,31,99,31,224,31,55,31,148,31,148,30,148,29,81,31,139,31,39,31,150,31,29,31,29,30,29,29,146,31,214,31,214,30,214,29,54,31,60,31,114,31,35,31,12,31,101,31,101,30,150,31,124,31,124,30,5,31,5,30,205,31,166,31,213,31,52,31,215,31,150,31,225,31,221,31,221,30,38,31,38,30,127,31,204,31,52,31,179,31,19,31,25,31,159,31,159,30,62,31,153,31,230,31,123,31,123,30,67,31,67,30,67,29,161,31,161,30,161,29,214,31,33,31,33,31,84,31,116,31,178,31,7,31,7,30,3,31,144,31,223,31,223,30,22,31,121,31,48,31,254,31,184,31,192,31,228,31,228,30,127,31,243,31,79,31,236,31,100,31,59,31,177,31,32,31,220,31,201,31,48,31,245,31,44,31,105,31,105,30,105,29,15,31,96,31,76,31,114,31,160,31,176,31,232,31,49,31,116,31,110,31,3,31,71,31,1,31,51,31,51,30,51,29,8,31,60,31,169,31,87,31,42,31,42,30,42,29,55,31,225,31,245,31,245,30,100,31,245,31,245,30,208,31,145,31,140,31,218,31,104,31,244,31,154,31,55,31,108,31,122,31,47,31,125,31,146,31,57,31,154,31,198,31,134,31,159,31,38,31,8,31,25,31,25,30,68,31,25,31,25,30,200,31,97,31,101,31,101,30,226,31,81,31,67,31,195,31,195,30,150,31,75,31,217,31,165,31,164,31,56,31,142,31,142,30,159,31,156,31,183,31,172,31,127,31,200,31,130,31,130,30,92,31,4,31,166,31,254,31,32,31,228,31,130,31,110,31,69,31,116,31,210,31,210,30,16,31,153,31,63,31,80,31,118,31,178,31,72,31,59,31,234,31,234,30,158,31,94,31,99,31,112,31,90,31,146,31,146,30,112,31,105,31,97,31,195,31,46,31,46,30,246,31,246,30,50,31,176,31,201,31,252,31,65,31,66,31,22,31,80,31,111,31,241,31,226,31,5,31,188,31,234,31,234,30,226,31,107,31,127,31,199,31,148,31,148,30,129,31,27,31,99,31,104,31,104,30,58,31,38,31,38,30,58,31,226,31,205,31,84,31,48,31,104,31,123,31,214,31,167,31,167,30,221,31,194,31,152,31,29,31,29,30,21,31,158,31,193,31,169,31,60,31,60,30,29,31,115,31,228,31,228,30,254,31,19,31,173,31,173,30,59,31,59,30,211,31,227,31,118,31,88,31,251,31,50,31,85,31,191,31,191,30,60,31,85,31,92,31,48,31,48,30,252,31,223,31,90,31,90,30,51,31,9,31,65,31,237,31,124,31,198,31,198,30,230,31,69,31,19,31,178,31,17,31,121,31,162,31,80,31,80,30,236,31,236,30,29,31,201,31,201,30,92,31,97,31,98,31,98,30,143,31,123,31,207,31,193,31,193,30,106,31,36,31,144,31,52,31,41,31,56,31,188,31,143,31,143,30,143,29,240,31,240,30,13,31,13,30,227,31,182,31,63,31,28,31,68,31,202,31,164,31,164,30,53,31,53,30,169,31,199,31,199,30,13,31,129,31,178,31,137,31,196,31,175,31,128,31,229,31,122,31,166,31,197,31,246,31,42,31,148,31,65,31,184,31,95,31,196,31,196,30,216,31,185,31,141,31,69,31,41,31,41,30,89,31,186,31,115,31,127,31,254,31,38,31,60,31,122,31,42,31,42,30,250,31,250,30,132,31,82,31,170,31,171,31,227,31,161,31,198,31,146,31,194,31,40,31,58,31,60,31,60,30,60,29,13,31,234,31,154,31,83,31,83,30,66,31,135,31,213,31,169,31,168,31,247,31,157,31,101,31,132,31,241,31,241,30,35,31,253,31,231,31,175,31,202,31,215,31,42,31,57,31,130,31,148,31,104,31,194,31,188,31,196,31,44,31,255,31,84,31,210,31,111,31,111,30,111,29,104,31,147,31,145,31,145,30,145,29,80,31,227,31,203,31,160,31,53,31,73,31,201,31,34,31,171,31,38,31,69,31,69,30,17,31,17,30,131,31,254,31,68,31,119,31,13,31,13,30,140,31,69,31,193,31,77,31,65,31,33,31,165,31,201,31,150,31,101,31,87,31,165,31,215,31,223,31,223,30,223,29,81,31,81,30,169,31,169,30,193,31,180,31,180,30,1,31,1,30,166,31,30,31,30,30,30,29,210,31,79,31,17,31,62,31,92,31,252,31,252,30,252,29,252,28,252,27,96,31,96,30,226,31,137,31,58,31,205,31,232,31,232,30,60,31,77,31,32,31,32,30,32,29,32,31,32,30,64,31,57,31,112,31,123,31,123,30,239,31,207,31,74,31,100,31,202,31,202,30,202,29,45,31,45,30,80,31,80,30,80,29,119,31,63,31,186,31,186,30,92,31,50,31,58,31,179,31,179,30,228,31,228,30,228,29,228,28,125,31,125,30,187,31,144,31,105,31,232,31,232,30,112,31,224,31,224,30,148,31,238,31,19,31,19,30,32,31,163,31,136,31,119,31,102,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
