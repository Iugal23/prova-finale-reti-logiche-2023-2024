-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_345 is
end project_tb_345;

architecture project_tb_arch_345 of project_tb_345 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 670;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (137,0,0,0,38,0,0,0,185,0,190,0,100,0,171,0,156,0,200,0,0,0,95,0,246,0,52,0,0,0,1,0,215,0,91,0,144,0,62,0,154,0,119,0,112,0,0,0,11,0,139,0,237,0,253,0,0,0,159,0,73,0,206,0,104,0,0,0,0,0,66,0,214,0,0,0,68,0,106,0,27,0,0,0,93,0,31,0,78,0,240,0,0,0,252,0,43,0,235,0,206,0,20,0,255,0,0,0,113,0,230,0,121,0,139,0,161,0,0,0,253,0,0,0,154,0,202,0,0,0,237,0,77,0,0,0,104,0,33,0,0,0,232,0,123,0,85,0,216,0,146,0,47,0,62,0,152,0,137,0,19,0,200,0,119,0,165,0,170,0,34,0,51,0,92,0,0,0,250,0,2,0,0,0,25,0,0,0,68,0,88,0,127,0,0,0,0,0,67,0,111,0,51,0,0,0,57,0,129,0,254,0,239,0,74,0,44,0,110,0,38,0,63,0,214,0,0,0,80,0,217,0,142,0,19,0,185,0,91,0,164,0,172,0,0,0,0,0,0,0,225,0,104,0,56,0,35,0,164,0,236,0,149,0,186,0,217,0,44,0,0,0,101,0,2,0,120,0,241,0,0,0,56,0,153,0,248,0,162,0,211,0,188,0,244,0,183,0,71,0,5,0,57,0,0,0,0,0,171,0,195,0,220,0,118,0,165,0,79,0,0,0,134,0,9,0,58,0,0,0,0,0,0,0,117,0,99,0,47,0,246,0,29,0,171,0,0,0,89,0,0,0,70,0,250,0,101,0,230,0,139,0,59,0,248,0,0,0,0,0,179,0,93,0,0,0,0,0,98,0,0,0,144,0,46,0,29,0,223,0,0,0,65,0,0,0,110,0,0,0,0,0,110,0,184,0,22,0,152,0,249,0,84,0,36,0,214,0,59,0,193,0,0,0,190,0,0,0,217,0,0,0,96,0,0,0,227,0,49,0,88,0,12,0,0,0,0,0,0,0,2,0,62,0,0,0,16,0,53,0,140,0,73,0,150,0,171,0,141,0,98,0,0,0,0,0,89,0,140,0,77,0,179,0,6,0,200,0,204,0,233,0,0,0,129,0,0,0,143,0,234,0,80,0,236,0,120,0,55,0,137,0,0,0,249,0,9,0,174,0,159,0,120,0,0,0,0,0,160,0,9,0,0,0,77,0,0,0,190,0,104,0,248,0,253,0,190,0,0,0,0,0,19,0,22,0,191,0,243,0,84,0,48,0,145,0,82,0,32,0,243,0,252,0,85,0,97,0,186,0,58,0,69,0,77,0,62,0,204,0,168,0,157,0,0,0,10,0,58,0,59,0,0,0,181,0,97,0,0,0,0,0,204,0,40,0,0,0,30,0,2,0,126,0,186,0,18,0,232,0,181,0,161,0,2,0,185,0,9,0,219,0,79,0,0,0,0,0,172,0,86,0,140,0,136,0,0,0,56,0,0,0,119,0,70,0,81,0,52,0,114,0,0,0,80,0,82,0,0,0,0,0,162,0,214,0,104,0,0,0,77,0,246,0,19,0,101,0,20,0,32,0,229,0,209,0,224,0,120,0,74,0,74,0,250,0,0,0,0,0,0,0,140,0,0,0,45,0,19,0,237,0,25,0,0,0,186,0,208,0,57,0,54,0,52,0,62,0,165,0,180,0,0,0,249,0,21,0,217,0,117,0,100,0,0,0,176,0,70,0,18,0,59,0,84,0,63,0,66,0,0,0,76,0,5,0,240,0,224,0,187,0,187,0,147,0,133,0,199,0,113,0,0,0,141,0,60,0,0,0,5,0,179,0,21,0,167,0,5,0,106,0,148,0,7,0,4,0,0,0,26,0,0,0,130,0,169,0,169,0,137,0,0,0,78,0,97,0,96,0,143,0,0,0,0,0,77,0,129,0,0,0,158,0,106,0,145,0,234,0,77,0,162,0,224,0,0,0,0,0,208,0,165,0,217,0,0,0,198,0,50,0,52,0,181,0,64,0,103,0,0,0,60,0,22,0,211,0,0,0,117,0,175,0,151,0,0,0,151,0,247,0,0,0,72,0,49,0,0,0,0,0,144,0,163,0,175,0,37,0,155,0,40,0,196,0,123,0,130,0,181,0,0,0,139,0,186,0,145,0,112,0,158,0,161,0,251,0,166,0,0,0,58,0,39,0,53,0,0,0,5,0,0,0,182,0,248,0,0,0,124,0,163,0,0,0,114,0,0,0,0,0,100,0,0,0,0,0,0,0,231,0,142,0,201,0,249,0,0,0,68,0,171,0,94,0,161,0,154,0,217,0,0,0,69,0,242,0,178,0,253,0,144,0,126,0,255,0,107,0,28,0,191,0,146,0,123,0,188,0,77,0,74,0,88,0,19,0,5,0,0,0,0,0,16,0,123,0,0,0,0,0,0,0,28,0,119,0,0,0,154,0,182,0,92,0,0,0,199,0,4,0,27,0,161,0,39,0,5,0,85,0,166,0,254,0,77,0,113,0,236,0,33,0,189,0,90,0,214,0,208,0,45,0,123,0,101,0,243,0,53,0,115,0,190,0,228,0,0,0,0,0,0,0,77,0,136,0,1,0,0,0,60,0,254,0,0,0,103,0,193,0,177,0,0,0,0,0,210,0,104,0,198,0,0,0,58,0,15,0,22,0,213,0,14,0,81,0,0,0,0,0,58,0,61,0,32,0,219,0,134,0,244,0,189,0,188,0,87,0,226,0,132,0,0,0,0,0,100,0,2,0,79,0,0,0,209,0,106,0,46,0,6,0,100,0,105,0,0,0,10,0,0,0,193,0,54,0,95,0,239,0,85,0,91,0,63,0,29,0,0,0,0,0,117,0,205,0,8,0,0,0,0,0,34,0,143,0,100,0,230,0,107,0,193,0,132,0,209,0,0,0,0,0,0,0,31,0,47,0,93,0,115,0,53,0,243,0,50,0,187,0,67,0,192,0,184,0,15,0,71,0,108,0,157,0,124,0,122,0);
signal scenario_full  : scenario_type := (137,31,137,30,38,31,38,30,185,31,190,31,100,31,171,31,156,31,200,31,200,30,95,31,246,31,52,31,52,30,1,31,215,31,91,31,144,31,62,31,154,31,119,31,112,31,112,30,11,31,139,31,237,31,253,31,253,30,159,31,73,31,206,31,104,31,104,30,104,29,66,31,214,31,214,30,68,31,106,31,27,31,27,30,93,31,31,31,78,31,240,31,240,30,252,31,43,31,235,31,206,31,20,31,255,31,255,30,113,31,230,31,121,31,139,31,161,31,161,30,253,31,253,30,154,31,202,31,202,30,237,31,77,31,77,30,104,31,33,31,33,30,232,31,123,31,85,31,216,31,146,31,47,31,62,31,152,31,137,31,19,31,200,31,119,31,165,31,170,31,34,31,51,31,92,31,92,30,250,31,2,31,2,30,25,31,25,30,68,31,88,31,127,31,127,30,127,29,67,31,111,31,51,31,51,30,57,31,129,31,254,31,239,31,74,31,44,31,110,31,38,31,63,31,214,31,214,30,80,31,217,31,142,31,19,31,185,31,91,31,164,31,172,31,172,30,172,29,172,28,225,31,104,31,56,31,35,31,164,31,236,31,149,31,186,31,217,31,44,31,44,30,101,31,2,31,120,31,241,31,241,30,56,31,153,31,248,31,162,31,211,31,188,31,244,31,183,31,71,31,5,31,57,31,57,30,57,29,171,31,195,31,220,31,118,31,165,31,79,31,79,30,134,31,9,31,58,31,58,30,58,29,58,28,117,31,99,31,47,31,246,31,29,31,171,31,171,30,89,31,89,30,70,31,250,31,101,31,230,31,139,31,59,31,248,31,248,30,248,29,179,31,93,31,93,30,93,29,98,31,98,30,144,31,46,31,29,31,223,31,223,30,65,31,65,30,110,31,110,30,110,29,110,31,184,31,22,31,152,31,249,31,84,31,36,31,214,31,59,31,193,31,193,30,190,31,190,30,217,31,217,30,96,31,96,30,227,31,49,31,88,31,12,31,12,30,12,29,12,28,2,31,62,31,62,30,16,31,53,31,140,31,73,31,150,31,171,31,141,31,98,31,98,30,98,29,89,31,140,31,77,31,179,31,6,31,200,31,204,31,233,31,233,30,129,31,129,30,143,31,234,31,80,31,236,31,120,31,55,31,137,31,137,30,249,31,9,31,174,31,159,31,120,31,120,30,120,29,160,31,9,31,9,30,77,31,77,30,190,31,104,31,248,31,253,31,190,31,190,30,190,29,19,31,22,31,191,31,243,31,84,31,48,31,145,31,82,31,32,31,243,31,252,31,85,31,97,31,186,31,58,31,69,31,77,31,62,31,204,31,168,31,157,31,157,30,10,31,58,31,59,31,59,30,181,31,97,31,97,30,97,29,204,31,40,31,40,30,30,31,2,31,126,31,186,31,18,31,232,31,181,31,161,31,2,31,185,31,9,31,219,31,79,31,79,30,79,29,172,31,86,31,140,31,136,31,136,30,56,31,56,30,119,31,70,31,81,31,52,31,114,31,114,30,80,31,82,31,82,30,82,29,162,31,214,31,104,31,104,30,77,31,246,31,19,31,101,31,20,31,32,31,229,31,209,31,224,31,120,31,74,31,74,31,250,31,250,30,250,29,250,28,140,31,140,30,45,31,19,31,237,31,25,31,25,30,186,31,208,31,57,31,54,31,52,31,62,31,165,31,180,31,180,30,249,31,21,31,217,31,117,31,100,31,100,30,176,31,70,31,18,31,59,31,84,31,63,31,66,31,66,30,76,31,5,31,240,31,224,31,187,31,187,31,147,31,133,31,199,31,113,31,113,30,141,31,60,31,60,30,5,31,179,31,21,31,167,31,5,31,106,31,148,31,7,31,4,31,4,30,26,31,26,30,130,31,169,31,169,31,137,31,137,30,78,31,97,31,96,31,143,31,143,30,143,29,77,31,129,31,129,30,158,31,106,31,145,31,234,31,77,31,162,31,224,31,224,30,224,29,208,31,165,31,217,31,217,30,198,31,50,31,52,31,181,31,64,31,103,31,103,30,60,31,22,31,211,31,211,30,117,31,175,31,151,31,151,30,151,31,247,31,247,30,72,31,49,31,49,30,49,29,144,31,163,31,175,31,37,31,155,31,40,31,196,31,123,31,130,31,181,31,181,30,139,31,186,31,145,31,112,31,158,31,161,31,251,31,166,31,166,30,58,31,39,31,53,31,53,30,5,31,5,30,182,31,248,31,248,30,124,31,163,31,163,30,114,31,114,30,114,29,100,31,100,30,100,29,100,28,231,31,142,31,201,31,249,31,249,30,68,31,171,31,94,31,161,31,154,31,217,31,217,30,69,31,242,31,178,31,253,31,144,31,126,31,255,31,107,31,28,31,191,31,146,31,123,31,188,31,77,31,74,31,88,31,19,31,5,31,5,30,5,29,16,31,123,31,123,30,123,29,123,28,28,31,119,31,119,30,154,31,182,31,92,31,92,30,199,31,4,31,27,31,161,31,39,31,5,31,85,31,166,31,254,31,77,31,113,31,236,31,33,31,189,31,90,31,214,31,208,31,45,31,123,31,101,31,243,31,53,31,115,31,190,31,228,31,228,30,228,29,228,28,77,31,136,31,1,31,1,30,60,31,254,31,254,30,103,31,193,31,177,31,177,30,177,29,210,31,104,31,198,31,198,30,58,31,15,31,22,31,213,31,14,31,81,31,81,30,81,29,58,31,61,31,32,31,219,31,134,31,244,31,189,31,188,31,87,31,226,31,132,31,132,30,132,29,100,31,2,31,79,31,79,30,209,31,106,31,46,31,6,31,100,31,105,31,105,30,10,31,10,30,193,31,54,31,95,31,239,31,85,31,91,31,63,31,29,31,29,30,29,29,117,31,205,31,8,31,8,30,8,29,34,31,143,31,100,31,230,31,107,31,193,31,132,31,209,31,209,30,209,29,209,28,31,31,47,31,93,31,115,31,53,31,243,31,50,31,187,31,67,31,192,31,184,31,15,31,71,31,108,31,157,31,124,31,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
