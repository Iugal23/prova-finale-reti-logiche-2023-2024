-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 273;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,177,0,114,0,54,0,176,0,176,0,5,0,0,0,110,0,177,0,0,0,164,0,91,0,67,0,252,0,0,0,73,0,70,0,192,0,239,0,88,0,121,0,144,0,197,0,85,0,88,0,139,0,81,0,0,0,50,0,116,0,0,0,0,0,80,0,38,0,0,0,242,0,252,0,177,0,94,0,200,0,0,0,60,0,247,0,52,0,180,0,245,0,243,0,238,0,254,0,31,0,48,0,121,0,241,0,234,0,0,0,0,0,220,0,81,0,33,0,102,0,176,0,138,0,115,0,246,0,15,0,55,0,118,0,0,0,206,0,0,0,242,0,0,0,38,0,0,0,146,0,150,0,102,0,206,0,27,0,0,0,214,0,15,0,108,0,92,0,37,0,0,0,0,0,0,0,0,0,40,0,186,0,189,0,251,0,0,0,232,0,0,0,222,0,84,0,90,0,0,0,251,0,93,0,171,0,145,0,0,0,0,0,0,0,0,0,60,0,85,0,231,0,57,0,182,0,17,0,77,0,43,0,0,0,0,0,87,0,0,0,97,0,0,0,180,0,160,0,231,0,158,0,38,0,0,0,164,0,137,0,176,0,59,0,0,0,99,0,254,0,173,0,21,0,214,0,31,0,0,0,89,0,112,0,0,0,210,0,18,0,214,0,81,0,192,0,0,0,83,0,0,0,123,0,53,0,226,0,0,0,139,0,26,0,0,0,26,0,0,0,57,0,187,0,0,0,178,0,152,0,253,0,181,0,159,0,245,0,83,0,0,0,162,0,240,0,36,0,0,0,0,0,141,0,0,0,88,0,38,0,147,0,112,0,58,0,146,0,109,0,84,0,155,0,0,0,207,0,250,0,135,0,240,0,205,0,30,0,159,0,134,0,64,0,61,0,0,0,237,0,246,0,60,0,27,0,3,0,63,0,131,0,3,0,165,0,103,0,64,0,186,0,245,0,24,0,229,0,0,0,6,0,21,0,188,0,8,0,120,0,105,0,207,0,232,0,250,0,95,0,195,0,200,0,135,0,146,0,0,0,53,0,171,0,46,0,0,0,210,0,167,0,223,0,198,0,117,0,9,0,87,0,0,0,186,0,125,0,213,0,100,0,38,0,230,0,254,0,32,0,0,0,166,0,0,0,11,0,138,0,0,0,0,0,168,0,109,0,246,0,222,0,122,0,193,0,0,0,114,0,4,0,82,0,37,0,0,0,135,0,180,0,130,0);
signal scenario_full  : scenario_type := (135,31,177,31,114,31,54,31,176,31,176,31,5,31,5,30,110,31,177,31,177,30,164,31,91,31,67,31,252,31,252,30,73,31,70,31,192,31,239,31,88,31,121,31,144,31,197,31,85,31,88,31,139,31,81,31,81,30,50,31,116,31,116,30,116,29,80,31,38,31,38,30,242,31,252,31,177,31,94,31,200,31,200,30,60,31,247,31,52,31,180,31,245,31,243,31,238,31,254,31,31,31,48,31,121,31,241,31,234,31,234,30,234,29,220,31,81,31,33,31,102,31,176,31,138,31,115,31,246,31,15,31,55,31,118,31,118,30,206,31,206,30,242,31,242,30,38,31,38,30,146,31,150,31,102,31,206,31,27,31,27,30,214,31,15,31,108,31,92,31,37,31,37,30,37,29,37,28,37,27,40,31,186,31,189,31,251,31,251,30,232,31,232,30,222,31,84,31,90,31,90,30,251,31,93,31,171,31,145,31,145,30,145,29,145,28,145,27,60,31,85,31,231,31,57,31,182,31,17,31,77,31,43,31,43,30,43,29,87,31,87,30,97,31,97,30,180,31,160,31,231,31,158,31,38,31,38,30,164,31,137,31,176,31,59,31,59,30,99,31,254,31,173,31,21,31,214,31,31,31,31,30,89,31,112,31,112,30,210,31,18,31,214,31,81,31,192,31,192,30,83,31,83,30,123,31,53,31,226,31,226,30,139,31,26,31,26,30,26,31,26,30,57,31,187,31,187,30,178,31,152,31,253,31,181,31,159,31,245,31,83,31,83,30,162,31,240,31,36,31,36,30,36,29,141,31,141,30,88,31,38,31,147,31,112,31,58,31,146,31,109,31,84,31,155,31,155,30,207,31,250,31,135,31,240,31,205,31,30,31,159,31,134,31,64,31,61,31,61,30,237,31,246,31,60,31,27,31,3,31,63,31,131,31,3,31,165,31,103,31,64,31,186,31,245,31,24,31,229,31,229,30,6,31,21,31,188,31,8,31,120,31,105,31,207,31,232,31,250,31,95,31,195,31,200,31,135,31,146,31,146,30,53,31,171,31,46,31,46,30,210,31,167,31,223,31,198,31,117,31,9,31,87,31,87,30,186,31,125,31,213,31,100,31,38,31,230,31,254,31,32,31,32,30,166,31,166,30,11,31,138,31,138,30,138,29,168,31,109,31,246,31,222,31,122,31,193,31,193,30,114,31,4,31,82,31,37,31,37,30,135,31,180,31,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
