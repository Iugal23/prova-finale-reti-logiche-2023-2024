-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_462 is
end project_tb_462;

architecture project_tb_arch_462 of project_tb_462 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 348;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,99,0,163,0,108,0,1,0,113,0,141,0,128,0,228,0,52,0,0,0,211,0,40,0,0,0,179,0,0,0,89,0,221,0,122,0,235,0,239,0,254,0,25,0,40,0,200,0,50,0,63,0,225,0,57,0,74,0,0,0,60,0,0,0,29,0,159,0,0,0,0,0,1,0,206,0,0,0,66,0,192,0,159,0,138,0,250,0,145,0,149,0,186,0,94,0,0,0,173,0,43,0,141,0,81,0,99,0,0,0,212,0,59,0,52,0,58,0,144,0,82,0,76,0,220,0,111,0,85,0,118,0,145,0,178,0,53,0,215,0,245,0,240,0,6,0,103,0,0,0,152,0,0,0,57,0,207,0,252,0,216,0,220,0,162,0,179,0,66,0,179,0,229,0,200,0,240,0,0,0,0,0,0,0,112,0,163,0,135,0,101,0,0,0,0,0,0,0,25,0,37,0,91,0,173,0,0,0,83,0,70,0,74,0,246,0,140,0,0,0,39,0,0,0,15,0,102,0,87,0,219,0,90,0,0,0,63,0,120,0,0,0,75,0,175,0,28,0,79,0,0,0,0,0,75,0,80,0,205,0,68,0,1,0,225,0,155,0,181,0,136,0,221,0,62,0,125,0,154,0,174,0,160,0,74,0,188,0,192,0,155,0,157,0,203,0,112,0,0,0,179,0,186,0,117,0,0,0,4,0,167,0,14,0,176,0,225,0,0,0,125,0,240,0,175,0,25,0,0,0,192,0,194,0,162,0,168,0,109,0,43,0,161,0,66,0,9,0,59,0,195,0,233,0,44,0,92,0,131,0,92,0,155,0,43,0,44,0,186,0,113,0,0,0,169,0,172,0,116,0,43,0,186,0,132,0,251,0,0,0,175,0,136,0,134,0,218,0,163,0,184,0,216,0,209,0,0,0,32,0,163,0,37,0,72,0,22,0,64,0,0,0,0,0,240,0,154,0,155,0,0,0,0,0,91,0,72,0,106,0,112,0,198,0,0,0,94,0,182,0,70,0,117,0,183,0,66,0,29,0,130,0,232,0,194,0,0,0,177,0,204,0,109,0,130,0,0,0,124,0,9,0,0,0,146,0,112,0,0,0,119,0,115,0,179,0,0,0,145,0,219,0,22,0,96,0,123,0,201,0,126,0,186,0,110,0,79,0,0,0,0,0,165,0,13,0,58,0,199,0,0,0,0,0,0,0,0,0,194,0,0,0,0,0,83,0,90,0,174,0,76,0,49,0,245,0,0,0,40,0,103,0,0,0,0,0,0,0,156,0,151,0,92,0,227,0,0,0,229,0,139,0,92,0,162,0,0,0,4,0,104,0,163,0,0,0,3,0,228,0,150,0,0,0,213,0,20,0,6,0,159,0,0,0,181,0,51,0,0,0,52,0,42,0,30,0,49,0,15,0,235,0,17,0,39,0,229,0,140,0,101,0,107,0,0,0,232,0,100,0,0,0,57,0,0,0,121,0,210,0,76,0,168,0,225,0,107,0,190,0,10,0,115,0,74,0,248,0,152,0,45,0,121,0,0,0,0,0,187,0,4,0,75,0);
signal scenario_full  : scenario_type := (0,0,99,31,163,31,108,31,1,31,113,31,141,31,128,31,228,31,52,31,52,30,211,31,40,31,40,30,179,31,179,30,89,31,221,31,122,31,235,31,239,31,254,31,25,31,40,31,200,31,50,31,63,31,225,31,57,31,74,31,74,30,60,31,60,30,29,31,159,31,159,30,159,29,1,31,206,31,206,30,66,31,192,31,159,31,138,31,250,31,145,31,149,31,186,31,94,31,94,30,173,31,43,31,141,31,81,31,99,31,99,30,212,31,59,31,52,31,58,31,144,31,82,31,76,31,220,31,111,31,85,31,118,31,145,31,178,31,53,31,215,31,245,31,240,31,6,31,103,31,103,30,152,31,152,30,57,31,207,31,252,31,216,31,220,31,162,31,179,31,66,31,179,31,229,31,200,31,240,31,240,30,240,29,240,28,112,31,163,31,135,31,101,31,101,30,101,29,101,28,25,31,37,31,91,31,173,31,173,30,83,31,70,31,74,31,246,31,140,31,140,30,39,31,39,30,15,31,102,31,87,31,219,31,90,31,90,30,63,31,120,31,120,30,75,31,175,31,28,31,79,31,79,30,79,29,75,31,80,31,205,31,68,31,1,31,225,31,155,31,181,31,136,31,221,31,62,31,125,31,154,31,174,31,160,31,74,31,188,31,192,31,155,31,157,31,203,31,112,31,112,30,179,31,186,31,117,31,117,30,4,31,167,31,14,31,176,31,225,31,225,30,125,31,240,31,175,31,25,31,25,30,192,31,194,31,162,31,168,31,109,31,43,31,161,31,66,31,9,31,59,31,195,31,233,31,44,31,92,31,131,31,92,31,155,31,43,31,44,31,186,31,113,31,113,30,169,31,172,31,116,31,43,31,186,31,132,31,251,31,251,30,175,31,136,31,134,31,218,31,163,31,184,31,216,31,209,31,209,30,32,31,163,31,37,31,72,31,22,31,64,31,64,30,64,29,240,31,154,31,155,31,155,30,155,29,91,31,72,31,106,31,112,31,198,31,198,30,94,31,182,31,70,31,117,31,183,31,66,31,29,31,130,31,232,31,194,31,194,30,177,31,204,31,109,31,130,31,130,30,124,31,9,31,9,30,146,31,112,31,112,30,119,31,115,31,179,31,179,30,145,31,219,31,22,31,96,31,123,31,201,31,126,31,186,31,110,31,79,31,79,30,79,29,165,31,13,31,58,31,199,31,199,30,199,29,199,28,199,27,194,31,194,30,194,29,83,31,90,31,174,31,76,31,49,31,245,31,245,30,40,31,103,31,103,30,103,29,103,28,156,31,151,31,92,31,227,31,227,30,229,31,139,31,92,31,162,31,162,30,4,31,104,31,163,31,163,30,3,31,228,31,150,31,150,30,213,31,20,31,6,31,159,31,159,30,181,31,51,31,51,30,52,31,42,31,30,31,49,31,15,31,235,31,17,31,39,31,229,31,140,31,101,31,107,31,107,30,232,31,100,31,100,30,57,31,57,30,121,31,210,31,76,31,168,31,225,31,107,31,190,31,10,31,115,31,74,31,248,31,152,31,45,31,121,31,121,30,121,29,187,31,4,31,75,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
