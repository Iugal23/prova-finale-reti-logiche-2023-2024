-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_85 is
end project_tb_85;

architecture project_tb_arch_85 of project_tb_85 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 745;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (108,0,250,0,96,0,191,0,196,0,106,0,0,0,225,0,158,0,0,0,139,0,24,0,0,0,80,0,154,0,212,0,177,0,16,0,0,0,230,0,19,0,123,0,65,0,253,0,14,0,0,0,0,0,211,0,243,0,64,0,3,0,133,0,41,0,6,0,68,0,126,0,81,0,40,0,0,0,72,0,240,0,193,0,179,0,95,0,0,0,137,0,38,0,198,0,25,0,112,0,230,0,104,0,115,0,0,0,48,0,0,0,226,0,0,0,229,0,254,0,106,0,0,0,19,0,207,0,3,0,6,0,0,0,26,0,17,0,137,0,104,0,57,0,170,0,90,0,0,0,188,0,244,0,207,0,0,0,87,0,0,0,103,0,244,0,91,0,80,0,245,0,228,0,17,0,113,0,78,0,127,0,73,0,150,0,199,0,42,0,192,0,66,0,129,0,0,0,214,0,205,0,152,0,62,0,149,0,169,0,97,0,0,0,0,0,179,0,179,0,147,0,175,0,138,0,231,0,73,0,242,0,52,0,0,0,0,0,254,0,0,0,144,0,0,0,0,0,192,0,35,0,212,0,0,0,0,0,27,0,107,0,175,0,67,0,0,0,223,0,0,0,74,0,83,0,97,0,25,0,62,0,110,0,0,0,60,0,212,0,103,0,203,0,69,0,72,0,162,0,0,0,169,0,214,0,211,0,138,0,218,0,193,0,205,0,0,0,159,0,104,0,107,0,149,0,10,0,250,0,29,0,241,0,243,0,5,0,8,0,0,0,7,0,87,0,0,0,122,0,142,0,139,0,142,0,252,0,238,0,193,0,116,0,15,0,47,0,151,0,0,0,213,0,22,0,193,0,205,0,67,0,57,0,71,0,8,0,59,0,0,0,0,0,212,0,168,0,253,0,186,0,29,0,0,0,127,0,178,0,1,0,199,0,103,0,0,0,132,0,0,0,157,0,0,0,3,0,233,0,134,0,228,0,0,0,161,0,164,0,104,0,233,0,244,0,89,0,219,0,233,0,35,0,183,0,94,0,74,0,154,0,0,0,0,0,0,0,56,0,230,0,5,0,203,0,185,0,27,0,37,0,0,0,171,0,0,0,53,0,0,0,24,0,217,0,35,0,25,0,136,0,35,0,167,0,21,0,209,0,238,0,34,0,188,0,148,0,0,0,0,0,233,0,175,0,0,0,103,0,0,0,22,0,111,0,139,0,188,0,50,0,202,0,163,0,69,0,29,0,234,0,91,0,129,0,243,0,0,0,128,0,80,0,137,0,57,0,201,0,154,0,183,0,31,0,0,0,0,0,114,0,163,0,107,0,230,0,0,0,236,0,158,0,0,0,47,0,166,0,0,0,12,0,52,0,103,0,194,0,0,0,61,0,0,0,162,0,185,0,29,0,0,0,56,0,205,0,17,0,241,0,5,0,88,0,71,0,0,0,156,0,255,0,0,0,20,0,105,0,0,0,0,0,254,0,7,0,69,0,33,0,218,0,9,0,132,0,110,0,0,0,59,0,71,0,234,0,240,0,218,0,46,0,0,0,182,0,0,0,249,0,209,0,244,0,172,0,18,0,0,0,11,0,105,0,48,0,0,0,108,0,75,0,176,0,231,0,128,0,0,0,141,0,212,0,106,0,200,0,40,0,219,0,180,0,169,0,122,0,79,0,57,0,204,0,25,0,171,0,0,0,223,0,0,0,74,0,57,0,119,0,63,0,50,0,26,0,28,0,81,0,130,0,127,0,130,0,214,0,134,0,134,0,165,0,176,0,0,0,151,0,148,0,0,0,0,0,111,0,210,0,68,0,0,0,131,0,243,0,99,0,0,0,0,0,183,0,68,0,140,0,52,0,230,0,0,0,107,0,0,0,79,0,52,0,194,0,189,0,0,0,149,0,113,0,193,0,0,0,211,0,183,0,98,0,55,0,170,0,8,0,93,0,53,0,238,0,79,0,135,0,127,0,95,0,114,0,206,0,0,0,0,0,0,0,0,0,191,0,135,0,148,0,150,0,189,0,76,0,205,0,131,0,62,0,196,0,196,0,0,0,83,0,157,0,54,0,20,0,29,0,197,0,108,0,255,0,33,0,198,0,136,0,179,0,0,0,20,0,76,0,195,0,233,0,93,0,203,0,0,0,176,0,21,0,0,0,222,0,66,0,236,0,253,0,204,0,198,0,42,0,0,0,91,0,194,0,113,0,143,0,46,0,71,0,135,0,222,0,103,0,39,0,32,0,133,0,197,0,226,0,0,0,0,0,236,0,0,0,0,0,0,0,114,0,0,0,245,0,199,0,31,0,212,0,152,0,204,0,110,0,138,0,0,0,162,0,220,0,36,0,96,0,115,0,94,0,0,0,72,0,35,0,0,0,119,0,100,0,235,0,209,0,233,0,0,0,11,0,0,0,0,0,150,0,231,0,161,0,0,0,0,0,71,0,207,0,221,0,195,0,216,0,242,0,87,0,141,0,162,0,0,0,89,0,0,0,30,0,87,0,2,0,0,0,212,0,179,0,216,0,90,0,47,0,214,0,111,0,144,0,0,0,75,0,67,0,135,0,88,0,2,0,219,0,60,0,118,0,123,0,230,0,169,0,235,0,0,0,241,0,173,0,238,0,218,0,138,0,172,0,92,0,255,0,0,0,191,0,0,0,0,0,0,0,0,0,0,0,35,0,140,0,3,0,152,0,17,0,0,0,169,0,67,0,139,0,191,0,249,0,169,0,0,0,192,0,38,0,65,0,201,0,100,0,11,0,85,0,28,0,34,0,180,0,190,0,235,0,134,0,124,0,0,0,177,0,236,0,52,0,93,0,227,0,187,0,127,0,64,0,155,0,0,0,35,0,131,0,195,0,7,0,51,0,241,0,27,0,0,0,158,0,174,0,21,0,234,0,13,0,112,0,181,0,3,0,0,0,44,0,13,0,0,0,0,0,0,0,211,0,176,0,0,0,175,0,253,0,212,0,30,0,169,0,2,0,65,0,109,0,239,0,0,0,114,0,70,0,26,0,184,0,245,0,0,0,147,0,136,0,168,0,24,0,221,0,208,0,39,0,77,0,98,0,176,0,100,0,197,0,10,0,179,0,226,0,145,0,7,0,0,0,216,0,62,0,103,0,110,0,0,0,2,0,119,0,118,0,173,0,76,0,200,0,6,0,28,0,0,0,199,0,0,0,28,0,25,0,26,0,194,0,64,0,0,0,195,0,86,0,83,0,134,0,17,0,221,0,179,0,156,0,248,0,26,0,201,0,182,0,150,0,179,0,50,0,140,0,0,0,81,0,56,0,202,0,241,0,85,0,0,0,232,0,233,0,59,0,153,0,0,0,200,0,106,0,0,0);
signal scenario_full  : scenario_type := (108,31,250,31,96,31,191,31,196,31,106,31,106,30,225,31,158,31,158,30,139,31,24,31,24,30,80,31,154,31,212,31,177,31,16,31,16,30,230,31,19,31,123,31,65,31,253,31,14,31,14,30,14,29,211,31,243,31,64,31,3,31,133,31,41,31,6,31,68,31,126,31,81,31,40,31,40,30,72,31,240,31,193,31,179,31,95,31,95,30,137,31,38,31,198,31,25,31,112,31,230,31,104,31,115,31,115,30,48,31,48,30,226,31,226,30,229,31,254,31,106,31,106,30,19,31,207,31,3,31,6,31,6,30,26,31,17,31,137,31,104,31,57,31,170,31,90,31,90,30,188,31,244,31,207,31,207,30,87,31,87,30,103,31,244,31,91,31,80,31,245,31,228,31,17,31,113,31,78,31,127,31,73,31,150,31,199,31,42,31,192,31,66,31,129,31,129,30,214,31,205,31,152,31,62,31,149,31,169,31,97,31,97,30,97,29,179,31,179,31,147,31,175,31,138,31,231,31,73,31,242,31,52,31,52,30,52,29,254,31,254,30,144,31,144,30,144,29,192,31,35,31,212,31,212,30,212,29,27,31,107,31,175,31,67,31,67,30,223,31,223,30,74,31,83,31,97,31,25,31,62,31,110,31,110,30,60,31,212,31,103,31,203,31,69,31,72,31,162,31,162,30,169,31,214,31,211,31,138,31,218,31,193,31,205,31,205,30,159,31,104,31,107,31,149,31,10,31,250,31,29,31,241,31,243,31,5,31,8,31,8,30,7,31,87,31,87,30,122,31,142,31,139,31,142,31,252,31,238,31,193,31,116,31,15,31,47,31,151,31,151,30,213,31,22,31,193,31,205,31,67,31,57,31,71,31,8,31,59,31,59,30,59,29,212,31,168,31,253,31,186,31,29,31,29,30,127,31,178,31,1,31,199,31,103,31,103,30,132,31,132,30,157,31,157,30,3,31,233,31,134,31,228,31,228,30,161,31,164,31,104,31,233,31,244,31,89,31,219,31,233,31,35,31,183,31,94,31,74,31,154,31,154,30,154,29,154,28,56,31,230,31,5,31,203,31,185,31,27,31,37,31,37,30,171,31,171,30,53,31,53,30,24,31,217,31,35,31,25,31,136,31,35,31,167,31,21,31,209,31,238,31,34,31,188,31,148,31,148,30,148,29,233,31,175,31,175,30,103,31,103,30,22,31,111,31,139,31,188,31,50,31,202,31,163,31,69,31,29,31,234,31,91,31,129,31,243,31,243,30,128,31,80,31,137,31,57,31,201,31,154,31,183,31,31,31,31,30,31,29,114,31,163,31,107,31,230,31,230,30,236,31,158,31,158,30,47,31,166,31,166,30,12,31,52,31,103,31,194,31,194,30,61,31,61,30,162,31,185,31,29,31,29,30,56,31,205,31,17,31,241,31,5,31,88,31,71,31,71,30,156,31,255,31,255,30,20,31,105,31,105,30,105,29,254,31,7,31,69,31,33,31,218,31,9,31,132,31,110,31,110,30,59,31,71,31,234,31,240,31,218,31,46,31,46,30,182,31,182,30,249,31,209,31,244,31,172,31,18,31,18,30,11,31,105,31,48,31,48,30,108,31,75,31,176,31,231,31,128,31,128,30,141,31,212,31,106,31,200,31,40,31,219,31,180,31,169,31,122,31,79,31,57,31,204,31,25,31,171,31,171,30,223,31,223,30,74,31,57,31,119,31,63,31,50,31,26,31,28,31,81,31,130,31,127,31,130,31,214,31,134,31,134,31,165,31,176,31,176,30,151,31,148,31,148,30,148,29,111,31,210,31,68,31,68,30,131,31,243,31,99,31,99,30,99,29,183,31,68,31,140,31,52,31,230,31,230,30,107,31,107,30,79,31,52,31,194,31,189,31,189,30,149,31,113,31,193,31,193,30,211,31,183,31,98,31,55,31,170,31,8,31,93,31,53,31,238,31,79,31,135,31,127,31,95,31,114,31,206,31,206,30,206,29,206,28,206,27,191,31,135,31,148,31,150,31,189,31,76,31,205,31,131,31,62,31,196,31,196,31,196,30,83,31,157,31,54,31,20,31,29,31,197,31,108,31,255,31,33,31,198,31,136,31,179,31,179,30,20,31,76,31,195,31,233,31,93,31,203,31,203,30,176,31,21,31,21,30,222,31,66,31,236,31,253,31,204,31,198,31,42,31,42,30,91,31,194,31,113,31,143,31,46,31,71,31,135,31,222,31,103,31,39,31,32,31,133,31,197,31,226,31,226,30,226,29,236,31,236,30,236,29,236,28,114,31,114,30,245,31,199,31,31,31,212,31,152,31,204,31,110,31,138,31,138,30,162,31,220,31,36,31,96,31,115,31,94,31,94,30,72,31,35,31,35,30,119,31,100,31,235,31,209,31,233,31,233,30,11,31,11,30,11,29,150,31,231,31,161,31,161,30,161,29,71,31,207,31,221,31,195,31,216,31,242,31,87,31,141,31,162,31,162,30,89,31,89,30,30,31,87,31,2,31,2,30,212,31,179,31,216,31,90,31,47,31,214,31,111,31,144,31,144,30,75,31,67,31,135,31,88,31,2,31,219,31,60,31,118,31,123,31,230,31,169,31,235,31,235,30,241,31,173,31,238,31,218,31,138,31,172,31,92,31,255,31,255,30,191,31,191,30,191,29,191,28,191,27,191,26,35,31,140,31,3,31,152,31,17,31,17,30,169,31,67,31,139,31,191,31,249,31,169,31,169,30,192,31,38,31,65,31,201,31,100,31,11,31,85,31,28,31,34,31,180,31,190,31,235,31,134,31,124,31,124,30,177,31,236,31,52,31,93,31,227,31,187,31,127,31,64,31,155,31,155,30,35,31,131,31,195,31,7,31,51,31,241,31,27,31,27,30,158,31,174,31,21,31,234,31,13,31,112,31,181,31,3,31,3,30,44,31,13,31,13,30,13,29,13,28,211,31,176,31,176,30,175,31,253,31,212,31,30,31,169,31,2,31,65,31,109,31,239,31,239,30,114,31,70,31,26,31,184,31,245,31,245,30,147,31,136,31,168,31,24,31,221,31,208,31,39,31,77,31,98,31,176,31,100,31,197,31,10,31,179,31,226,31,145,31,7,31,7,30,216,31,62,31,103,31,110,31,110,30,2,31,119,31,118,31,173,31,76,31,200,31,6,31,28,31,28,30,199,31,199,30,28,31,25,31,26,31,194,31,64,31,64,30,195,31,86,31,83,31,134,31,17,31,221,31,179,31,156,31,248,31,26,31,201,31,182,31,150,31,179,31,50,31,140,31,140,30,81,31,56,31,202,31,241,31,85,31,85,30,232,31,233,31,59,31,153,31,153,30,200,31,106,31,106,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
