-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 732;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (141,0,61,0,223,0,63,0,47,0,199,0,151,0,0,0,50,0,151,0,33,0,50,0,59,0,104,0,156,0,143,0,12,0,215,0,121,0,0,0,0,0,61,0,187,0,42,0,242,0,0,0,202,0,0,0,254,0,0,0,0,0,19,0,151,0,245,0,0,0,126,0,64,0,28,0,0,0,11,0,138,0,212,0,202,0,173,0,104,0,153,0,213,0,0,0,225,0,116,0,173,0,16,0,1,0,69,0,227,0,176,0,113,0,0,0,177,0,208,0,228,0,96,0,168,0,112,0,32,0,19,0,100,0,83,0,140,0,149,0,51,0,0,0,0,0,161,0,121,0,50,0,107,0,0,0,185,0,0,0,165,0,0,0,164,0,165,0,0,0,16,0,11,0,176,0,81,0,78,0,0,0,199,0,191,0,0,0,0,0,0,0,0,0,0,0,140,0,0,0,40,0,14,0,182,0,142,0,0,0,37,0,187,0,196,0,174,0,12,0,209,0,0,0,103,0,170,0,173,0,205,0,53,0,0,0,227,0,86,0,247,0,170,0,116,0,232,0,138,0,253,0,74,0,0,0,195,0,240,0,104,0,0,0,192,0,1,0,92,0,174,0,0,0,92,0,55,0,0,0,54,0,0,0,0,0,0,0,36,0,46,0,0,0,72,0,65,0,0,0,0,0,0,0,167,0,5,0,130,0,188,0,115,0,190,0,150,0,188,0,194,0,50,0,99,0,242,0,46,0,0,0,16,0,0,0,0,0,167,0,198,0,182,0,15,0,245,0,65,0,155,0,113,0,0,0,86,0,83,0,173,0,0,0,39,0,188,0,95,0,91,0,81,0,155,0,194,0,133,0,34,0,245,0,0,0,80,0,200,0,167,0,248,0,0,0,0,0,0,0,50,0,115,0,64,0,232,0,192,0,137,0,129,0,0,0,0,0,0,0,42,0,62,0,0,0,0,0,158,0,216,0,90,0,238,0,0,0,225,0,217,0,0,0,0,0,8,0,161,0,102,0,108,0,172,0,0,0,109,0,100,0,46,0,90,0,200,0,29,0,254,0,0,0,65,0,28,0,140,0,101,0,143,0,0,0,32,0,57,0,254,0,49,0,192,0,148,0,0,0,86,0,0,0,0,0,171,0,70,0,51,0,59,0,76,0,216,0,162,0,0,0,187,0,0,0,225,0,37,0,216,0,176,0,0,0,217,0,123,0,0,0,0,0,78,0,0,0,133,0,125,0,34,0,217,0,0,0,246,0,63,0,222,0,244,0,0,0,0,0,0,0,0,0,105,0,136,0,0,0,135,0,155,0,0,0,175,0,143,0,67,0,192,0,0,0,119,0,168,0,0,0,17,0,9,0,205,0,0,0,143,0,134,0,100,0,46,0,252,0,10,0,227,0,115,0,251,0,127,0,144,0,39,0,129,0,90,0,22,0,0,0,108,0,68,0,233,0,249,0,156,0,250,0,235,0,12,0,47,0,0,0,140,0,162,0,96,0,54,0,83,0,47,0,247,0,169,0,150,0,233,0,223,0,104,0,47,0,50,0,43,0,156,0,13,0,106,0,0,0,186,0,200,0,92,0,153,0,0,0,231,0,140,0,0,0,102,0,37,0,0,0,0,0,0,0,0,0,9,0,86,0,244,0,128,0,201,0,0,0,151,0,26,0,39,0,138,0,212,0,38,0,143,0,51,0,0,0,98,0,63,0,101,0,12,0,0,0,0,0,255,0,201,0,25,0,125,0,0,0,0,0,110,0,140,0,6,0,58,0,0,0,60,0,114,0,227,0,221,0,205,0,59,0,148,0,70,0,140,0,215,0,148,0,0,0,255,0,0,0,103,0,145,0,58,0,176,0,2,0,85,0,212,0,174,0,34,0,77,0,33,0,20,0,137,0,193,0,136,0,250,0,171,0,117,0,0,0,212,0,0,0,0,0,0,0,16,0,129,0,41,0,194,0,40,0,0,0,204,0,167,0,196,0,0,0,49,0,0,0,0,0,44,0,31,0,0,0,129,0,176,0,223,0,208,0,63,0,249,0,0,0,28,0,222,0,186,0,27,0,207,0,0,0,0,0,230,0,0,0,59,0,248,0,158,0,108,0,28,0,154,0,43,0,96,0,101,0,0,0,212,0,6,0,158,0,180,0,140,0,38,0,0,0,125,0,45,0,0,0,214,0,239,0,157,0,11,0,193,0,0,0,0,0,196,0,87,0,185,0,0,0,27,0,213,0,35,0,130,0,20,0,237,0,179,0,254,0,0,0,160,0,0,0,158,0,148,0,142,0,148,0,0,0,75,0,221,0,72,0,194,0,234,0,86,0,51,0,0,0,27,0,40,0,204,0,225,0,91,0,75,0,44,0,196,0,0,0,96,0,42,0,101,0,197,0,117,0,197,0,146,0,224,0,0,0,17,0,137,0,63,0,110,0,29,0,142,0,228,0,242,0,0,0,0,0,198,0,157,0,193,0,54,0,138,0,0,0,123,0,135,0,237,0,121,0,182,0,187,0,249,0,0,0,102,0,0,0,108,0,0,0,0,0,47,0,17,0,0,0,147,0,0,0,3,0,0,0,195,0,76,0,189,0,201,0,0,0,213,0,243,0,39,0,94,0,39,0,59,0,231,0,0,0,135,0,80,0,0,0,59,0,123,0,149,0,0,0,252,0,0,0,0,0,76,0,103,0,39,0,0,0,105,0,26,0,104,0,145,0,251,0,116,0,129,0,71,0,69,0,250,0,40,0,71,0,125,0,0,0,50,0,0,0,247,0,89,0,142,0,10,0,240,0,0,0,0,0,56,0,0,0,125,0,15,0,137,0,0,0,1,0,232,0,0,0,0,0,186,0,0,0,42,0,0,0,40,0,0,0,216,0,223,0,234,0,214,0,176,0,0,0,6,0,227,0,229,0,126,0,0,0,50,0,0,0,0,0,200,0,0,0,107,0,208,0,53,0,151,0,139,0,0,0,0,0,41,0,9,0,40,0,0,0,0,0,64,0,32,0,237,0,117,0,238,0,135,0,35,0,88,0,0,0,28,0,224,0,5,0,79,0,203,0,169,0,10,0,20,0,121,0,116,0,64,0,161,0,37,0,119,0,167,0,226,0,122,0,0,0,65,0,209,0,47,0,56,0,63,0,0,0,80,0,127,0,148,0,0,0,0,0,26,0,41,0,195,0,11,0,181,0,0,0,170,0,138,0,247,0,45,0,0,0,0,0,0,0,190,0,0,0,82,0,0,0,158,0,240,0,167,0,106,0,92,0,92,0,0,0,0,0,173,0);
signal scenario_full  : scenario_type := (141,31,61,31,223,31,63,31,47,31,199,31,151,31,151,30,50,31,151,31,33,31,50,31,59,31,104,31,156,31,143,31,12,31,215,31,121,31,121,30,121,29,61,31,187,31,42,31,242,31,242,30,202,31,202,30,254,31,254,30,254,29,19,31,151,31,245,31,245,30,126,31,64,31,28,31,28,30,11,31,138,31,212,31,202,31,173,31,104,31,153,31,213,31,213,30,225,31,116,31,173,31,16,31,1,31,69,31,227,31,176,31,113,31,113,30,177,31,208,31,228,31,96,31,168,31,112,31,32,31,19,31,100,31,83,31,140,31,149,31,51,31,51,30,51,29,161,31,121,31,50,31,107,31,107,30,185,31,185,30,165,31,165,30,164,31,165,31,165,30,16,31,11,31,176,31,81,31,78,31,78,30,199,31,191,31,191,30,191,29,191,28,191,27,191,26,140,31,140,30,40,31,14,31,182,31,142,31,142,30,37,31,187,31,196,31,174,31,12,31,209,31,209,30,103,31,170,31,173,31,205,31,53,31,53,30,227,31,86,31,247,31,170,31,116,31,232,31,138,31,253,31,74,31,74,30,195,31,240,31,104,31,104,30,192,31,1,31,92,31,174,31,174,30,92,31,55,31,55,30,54,31,54,30,54,29,54,28,36,31,46,31,46,30,72,31,65,31,65,30,65,29,65,28,167,31,5,31,130,31,188,31,115,31,190,31,150,31,188,31,194,31,50,31,99,31,242,31,46,31,46,30,16,31,16,30,16,29,167,31,198,31,182,31,15,31,245,31,65,31,155,31,113,31,113,30,86,31,83,31,173,31,173,30,39,31,188,31,95,31,91,31,81,31,155,31,194,31,133,31,34,31,245,31,245,30,80,31,200,31,167,31,248,31,248,30,248,29,248,28,50,31,115,31,64,31,232,31,192,31,137,31,129,31,129,30,129,29,129,28,42,31,62,31,62,30,62,29,158,31,216,31,90,31,238,31,238,30,225,31,217,31,217,30,217,29,8,31,161,31,102,31,108,31,172,31,172,30,109,31,100,31,46,31,90,31,200,31,29,31,254,31,254,30,65,31,28,31,140,31,101,31,143,31,143,30,32,31,57,31,254,31,49,31,192,31,148,31,148,30,86,31,86,30,86,29,171,31,70,31,51,31,59,31,76,31,216,31,162,31,162,30,187,31,187,30,225,31,37,31,216,31,176,31,176,30,217,31,123,31,123,30,123,29,78,31,78,30,133,31,125,31,34,31,217,31,217,30,246,31,63,31,222,31,244,31,244,30,244,29,244,28,244,27,105,31,136,31,136,30,135,31,155,31,155,30,175,31,143,31,67,31,192,31,192,30,119,31,168,31,168,30,17,31,9,31,205,31,205,30,143,31,134,31,100,31,46,31,252,31,10,31,227,31,115,31,251,31,127,31,144,31,39,31,129,31,90,31,22,31,22,30,108,31,68,31,233,31,249,31,156,31,250,31,235,31,12,31,47,31,47,30,140,31,162,31,96,31,54,31,83,31,47,31,247,31,169,31,150,31,233,31,223,31,104,31,47,31,50,31,43,31,156,31,13,31,106,31,106,30,186,31,200,31,92,31,153,31,153,30,231,31,140,31,140,30,102,31,37,31,37,30,37,29,37,28,37,27,9,31,86,31,244,31,128,31,201,31,201,30,151,31,26,31,39,31,138,31,212,31,38,31,143,31,51,31,51,30,98,31,63,31,101,31,12,31,12,30,12,29,255,31,201,31,25,31,125,31,125,30,125,29,110,31,140,31,6,31,58,31,58,30,60,31,114,31,227,31,221,31,205,31,59,31,148,31,70,31,140,31,215,31,148,31,148,30,255,31,255,30,103,31,145,31,58,31,176,31,2,31,85,31,212,31,174,31,34,31,77,31,33,31,20,31,137,31,193,31,136,31,250,31,171,31,117,31,117,30,212,31,212,30,212,29,212,28,16,31,129,31,41,31,194,31,40,31,40,30,204,31,167,31,196,31,196,30,49,31,49,30,49,29,44,31,31,31,31,30,129,31,176,31,223,31,208,31,63,31,249,31,249,30,28,31,222,31,186,31,27,31,207,31,207,30,207,29,230,31,230,30,59,31,248,31,158,31,108,31,28,31,154,31,43,31,96,31,101,31,101,30,212,31,6,31,158,31,180,31,140,31,38,31,38,30,125,31,45,31,45,30,214,31,239,31,157,31,11,31,193,31,193,30,193,29,196,31,87,31,185,31,185,30,27,31,213,31,35,31,130,31,20,31,237,31,179,31,254,31,254,30,160,31,160,30,158,31,148,31,142,31,148,31,148,30,75,31,221,31,72,31,194,31,234,31,86,31,51,31,51,30,27,31,40,31,204,31,225,31,91,31,75,31,44,31,196,31,196,30,96,31,42,31,101,31,197,31,117,31,197,31,146,31,224,31,224,30,17,31,137,31,63,31,110,31,29,31,142,31,228,31,242,31,242,30,242,29,198,31,157,31,193,31,54,31,138,31,138,30,123,31,135,31,237,31,121,31,182,31,187,31,249,31,249,30,102,31,102,30,108,31,108,30,108,29,47,31,17,31,17,30,147,31,147,30,3,31,3,30,195,31,76,31,189,31,201,31,201,30,213,31,243,31,39,31,94,31,39,31,59,31,231,31,231,30,135,31,80,31,80,30,59,31,123,31,149,31,149,30,252,31,252,30,252,29,76,31,103,31,39,31,39,30,105,31,26,31,104,31,145,31,251,31,116,31,129,31,71,31,69,31,250,31,40,31,71,31,125,31,125,30,50,31,50,30,247,31,89,31,142,31,10,31,240,31,240,30,240,29,56,31,56,30,125,31,15,31,137,31,137,30,1,31,232,31,232,30,232,29,186,31,186,30,42,31,42,30,40,31,40,30,216,31,223,31,234,31,214,31,176,31,176,30,6,31,227,31,229,31,126,31,126,30,50,31,50,30,50,29,200,31,200,30,107,31,208,31,53,31,151,31,139,31,139,30,139,29,41,31,9,31,40,31,40,30,40,29,64,31,32,31,237,31,117,31,238,31,135,31,35,31,88,31,88,30,28,31,224,31,5,31,79,31,203,31,169,31,10,31,20,31,121,31,116,31,64,31,161,31,37,31,119,31,167,31,226,31,122,31,122,30,65,31,209,31,47,31,56,31,63,31,63,30,80,31,127,31,148,31,148,30,148,29,26,31,41,31,195,31,11,31,181,31,181,30,170,31,138,31,247,31,45,31,45,30,45,29,45,28,190,31,190,30,82,31,82,30,158,31,240,31,167,31,106,31,92,31,92,31,92,30,92,29,173,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
