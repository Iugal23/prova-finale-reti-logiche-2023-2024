-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_0 is
end project_tb_0;

architecture project_tb_arch_0 of project_tb_0 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 877;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,112,0,74,0,175,0,195,0,134,0,252,0,179,0,143,0,0,0,243,0,166,0,0,0,217,0,228,0,0,0,36,0,103,0,0,0,0,0,83,0,1,0,33,0,46,0,245,0,0,0,0,0,0,0,150,0,209,0,0,0,70,0,0,0,54,0,133,0,30,0,218,0,81,0,170,0,242,0,218,0,100,0,185,0,204,0,251,0,212,0,206,0,251,0,0,0,238,0,180,0,227,0,0,0,93,0,239,0,0,0,26,0,225,0,161,0,119,0,140,0,50,0,0,0,139,0,0,0,242,0,0,0,152,0,0,0,137,0,33,0,150,0,0,0,154,0,52,0,27,0,135,0,214,0,0,0,0,0,188,0,249,0,0,0,166,0,0,0,161,0,7,0,172,0,172,0,127,0,98,0,26,0,193,0,0,0,182,0,0,0,100,0,250,0,247,0,34,0,0,0,120,0,221,0,28,0,31,0,63,0,91,0,234,0,112,0,0,0,90,0,54,0,158,0,199,0,170,0,0,0,115,0,166,0,172,0,0,0,10,0,41,0,56,0,211,0,212,0,187,0,0,0,162,0,142,0,119,0,52,0,0,0,23,0,181,0,42,0,174,0,0,0,218,0,0,0,119,0,140,0,103,0,36,0,0,0,47,0,0,0,0,0,125,0,235,0,16,0,47,0,0,0,10,0,76,0,0,0,13,0,155,0,0,0,96,0,120,0,232,0,59,0,0,0,214,0,116,0,46,0,64,0,119,0,66,0,208,0,0,0,11,0,252,0,160,0,0,0,94,0,56,0,0,0,0,0,193,0,0,0,0,0,0,0,214,0,0,0,168,0,49,0,21,0,197,0,0,0,157,0,21,0,0,0,253,0,113,0,17,0,222,0,65,0,154,0,116,0,157,0,170,0,18,0,0,0,0,0,109,0,248,0,237,0,151,0,0,0,72,0,154,0,102,0,131,0,0,0,178,0,13,0,174,0,124,0,0,0,117,0,208,0,253,0,5,0,6,0,46,0,0,0,115,0,222,0,0,0,42,0,21,0,75,0,207,0,115,0,107,0,19,0,0,0,241,0,105,0,103,0,12,0,158,0,0,0,96,0,0,0,3,0,62,0,232,0,32,0,77,0,0,0,0,0,169,0,85,0,0,0,144,0,200,0,56,0,0,0,115,0,232,0,89,0,43,0,7,0,109,0,199,0,116,0,145,0,70,0,94,0,164,0,96,0,246,0,249,0,108,0,0,0,123,0,152,0,19,0,129,0,204,0,250,0,24,0,240,0,148,0,5,0,148,0,27,0,0,0,0,0,134,0,45,0,146,0,0,0,163,0,0,0,0,0,159,0,144,0,255,0,100,0,135,0,252,0,86,0,0,0,0,0,0,0,0,0,20,0,54,0,45,0,151,0,161,0,105,0,154,0,203,0,253,0,0,0,0,0,76,0,197,0,0,0,227,0,163,0,203,0,140,0,12,0,181,0,1,0,195,0,155,0,0,0,57,0,134,0,65,0,0,0,234,0,83,0,229,0,47,0,137,0,241,0,0,0,114,0,0,0,66,0,70,0,146,0,174,0,211,0,0,0,136,0,0,0,0,0,211,0,0,0,0,0,166,0,188,0,213,0,23,0,49,0,155,0,194,0,64,0,0,0,133,0,223,0,253,0,119,0,105,0,0,0,155,0,220,0,106,0,152,0,31,0,130,0,7,0,245,0,0,0,0,0,0,0,229,0,0,0,135,0,92,0,0,0,109,0,251,0,243,0,155,0,122,0,167,0,252,0,49,0,102,0,84,0,86,0,241,0,238,0,0,0,47,0,54,0,205,0,0,0,13,0,222,0,0,0,195,0,104,0,116,0,75,0,0,0,93,0,214,0,76,0,223,0,115,0,69,0,143,0,236,0,0,0,0,0,0,0,179,0,146,0,102,0,0,0,222,0,73,0,228,0,15,0,87,0,3,0,80,0,215,0,76,0,248,0,0,0,161,0,233,0,1,0,249,0,0,0,195,0,0,0,9,0,185,0,33,0,0,0,203,0,0,0,233,0,44,0,216,0,29,0,150,0,158,0,212,0,0,0,26,0,42,0,0,0,9,0,157,0,0,0,146,0,42,0,43,0,250,0,5,0,0,0,35,0,0,0,202,0,147,0,209,0,174,0,130,0,130,0,227,0,120,0,198,0,133,0,112,0,0,0,16,0,183,0,236,0,157,0,249,0,183,0,142,0,80,0,0,0,44,0,0,0,0,0,97,0,0,0,0,0,0,0,35,0,66,0,88,0,0,0,70,0,165,0,104,0,104,0,198,0,0,0,138,0,158,0,104,0,0,0,0,0,0,0,172,0,0,0,14,0,83,0,0,0,176,0,193,0,0,0,0,0,109,0,19,0,163,0,0,0,40,0,242,0,3,0,54,0,52,0,41,0,231,0,243,0,178,0,157,0,0,0,98,0,127,0,225,0,149,0,0,0,223,0,153,0,46,0,204,0,0,0,221,0,40,0,128,0,82,0,0,0,54,0,0,0,79,0,0,0,69,0,126,0,221,0,115,0,52,0,113,0,165,0,42,0,107,0,114,0,239,0,240,0,157,0,0,0,88,0,0,0,19,0,37,0,0,0,154,0,127,0,163,0,172,0,172,0,0,0,0,0,151,0,163,0,137,0,231,0,0,0,226,0,0,0,137,0,15,0,0,0,255,0,0,0,85,0,22,0,205,0,195,0,8,0,228,0,52,0,48,0,233,0,0,0,91,0,253,0,0,0,46,0,0,0,33,0,0,0,44,0,4,0,0,0,0,0,83,0,142,0,76,0,0,0,0,0,0,0,0,0,196,0,0,0,245,0,93,0,97,0,32,0,37,0,0,0,126,0,212,0,249,0,21,0,84,0,123,0,228,0,219,0,0,0,172,0,75,0,12,0,118,0,0,0,49,0,103,0,0,0,0,0,187,0,250,0,227,0,0,0,16,0,57,0,12,0,0,0,91,0,70,0,170,0,229,0,243,0,142,0,0,0,64,0,97,0,104,0,87,0,150,0,25,0,109,0,119,0,0,0,233,0,145,0,0,0,0,0,227,0,44,0,207,0,225,0,74,0,0,0,194,0,0,0,0,0,64,0,104,0,158,0,67,0,29,0,218,0,7,0,42,0,0,0,25,0,155,0,222,0,128,0,221,0,79,0,91,0,0,0,0,0,255,0,91,0,10,0,178,0,150,0,37,0,0,0,153,0,49,0,182,0,70,0,67,0,0,0,151,0,237,0,127,0,1,0,91,0,28,0,42,0,60,0,145,0,157,0,95,0,140,0,15,0,221,0,137,0,255,0,232,0,120,0,36,0,93,0,133,0,28,0,82,0,193,0,45,0,97,0,162,0,0,0,155,0,253,0,124,0,232,0,57,0,0,0,65,0,36,0,248,0,125,0,154,0,149,0,204,0,0,0,252,0,157,0,232,0,150,0,6,0,0,0,0,0,115,0,155,0,118,0,89,0,155,0,145,0,242,0,193,0,174,0,156,0,196,0,26,0,249,0,0,0,26,0,104,0,0,0,28,0,0,0,155,0,164,0,128,0,252,0,100,0,209,0,0,0,194,0,135,0,247,0,247,0,49,0,186,0,121,0,100,0,63,0,0,0,15,0,175,0,0,0,78,0,229,0,113,0,156,0,48,0,65,0,0,0,99,0,241,0,178,0,0,0,218,0,41,0,85,0,0,0,0,0,0,0,165,0,0,0,158,0,141,0,0,0,18,0,231,0,0,0,186,0,0,0,0,0,69,0,232,0,0,0,188,0,93,0,2,0,94,0,0,0,72,0,254,0,0,0,247,0,53,0,76,0,109,0,107,0,0,0,120,0,175,0,0,0,231,0,71,0,3,0,0,0,175,0,174,0,134,0,139,0,12,0,30,0,99,0,49,0,249,0,0,0,150,0,163,0,27,0,43,0);
signal scenario_full  : scenario_type := (6,31,112,31,74,31,175,31,195,31,134,31,252,31,179,31,143,31,143,30,243,31,166,31,166,30,217,31,228,31,228,30,36,31,103,31,103,30,103,29,83,31,1,31,33,31,46,31,245,31,245,30,245,29,245,28,150,31,209,31,209,30,70,31,70,30,54,31,133,31,30,31,218,31,81,31,170,31,242,31,218,31,100,31,185,31,204,31,251,31,212,31,206,31,251,31,251,30,238,31,180,31,227,31,227,30,93,31,239,31,239,30,26,31,225,31,161,31,119,31,140,31,50,31,50,30,139,31,139,30,242,31,242,30,152,31,152,30,137,31,33,31,150,31,150,30,154,31,52,31,27,31,135,31,214,31,214,30,214,29,188,31,249,31,249,30,166,31,166,30,161,31,7,31,172,31,172,31,127,31,98,31,26,31,193,31,193,30,182,31,182,30,100,31,250,31,247,31,34,31,34,30,120,31,221,31,28,31,31,31,63,31,91,31,234,31,112,31,112,30,90,31,54,31,158,31,199,31,170,31,170,30,115,31,166,31,172,31,172,30,10,31,41,31,56,31,211,31,212,31,187,31,187,30,162,31,142,31,119,31,52,31,52,30,23,31,181,31,42,31,174,31,174,30,218,31,218,30,119,31,140,31,103,31,36,31,36,30,47,31,47,30,47,29,125,31,235,31,16,31,47,31,47,30,10,31,76,31,76,30,13,31,155,31,155,30,96,31,120,31,232,31,59,31,59,30,214,31,116,31,46,31,64,31,119,31,66,31,208,31,208,30,11,31,252,31,160,31,160,30,94,31,56,31,56,30,56,29,193,31,193,30,193,29,193,28,214,31,214,30,168,31,49,31,21,31,197,31,197,30,157,31,21,31,21,30,253,31,113,31,17,31,222,31,65,31,154,31,116,31,157,31,170,31,18,31,18,30,18,29,109,31,248,31,237,31,151,31,151,30,72,31,154,31,102,31,131,31,131,30,178,31,13,31,174,31,124,31,124,30,117,31,208,31,253,31,5,31,6,31,46,31,46,30,115,31,222,31,222,30,42,31,21,31,75,31,207,31,115,31,107,31,19,31,19,30,241,31,105,31,103,31,12,31,158,31,158,30,96,31,96,30,3,31,62,31,232,31,32,31,77,31,77,30,77,29,169,31,85,31,85,30,144,31,200,31,56,31,56,30,115,31,232,31,89,31,43,31,7,31,109,31,199,31,116,31,145,31,70,31,94,31,164,31,96,31,246,31,249,31,108,31,108,30,123,31,152,31,19,31,129,31,204,31,250,31,24,31,240,31,148,31,5,31,148,31,27,31,27,30,27,29,134,31,45,31,146,31,146,30,163,31,163,30,163,29,159,31,144,31,255,31,100,31,135,31,252,31,86,31,86,30,86,29,86,28,86,27,20,31,54,31,45,31,151,31,161,31,105,31,154,31,203,31,253,31,253,30,253,29,76,31,197,31,197,30,227,31,163,31,203,31,140,31,12,31,181,31,1,31,195,31,155,31,155,30,57,31,134,31,65,31,65,30,234,31,83,31,229,31,47,31,137,31,241,31,241,30,114,31,114,30,66,31,70,31,146,31,174,31,211,31,211,30,136,31,136,30,136,29,211,31,211,30,211,29,166,31,188,31,213,31,23,31,49,31,155,31,194,31,64,31,64,30,133,31,223,31,253,31,119,31,105,31,105,30,155,31,220,31,106,31,152,31,31,31,130,31,7,31,245,31,245,30,245,29,245,28,229,31,229,30,135,31,92,31,92,30,109,31,251,31,243,31,155,31,122,31,167,31,252,31,49,31,102,31,84,31,86,31,241,31,238,31,238,30,47,31,54,31,205,31,205,30,13,31,222,31,222,30,195,31,104,31,116,31,75,31,75,30,93,31,214,31,76,31,223,31,115,31,69,31,143,31,236,31,236,30,236,29,236,28,179,31,146,31,102,31,102,30,222,31,73,31,228,31,15,31,87,31,3,31,80,31,215,31,76,31,248,31,248,30,161,31,233,31,1,31,249,31,249,30,195,31,195,30,9,31,185,31,33,31,33,30,203,31,203,30,233,31,44,31,216,31,29,31,150,31,158,31,212,31,212,30,26,31,42,31,42,30,9,31,157,31,157,30,146,31,42,31,43,31,250,31,5,31,5,30,35,31,35,30,202,31,147,31,209,31,174,31,130,31,130,31,227,31,120,31,198,31,133,31,112,31,112,30,16,31,183,31,236,31,157,31,249,31,183,31,142,31,80,31,80,30,44,31,44,30,44,29,97,31,97,30,97,29,97,28,35,31,66,31,88,31,88,30,70,31,165,31,104,31,104,31,198,31,198,30,138,31,158,31,104,31,104,30,104,29,104,28,172,31,172,30,14,31,83,31,83,30,176,31,193,31,193,30,193,29,109,31,19,31,163,31,163,30,40,31,242,31,3,31,54,31,52,31,41,31,231,31,243,31,178,31,157,31,157,30,98,31,127,31,225,31,149,31,149,30,223,31,153,31,46,31,204,31,204,30,221,31,40,31,128,31,82,31,82,30,54,31,54,30,79,31,79,30,69,31,126,31,221,31,115,31,52,31,113,31,165,31,42,31,107,31,114,31,239,31,240,31,157,31,157,30,88,31,88,30,19,31,37,31,37,30,154,31,127,31,163,31,172,31,172,31,172,30,172,29,151,31,163,31,137,31,231,31,231,30,226,31,226,30,137,31,15,31,15,30,255,31,255,30,85,31,22,31,205,31,195,31,8,31,228,31,52,31,48,31,233,31,233,30,91,31,253,31,253,30,46,31,46,30,33,31,33,30,44,31,4,31,4,30,4,29,83,31,142,31,76,31,76,30,76,29,76,28,76,27,196,31,196,30,245,31,93,31,97,31,32,31,37,31,37,30,126,31,212,31,249,31,21,31,84,31,123,31,228,31,219,31,219,30,172,31,75,31,12,31,118,31,118,30,49,31,103,31,103,30,103,29,187,31,250,31,227,31,227,30,16,31,57,31,12,31,12,30,91,31,70,31,170,31,229,31,243,31,142,31,142,30,64,31,97,31,104,31,87,31,150,31,25,31,109,31,119,31,119,30,233,31,145,31,145,30,145,29,227,31,44,31,207,31,225,31,74,31,74,30,194,31,194,30,194,29,64,31,104,31,158,31,67,31,29,31,218,31,7,31,42,31,42,30,25,31,155,31,222,31,128,31,221,31,79,31,91,31,91,30,91,29,255,31,91,31,10,31,178,31,150,31,37,31,37,30,153,31,49,31,182,31,70,31,67,31,67,30,151,31,237,31,127,31,1,31,91,31,28,31,42,31,60,31,145,31,157,31,95,31,140,31,15,31,221,31,137,31,255,31,232,31,120,31,36,31,93,31,133,31,28,31,82,31,193,31,45,31,97,31,162,31,162,30,155,31,253,31,124,31,232,31,57,31,57,30,65,31,36,31,248,31,125,31,154,31,149,31,204,31,204,30,252,31,157,31,232,31,150,31,6,31,6,30,6,29,115,31,155,31,118,31,89,31,155,31,145,31,242,31,193,31,174,31,156,31,196,31,26,31,249,31,249,30,26,31,104,31,104,30,28,31,28,30,155,31,164,31,128,31,252,31,100,31,209,31,209,30,194,31,135,31,247,31,247,31,49,31,186,31,121,31,100,31,63,31,63,30,15,31,175,31,175,30,78,31,229,31,113,31,156,31,48,31,65,31,65,30,99,31,241,31,178,31,178,30,218,31,41,31,85,31,85,30,85,29,85,28,165,31,165,30,158,31,141,31,141,30,18,31,231,31,231,30,186,31,186,30,186,29,69,31,232,31,232,30,188,31,93,31,2,31,94,31,94,30,72,31,254,31,254,30,247,31,53,31,76,31,109,31,107,31,107,30,120,31,175,31,175,30,231,31,71,31,3,31,3,30,175,31,174,31,134,31,139,31,12,31,30,31,99,31,49,31,249,31,249,30,150,31,163,31,27,31,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
