-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_196 is
end project_tb_196;

architecture project_tb_arch_196 of project_tb_196 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 812;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (47,0,157,0,69,0,232,0,0,0,37,0,156,0,19,0,11,0,57,0,0,0,1,0,0,0,136,0,226,0,167,0,178,0,108,0,11,0,0,0,0,0,0,0,27,0,74,0,186,0,0,0,109,0,108,0,235,0,103,0,120,0,8,0,49,0,0,0,191,0,164,0,138,0,212,0,147,0,154,0,239,0,150,0,131,0,96,0,14,0,211,0,113,0,162,0,21,0,130,0,250,0,0,0,107,0,12,0,182,0,190,0,202,0,97,0,174,0,79,0,62,0,94,0,0,0,121,0,218,0,226,0,204,0,184,0,183,0,0,0,128,0,120,0,148,0,228,0,29,0,193,0,0,0,139,0,181,0,16,0,36,0,247,0,0,0,172,0,0,0,66,0,40,0,174,0,0,0,230,0,49,0,94,0,199,0,51,0,210,0,27,0,128,0,56,0,113,0,53,0,0,0,16,0,92,0,86,0,94,0,31,0,0,0,32,0,196,0,178,0,123,0,71,0,0,0,125,0,30,0,234,0,202,0,218,0,0,0,251,0,186,0,120,0,191,0,121,0,0,0,171,0,121,0,0,0,170,0,241,0,42,0,18,0,137,0,59,0,246,0,46,0,131,0,77,0,58,0,177,0,0,0,59,0,50,0,220,0,18,0,67,0,110,0,178,0,146,0,46,0,167,0,34,0,0,0,146,0,116,0,58,0,104,0,209,0,0,0,203,0,214,0,95,0,0,0,227,0,0,0,17,0,83,0,184,0,183,0,0,0,0,0,120,0,27,0,229,0,0,0,95,0,0,0,49,0,206,0,161,0,0,0,144,0,82,0,77,0,0,0,0,0,199,0,13,0,192,0,226,0,65,0,0,0,94,0,56,0,222,0,63,0,73,0,0,0,0,0,203,0,218,0,67,0,190,0,61,0,110,0,106,0,189,0,209,0,181,0,197,0,4,0,42,0,0,0,16,0,237,0,125,0,251,0,0,0,162,0,33,0,0,0,0,0,225,0,71,0,60,0,6,0,241,0,105,0,66,0,0,0,226,0,56,0,137,0,0,0,0,0,170,0,28,0,210,0,92,0,83,0,0,0,146,0,214,0,0,0,161,0,1,0,67,0,219,0,122,0,204,0,116,0,14,0,46,0,113,0,0,0,237,0,25,0,18,0,225,0,241,0,31,0,112,0,0,0,16,0,45,0,23,0,92,0,168,0,248,0,30,0,14,0,45,0,159,0,126,0,88,0,150,0,226,0,175,0,14,0,45,0,143,0,0,0,234,0,205,0,56,0,197,0,17,0,49,0,0,0,223,0,85,0,236,0,94,0,158,0,44,0,167,0,28,0,0,0,4,0,168,0,43,0,138,0,231,0,0,0,0,0,68,0,164,0,132,0,0,0,0,0,0,0,77,0,70,0,224,0,99,0,69,0,145,0,156,0,0,0,0,0,15,0,89,0,175,0,0,0,76,0,192,0,0,0,0,0,201,0,31,0,74,0,175,0,214,0,147,0,0,0,199,0,75,0,43,0,102,0,0,0,79,0,69,0,141,0,207,0,65,0,0,0,61,0,26,0,231,0,0,0,0,0,142,0,220,0,164,0,134,0,237,0,175,0,144,0,32,0,91,0,0,0,3,0,246,0,229,0,148,0,75,0,0,0,0,0,149,0,0,0,196,0,178,0,251,0,115,0,221,0,180,0,227,0,106,0,107,0,179,0,38,0,0,0,171,0,77,0,23,0,0,0,0,0,177,0,118,0,117,0,156,0,163,0,58,0,196,0,41,0,36,0,93,0,255,0,94,0,0,0,125,0,60,0,118,0,64,0,86,0,100,0,0,0,30,0,15,0,22,0,5,0,188,0,45,0,0,0,8,0,236,0,0,0,206,0,55,0,73,0,13,0,0,0,65,0,0,0,153,0,39,0,96,0,136,0,36,0,44,0,127,0,122,0,86,0,224,0,161,0,181,0,110,0,0,0,152,0,110,0,246,0,253,0,226,0,0,0,54,0,175,0,49,0,85,0,195,0,191,0,0,0,172,0,210,0,239,0,0,0,74,0,187,0,0,0,7,0,195,0,45,0,204,0,64,0,163,0,178,0,137,0,93,0,0,0,0,0,11,0,71,0,242,0,226,0,214,0,0,0,209,0,196,0,221,0,195,0,71,0,179,0,81,0,166,0,14,0,207,0,6,0,174,0,159,0,86,0,214,0,64,0,137,0,191,0,226,0,154,0,0,0,91,0,108,0,3,0,157,0,9,0,102,0,0,0,95,0,130,0,194,0,41,0,16,0,0,0,42,0,161,0,0,0,87,0,144,0,73,0,179,0,223,0,96,0,195,0,90,0,131,0,0,0,146,0,0,0,129,0,107,0,91,0,179,0,0,0,0,0,229,0,212,0,1,0,223,0,0,0,182,0,234,0,0,0,0,0,103,0,45,0,112,0,244,0,227,0,9,0,232,0,183,0,152,0,45,0,0,0,36,0,0,0,99,0,254,0,241,0,84,0,179,0,247,0,168,0,253,0,163,0,0,0,248,0,224,0,116,0,130,0,158,0,60,0,129,0,110,0,75,0,75,0,171,0,0,0,253,0,64,0,0,0,110,0,0,0,55,0,57,0,155,0,0,0,0,0,159,0,78,0,104,0,224,0,0,0,0,0,130,0,0,0,141,0,34,0,172,0,77,0,38,0,0,0,100,0,142,0,1,0,43,0,90,0,51,0,42,0,249,0,115,0,165,0,127,0,0,0,199,0,0,0,195,0,179,0,255,0,123,0,0,0,198,0,235,0,0,0,47,0,38,0,0,0,116,0,0,0,121,0,71,0,206,0,199,0,0,0,30,0,181,0,232,0,3,0,201,0,53,0,16,0,0,0,96,0,152,0,145,0,187,0,184,0,100,0,153,0,66,0,180,0,218,0,126,0,0,0,232,0,73,0,156,0,0,0,37,0,153,0,0,0,0,0,10,0,0,0,0,0,226,0,0,0,54,0,168,0,247,0,217,0,114,0,107,0,249,0,8,0,233,0,152,0,47,0,0,0,162,0,0,0,55,0,105,0,72,0,119,0,24,0,26,0,140,0,169,0,3,0,37,0,199,0,54,0,103,0,218,0,188,0,114,0,125,0,0,0,219,0,0,0,203,0,97,0,160,0,53,0,134,0,0,0,47,0,190,0,168,0,139,0,25,0,0,0,0,0,86,0,168,0,0,0,106,0,130,0,83,0,158,0,106,0,0,0,128,0,46,0,204,0,89,0,13,0,104,0,113,0,242,0,123,0,214,0,0,0,250,0,0,0,145,0,42,0,210,0,146,0,198,0,80,0,6,0,2,0,0,0,116,0,33,0,151,0,0,0,252,0,151,0,97,0,141,0,0,0,41,0,25,0,84,0,134,0,118,0,4,0,24,0,164,0,0,0,80,0,0,0,0,0,241,0,112,0,158,0,73,0,0,0,130,0,80,0,44,0,145,0,115,0,212,0,0,0,89,0,209,0,104,0,185,0,158,0,35,0,50,0,212,0,58,0,0,0,0,0,0,0,252,0,96,0,86,0,59,0,121,0,0,0,145,0,0,0,25,0,0,0,24,0,116,0,0,0,0,0,0,0,19,0,247,0,194,0,65,0,56,0,126,0,192,0,193,0,0,0,191,0,130,0);
signal scenario_full  : scenario_type := (47,31,157,31,69,31,232,31,232,30,37,31,156,31,19,31,11,31,57,31,57,30,1,31,1,30,136,31,226,31,167,31,178,31,108,31,11,31,11,30,11,29,11,28,27,31,74,31,186,31,186,30,109,31,108,31,235,31,103,31,120,31,8,31,49,31,49,30,191,31,164,31,138,31,212,31,147,31,154,31,239,31,150,31,131,31,96,31,14,31,211,31,113,31,162,31,21,31,130,31,250,31,250,30,107,31,12,31,182,31,190,31,202,31,97,31,174,31,79,31,62,31,94,31,94,30,121,31,218,31,226,31,204,31,184,31,183,31,183,30,128,31,120,31,148,31,228,31,29,31,193,31,193,30,139,31,181,31,16,31,36,31,247,31,247,30,172,31,172,30,66,31,40,31,174,31,174,30,230,31,49,31,94,31,199,31,51,31,210,31,27,31,128,31,56,31,113,31,53,31,53,30,16,31,92,31,86,31,94,31,31,31,31,30,32,31,196,31,178,31,123,31,71,31,71,30,125,31,30,31,234,31,202,31,218,31,218,30,251,31,186,31,120,31,191,31,121,31,121,30,171,31,121,31,121,30,170,31,241,31,42,31,18,31,137,31,59,31,246,31,46,31,131,31,77,31,58,31,177,31,177,30,59,31,50,31,220,31,18,31,67,31,110,31,178,31,146,31,46,31,167,31,34,31,34,30,146,31,116,31,58,31,104,31,209,31,209,30,203,31,214,31,95,31,95,30,227,31,227,30,17,31,83,31,184,31,183,31,183,30,183,29,120,31,27,31,229,31,229,30,95,31,95,30,49,31,206,31,161,31,161,30,144,31,82,31,77,31,77,30,77,29,199,31,13,31,192,31,226,31,65,31,65,30,94,31,56,31,222,31,63,31,73,31,73,30,73,29,203,31,218,31,67,31,190,31,61,31,110,31,106,31,189,31,209,31,181,31,197,31,4,31,42,31,42,30,16,31,237,31,125,31,251,31,251,30,162,31,33,31,33,30,33,29,225,31,71,31,60,31,6,31,241,31,105,31,66,31,66,30,226,31,56,31,137,31,137,30,137,29,170,31,28,31,210,31,92,31,83,31,83,30,146,31,214,31,214,30,161,31,1,31,67,31,219,31,122,31,204,31,116,31,14,31,46,31,113,31,113,30,237,31,25,31,18,31,225,31,241,31,31,31,112,31,112,30,16,31,45,31,23,31,92,31,168,31,248,31,30,31,14,31,45,31,159,31,126,31,88,31,150,31,226,31,175,31,14,31,45,31,143,31,143,30,234,31,205,31,56,31,197,31,17,31,49,31,49,30,223,31,85,31,236,31,94,31,158,31,44,31,167,31,28,31,28,30,4,31,168,31,43,31,138,31,231,31,231,30,231,29,68,31,164,31,132,31,132,30,132,29,132,28,77,31,70,31,224,31,99,31,69,31,145,31,156,31,156,30,156,29,15,31,89,31,175,31,175,30,76,31,192,31,192,30,192,29,201,31,31,31,74,31,175,31,214,31,147,31,147,30,199,31,75,31,43,31,102,31,102,30,79,31,69,31,141,31,207,31,65,31,65,30,61,31,26,31,231,31,231,30,231,29,142,31,220,31,164,31,134,31,237,31,175,31,144,31,32,31,91,31,91,30,3,31,246,31,229,31,148,31,75,31,75,30,75,29,149,31,149,30,196,31,178,31,251,31,115,31,221,31,180,31,227,31,106,31,107,31,179,31,38,31,38,30,171,31,77,31,23,31,23,30,23,29,177,31,118,31,117,31,156,31,163,31,58,31,196,31,41,31,36,31,93,31,255,31,94,31,94,30,125,31,60,31,118,31,64,31,86,31,100,31,100,30,30,31,15,31,22,31,5,31,188,31,45,31,45,30,8,31,236,31,236,30,206,31,55,31,73,31,13,31,13,30,65,31,65,30,153,31,39,31,96,31,136,31,36,31,44,31,127,31,122,31,86,31,224,31,161,31,181,31,110,31,110,30,152,31,110,31,246,31,253,31,226,31,226,30,54,31,175,31,49,31,85,31,195,31,191,31,191,30,172,31,210,31,239,31,239,30,74,31,187,31,187,30,7,31,195,31,45,31,204,31,64,31,163,31,178,31,137,31,93,31,93,30,93,29,11,31,71,31,242,31,226,31,214,31,214,30,209,31,196,31,221,31,195,31,71,31,179,31,81,31,166,31,14,31,207,31,6,31,174,31,159,31,86,31,214,31,64,31,137,31,191,31,226,31,154,31,154,30,91,31,108,31,3,31,157,31,9,31,102,31,102,30,95,31,130,31,194,31,41,31,16,31,16,30,42,31,161,31,161,30,87,31,144,31,73,31,179,31,223,31,96,31,195,31,90,31,131,31,131,30,146,31,146,30,129,31,107,31,91,31,179,31,179,30,179,29,229,31,212,31,1,31,223,31,223,30,182,31,234,31,234,30,234,29,103,31,45,31,112,31,244,31,227,31,9,31,232,31,183,31,152,31,45,31,45,30,36,31,36,30,99,31,254,31,241,31,84,31,179,31,247,31,168,31,253,31,163,31,163,30,248,31,224,31,116,31,130,31,158,31,60,31,129,31,110,31,75,31,75,31,171,31,171,30,253,31,64,31,64,30,110,31,110,30,55,31,57,31,155,31,155,30,155,29,159,31,78,31,104,31,224,31,224,30,224,29,130,31,130,30,141,31,34,31,172,31,77,31,38,31,38,30,100,31,142,31,1,31,43,31,90,31,51,31,42,31,249,31,115,31,165,31,127,31,127,30,199,31,199,30,195,31,179,31,255,31,123,31,123,30,198,31,235,31,235,30,47,31,38,31,38,30,116,31,116,30,121,31,71,31,206,31,199,31,199,30,30,31,181,31,232,31,3,31,201,31,53,31,16,31,16,30,96,31,152,31,145,31,187,31,184,31,100,31,153,31,66,31,180,31,218,31,126,31,126,30,232,31,73,31,156,31,156,30,37,31,153,31,153,30,153,29,10,31,10,30,10,29,226,31,226,30,54,31,168,31,247,31,217,31,114,31,107,31,249,31,8,31,233,31,152,31,47,31,47,30,162,31,162,30,55,31,105,31,72,31,119,31,24,31,26,31,140,31,169,31,3,31,37,31,199,31,54,31,103,31,218,31,188,31,114,31,125,31,125,30,219,31,219,30,203,31,97,31,160,31,53,31,134,31,134,30,47,31,190,31,168,31,139,31,25,31,25,30,25,29,86,31,168,31,168,30,106,31,130,31,83,31,158,31,106,31,106,30,128,31,46,31,204,31,89,31,13,31,104,31,113,31,242,31,123,31,214,31,214,30,250,31,250,30,145,31,42,31,210,31,146,31,198,31,80,31,6,31,2,31,2,30,116,31,33,31,151,31,151,30,252,31,151,31,97,31,141,31,141,30,41,31,25,31,84,31,134,31,118,31,4,31,24,31,164,31,164,30,80,31,80,30,80,29,241,31,112,31,158,31,73,31,73,30,130,31,80,31,44,31,145,31,115,31,212,31,212,30,89,31,209,31,104,31,185,31,158,31,35,31,50,31,212,31,58,31,58,30,58,29,58,28,252,31,96,31,86,31,59,31,121,31,121,30,145,31,145,30,25,31,25,30,24,31,116,31,116,30,116,29,116,28,19,31,247,31,194,31,65,31,56,31,126,31,192,31,193,31,193,30,191,31,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
