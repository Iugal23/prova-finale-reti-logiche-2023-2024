-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_817 is
end project_tb_817;

architecture project_tb_arch_817 of project_tb_817 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,148,0,98,0,116,0,0,0,113,0,98,0,46,0,0,0,46,0,145,0,10,0,183,0,0,0,0,0,86,0,77,0,0,0,0,0,54,0,213,0,54,0,20,0,41,0,6,0,250,0,147,0,0,0,35,0,177,0,29,0,231,0,234,0,184,0,43,0,13,0,71,0,156,0,0,0,136,0,0,0,60,0,199,0,149,0,52,0,73,0,0,0,110,0,0,0,186,0,0,0,152,0,19,0,167,0,35,0,161,0,89,0,231,0,90,0,64,0,160,0,237,0,124,0,203,0,53,0,0,0,114,0,215,0,0,0,68,0,135,0,5,0,251,0,90,0,74,0,221,0,0,0,213,0,39,0,47,0,191,0,78,0,194,0,82,0,0,0,234,0,36,0,114,0,160,0,205,0,0,0,235,0,117,0,1,0,159,0,0,0,177,0,146,0,59,0,95,0,0,0,140,0,133,0,149,0,150,0,131,0,206,0,192,0,215,0,218,0,142,0,0,0,177,0,232,0,151,0,93,0,0,0,197,0,149,0,254,0,83,0,172,0,0,0,119,0,82,0,41,0,221,0,104,0,172,0,29,0,0,0,0,0,174,0,153,0,37,0,98,0,8,0,105,0,42,0,0,0,51,0,124,0,64,0,149,0,170,0,1,0,88,0,121,0,177,0,61,0,16,0,238,0,229,0,111,0,29,0,51,0,98,0,34,0,38,0,37,0,7,0,130,0,129,0,247,0,87,0,0,0,82,0,51,0,186,0,0,0,34,0,158,0,143,0,46,0,128,0,131,0,0,0,35,0,181,0,204,0,169,0,0,0,49,0,23,0,0,0,72,0,207,0,162,0,132,0,69,0,0,0,0,0,40,0,86,0,19,0,0,0,0,0,99,0,131,0,91,0,154,0,236,0,11,0,114,0,0,0,113,0,208,0,0,0,0,0,0,0,0,0,31,0,51,0,130,0,3,0,181,0,180,0,78,0,114,0,226,0,63,0,250,0,6,0,198,0,0,0,245,0,5,0,3,0,253,0,104,0,38,0,215,0,184,0,49,0,59,0,0,0,72,0,105,0,250,0,185,0,100,0,0,0,142,0,0,0,1,0,152,0,0,0,162,0,0,0,0,0,0,0,74,0,0,0,109,0,126,0,60,0,172,0,141,0,148,0,159,0,227,0,0,0,33,0,138,0,59,0,245,0,169,0,242,0,12,0,170,0,0,0,185,0,0,0,236,0,224,0,0,0,121,0,205,0,41,0,0,0,92,0,98,0,231,0,244,0,42,0,50,0,129,0,68,0,0,0,0,0,0,0,7,0,73,0,32,0,90,0,0,0,195,0,0,0,20,0,79,0,72,0,184,0,179,0,212,0,56,0,164,0,47,0,38,0,34,0,246,0,0,0,57,0,127,0,199,0,216,0,222,0,111,0,0,0,0,0,218,0,187,0,97,0,0,0,57,0,255,0,183,0,13,0,112,0,126,0,170,0,189,0,45,0,118,0,71,0,0,0,20,0,97,0,94,0,202,0,227,0,46,0,158,0,0,0,105,0,89,0,33,0,1,0,144,0,99,0,173,0,0,0,195,0,0,0,0,0,125,0,170,0,41,0,182,0,110,0,8,0,0,0,160,0,16,0,236,0,23,0,0,0,110,0,75,0,159,0,25,0,2,0,126,0,200,0,30,0,44,0,50,0,0,0,7,0,17,0,42,0,111,0,155,0,102,0,121,0,0,0,133,0,101,0,70,0,207,0,152,0,197,0,154,0,154,0,176,0,163,0,80,0,181,0,0,0,136,0,75,0,0,0,0,0,225,0,73,0,0,0,198,0,149,0,192,0,0,0,84,0,0,0,67,0,0,0,104,0,118,0,158,0,200,0,248,0,102,0,132,0,230,0,91,0,237,0,250,0,53,0,0,0,53,0,60,0,126,0,38,0,58,0,151,0,209,0,158,0,42,0,17,0,0,0,0,0,198,0,113,0,202,0,12,0,208,0,0,0,0,0,136,0,248,0,0,0,181,0,19,0,223,0,140,0,67,0,104,0,251,0,16,0,155,0,191,0,138,0,0,0,53,0,184,0,231,0,196,0,69,0,128,0,0,0,135,0,99,0,188,0,158,0,36,0,239,0,183,0,12,0,0,0,69,0,205,0,0,0,111,0,188,0,0,0,35,0,143,0,201,0,231,0,252,0,2,0,108,0,86,0,57,0,118,0,191,0,182,0,200,0,137,0,232,0,97,0,0,0,114,0,0,0,0,0,95,0,130,0,122,0,0,0,100,0,196,0,0,0,171,0,223,0,88,0,185,0,1,0,180,0,0,0,0,0,204,0,240,0,235,0,95,0,0,0,0,0,250,0,0,0,49,0,151,0,0,0,156,0,198,0,147,0,71,0,94,0,4,0,131,0,44,0,191,0,13,0,0,0,207,0,76,0,221,0,113,0,0,0,105,0,76,0,63,0,195,0,111,0,245,0,133,0,122,0,209,0,227,0,86,0,245,0,141,0,0,0,30,0,0,0,194,0,0,0,39,0,0,0,0,0,197,0,194,0,64,0,13,0,132,0,179,0,177,0,234,0,3,0,244,0,185,0,0,0,12,0,110,0,2,0,85,0,160,0,96,0,0,0,0,0,235,0,16,0,0,0,0,0,169,0,0,0,226,0,0,0,246,0,162,0,89,0,77,0,0,0,217,0,82,0,187,0,20,0,181,0,0,0,227,0,2,0,137,0,0,0,20,0,224,0,188,0,0,0,47,0,0,0,82,0,28,0,127,0,249,0,0,0,210,0,89,0,144,0,76,0,0,0,105,0,102,0,145,0,104,0,47,0,0,0,207,0,254,0,61,0,6,0,196,0,203,0,6,0,183,0,0,0,195,0,8,0,165,0,0,0,55,0,0,0,0,0,98,0,164,0,111,0,112,0,242,0,0,0,33,0,14,0,48,0,41,0,235,0,0,0,138,0,83,0,248,0,3,0,112,0,18,0,18,0,0,0,235,0,224,0,185,0,167,0,211,0,99,0,219,0,108,0,82,0,202,0,0,0,214,0,112,0,0,0,51,0,203,0,108,0,2,0,72,0,0,0,30,0,78,0,182,0,0,0,228,0,205,0,157,0,17,0,236,0,133,0,0,0,0,0,10,0,159,0,8,0,0,0,202,0,146,0,19,0,255,0,0,0,128,0,165,0,206,0,237,0,191,0,220,0,138,0,134,0,0,0,232,0,118,0,88,0,204,0,219,0,0,0,212,0,225,0,133,0,149,0,76,0,1,0,43,0,138,0,198,0,188,0,84,0,124,0,161,0,245,0,0,0,205,0,9,0,90,0,91,0,166,0,113,0,197,0,138,0,0,0,204,0,0,0,0,0,14,0,75,0,67,0,0,0,127,0,131,0,232,0,21,0,8,0,0,0,14,0,0,0,253,0,249,0,16,0,83,0,84,0,225,0,97,0,150,0,24,0,133,0,3,0,0,0,242,0,0,0,42,0,239,0,0,0,58,0,147,0,16,0,0,0,239,0,143,0,0,0,221,0,231,0,0,0,52,0,195,0,130,0,223,0,0,0,0,0,211,0,0,0,209,0,170,0,0,0,223,0,100,0,0,0,62,0,0,0,11,0,0,0,94,0,0,0,0,0,0,0,201,0,254,0,122,0,11,0,0,0,0,0,211,0,0,0,0,0,8,0,32,0,94,0,141,0,0,0,0,0,148,0,0,0,38,0,115,0,0,0,152,0,0,0,166,0,189,0,0,0,0,0,7,0,0,0,17,0,29,0,0,0,88,0,0,0,237,0,131,0,95,0,0,0,49,0,71,0,236,0,0,0,244,0,248,0,0,0,123,0,183,0,176,0,136,0,124,0,15,0,155,0,118,0,119,0,217,0,20,0,71,0,72,0,65,0,0,0,214,0,166,0,90,0,125,0,229,0,149,0,51,0,95,0,158,0,205,0,251,0,169,0,154,0,126,0,195,0,189,0,186,0,176,0,168,0,0,0,125,0,222,0,117,0,70,0,126,0,161,0,115,0,253,0,49,0,12,0,131,0,0,0,220,0,108,0,13,0,0,0,17,0,241,0,223,0,118,0,203,0,27,0,47,0,0,0,42,0,195,0,0,0,146,0,247,0,0,0,81,0,0,0,200,0,0,0,134,0,0,0,122,0,227,0,48,0,138,0,0,0,194,0,46,0,16,0,124,0,14,0,179,0,0,0,255,0,0,0,227,0,99,0,80,0,137,0,68,0,122,0,97,0,186,0,109,0,249,0,58,0,46,0,169,0,153,0,211,0,126,0,0,0,158,0,63,0,124,0,180,0,90,0,46,0,0,0,214,0,0,0,232,0,0,0,189,0,84,0,84,0,79,0,18,0,139,0,0,0,129,0);
signal scenario_full  : scenario_type := (0,0,148,31,98,31,116,31,116,30,113,31,98,31,46,31,46,30,46,31,145,31,10,31,183,31,183,30,183,29,86,31,77,31,77,30,77,29,54,31,213,31,54,31,20,31,41,31,6,31,250,31,147,31,147,30,35,31,177,31,29,31,231,31,234,31,184,31,43,31,13,31,71,31,156,31,156,30,136,31,136,30,60,31,199,31,149,31,52,31,73,31,73,30,110,31,110,30,186,31,186,30,152,31,19,31,167,31,35,31,161,31,89,31,231,31,90,31,64,31,160,31,237,31,124,31,203,31,53,31,53,30,114,31,215,31,215,30,68,31,135,31,5,31,251,31,90,31,74,31,221,31,221,30,213,31,39,31,47,31,191,31,78,31,194,31,82,31,82,30,234,31,36,31,114,31,160,31,205,31,205,30,235,31,117,31,1,31,159,31,159,30,177,31,146,31,59,31,95,31,95,30,140,31,133,31,149,31,150,31,131,31,206,31,192,31,215,31,218,31,142,31,142,30,177,31,232,31,151,31,93,31,93,30,197,31,149,31,254,31,83,31,172,31,172,30,119,31,82,31,41,31,221,31,104,31,172,31,29,31,29,30,29,29,174,31,153,31,37,31,98,31,8,31,105,31,42,31,42,30,51,31,124,31,64,31,149,31,170,31,1,31,88,31,121,31,177,31,61,31,16,31,238,31,229,31,111,31,29,31,51,31,98,31,34,31,38,31,37,31,7,31,130,31,129,31,247,31,87,31,87,30,82,31,51,31,186,31,186,30,34,31,158,31,143,31,46,31,128,31,131,31,131,30,35,31,181,31,204,31,169,31,169,30,49,31,23,31,23,30,72,31,207,31,162,31,132,31,69,31,69,30,69,29,40,31,86,31,19,31,19,30,19,29,99,31,131,31,91,31,154,31,236,31,11,31,114,31,114,30,113,31,208,31,208,30,208,29,208,28,208,27,31,31,51,31,130,31,3,31,181,31,180,31,78,31,114,31,226,31,63,31,250,31,6,31,198,31,198,30,245,31,5,31,3,31,253,31,104,31,38,31,215,31,184,31,49,31,59,31,59,30,72,31,105,31,250,31,185,31,100,31,100,30,142,31,142,30,1,31,152,31,152,30,162,31,162,30,162,29,162,28,74,31,74,30,109,31,126,31,60,31,172,31,141,31,148,31,159,31,227,31,227,30,33,31,138,31,59,31,245,31,169,31,242,31,12,31,170,31,170,30,185,31,185,30,236,31,224,31,224,30,121,31,205,31,41,31,41,30,92,31,98,31,231,31,244,31,42,31,50,31,129,31,68,31,68,30,68,29,68,28,7,31,73,31,32,31,90,31,90,30,195,31,195,30,20,31,79,31,72,31,184,31,179,31,212,31,56,31,164,31,47,31,38,31,34,31,246,31,246,30,57,31,127,31,199,31,216,31,222,31,111,31,111,30,111,29,218,31,187,31,97,31,97,30,57,31,255,31,183,31,13,31,112,31,126,31,170,31,189,31,45,31,118,31,71,31,71,30,20,31,97,31,94,31,202,31,227,31,46,31,158,31,158,30,105,31,89,31,33,31,1,31,144,31,99,31,173,31,173,30,195,31,195,30,195,29,125,31,170,31,41,31,182,31,110,31,8,31,8,30,160,31,16,31,236,31,23,31,23,30,110,31,75,31,159,31,25,31,2,31,126,31,200,31,30,31,44,31,50,31,50,30,7,31,17,31,42,31,111,31,155,31,102,31,121,31,121,30,133,31,101,31,70,31,207,31,152,31,197,31,154,31,154,31,176,31,163,31,80,31,181,31,181,30,136,31,75,31,75,30,75,29,225,31,73,31,73,30,198,31,149,31,192,31,192,30,84,31,84,30,67,31,67,30,104,31,118,31,158,31,200,31,248,31,102,31,132,31,230,31,91,31,237,31,250,31,53,31,53,30,53,31,60,31,126,31,38,31,58,31,151,31,209,31,158,31,42,31,17,31,17,30,17,29,198,31,113,31,202,31,12,31,208,31,208,30,208,29,136,31,248,31,248,30,181,31,19,31,223,31,140,31,67,31,104,31,251,31,16,31,155,31,191,31,138,31,138,30,53,31,184,31,231,31,196,31,69,31,128,31,128,30,135,31,99,31,188,31,158,31,36,31,239,31,183,31,12,31,12,30,69,31,205,31,205,30,111,31,188,31,188,30,35,31,143,31,201,31,231,31,252,31,2,31,108,31,86,31,57,31,118,31,191,31,182,31,200,31,137,31,232,31,97,31,97,30,114,31,114,30,114,29,95,31,130,31,122,31,122,30,100,31,196,31,196,30,171,31,223,31,88,31,185,31,1,31,180,31,180,30,180,29,204,31,240,31,235,31,95,31,95,30,95,29,250,31,250,30,49,31,151,31,151,30,156,31,198,31,147,31,71,31,94,31,4,31,131,31,44,31,191,31,13,31,13,30,207,31,76,31,221,31,113,31,113,30,105,31,76,31,63,31,195,31,111,31,245,31,133,31,122,31,209,31,227,31,86,31,245,31,141,31,141,30,30,31,30,30,194,31,194,30,39,31,39,30,39,29,197,31,194,31,64,31,13,31,132,31,179,31,177,31,234,31,3,31,244,31,185,31,185,30,12,31,110,31,2,31,85,31,160,31,96,31,96,30,96,29,235,31,16,31,16,30,16,29,169,31,169,30,226,31,226,30,246,31,162,31,89,31,77,31,77,30,217,31,82,31,187,31,20,31,181,31,181,30,227,31,2,31,137,31,137,30,20,31,224,31,188,31,188,30,47,31,47,30,82,31,28,31,127,31,249,31,249,30,210,31,89,31,144,31,76,31,76,30,105,31,102,31,145,31,104,31,47,31,47,30,207,31,254,31,61,31,6,31,196,31,203,31,6,31,183,31,183,30,195,31,8,31,165,31,165,30,55,31,55,30,55,29,98,31,164,31,111,31,112,31,242,31,242,30,33,31,14,31,48,31,41,31,235,31,235,30,138,31,83,31,248,31,3,31,112,31,18,31,18,31,18,30,235,31,224,31,185,31,167,31,211,31,99,31,219,31,108,31,82,31,202,31,202,30,214,31,112,31,112,30,51,31,203,31,108,31,2,31,72,31,72,30,30,31,78,31,182,31,182,30,228,31,205,31,157,31,17,31,236,31,133,31,133,30,133,29,10,31,159,31,8,31,8,30,202,31,146,31,19,31,255,31,255,30,128,31,165,31,206,31,237,31,191,31,220,31,138,31,134,31,134,30,232,31,118,31,88,31,204,31,219,31,219,30,212,31,225,31,133,31,149,31,76,31,1,31,43,31,138,31,198,31,188,31,84,31,124,31,161,31,245,31,245,30,205,31,9,31,90,31,91,31,166,31,113,31,197,31,138,31,138,30,204,31,204,30,204,29,14,31,75,31,67,31,67,30,127,31,131,31,232,31,21,31,8,31,8,30,14,31,14,30,253,31,249,31,16,31,83,31,84,31,225,31,97,31,150,31,24,31,133,31,3,31,3,30,242,31,242,30,42,31,239,31,239,30,58,31,147,31,16,31,16,30,239,31,143,31,143,30,221,31,231,31,231,30,52,31,195,31,130,31,223,31,223,30,223,29,211,31,211,30,209,31,170,31,170,30,223,31,100,31,100,30,62,31,62,30,11,31,11,30,94,31,94,30,94,29,94,28,201,31,254,31,122,31,11,31,11,30,11,29,211,31,211,30,211,29,8,31,32,31,94,31,141,31,141,30,141,29,148,31,148,30,38,31,115,31,115,30,152,31,152,30,166,31,189,31,189,30,189,29,7,31,7,30,17,31,29,31,29,30,88,31,88,30,237,31,131,31,95,31,95,30,49,31,71,31,236,31,236,30,244,31,248,31,248,30,123,31,183,31,176,31,136,31,124,31,15,31,155,31,118,31,119,31,217,31,20,31,71,31,72,31,65,31,65,30,214,31,166,31,90,31,125,31,229,31,149,31,51,31,95,31,158,31,205,31,251,31,169,31,154,31,126,31,195,31,189,31,186,31,176,31,168,31,168,30,125,31,222,31,117,31,70,31,126,31,161,31,115,31,253,31,49,31,12,31,131,31,131,30,220,31,108,31,13,31,13,30,17,31,241,31,223,31,118,31,203,31,27,31,47,31,47,30,42,31,195,31,195,30,146,31,247,31,247,30,81,31,81,30,200,31,200,30,134,31,134,30,122,31,227,31,48,31,138,31,138,30,194,31,46,31,16,31,124,31,14,31,179,31,179,30,255,31,255,30,227,31,99,31,80,31,137,31,68,31,122,31,97,31,186,31,109,31,249,31,58,31,46,31,169,31,153,31,211,31,126,31,126,30,158,31,63,31,124,31,180,31,90,31,46,31,46,30,214,31,214,30,232,31,232,30,189,31,84,31,84,31,79,31,18,31,139,31,139,30,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
