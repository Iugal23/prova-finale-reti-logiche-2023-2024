-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 252;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,185,0,0,0,184,0,149,0,12,0,102,0,37,0,134,0,101,0,150,0,0,0,59,0,52,0,183,0,104,0,251,0,191,0,2,0,183,0,0,0,201,0,158,0,6,0,215,0,228,0,73,0,99,0,0,0,253,0,39,0,208,0,255,0,103,0,193,0,166,0,231,0,153,0,115,0,119,0,0,0,0,0,162,0,103,0,0,0,150,0,177,0,155,0,0,0,162,0,0,0,211,0,244,0,171,0,156,0,0,0,45,0,0,0,244,0,235,0,138,0,196,0,22,0,159,0,0,0,0,0,125,0,37,0,182,0,121,0,41,0,167,0,95,0,81,0,13,0,0,0,210,0,0,0,0,0,184,0,181,0,243,0,191,0,177,0,185,0,127,0,150,0,82,0,249,0,77,0,245,0,0,0,152,0,105,0,39,0,0,0,0,0,0,0,80,0,0,0,232,0,0,0,118,0,169,0,176,0,106,0,121,0,34,0,250,0,90,0,107,0,178,0,196,0,239,0,147,0,185,0,223,0,147,0,71,0,0,0,0,0,166,0,20,0,196,0,223,0,0,0,16,0,192,0,37,0,118,0,104,0,0,0,42,0,222,0,232,0,99,0,11,0,191,0,0,0,136,0,0,0,104,0,191,0,121,0,0,0,100,0,190,0,0,0,164,0,131,0,119,0,103,0,0,0,0,0,113,0,119,0,22,0,212,0,0,0,112,0,188,0,125,0,129,0,208,0,96,0,63,0,0,0,0,0,238,0,85,0,0,0,238,0,17,0,79,0,217,0,243,0,0,0,106,0,94,0,220,0,68,0,0,0,199,0,234,0,64,0,0,0,238,0,0,0,253,0,153,0,164,0,52,0,183,0,221,0,118,0,187,0,147,0,0,0,112,0,0,0,142,0,0,0,57,0,0,0,5,0,93,0,86,0,0,0,131,0,45,0,0,0,0,0,2,0,24,0,30,0,0,0,162,0,124,0,0,0,0,0,212,0,0,0,0,0,48,0,96,0,189,0,203,0,90,0,152,0,0,0,232,0,38,0,85,0,0,0,189,0,223,0,0,0,240,0,240,0,0,0,99,0,0,0,199,0,201,0,140,0,76,0,19,0,166,0,176,0,173,0,191,0,2,0);
signal scenario_full  : scenario_type := (87,31,185,31,185,30,184,31,149,31,12,31,102,31,37,31,134,31,101,31,150,31,150,30,59,31,52,31,183,31,104,31,251,31,191,31,2,31,183,31,183,30,201,31,158,31,6,31,215,31,228,31,73,31,99,31,99,30,253,31,39,31,208,31,255,31,103,31,193,31,166,31,231,31,153,31,115,31,119,31,119,30,119,29,162,31,103,31,103,30,150,31,177,31,155,31,155,30,162,31,162,30,211,31,244,31,171,31,156,31,156,30,45,31,45,30,244,31,235,31,138,31,196,31,22,31,159,31,159,30,159,29,125,31,37,31,182,31,121,31,41,31,167,31,95,31,81,31,13,31,13,30,210,31,210,30,210,29,184,31,181,31,243,31,191,31,177,31,185,31,127,31,150,31,82,31,249,31,77,31,245,31,245,30,152,31,105,31,39,31,39,30,39,29,39,28,80,31,80,30,232,31,232,30,118,31,169,31,176,31,106,31,121,31,34,31,250,31,90,31,107,31,178,31,196,31,239,31,147,31,185,31,223,31,147,31,71,31,71,30,71,29,166,31,20,31,196,31,223,31,223,30,16,31,192,31,37,31,118,31,104,31,104,30,42,31,222,31,232,31,99,31,11,31,191,31,191,30,136,31,136,30,104,31,191,31,121,31,121,30,100,31,190,31,190,30,164,31,131,31,119,31,103,31,103,30,103,29,113,31,119,31,22,31,212,31,212,30,112,31,188,31,125,31,129,31,208,31,96,31,63,31,63,30,63,29,238,31,85,31,85,30,238,31,17,31,79,31,217,31,243,31,243,30,106,31,94,31,220,31,68,31,68,30,199,31,234,31,64,31,64,30,238,31,238,30,253,31,153,31,164,31,52,31,183,31,221,31,118,31,187,31,147,31,147,30,112,31,112,30,142,31,142,30,57,31,57,30,5,31,93,31,86,31,86,30,131,31,45,31,45,30,45,29,2,31,24,31,30,31,30,30,162,31,124,31,124,30,124,29,212,31,212,30,212,29,48,31,96,31,189,31,203,31,90,31,152,31,152,30,232,31,38,31,85,31,85,30,189,31,223,31,223,30,240,31,240,31,240,30,99,31,99,30,199,31,201,31,140,31,76,31,19,31,166,31,176,31,173,31,191,31,2,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
