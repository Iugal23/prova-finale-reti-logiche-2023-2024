-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 989;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,132,0,173,0,200,0,0,0,162,0,167,0,219,0,222,0,230,0,235,0,206,0,0,0,142,0,77,0,32,0,124,0,106,0,121,0,0,0,109,0,106,0,221,0,163,0,171,0,60,0,241,0,139,0,58,0,120,0,211,0,0,0,0,0,60,0,0,0,225,0,0,0,136,0,181,0,46,0,126,0,0,0,43,0,58,0,246,0,254,0,216,0,98,0,77,0,150,0,66,0,47,0,112,0,0,0,10,0,0,0,0,0,255,0,233,0,83,0,95,0,149,0,0,0,171,0,154,0,0,0,215,0,23,0,0,0,72,0,89,0,41,0,101,0,0,0,23,0,185,0,58,0,245,0,0,0,189,0,251,0,22,0,78,0,139,0,142,0,16,0,250,0,68,0,41,0,0,0,98,0,127,0,94,0,0,0,100,0,0,0,0,0,0,0,227,0,17,0,176,0,104,0,136,0,216,0,236,0,238,0,86,0,15,0,93,0,57,0,31,0,175,0,56,0,0,0,216,0,177,0,31,0,183,0,190,0,205,0,0,0,253,0,251,0,243,0,77,0,208,0,0,0,93,0,179,0,175,0,8,0,0,0,240,0,17,0,102,0,109,0,68,0,0,0,209,0,78,0,108,0,41,0,0,0,0,0,186,0,235,0,183,0,224,0,0,0,118,0,0,0,96,0,77,0,111,0,34,0,171,0,175,0,241,0,190,0,246,0,0,0,216,0,83,0,0,0,0,0,164,0,216,0,178,0,200,0,219,0,30,0,0,0,39,0,139,0,57,0,121,0,80,0,6,0,244,0,0,0,96,0,0,0,26,0,203,0,16,0,79,0,15,0,195,0,0,0,0,0,0,0,243,0,109,0,179,0,144,0,76,0,0,0,254,0,61,0,84,0,0,0,168,0,150,0,14,0,165,0,138,0,65,0,218,0,34,0,230,0,19,0,4,0,0,0,14,0,12,0,104,0,54,0,225,0,180,0,0,0,0,0,89,0,158,0,219,0,55,0,29,0,19,0,96,0,144,0,186,0,102,0,175,0,37,0,182,0,0,0,0,0,0,0,0,0,14,0,3,0,155,0,240,0,95,0,199,0,104,0,247,0,36,0,222,0,153,0,0,0,129,0,0,0,106,0,64,0,0,0,169,0,236,0,69,0,100,0,9,0,101,0,102,0,239,0,0,0,166,0,0,0,160,0,149,0,135,0,58,0,0,0,191,0,28,0,77,0,192,0,231,0,234,0,214,0,217,0,156,0,79,0,33,0,86,0,165,0,77,0,210,0,163,0,241,0,0,0,85,0,249,0,7,0,252,0,66,0,216,0,2,0,248,0,244,0,250,0,253,0,133,0,88,0,91,0,0,0,104,0,0,0,148,0,172,0,227,0,219,0,0,0,133,0,73,0,0,0,85,0,177,0,35,0,111,0,68,0,175,0,42,0,138,0,33,0,95,0,12,0,61,0,122,0,133,0,0,0,151,0,0,0,167,0,0,0,117,0,85,0,0,0,114,0,54,0,230,0,97,0,71,0,121,0,39,0,8,0,254,0,194,0,238,0,20,0,239,0,185,0,148,0,179,0,228,0,168,0,2,0,0,0,188,0,0,0,110,0,153,0,87,0,0,0,120,0,142,0,62,0,224,0,44,0,245,0,137,0,133,0,72,0,17,0,155,0,233,0,79,0,17,0,31,0,223,0,143,0,222,0,0,0,0,0,15,0,0,0,37,0,249,0,121,0,0,0,82,0,223,0,48,0,245,0,0,0,7,0,22,0,32,0,129,0,95,0,13,0,0,0,50,0,196,0,0,0,157,0,75,0,0,0,4,0,27,0,61,0,146,0,83,0,246,0,52,0,254,0,144,0,212,0,239,0,186,0,48,0,176,0,19,0,213,0,0,0,115,0,164,0,148,0,115,0,0,0,233,0,145,0,189,0,195,0,67,0,95,0,105,0,207,0,24,0,91,0,239,0,98,0,90,0,14,0,164,0,72,0,181,0,249,0,210,0,0,0,233,0,107,0,94,0,0,0,138,0,198,0,134,0,2,0,231,0,144,0,26,0,27,0,43,0,142,0,225,0,34,0,42,0,241,0,140,0,115,0,139,0,160,0,117,0,127,0,230,0,109,0,173,0,51,0,51,0,116,0,174,0,67,0,208,0,14,0,0,0,194,0,110,0,0,0,158,0,165,0,5,0,160,0,134,0,0,0,137,0,186,0,199,0,253,0,0,0,114,0,35,0,220,0,114,0,187,0,19,0,98,0,132,0,39,0,176,0,208,0,186,0,250,0,162,0,35,0,161,0,168,0,0,0,29,0,0,0,62,0,164,0,0,0,205,0,249,0,34,0,159,0,150,0,28,0,91,0,9,0,102,0,28,0,86,0,48,0,7,0,0,0,166,0,187,0,0,0,116,0,44,0,171,0,77,0,169,0,0,0,145,0,145,0,190,0,107,0,16,0,89,0,180,0,68,0,82,0,19,0,7,0,148,0,40,0,86,0,120,0,0,0,139,0,6,0,43,0,126,0,4,0,186,0,111,0,0,0,77,0,143,0,27,0,137,0,0,0,82,0,49,0,225,0,34,0,88,0,81,0,203,0,18,0,171,0,95,0,69,0,68,0,0,0,148,0,0,0,52,0,0,0,114,0,211,0,44,0,128,0,160,0,114,0,107,0,229,0,0,0,159,0,0,0,37,0,0,0,148,0,215,0,253,0,122,0,170,0,144,0,207,0,183,0,230,0,226,0,159,0,83,0,142,0,131,0,240,0,174,0,72,0,247,0,191,0,64,0,72,0,131,0,0,0,41,0,255,0,254,0,170,0,13,0,150,0,188,0,138,0,218,0,0,0,237,0,96,0,230,0,22,0,44,0,160,0,239,0,51,0,207,0,201,0,122,0,186,0,155,0,59,0,28,0,112,0,53,0,0,0,36,0,67,0,109,0,0,0,49,0,176,0,0,0,4,0,222,0,229,0,85,0,231,0,148,0,233,0,179,0,47,0,64,0,139,0,89,0,79,0,19,0,241,0,204,0,86,0,124,0,0,0,0,0,20,0,91,0,43,0,0,0,138,0,0,0,36,0,0,0,159,0,97,0,237,0,0,0,53,0,147,0,148,0,215,0,149,0,191,0,211,0,0,0,191,0,139,0,27,0,210,0,25,0,191,0,102,0,0,0,227,0,173,0,231,0,172,0,249,0,218,0,145,0,217,0,0,0,156,0,0,0,29,0,180,0,192,0,204,0,21,0,223,0,236,0,0,0,102,0,84,0,79,0,247,0,12,0,182,0,231,0,0,0,128,0,236,0,157,0,250,0,181,0,189,0,147,0,7,0,130,0,136,0,116,0,163,0,179,0,73,0,123,0,73,0,97,0,231,0,85,0,90,0,78,0,0,0,18,0,94,0,165,0,0,0,0,0,24,0,36,0,0,0,6,0,141,0,8,0,243,0,125,0,250,0,83,0,221,0,32,0,164,0,141,0,143,0,0,0,166,0,9,0,112,0,0,0,196,0,62,0,247,0,213,0,8,0,84,0,212,0,0,0,0,0,66,0,121,0,24,0,18,0,0,0,206,0,199,0,0,0,0,0,136,0,0,0,0,0,132,0,113,0,99,0,178,0,153,0,225,0,8,0,151,0,148,0,189,0,5,0,93,0,0,0,230,0,136,0,59,0,0,0,247,0,0,0,191,0,133,0,243,0,116,0,218,0,190,0,222,0,246,0,232,0,135,0,41,0,161,0,0,0,240,0,121,0,81,0,213,0,30,0,0,0,103,0,174,0,160,0,0,0,3,0,30,0,0,0,239,0,199,0,121,0,0,0,0,0,0,0,255,0,164,0,29,0,100,0,98,0,172,0,37,0,178,0,222,0,239,0,168,0,0,0,104,0,16,0,231,0,203,0,132,0,0,0,128,0,23,0,165,0,39,0,154,0,59,0,13,0,91,0,0,0,54,0,214,0,211,0,8,0,151,0,31,0,109,0,0,0,0,0,69,0,48,0,84,0,250,0,142,0,157,0,84,0,149,0,88,0,113,0,0,0,57,0,132,0,251,0,87,0,0,0,25,0,134,0,10,0,141,0,31,0,0,0,255,0,0,0,166,0,0,0,229,0,0,0,124,0,0,0,198,0,0,0,193,0,9,0,189,0,60,0,0,0,206,0,68,0,89,0,53,0,6,0,147,0,0,0,170,0,94,0,91,0,70,0,147,0,216,0,69,0,7,0,159,0,54,0,133,0,0,0,133,0,0,0,0,0,235,0,13,0,112,0,158,0,35,0,72,0,251,0,130,0,0,0,23,0,115,0,0,0,39,0,117,0,103,0,234,0,41,0,0,0,127,0,205,0,187,0,72,0,66,0,21,0,0,0,97,0,107,0,180,0,0,0,26,0,2,0,25,0,25,0,66,0,179,0,191,0,0,0,118,0,168,0,83,0);
signal scenario_full  : scenario_type := (0,0,132,31,173,31,200,31,200,30,162,31,167,31,219,31,222,31,230,31,235,31,206,31,206,30,142,31,77,31,32,31,124,31,106,31,121,31,121,30,109,31,106,31,221,31,163,31,171,31,60,31,241,31,139,31,58,31,120,31,211,31,211,30,211,29,60,31,60,30,225,31,225,30,136,31,181,31,46,31,126,31,126,30,43,31,58,31,246,31,254,31,216,31,98,31,77,31,150,31,66,31,47,31,112,31,112,30,10,31,10,30,10,29,255,31,233,31,83,31,95,31,149,31,149,30,171,31,154,31,154,30,215,31,23,31,23,30,72,31,89,31,41,31,101,31,101,30,23,31,185,31,58,31,245,31,245,30,189,31,251,31,22,31,78,31,139,31,142,31,16,31,250,31,68,31,41,31,41,30,98,31,127,31,94,31,94,30,100,31,100,30,100,29,100,28,227,31,17,31,176,31,104,31,136,31,216,31,236,31,238,31,86,31,15,31,93,31,57,31,31,31,175,31,56,31,56,30,216,31,177,31,31,31,183,31,190,31,205,31,205,30,253,31,251,31,243,31,77,31,208,31,208,30,93,31,179,31,175,31,8,31,8,30,240,31,17,31,102,31,109,31,68,31,68,30,209,31,78,31,108,31,41,31,41,30,41,29,186,31,235,31,183,31,224,31,224,30,118,31,118,30,96,31,77,31,111,31,34,31,171,31,175,31,241,31,190,31,246,31,246,30,216,31,83,31,83,30,83,29,164,31,216,31,178,31,200,31,219,31,30,31,30,30,39,31,139,31,57,31,121,31,80,31,6,31,244,31,244,30,96,31,96,30,26,31,203,31,16,31,79,31,15,31,195,31,195,30,195,29,195,28,243,31,109,31,179,31,144,31,76,31,76,30,254,31,61,31,84,31,84,30,168,31,150,31,14,31,165,31,138,31,65,31,218,31,34,31,230,31,19,31,4,31,4,30,14,31,12,31,104,31,54,31,225,31,180,31,180,30,180,29,89,31,158,31,219,31,55,31,29,31,19,31,96,31,144,31,186,31,102,31,175,31,37,31,182,31,182,30,182,29,182,28,182,27,14,31,3,31,155,31,240,31,95,31,199,31,104,31,247,31,36,31,222,31,153,31,153,30,129,31,129,30,106,31,64,31,64,30,169,31,236,31,69,31,100,31,9,31,101,31,102,31,239,31,239,30,166,31,166,30,160,31,149,31,135,31,58,31,58,30,191,31,28,31,77,31,192,31,231,31,234,31,214,31,217,31,156,31,79,31,33,31,86,31,165,31,77,31,210,31,163,31,241,31,241,30,85,31,249,31,7,31,252,31,66,31,216,31,2,31,248,31,244,31,250,31,253,31,133,31,88,31,91,31,91,30,104,31,104,30,148,31,172,31,227,31,219,31,219,30,133,31,73,31,73,30,85,31,177,31,35,31,111,31,68,31,175,31,42,31,138,31,33,31,95,31,12,31,61,31,122,31,133,31,133,30,151,31,151,30,167,31,167,30,117,31,85,31,85,30,114,31,54,31,230,31,97,31,71,31,121,31,39,31,8,31,254,31,194,31,238,31,20,31,239,31,185,31,148,31,179,31,228,31,168,31,2,31,2,30,188,31,188,30,110,31,153,31,87,31,87,30,120,31,142,31,62,31,224,31,44,31,245,31,137,31,133,31,72,31,17,31,155,31,233,31,79,31,17,31,31,31,223,31,143,31,222,31,222,30,222,29,15,31,15,30,37,31,249,31,121,31,121,30,82,31,223,31,48,31,245,31,245,30,7,31,22,31,32,31,129,31,95,31,13,31,13,30,50,31,196,31,196,30,157,31,75,31,75,30,4,31,27,31,61,31,146,31,83,31,246,31,52,31,254,31,144,31,212,31,239,31,186,31,48,31,176,31,19,31,213,31,213,30,115,31,164,31,148,31,115,31,115,30,233,31,145,31,189,31,195,31,67,31,95,31,105,31,207,31,24,31,91,31,239,31,98,31,90,31,14,31,164,31,72,31,181,31,249,31,210,31,210,30,233,31,107,31,94,31,94,30,138,31,198,31,134,31,2,31,231,31,144,31,26,31,27,31,43,31,142,31,225,31,34,31,42,31,241,31,140,31,115,31,139,31,160,31,117,31,127,31,230,31,109,31,173,31,51,31,51,31,116,31,174,31,67,31,208,31,14,31,14,30,194,31,110,31,110,30,158,31,165,31,5,31,160,31,134,31,134,30,137,31,186,31,199,31,253,31,253,30,114,31,35,31,220,31,114,31,187,31,19,31,98,31,132,31,39,31,176,31,208,31,186,31,250,31,162,31,35,31,161,31,168,31,168,30,29,31,29,30,62,31,164,31,164,30,205,31,249,31,34,31,159,31,150,31,28,31,91,31,9,31,102,31,28,31,86,31,48,31,7,31,7,30,166,31,187,31,187,30,116,31,44,31,171,31,77,31,169,31,169,30,145,31,145,31,190,31,107,31,16,31,89,31,180,31,68,31,82,31,19,31,7,31,148,31,40,31,86,31,120,31,120,30,139,31,6,31,43,31,126,31,4,31,186,31,111,31,111,30,77,31,143,31,27,31,137,31,137,30,82,31,49,31,225,31,34,31,88,31,81,31,203,31,18,31,171,31,95,31,69,31,68,31,68,30,148,31,148,30,52,31,52,30,114,31,211,31,44,31,128,31,160,31,114,31,107,31,229,31,229,30,159,31,159,30,37,31,37,30,148,31,215,31,253,31,122,31,170,31,144,31,207,31,183,31,230,31,226,31,159,31,83,31,142,31,131,31,240,31,174,31,72,31,247,31,191,31,64,31,72,31,131,31,131,30,41,31,255,31,254,31,170,31,13,31,150,31,188,31,138,31,218,31,218,30,237,31,96,31,230,31,22,31,44,31,160,31,239,31,51,31,207,31,201,31,122,31,186,31,155,31,59,31,28,31,112,31,53,31,53,30,36,31,67,31,109,31,109,30,49,31,176,31,176,30,4,31,222,31,229,31,85,31,231,31,148,31,233,31,179,31,47,31,64,31,139,31,89,31,79,31,19,31,241,31,204,31,86,31,124,31,124,30,124,29,20,31,91,31,43,31,43,30,138,31,138,30,36,31,36,30,159,31,97,31,237,31,237,30,53,31,147,31,148,31,215,31,149,31,191,31,211,31,211,30,191,31,139,31,27,31,210,31,25,31,191,31,102,31,102,30,227,31,173,31,231,31,172,31,249,31,218,31,145,31,217,31,217,30,156,31,156,30,29,31,180,31,192,31,204,31,21,31,223,31,236,31,236,30,102,31,84,31,79,31,247,31,12,31,182,31,231,31,231,30,128,31,236,31,157,31,250,31,181,31,189,31,147,31,7,31,130,31,136,31,116,31,163,31,179,31,73,31,123,31,73,31,97,31,231,31,85,31,90,31,78,31,78,30,18,31,94,31,165,31,165,30,165,29,24,31,36,31,36,30,6,31,141,31,8,31,243,31,125,31,250,31,83,31,221,31,32,31,164,31,141,31,143,31,143,30,166,31,9,31,112,31,112,30,196,31,62,31,247,31,213,31,8,31,84,31,212,31,212,30,212,29,66,31,121,31,24,31,18,31,18,30,206,31,199,31,199,30,199,29,136,31,136,30,136,29,132,31,113,31,99,31,178,31,153,31,225,31,8,31,151,31,148,31,189,31,5,31,93,31,93,30,230,31,136,31,59,31,59,30,247,31,247,30,191,31,133,31,243,31,116,31,218,31,190,31,222,31,246,31,232,31,135,31,41,31,161,31,161,30,240,31,121,31,81,31,213,31,30,31,30,30,103,31,174,31,160,31,160,30,3,31,30,31,30,30,239,31,199,31,121,31,121,30,121,29,121,28,255,31,164,31,29,31,100,31,98,31,172,31,37,31,178,31,222,31,239,31,168,31,168,30,104,31,16,31,231,31,203,31,132,31,132,30,128,31,23,31,165,31,39,31,154,31,59,31,13,31,91,31,91,30,54,31,214,31,211,31,8,31,151,31,31,31,109,31,109,30,109,29,69,31,48,31,84,31,250,31,142,31,157,31,84,31,149,31,88,31,113,31,113,30,57,31,132,31,251,31,87,31,87,30,25,31,134,31,10,31,141,31,31,31,31,30,255,31,255,30,166,31,166,30,229,31,229,30,124,31,124,30,198,31,198,30,193,31,9,31,189,31,60,31,60,30,206,31,68,31,89,31,53,31,6,31,147,31,147,30,170,31,94,31,91,31,70,31,147,31,216,31,69,31,7,31,159,31,54,31,133,31,133,30,133,31,133,30,133,29,235,31,13,31,112,31,158,31,35,31,72,31,251,31,130,31,130,30,23,31,115,31,115,30,39,31,117,31,103,31,234,31,41,31,41,30,127,31,205,31,187,31,72,31,66,31,21,31,21,30,97,31,107,31,180,31,180,30,26,31,2,31,25,31,25,31,66,31,179,31,191,31,191,30,118,31,168,31,83,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
