-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1017;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,232,0,229,0,69,0,235,0,251,0,14,0,175,0,167,0,0,0,23,0,80,0,80,0,0,0,0,0,184,0,0,0,178,0,233,0,115,0,181,0,25,0,71,0,230,0,206,0,215,0,0,0,169,0,255,0,0,0,165,0,0,0,145,0,47,0,15,0,76,0,238,0,5,0,98,0,0,0,145,0,13,0,0,0,240,0,0,0,0,0,0,0,170,0,120,0,102,0,110,0,0,0,217,0,134,0,0,0,123,0,199,0,0,0,81,0,81,0,178,0,98,0,58,0,140,0,77,0,96,0,25,0,132,0,253,0,208,0,89,0,88,0,84,0,243,0,0,0,213,0,0,0,183,0,0,0,51,0,109,0,0,0,146,0,59,0,199,0,195,0,50,0,199,0,241,0,0,0,129,0,5,0,40,0,121,0,183,0,83,0,28,0,127,0,0,0,27,0,98,0,107,0,175,0,59,0,0,0,0,0,140,0,0,0,139,0,0,0,45,0,1,0,175,0,109,0,220,0,194,0,186,0,204,0,5,0,0,0,98,0,223,0,70,0,96,0,162,0,0,0,0,0,187,0,151,0,31,0,9,0,23,0,40,0,229,0,52,0,34,0,0,0,0,0,184,0,174,0,221,0,1,0,135,0,89,0,11,0,176,0,71,0,161,0,243,0,254,0,143,0,41,0,79,0,177,0,48,0,132,0,219,0,0,0,229,0,3,0,84,0,212,0,229,0,214,0,191,0,21,0,0,0,205,0,154,0,0,0,12,0,63,0,208,0,89,0,223,0,80,0,0,0,0,0,220,0,197,0,98,0,95,0,173,0,26,0,188,0,59,0,220,0,232,0,139,0,185,0,132,0,0,0,34,0,0,0,150,0,0,0,0,0,0,0,0,0,68,0,112,0,17,0,95,0,184,0,242,0,0,0,0,0,0,0,211,0,161,0,31,0,0,0,145,0,0,0,40,0,240,0,0,0,146,0,90,0,0,0,177,0,11,0,41,0,24,0,0,0,179,0,244,0,137,0,0,0,0,0,0,0,0,0,151,0,14,0,80,0,73,0,240,0,0,0,71,0,159,0,0,0,206,0,0,0,13,0,2,0,167,0,0,0,0,0,241,0,85,0,0,0,236,0,163,0,0,0,0,0,51,0,0,0,114,0,173,0,146,0,139,0,145,0,79,0,151,0,191,0,53,0,108,0,0,0,82,0,0,0,183,0,20,0,176,0,231,0,133,0,158,0,0,0,62,0,247,0,171,0,246,0,61,0,181,0,0,0,15,0,31,0,138,0,146,0,123,0,175,0,0,0,53,0,116,0,205,0,0,0,44,0,0,0,124,0,0,0,121,0,66,0,234,0,0,0,50,0,176,0,95,0,0,0,70,0,215,0,184,0,0,0,0,0,199,0,37,0,208,0,0,0,60,0,0,0,119,0,148,0,0,0,57,0,141,0,228,0,0,0,177,0,121,0,90,0,0,0,26,0,0,0,0,0,28,0,58,0,154,0,0,0,82,0,0,0,0,0,221,0,28,0,38,0,89,0,44,0,69,0,111,0,180,0,13,0,94,0,70,0,233,0,207,0,115,0,131,0,57,0,60,0,45,0,0,0,143,0,179,0,77,0,144,0,10,0,248,0,35,0,0,0,0,0,254,0,39,0,0,0,242,0,30,0,127,0,138,0,134,0,67,0,84,0,0,0,42,0,231,0,174,0,0,0,116,0,189,0,25,0,109,0,219,0,0,0,0,0,206,0,234,0,116,0,212,0,43,0,93,0,141,0,242,0,238,0,62,0,208,0,0,0,89,0,233,0,0,0,9,0,0,0,210,0,79,0,0,0,0,0,51,0,33,0,129,0,0,0,16,0,234,0,92,0,34,0,0,0,245,0,197,0,25,0,195,0,0,0,158,0,16,0,20,0,0,0,223,0,25,0,0,0,179,0,163,0,240,0,8,0,237,0,23,0,0,0,221,0,0,0,194,0,199,0,199,0,132,0,192,0,80,0,0,0,40,0,100,0,45,0,150,0,0,0,104,0,57,0,250,0,58,0,91,0,159,0,236,0,183,0,131,0,51,0,225,0,58,0,80,0,0,0,208,0,76,0,90,0,222,0,0,0,142,0,48,0,59,0,15,0,1,0,195,0,38,0,101,0,0,0,45,0,95,0,0,0,235,0,131,0,206,0,218,0,148,0,34,0,38,0,244,0,214,0,0,0,152,0,126,0,42,0,3,0,132,0,23,0,103,0,43,0,227,0,37,0,66,0,60,0,49,0,174,0,235,0,0,0,207,0,17,0,114,0,82,0,0,0,215,0,0,0,67,0,0,0,3,0,40,0,40,0,0,0,31,0,159,0,60,0,190,0,238,0,243,0,118,0,30,0,197,0,0,0,34,0,0,0,25,0,132,0,51,0,22,0,196,0,239,0,0,0,168,0,169,0,144,0,0,0,0,0,78,0,0,0,0,0,248,0,204,0,8,0,237,0,125,0,37,0,198,0,15,0,0,0,0,0,140,0,54,0,198,0,38,0,98,0,111,0,239,0,0,0,138,0,31,0,68,0,190,0,0,0,0,0,172,0,189,0,84,0,21,0,2,0,0,0,40,0,232,0,89,0,0,0,73,0,0,0,75,0,216,0,51,0,28,0,0,0,0,0,0,0,142,0,95,0,104,0,35,0,0,0,166,0,241,0,4,0,131,0,20,0,241,0,247,0,56,0,48,0,168,0,237,0,21,0,200,0,101,0,11,0,118,0,13,0,217,0,250,0,0,0,140,0,7,0,154,0,0,0,79,0,92,0,0,0,101,0,180,0,135,0,7,0,48,0,35,0,222,0,141,0,136,0,5,0,110,0,0,0,0,0,0,0,159,0,78,0,50,0,68,0,35,0,0,0,7,0,146,0,239,0,94,0,0,0,25,0,237,0,42,0,85,0,203,0,145,0,243,0,174,0,240,0,79,0,35,0,184,0,0,0,0,0,155,0,126,0,228,0,95,0,92,0,229,0,216,0,151,0,210,0,213,0,68,0,3,0,182,0,0,0,34,0,208,0,217,0,17,0,236,0,127,0,0,0,2,0,42,0,189,0,242,0,97,0,245,0,106,0,5,0,25,0,94,0,114,0,197,0,0,0,0,0,248,0,77,0,60,0,116,0,222,0,37,0,182,0,199,0,125,0,222,0,0,0,151,0,211,0,205,0,7,0,228,0,0,0,0,0,1,0,83,0,244,0,8,0,194,0,21,0,178,0,0,0,20,0,101,0,194,0,0,0,244,0,176,0,95,0,240,0,183,0,128,0,26,0,40,0,243,0,94,0,51,0,0,0,6,0,244,0,237,0,19,0,0,0,242,0,221,0,4,0,9,0,168,0,142,0,208,0,0,0,112,0,0,0,0,0,187,0,177,0,134,0,178,0,92,0,0,0,0,0,183,0,144,0,123,0,84,0,0,0,0,0,95,0,88,0,24,0,143,0,51,0,151,0,214,0,66,0,114,0,142,0,0,0,73,0,41,0,44,0,0,0,52,0,102,0,198,0,197,0,17,0,126,0,51,0,4,0,230,0,81,0,25,0,102,0,233,0,141,0,53,0,209,0,65,0,114,0,204,0,0,0,101,0,205,0,160,0,0,0,193,0,183,0,181,0,122,0,91,0,0,0,0,0,238,0,162,0,128,0,0,0,107,0,101,0,210,0,90,0,241,0,0,0,122,0,167,0,161,0,166,0,170,0,16,0,0,0,218,0,0,0,0,0,157,0,0,0,239,0,243,0,0,0,227,0,176,0,145,0,0,0,210,0,128,0,8,0,230,0,190,0,57,0,4,0,114,0,27,0,126,0,3,0,220,0,114,0,100,0,0,0,9,0,212,0,34,0,209,0,248,0,62,0,67,0,90,0,136,0,10,0,185,0,7,0,0,0,177,0,236,0,192,0,75,0,12,0,0,0,35,0,0,0,23,0,0,0,143,0,0,0,0,0,29,0,0,0,217,0,154,0,105,0,24,0,0,0,248,0,21,0,76,0,29,0,176,0,5,0,0,0,167,0,209,0,155,0,0,0,64,0,136,0,29,0,0,0,106,0,4,0,65,0,101,0,191,0,246,0,229,0,89,0,57,0,194,0,146,0,0,0,247,0,67,0,31,0,109,0,98,0,151,0,215,0,79,0,25,0,64,0,169,0,230,0,55,0,86,0,88,0,5,0,117,0,1,0,223,0,138,0,254,0,143,0,0,0,202,0,158,0,189,0,0,0,0,0,99,0,200,0,241,0,159,0,0,0,127,0,0,0,195,0,217,0,167,0,162,0,142,0,177,0,0,0,202,0,94,0,0,0,0,0,83,0,253,0,6,0,105,0,0,0,250,0,0,0,131,0,168,0,24,0,150,0,6,0,34,0,228,0,214,0,92,0,144,0,166,0,0,0,0,0,151,0,0,0,0,0,55,0,0,0,182,0,159,0,226,0,160,0,175,0,145,0,0,0,245,0,22,0,0,0,40,0,163,0,141,0,0,0,104,0,1,0,82,0,202,0,138,0,149,0,202,0,123,0,0,0,50,0,82,0,3,0,49,0);
signal scenario_full  : scenario_type := (0,0,232,31,229,31,69,31,235,31,251,31,14,31,175,31,167,31,167,30,23,31,80,31,80,31,80,30,80,29,184,31,184,30,178,31,233,31,115,31,181,31,25,31,71,31,230,31,206,31,215,31,215,30,169,31,255,31,255,30,165,31,165,30,145,31,47,31,15,31,76,31,238,31,5,31,98,31,98,30,145,31,13,31,13,30,240,31,240,30,240,29,240,28,170,31,120,31,102,31,110,31,110,30,217,31,134,31,134,30,123,31,199,31,199,30,81,31,81,31,178,31,98,31,58,31,140,31,77,31,96,31,25,31,132,31,253,31,208,31,89,31,88,31,84,31,243,31,243,30,213,31,213,30,183,31,183,30,51,31,109,31,109,30,146,31,59,31,199,31,195,31,50,31,199,31,241,31,241,30,129,31,5,31,40,31,121,31,183,31,83,31,28,31,127,31,127,30,27,31,98,31,107,31,175,31,59,31,59,30,59,29,140,31,140,30,139,31,139,30,45,31,1,31,175,31,109,31,220,31,194,31,186,31,204,31,5,31,5,30,98,31,223,31,70,31,96,31,162,31,162,30,162,29,187,31,151,31,31,31,9,31,23,31,40,31,229,31,52,31,34,31,34,30,34,29,184,31,174,31,221,31,1,31,135,31,89,31,11,31,176,31,71,31,161,31,243,31,254,31,143,31,41,31,79,31,177,31,48,31,132,31,219,31,219,30,229,31,3,31,84,31,212,31,229,31,214,31,191,31,21,31,21,30,205,31,154,31,154,30,12,31,63,31,208,31,89,31,223,31,80,31,80,30,80,29,220,31,197,31,98,31,95,31,173,31,26,31,188,31,59,31,220,31,232,31,139,31,185,31,132,31,132,30,34,31,34,30,150,31,150,30,150,29,150,28,150,27,68,31,112,31,17,31,95,31,184,31,242,31,242,30,242,29,242,28,211,31,161,31,31,31,31,30,145,31,145,30,40,31,240,31,240,30,146,31,90,31,90,30,177,31,11,31,41,31,24,31,24,30,179,31,244,31,137,31,137,30,137,29,137,28,137,27,151,31,14,31,80,31,73,31,240,31,240,30,71,31,159,31,159,30,206,31,206,30,13,31,2,31,167,31,167,30,167,29,241,31,85,31,85,30,236,31,163,31,163,30,163,29,51,31,51,30,114,31,173,31,146,31,139,31,145,31,79,31,151,31,191,31,53,31,108,31,108,30,82,31,82,30,183,31,20,31,176,31,231,31,133,31,158,31,158,30,62,31,247,31,171,31,246,31,61,31,181,31,181,30,15,31,31,31,138,31,146,31,123,31,175,31,175,30,53,31,116,31,205,31,205,30,44,31,44,30,124,31,124,30,121,31,66,31,234,31,234,30,50,31,176,31,95,31,95,30,70,31,215,31,184,31,184,30,184,29,199,31,37,31,208,31,208,30,60,31,60,30,119,31,148,31,148,30,57,31,141,31,228,31,228,30,177,31,121,31,90,31,90,30,26,31,26,30,26,29,28,31,58,31,154,31,154,30,82,31,82,30,82,29,221,31,28,31,38,31,89,31,44,31,69,31,111,31,180,31,13,31,94,31,70,31,233,31,207,31,115,31,131,31,57,31,60,31,45,31,45,30,143,31,179,31,77,31,144,31,10,31,248,31,35,31,35,30,35,29,254,31,39,31,39,30,242,31,30,31,127,31,138,31,134,31,67,31,84,31,84,30,42,31,231,31,174,31,174,30,116,31,189,31,25,31,109,31,219,31,219,30,219,29,206,31,234,31,116,31,212,31,43,31,93,31,141,31,242,31,238,31,62,31,208,31,208,30,89,31,233,31,233,30,9,31,9,30,210,31,79,31,79,30,79,29,51,31,33,31,129,31,129,30,16,31,234,31,92,31,34,31,34,30,245,31,197,31,25,31,195,31,195,30,158,31,16,31,20,31,20,30,223,31,25,31,25,30,179,31,163,31,240,31,8,31,237,31,23,31,23,30,221,31,221,30,194,31,199,31,199,31,132,31,192,31,80,31,80,30,40,31,100,31,45,31,150,31,150,30,104,31,57,31,250,31,58,31,91,31,159,31,236,31,183,31,131,31,51,31,225,31,58,31,80,31,80,30,208,31,76,31,90,31,222,31,222,30,142,31,48,31,59,31,15,31,1,31,195,31,38,31,101,31,101,30,45,31,95,31,95,30,235,31,131,31,206,31,218,31,148,31,34,31,38,31,244,31,214,31,214,30,152,31,126,31,42,31,3,31,132,31,23,31,103,31,43,31,227,31,37,31,66,31,60,31,49,31,174,31,235,31,235,30,207,31,17,31,114,31,82,31,82,30,215,31,215,30,67,31,67,30,3,31,40,31,40,31,40,30,31,31,159,31,60,31,190,31,238,31,243,31,118,31,30,31,197,31,197,30,34,31,34,30,25,31,132,31,51,31,22,31,196,31,239,31,239,30,168,31,169,31,144,31,144,30,144,29,78,31,78,30,78,29,248,31,204,31,8,31,237,31,125,31,37,31,198,31,15,31,15,30,15,29,140,31,54,31,198,31,38,31,98,31,111,31,239,31,239,30,138,31,31,31,68,31,190,31,190,30,190,29,172,31,189,31,84,31,21,31,2,31,2,30,40,31,232,31,89,31,89,30,73,31,73,30,75,31,216,31,51,31,28,31,28,30,28,29,28,28,142,31,95,31,104,31,35,31,35,30,166,31,241,31,4,31,131,31,20,31,241,31,247,31,56,31,48,31,168,31,237,31,21,31,200,31,101,31,11,31,118,31,13,31,217,31,250,31,250,30,140,31,7,31,154,31,154,30,79,31,92,31,92,30,101,31,180,31,135,31,7,31,48,31,35,31,222,31,141,31,136,31,5,31,110,31,110,30,110,29,110,28,159,31,78,31,50,31,68,31,35,31,35,30,7,31,146,31,239,31,94,31,94,30,25,31,237,31,42,31,85,31,203,31,145,31,243,31,174,31,240,31,79,31,35,31,184,31,184,30,184,29,155,31,126,31,228,31,95,31,92,31,229,31,216,31,151,31,210,31,213,31,68,31,3,31,182,31,182,30,34,31,208,31,217,31,17,31,236,31,127,31,127,30,2,31,42,31,189,31,242,31,97,31,245,31,106,31,5,31,25,31,94,31,114,31,197,31,197,30,197,29,248,31,77,31,60,31,116,31,222,31,37,31,182,31,199,31,125,31,222,31,222,30,151,31,211,31,205,31,7,31,228,31,228,30,228,29,1,31,83,31,244,31,8,31,194,31,21,31,178,31,178,30,20,31,101,31,194,31,194,30,244,31,176,31,95,31,240,31,183,31,128,31,26,31,40,31,243,31,94,31,51,31,51,30,6,31,244,31,237,31,19,31,19,30,242,31,221,31,4,31,9,31,168,31,142,31,208,31,208,30,112,31,112,30,112,29,187,31,177,31,134,31,178,31,92,31,92,30,92,29,183,31,144,31,123,31,84,31,84,30,84,29,95,31,88,31,24,31,143,31,51,31,151,31,214,31,66,31,114,31,142,31,142,30,73,31,41,31,44,31,44,30,52,31,102,31,198,31,197,31,17,31,126,31,51,31,4,31,230,31,81,31,25,31,102,31,233,31,141,31,53,31,209,31,65,31,114,31,204,31,204,30,101,31,205,31,160,31,160,30,193,31,183,31,181,31,122,31,91,31,91,30,91,29,238,31,162,31,128,31,128,30,107,31,101,31,210,31,90,31,241,31,241,30,122,31,167,31,161,31,166,31,170,31,16,31,16,30,218,31,218,30,218,29,157,31,157,30,239,31,243,31,243,30,227,31,176,31,145,31,145,30,210,31,128,31,8,31,230,31,190,31,57,31,4,31,114,31,27,31,126,31,3,31,220,31,114,31,100,31,100,30,9,31,212,31,34,31,209,31,248,31,62,31,67,31,90,31,136,31,10,31,185,31,7,31,7,30,177,31,236,31,192,31,75,31,12,31,12,30,35,31,35,30,23,31,23,30,143,31,143,30,143,29,29,31,29,30,217,31,154,31,105,31,24,31,24,30,248,31,21,31,76,31,29,31,176,31,5,31,5,30,167,31,209,31,155,31,155,30,64,31,136,31,29,31,29,30,106,31,4,31,65,31,101,31,191,31,246,31,229,31,89,31,57,31,194,31,146,31,146,30,247,31,67,31,31,31,109,31,98,31,151,31,215,31,79,31,25,31,64,31,169,31,230,31,55,31,86,31,88,31,5,31,117,31,1,31,223,31,138,31,254,31,143,31,143,30,202,31,158,31,189,31,189,30,189,29,99,31,200,31,241,31,159,31,159,30,127,31,127,30,195,31,217,31,167,31,162,31,142,31,177,31,177,30,202,31,94,31,94,30,94,29,83,31,253,31,6,31,105,31,105,30,250,31,250,30,131,31,168,31,24,31,150,31,6,31,34,31,228,31,214,31,92,31,144,31,166,31,166,30,166,29,151,31,151,30,151,29,55,31,55,30,182,31,159,31,226,31,160,31,175,31,145,31,145,30,245,31,22,31,22,30,40,31,163,31,141,31,141,30,104,31,1,31,82,31,202,31,138,31,149,31,202,31,123,31,123,30,50,31,82,31,3,31,49,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
