-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 358;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,205,0,19,0,229,0,132,0,0,0,82,0,0,0,116,0,157,0,197,0,112,0,0,0,10,0,159,0,6,0,165,0,70,0,46,0,139,0,129,0,199,0,228,0,15,0,4,0,22,0,13,0,33,0,100,0,156,0,113,0,180,0,0,0,0,0,180,0,217,0,254,0,130,0,197,0,15,0,0,0,30,0,0,0,201,0,118,0,21,0,45,0,0,0,208,0,2,0,0,0,67,0,176,0,202,0,44,0,0,0,33,0,182,0,0,0,0,0,250,0,0,0,64,0,126,0,18,0,6,0,114,0,234,0,28,0,215,0,1,0,234,0,220,0,188,0,190,0,232,0,252,0,117,0,176,0,181,0,114,0,89,0,0,0,6,0,84,0,10,0,72,0,123,0,55,0,205,0,0,0,155,0,106,0,174,0,41,0,27,0,85,0,147,0,39,0,38,0,26,0,0,0,114,0,0,0,25,0,0,0,102,0,30,0,226,0,123,0,215,0,194,0,2,0,49,0,32,0,162,0,89,0,166,0,164,0,218,0,146,0,190,0,110,0,22,0,0,0,244,0,1,0,142,0,47,0,137,0,0,0,0,0,127,0,101,0,205,0,0,0,0,0,230,0,100,0,0,0,181,0,0,0,56,0,183,0,43,0,193,0,117,0,53,0,110,0,192,0,0,0,45,0,57,0,172,0,59,0,167,0,0,0,203,0,198,0,162,0,118,0,228,0,140,0,0,0,112,0,236,0,132,0,193,0,60,0,0,0,208,0,105,0,0,0,5,0,217,0,228,0,165,0,101,0,252,0,251,0,99,0,174,0,95,0,110,0,96,0,0,0,136,0,227,0,51,0,91,0,0,0,0,0,92,0,0,0,156,0,82,0,146,0,0,0,228,0,202,0,55,0,155,0,100,0,60,0,100,0,79,0,56,0,32,0,207,0,186,0,0,0,179,0,175,0,231,0,125,0,68,0,114,0,76,0,226,0,127,0,0,0,130,0,234,0,91,0,148,0,0,0,94,0,87,0,0,0,26,0,0,0,0,0,124,0,156,0,64,0,14,0,173,0,124,0,85,0,169,0,51,0,249,0,195,0,0,0,137,0,9,0,183,0,207,0,13,0,40,0,93,0,254,0,0,0,246,0,101,0,217,0,138,0,215,0,147,0,0,0,51,0,14,0,243,0,40,0,88,0,22,0,229,0,127,0,109,0,12,0,223,0,195,0,197,0,138,0,0,0,58,0,94,0,254,0,4,0,100,0,180,0,0,0,53,0,52,0,215,0,159,0,0,0,202,0,129,0,0,0,24,0,175,0,0,0,0,0,44,0,165,0,71,0,0,0,72,0,137,0,0,0,3,0,0,0,0,0,46,0,10,0,154,0,82,0,213,0,21,0,47,0,230,0,249,0,99,0,219,0,229,0,214,0,46,0,249,0,47,0,75,0,102,0,56,0,77,0,0,0,26,0,161,0,10,0,189,0,20,0,40,0,148,0,241,0,128,0,162,0,17,0,183,0,63,0,102,0,17,0,0,0,202,0,8,0,98,0,189,0,110,0,0,0,141,0,154,0,193,0,117,0,115,0,0,0,86,0,117,0,218,0,0,0,81,0);
signal scenario_full  : scenario_type := (69,31,205,31,19,31,229,31,132,31,132,30,82,31,82,30,116,31,157,31,197,31,112,31,112,30,10,31,159,31,6,31,165,31,70,31,46,31,139,31,129,31,199,31,228,31,15,31,4,31,22,31,13,31,33,31,100,31,156,31,113,31,180,31,180,30,180,29,180,31,217,31,254,31,130,31,197,31,15,31,15,30,30,31,30,30,201,31,118,31,21,31,45,31,45,30,208,31,2,31,2,30,67,31,176,31,202,31,44,31,44,30,33,31,182,31,182,30,182,29,250,31,250,30,64,31,126,31,18,31,6,31,114,31,234,31,28,31,215,31,1,31,234,31,220,31,188,31,190,31,232,31,252,31,117,31,176,31,181,31,114,31,89,31,89,30,6,31,84,31,10,31,72,31,123,31,55,31,205,31,205,30,155,31,106,31,174,31,41,31,27,31,85,31,147,31,39,31,38,31,26,31,26,30,114,31,114,30,25,31,25,30,102,31,30,31,226,31,123,31,215,31,194,31,2,31,49,31,32,31,162,31,89,31,166,31,164,31,218,31,146,31,190,31,110,31,22,31,22,30,244,31,1,31,142,31,47,31,137,31,137,30,137,29,127,31,101,31,205,31,205,30,205,29,230,31,100,31,100,30,181,31,181,30,56,31,183,31,43,31,193,31,117,31,53,31,110,31,192,31,192,30,45,31,57,31,172,31,59,31,167,31,167,30,203,31,198,31,162,31,118,31,228,31,140,31,140,30,112,31,236,31,132,31,193,31,60,31,60,30,208,31,105,31,105,30,5,31,217,31,228,31,165,31,101,31,252,31,251,31,99,31,174,31,95,31,110,31,96,31,96,30,136,31,227,31,51,31,91,31,91,30,91,29,92,31,92,30,156,31,82,31,146,31,146,30,228,31,202,31,55,31,155,31,100,31,60,31,100,31,79,31,56,31,32,31,207,31,186,31,186,30,179,31,175,31,231,31,125,31,68,31,114,31,76,31,226,31,127,31,127,30,130,31,234,31,91,31,148,31,148,30,94,31,87,31,87,30,26,31,26,30,26,29,124,31,156,31,64,31,14,31,173,31,124,31,85,31,169,31,51,31,249,31,195,31,195,30,137,31,9,31,183,31,207,31,13,31,40,31,93,31,254,31,254,30,246,31,101,31,217,31,138,31,215,31,147,31,147,30,51,31,14,31,243,31,40,31,88,31,22,31,229,31,127,31,109,31,12,31,223,31,195,31,197,31,138,31,138,30,58,31,94,31,254,31,4,31,100,31,180,31,180,30,53,31,52,31,215,31,159,31,159,30,202,31,129,31,129,30,24,31,175,31,175,30,175,29,44,31,165,31,71,31,71,30,72,31,137,31,137,30,3,31,3,30,3,29,46,31,10,31,154,31,82,31,213,31,21,31,47,31,230,31,249,31,99,31,219,31,229,31,214,31,46,31,249,31,47,31,75,31,102,31,56,31,77,31,77,30,26,31,161,31,10,31,189,31,20,31,40,31,148,31,241,31,128,31,162,31,17,31,183,31,63,31,102,31,17,31,17,30,202,31,8,31,98,31,189,31,110,31,110,30,141,31,154,31,193,31,117,31,115,31,115,30,86,31,117,31,218,31,218,30,81,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
