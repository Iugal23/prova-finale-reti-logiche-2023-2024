-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 634;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (58,0,16,0,201,0,188,0,178,0,60,0,0,0,0,0,240,0,71,0,139,0,94,0,143,0,254,0,0,0,240,0,252,0,0,0,192,0,0,0,138,0,0,0,98,0,83,0,0,0,35,0,0,0,249,0,169,0,0,0,240,0,196,0,3,0,243,0,63,0,130,0,4,0,0,0,66,0,231,0,32,0,213,0,0,0,158,0,0,0,0,0,201,0,0,0,19,0,236,0,126,0,165,0,101,0,176,0,138,0,88,0,82,0,129,0,66,0,14,0,160,0,0,0,158,0,31,0,78,0,172,0,0,0,0,0,242,0,10,0,239,0,107,0,16,0,46,0,0,0,246,0,0,0,69,0,69,0,196,0,0,0,0,0,145,0,142,0,194,0,190,0,232,0,3,0,161,0,128,0,169,0,120,0,20,0,72,0,241,0,0,0,83,0,12,0,0,0,229,0,63,0,8,0,165,0,0,0,166,0,198,0,121,0,205,0,228,0,0,0,251,0,0,0,61,0,152,0,120,0,0,0,85,0,0,0,52,0,0,0,90,0,182,0,118,0,66,0,127,0,52,0,201,0,0,0,163,0,164,0,0,0,75,0,43,0,95,0,173,0,125,0,0,0,13,0,98,0,74,0,157,0,254,0,236,0,149,0,42,0,0,0,0,0,153,0,250,0,35,0,0,0,178,0,57,0,80,0,168,0,204,0,0,0,14,0,180,0,190,0,0,0,83,0,134,0,67,0,55,0,0,0,242,0,193,0,131,0,104,0,47,0,226,0,173,0,56,0,106,0,40,0,135,0,82,0,186,0,6,0,50,0,202,0,251,0,11,0,0,0,10,0,0,0,20,0,253,0,212,0,45,0,0,0,124,0,218,0,0,0,51,0,135,0,0,0,191,0,0,0,107,0,246,0,0,0,111,0,177,0,241,0,178,0,0,0,129,0,0,0,179,0,0,0,0,0,204,0,138,0,111,0,225,0,208,0,0,0,35,0,116,0,61,0,212,0,23,0,219,0,75,0,0,0,17,0,196,0,21,0,0,0,50,0,76,0,171,0,3,0,79,0,154,0,0,0,0,0,246,0,250,0,151,0,103,0,84,0,33,0,72,0,230,0,0,0,0,0,124,0,200,0,0,0,168,0,103,0,0,0,0,0,245,0,129,0,197,0,3,0,123,0,0,0,252,0,0,0,185,0,156,0,82,0,147,0,0,0,123,0,192,0,91,0,0,0,46,0,0,0,180,0,0,0,216,0,0,0,165,0,157,0,187,0,189,0,0,0,251,0,174,0,121,0,154,0,151,0,0,0,0,0,36,0,0,0,0,0,90,0,210,0,37,0,251,0,3,0,0,0,152,0,141,0,162,0,50,0,251,0,79,0,0,0,98,0,0,0,140,0,85,0,100,0,226,0,14,0,186,0,166,0,23,0,187,0,186,0,0,0,180,0,24,0,196,0,0,0,0,0,34,0,30,0,40,0,80,0,253,0,60,0,30,0,127,0,129,0,0,0,0,0,0,0,38,0,0,0,0,0,117,0,119,0,25,0,174,0,22,0,186,0,143,0,232,0,0,0,122,0,7,0,113,0,9,0,191,0,177,0,94,0,153,0,10,0,189,0,105,0,54,0,114,0,52,0,107,0,79,0,0,0,169,0,227,0,101,0,5,0,16,0,0,0,120,0,171,0,77,0,6,0,0,0,48,0,157,0,220,0,215,0,0,0,138,0,0,0,159,0,32,0,221,0,0,0,218,0,197,0,3,0,248,0,0,0,240,0,145,0,191,0,0,0,11,0,255,0,58,0,0,0,181,0,110,0,104,0,109,0,99,0,105,0,181,0,102,0,244,0,79,0,156,0,13,0,0,0,0,0,235,0,108,0,143,0,189,0,168,0,14,0,176,0,58,0,39,0,215,0,108,0,79,0,0,0,85,0,0,0,157,0,89,0,76,0,0,0,233,0,167,0,0,0,233,0,93,0,143,0,118,0,0,0,251,0,113,0,45,0,124,0,183,0,176,0,153,0,229,0,221,0,160,0,70,0,18,0,139,0,77,0,94,0,0,0,80,0,133,0,246,0,141,0,168,0,0,0,0,0,231,0,187,0,82,0,216,0,0,0,163,0,237,0,12,0,95,0,0,0,165,0,81,0,0,0,101,0,62,0,28,0,135,0,120,0,209,0,0,0,99,0,107,0,202,0,27,0,0,0,142,0,0,0,101,0,0,0,227,0,0,0,83,0,0,0,0,0,112,0,54,0,52,0,0,0,19,0,137,0,0,0,113,0,240,0,229,0,94,0,195,0,220,0,247,0,86,0,226,0,1,0,0,0,44,0,38,0,194,0,208,0,96,0,42,0,100,0,0,0,252,0,97,0,0,0,88,0,0,0,0,0,71,0,117,0,74,0,91,0,224,0,0,0,199,0,153,0,69,0,218,0,118,0,89,0,0,0,192,0,134,0,181,0,147,0,231,0,254,0,89,0,0,0,212,0,0,0,178,0,50,0,21,0,70,0,0,0,207,0,200,0,217,0,98,0,136,0,0,0,121,0,0,0,13,0,210,0,102,0,173,0,153,0,179,0,117,0,183,0,190,0,74,0,116,0,102,0,111,0,8,0,143,0,68,0,187,0,139,0,155,0,116,0,227,0,77,0,133,0,0,0,179,0,2,0,213,0,186,0,220,0,72,0,245,0,53,0,165,0,63,0,155,0,253,0,0,0,0,0,216,0,189,0,72,0,0,0,163,0,217,0,155,0,250,0,38,0,252,0,100,0,212,0,243,0,172,0,196,0,0,0,64,0,145,0,0,0,0,0,143,0,0,0,20,0,58,0,193,0,105,0,168,0,216,0,74,0);
signal scenario_full  : scenario_type := (58,31,16,31,201,31,188,31,178,31,60,31,60,30,60,29,240,31,71,31,139,31,94,31,143,31,254,31,254,30,240,31,252,31,252,30,192,31,192,30,138,31,138,30,98,31,83,31,83,30,35,31,35,30,249,31,169,31,169,30,240,31,196,31,3,31,243,31,63,31,130,31,4,31,4,30,66,31,231,31,32,31,213,31,213,30,158,31,158,30,158,29,201,31,201,30,19,31,236,31,126,31,165,31,101,31,176,31,138,31,88,31,82,31,129,31,66,31,14,31,160,31,160,30,158,31,31,31,78,31,172,31,172,30,172,29,242,31,10,31,239,31,107,31,16,31,46,31,46,30,246,31,246,30,69,31,69,31,196,31,196,30,196,29,145,31,142,31,194,31,190,31,232,31,3,31,161,31,128,31,169,31,120,31,20,31,72,31,241,31,241,30,83,31,12,31,12,30,229,31,63,31,8,31,165,31,165,30,166,31,198,31,121,31,205,31,228,31,228,30,251,31,251,30,61,31,152,31,120,31,120,30,85,31,85,30,52,31,52,30,90,31,182,31,118,31,66,31,127,31,52,31,201,31,201,30,163,31,164,31,164,30,75,31,43,31,95,31,173,31,125,31,125,30,13,31,98,31,74,31,157,31,254,31,236,31,149,31,42,31,42,30,42,29,153,31,250,31,35,31,35,30,178,31,57,31,80,31,168,31,204,31,204,30,14,31,180,31,190,31,190,30,83,31,134,31,67,31,55,31,55,30,242,31,193,31,131,31,104,31,47,31,226,31,173,31,56,31,106,31,40,31,135,31,82,31,186,31,6,31,50,31,202,31,251,31,11,31,11,30,10,31,10,30,20,31,253,31,212,31,45,31,45,30,124,31,218,31,218,30,51,31,135,31,135,30,191,31,191,30,107,31,246,31,246,30,111,31,177,31,241,31,178,31,178,30,129,31,129,30,179,31,179,30,179,29,204,31,138,31,111,31,225,31,208,31,208,30,35,31,116,31,61,31,212,31,23,31,219,31,75,31,75,30,17,31,196,31,21,31,21,30,50,31,76,31,171,31,3,31,79,31,154,31,154,30,154,29,246,31,250,31,151,31,103,31,84,31,33,31,72,31,230,31,230,30,230,29,124,31,200,31,200,30,168,31,103,31,103,30,103,29,245,31,129,31,197,31,3,31,123,31,123,30,252,31,252,30,185,31,156,31,82,31,147,31,147,30,123,31,192,31,91,31,91,30,46,31,46,30,180,31,180,30,216,31,216,30,165,31,157,31,187,31,189,31,189,30,251,31,174,31,121,31,154,31,151,31,151,30,151,29,36,31,36,30,36,29,90,31,210,31,37,31,251,31,3,31,3,30,152,31,141,31,162,31,50,31,251,31,79,31,79,30,98,31,98,30,140,31,85,31,100,31,226,31,14,31,186,31,166,31,23,31,187,31,186,31,186,30,180,31,24,31,196,31,196,30,196,29,34,31,30,31,40,31,80,31,253,31,60,31,30,31,127,31,129,31,129,30,129,29,129,28,38,31,38,30,38,29,117,31,119,31,25,31,174,31,22,31,186,31,143,31,232,31,232,30,122,31,7,31,113,31,9,31,191,31,177,31,94,31,153,31,10,31,189,31,105,31,54,31,114,31,52,31,107,31,79,31,79,30,169,31,227,31,101,31,5,31,16,31,16,30,120,31,171,31,77,31,6,31,6,30,48,31,157,31,220,31,215,31,215,30,138,31,138,30,159,31,32,31,221,31,221,30,218,31,197,31,3,31,248,31,248,30,240,31,145,31,191,31,191,30,11,31,255,31,58,31,58,30,181,31,110,31,104,31,109,31,99,31,105,31,181,31,102,31,244,31,79,31,156,31,13,31,13,30,13,29,235,31,108,31,143,31,189,31,168,31,14,31,176,31,58,31,39,31,215,31,108,31,79,31,79,30,85,31,85,30,157,31,89,31,76,31,76,30,233,31,167,31,167,30,233,31,93,31,143,31,118,31,118,30,251,31,113,31,45,31,124,31,183,31,176,31,153,31,229,31,221,31,160,31,70,31,18,31,139,31,77,31,94,31,94,30,80,31,133,31,246,31,141,31,168,31,168,30,168,29,231,31,187,31,82,31,216,31,216,30,163,31,237,31,12,31,95,31,95,30,165,31,81,31,81,30,101,31,62,31,28,31,135,31,120,31,209,31,209,30,99,31,107,31,202,31,27,31,27,30,142,31,142,30,101,31,101,30,227,31,227,30,83,31,83,30,83,29,112,31,54,31,52,31,52,30,19,31,137,31,137,30,113,31,240,31,229,31,94,31,195,31,220,31,247,31,86,31,226,31,1,31,1,30,44,31,38,31,194,31,208,31,96,31,42,31,100,31,100,30,252,31,97,31,97,30,88,31,88,30,88,29,71,31,117,31,74,31,91,31,224,31,224,30,199,31,153,31,69,31,218,31,118,31,89,31,89,30,192,31,134,31,181,31,147,31,231,31,254,31,89,31,89,30,212,31,212,30,178,31,50,31,21,31,70,31,70,30,207,31,200,31,217,31,98,31,136,31,136,30,121,31,121,30,13,31,210,31,102,31,173,31,153,31,179,31,117,31,183,31,190,31,74,31,116,31,102,31,111,31,8,31,143,31,68,31,187,31,139,31,155,31,116,31,227,31,77,31,133,31,133,30,179,31,2,31,213,31,186,31,220,31,72,31,245,31,53,31,165,31,63,31,155,31,253,31,253,30,253,29,216,31,189,31,72,31,72,30,163,31,217,31,155,31,250,31,38,31,252,31,100,31,212,31,243,31,172,31,196,31,196,30,64,31,145,31,145,30,145,29,143,31,143,30,20,31,58,31,193,31,105,31,168,31,216,31,74,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
