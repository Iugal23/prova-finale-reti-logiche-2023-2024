-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 415;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (65,0,0,0,70,0,165,0,17,0,216,0,136,0,100,0,6,0,251,0,0,0,0,0,40,0,0,0,137,0,231,0,239,0,0,0,251,0,128,0,0,0,238,0,194,0,164,0,0,0,223,0,221,0,48,0,0,0,93,0,0,0,210,0,15,0,160,0,144,0,54,0,5,0,0,0,50,0,78,0,177,0,138,0,239,0,203,0,45,0,113,0,0,0,71,0,184,0,193,0,0,0,216,0,228,0,107,0,227,0,67,0,0,0,86,0,0,0,28,0,157,0,194,0,204,0,198,0,156,0,0,0,236,0,169,0,87,0,146,0,143,0,198,0,243,0,0,0,0,0,223,0,82,0,0,0,230,0,86,0,89,0,77,0,70,0,244,0,214,0,178,0,0,0,13,0,73,0,227,0,189,0,121,0,221,0,34,0,242,0,239,0,53,0,118,0,245,0,182,0,78,0,5,0,0,0,126,0,136,0,213,0,32,0,0,0,0,0,246,0,167,0,46,0,0,0,0,0,0,0,171,0,151,0,254,0,0,0,0,0,250,0,0,0,45,0,28,0,123,0,0,0,219,0,174,0,57,0,0,0,219,0,0,0,0,0,5,0,58,0,194,0,99,0,139,0,123,0,68,0,0,0,186,0,122,0,85,0,19,0,100,0,28,0,0,0,229,0,217,0,93,0,0,0,0,0,0,0,4,0,2,0,0,0,15,0,0,0,22,0,90,0,215,0,226,0,111,0,113,0,0,0,0,0,235,0,79,0,0,0,36,0,94,0,164,0,188,0,201,0,0,0,245,0,167,0,172,0,0,0,0,0,0,0,191,0,172,0,147,0,124,0,235,0,54,0,0,0,82,0,176,0,202,0,0,0,48,0,189,0,18,0,195,0,4,0,24,0,30,0,183,0,222,0,90,0,197,0,233,0,201,0,117,0,34,0,112,0,0,0,158,0,186,0,0,0,44,0,183,0,248,0,10,0,63,0,227,0,39,0,120,0,181,0,116,0,37,0,0,0,175,0,175,0,212,0,71,0,232,0,166,0,108,0,139,0,74,0,0,0,83,0,0,0,0,0,0,0,127,0,100,0,59,0,137,0,70,0,175,0,0,0,25,0,88,0,187,0,163,0,64,0,115,0,243,0,16,0,126,0,74,0,219,0,194,0,120,0,30,0,122,0,242,0,50,0,38,0,0,0,0,0,0,0,13,0,82,0,0,0,250,0,195,0,34,0,56,0,213,0,189,0,0,0,49,0,179,0,35,0,121,0,241,0,95,0,219,0,0,0,100,0,238,0,239,0,0,0,0,0,85,0,118,0,176,0,238,0,61,0,137,0,0,0,12,0,114,0,181,0,131,0,21,0,30,0,167,0,0,0,28,0,71,0,170,0,50,0,183,0,135,0,92,0,199,0,184,0,23,0,237,0,0,0,22,0,0,0,0,0,36,0,116,0,0,0,140,0,119,0,87,0,239,0,132,0,193,0,250,0,0,0,117,0,201,0,235,0,82,0,0,0,31,0,0,0,0,0,112,0,1,0,104,0,166,0,0,0,0,0,0,0,113,0,0,0,0,0,189,0,96,0,149,0,95,0,62,0,211,0,169,0,10,0,135,0,0,0,246,0,159,0,94,0,240,0,51,0,138,0,19,0,171,0,66,0,131,0,0,0,233,0,67,0,138,0,117,0,128,0,0,0,0,0,127,0,1,0,245,0,127,0,71,0,0,0,0,0,39,0,0,0,8,0,0,0,97,0,61,0,25,0,0,0,66,0,168,0,148,0,16,0,183,0,0,0,190,0,4,0,98,0,0,0,109,0,54,0,34,0,135,0,148,0,0,0,159,0,235,0,164,0,101,0,170,0,86,0,0,0);
signal scenario_full  : scenario_type := (65,31,65,30,70,31,165,31,17,31,216,31,136,31,100,31,6,31,251,31,251,30,251,29,40,31,40,30,137,31,231,31,239,31,239,30,251,31,128,31,128,30,238,31,194,31,164,31,164,30,223,31,221,31,48,31,48,30,93,31,93,30,210,31,15,31,160,31,144,31,54,31,5,31,5,30,50,31,78,31,177,31,138,31,239,31,203,31,45,31,113,31,113,30,71,31,184,31,193,31,193,30,216,31,228,31,107,31,227,31,67,31,67,30,86,31,86,30,28,31,157,31,194,31,204,31,198,31,156,31,156,30,236,31,169,31,87,31,146,31,143,31,198,31,243,31,243,30,243,29,223,31,82,31,82,30,230,31,86,31,89,31,77,31,70,31,244,31,214,31,178,31,178,30,13,31,73,31,227,31,189,31,121,31,221,31,34,31,242,31,239,31,53,31,118,31,245,31,182,31,78,31,5,31,5,30,126,31,136,31,213,31,32,31,32,30,32,29,246,31,167,31,46,31,46,30,46,29,46,28,171,31,151,31,254,31,254,30,254,29,250,31,250,30,45,31,28,31,123,31,123,30,219,31,174,31,57,31,57,30,219,31,219,30,219,29,5,31,58,31,194,31,99,31,139,31,123,31,68,31,68,30,186,31,122,31,85,31,19,31,100,31,28,31,28,30,229,31,217,31,93,31,93,30,93,29,93,28,4,31,2,31,2,30,15,31,15,30,22,31,90,31,215,31,226,31,111,31,113,31,113,30,113,29,235,31,79,31,79,30,36,31,94,31,164,31,188,31,201,31,201,30,245,31,167,31,172,31,172,30,172,29,172,28,191,31,172,31,147,31,124,31,235,31,54,31,54,30,82,31,176,31,202,31,202,30,48,31,189,31,18,31,195,31,4,31,24,31,30,31,183,31,222,31,90,31,197,31,233,31,201,31,117,31,34,31,112,31,112,30,158,31,186,31,186,30,44,31,183,31,248,31,10,31,63,31,227,31,39,31,120,31,181,31,116,31,37,31,37,30,175,31,175,31,212,31,71,31,232,31,166,31,108,31,139,31,74,31,74,30,83,31,83,30,83,29,83,28,127,31,100,31,59,31,137,31,70,31,175,31,175,30,25,31,88,31,187,31,163,31,64,31,115,31,243,31,16,31,126,31,74,31,219,31,194,31,120,31,30,31,122,31,242,31,50,31,38,31,38,30,38,29,38,28,13,31,82,31,82,30,250,31,195,31,34,31,56,31,213,31,189,31,189,30,49,31,179,31,35,31,121,31,241,31,95,31,219,31,219,30,100,31,238,31,239,31,239,30,239,29,85,31,118,31,176,31,238,31,61,31,137,31,137,30,12,31,114,31,181,31,131,31,21,31,30,31,167,31,167,30,28,31,71,31,170,31,50,31,183,31,135,31,92,31,199,31,184,31,23,31,237,31,237,30,22,31,22,30,22,29,36,31,116,31,116,30,140,31,119,31,87,31,239,31,132,31,193,31,250,31,250,30,117,31,201,31,235,31,82,31,82,30,31,31,31,30,31,29,112,31,1,31,104,31,166,31,166,30,166,29,166,28,113,31,113,30,113,29,189,31,96,31,149,31,95,31,62,31,211,31,169,31,10,31,135,31,135,30,246,31,159,31,94,31,240,31,51,31,138,31,19,31,171,31,66,31,131,31,131,30,233,31,67,31,138,31,117,31,128,31,128,30,128,29,127,31,1,31,245,31,127,31,71,31,71,30,71,29,39,31,39,30,8,31,8,30,97,31,61,31,25,31,25,30,66,31,168,31,148,31,16,31,183,31,183,30,190,31,4,31,98,31,98,30,109,31,54,31,34,31,135,31,148,31,148,30,159,31,235,31,164,31,101,31,170,31,86,31,86,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
