-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_288 is
end project_tb_288;

architecture project_tb_arch_288 of project_tb_288 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 936;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,13,0,185,0,12,0,78,0,237,0,175,0,126,0,87,0,0,0,186,0,80,0,0,0,225,0,139,0,14,0,17,0,227,0,124,0,35,0,7,0,0,0,197,0,0,0,11,0,170,0,0,0,213,0,0,0,67,0,59,0,92,0,200,0,138,0,4,0,0,0,111,0,121,0,28,0,0,0,0,0,0,0,134,0,100,0,249,0,46,0,48,0,152,0,118,0,60,0,43,0,81,0,0,0,111,0,189,0,2,0,43,0,147,0,93,0,250,0,0,0,99,0,10,0,161,0,220,0,134,0,76,0,27,0,0,0,106,0,7,0,90,0,242,0,230,0,128,0,62,0,11,0,235,0,194,0,238,0,14,0,176,0,0,0,69,0,161,0,0,0,72,0,119,0,0,0,239,0,219,0,22,0,0,0,115,0,0,0,203,0,247,0,171,0,151,0,0,0,0,0,46,0,197,0,117,0,168,0,0,0,0,0,60,0,77,0,29,0,85,0,87,0,210,0,27,0,0,0,230,0,127,0,100,0,49,0,0,0,241,0,54,0,0,0,166,0,0,0,83,0,205,0,69,0,164,0,115,0,166,0,14,0,210,0,0,0,119,0,157,0,237,0,85,0,166,0,75,0,0,0,0,0,163,0,132,0,0,0,96,0,56,0,54,0,94,0,11,0,44,0,0,0,132,0,52,0,28,0,0,0,235,0,0,0,249,0,147,0,112,0,190,0,0,0,254,0,103,0,12,0,114,0,7,0,7,0,78,0,114,0,0,0,75,0,0,0,99,0,0,0,142,0,23,0,134,0,0,0,15,0,0,0,220,0,234,0,194,0,205,0,101,0,108,0,134,0,127,0,51,0,170,0,42,0,78,0,60,0,0,0,165,0,0,0,237,0,82,0,237,0,34,0,171,0,102,0,143,0,0,0,175,0,128,0,113,0,0,0,207,0,116,0,243,0,41,0,94,0,0,0,214,0,197,0,104,0,37,0,163,0,162,0,99,0,79,0,197,0,218,0,22,0,229,0,220,0,238,0,201,0,0,0,0,0,0,0,180,0,219,0,0,0,0,0,0,0,200,0,129,0,24,0,240,0,210,0,112,0,6,0,112,0,127,0,71,0,140,0,198,0,14,0,87,0,238,0,91,0,113,0,148,0,22,0,126,0,26,0,190,0,218,0,14,0,24,0,88,0,137,0,67,0,58,0,212,0,214,0,188,0,219,0,0,0,197,0,143,0,5,0,23,0,116,0,128,0,253,0,123,0,224,0,159,0,93,0,113,0,40,0,0,0,147,0,20,0,207,0,187,0,201,0,217,0,1,0,107,0,199,0,107,0,30,0,0,0,106,0,0,0,249,0,1,0,115,0,238,0,48,0,5,0,136,0,115,0,13,0,93,0,0,0,160,0,172,0,51,0,63,0,192,0,51,0,92,0,209,0,26,0,159,0,0,0,116,0,155,0,0,0,215,0,213,0,198,0,253,0,125,0,200,0,211,0,20,0,30,0,233,0,86,0,143,0,116,0,0,0,242,0,3,0,0,0,154,0,228,0,58,0,0,0,250,0,163,0,45,0,0,0,68,0,246,0,0,0,49,0,233,0,59,0,0,0,215,0,129,0,247,0,0,0,80,0,55,0,97,0,153,0,140,0,159,0,0,0,47,0,225,0,201,0,105,0,0,0,13,0,150,0,52,0,215,0,16,0,239,0,135,0,199,0,156,0,140,0,0,0,196,0,220,0,153,0,104,0,46,0,115,0,0,0,0,0,5,0,86,0,163,0,218,0,16,0,0,0,0,0,227,0,108,0,19,0,41,0,0,0,129,0,19,0,0,0,27,0,191,0,70,0,215,0,81,0,96,0,86,0,21,0,10,0,90,0,56,0,88,0,59,0,100,0,0,0,247,0,103,0,0,0,205,0,0,0,80,0,35,0,201,0,0,0,32,0,38,0,103,0,0,0,171,0,0,0,164,0,18,0,250,0,236,0,100,0,151,0,46,0,233,0,206,0,0,0,81,0,0,0,175,0,0,0,251,0,0,0,177,0,227,0,0,0,25,0,0,0,25,0,174,0,193,0,209,0,133,0,109,0,185,0,0,0,246,0,229,0,159,0,200,0,0,0,49,0,0,0,251,0,0,0,3,0,44,0,96,0,15,0,139,0,120,0,173,0,83,0,0,0,49,0,131,0,207,0,0,0,61,0,0,0,252,0,147,0,183,0,13,0,215,0,0,0,0,0,3,0,115,0,56,0,243,0,61,0,61,0,0,0,244,0,190,0,206,0,150,0,0,0,96,0,85,0,137,0,0,0,189,0,0,0,84,0,214,0,124,0,106,0,211,0,76,0,23,0,117,0,190,0,0,0,46,0,156,0,41,0,78,0,0,0,235,0,0,0,67,0,208,0,109,0,38,0,160,0,242,0,237,0,0,0,153,0,222,0,0,0,19,0,57,0,115,0,212,0,31,0,196,0,55,0,85,0,237,0,240,0,62,0,191,0,29,0,0,0,49,0,247,0,101,0,66,0,27,0,65,0,130,0,183,0,186,0,0,0,232,0,199,0,241,0,215,0,42,0,141,0,65,0,63,0,183,0,122,0,28,0,43,0,196,0,132,0,28,0,155,0,53,0,15,0,0,0,133,0,0,0,0,0,25,0,0,0,59,0,250,0,237,0,0,0,190,0,0,0,96,0,216,0,129,0,0,0,0,0,79,0,52,0,136,0,244,0,103,0,150,0,221,0,0,0,48,0,238,0,144,0,58,0,71,0,128,0,126,0,218,0,244,0,23,0,230,0,18,0,2,0,148,0,0,0,0,0,176,0,19,0,198,0,0,0,133,0,23,0,174,0,248,0,142,0,107,0,36,0,32,0,5,0,0,0,111,0,0,0,216,0,244,0,0,0,0,0,139,0,203,0,37,0,195,0,120,0,68,0,13,0,254,0,28,0,141,0,155,0,0,0,10,0,226,0,0,0,70,0,0,0,0,0,0,0,21,0,75,0,0,0,0,0,114,0,133,0,74,0,190,0,224,0,118,0,6,0,89,0,225,0,67,0,80,0,0,0,121,0,0,0,178,0,60,0,186,0,254,0,38,0,0,0,204,0,160,0,171,0,66,0,31,0,4,0,179,0,180,0,126,0,34,0,165,0,0,0,180,0,0,0,191,0,249,0,157,0,191,0,0,0,64,0,159,0,145,0,0,0,129,0,209,0,252,0,32,0,0,0,79,0,103,0,102,0,174,0,151,0,0,0,155,0,0,0,111,0,150,0,77,0,220,0,155,0,0,0,95,0,83,0,240,0,60,0,0,0,128,0,117,0,123,0,0,0,58,0,0,0,211,0,214,0,18,0,0,0,210,0,147,0,165,0,105,0,0,0,101,0,127,0,26,0,17,0,237,0,170,0,254,0,24,0,44,0,198,0,13,0,106,0,80,0,188,0,127,0,151,0,218,0,234,0,218,0,246,0,253,0,65,0,189,0,0,0,19,0,74,0,186,0,0,0,166,0,0,0,0,0,141,0,216,0,0,0,0,0,80,0,84,0,244,0,13,0,82,0,0,0,40,0,0,0,248,0,217,0,51,0,151,0,0,0,0,0,171,0,0,0,46,0,171,0,94,0,226,0,177,0,123,0,87,0,166,0,9,0,17,0,37,0,0,0,151,0,147,0,60,0,61,0,0,0,12,0,0,0,0,0,190,0,226,0,0,0,93,0,162,0,58,0,105,0,57,0,120,0,154,0,179,0,50,0,45,0,0,0,240,0,177,0,174,0,26,0,189,0,216,0,249,0,247,0,76,0,32,0,93,0,125,0,50,0,209,0,143,0,109,0,18,0,199,0,1,0,89,0,194,0,0,0,218,0,189,0,96,0,0,0,139,0,16,0,63,0,33,0,214,0,28,0,0,0,158,0,0,0,50,0,240,0,205,0,103,0,172,0,230,0,254,0,110,0,213,0,29,0,180,0,176,0,177,0,228,0,109,0,200,0,133,0,84,0,254,0,0,0,0,0,33,0,14,0,16,0,0,0,151,0,132,0,55,0,89,0,7,0,223,0,0,0,130,0,0,0,156,0,225,0,24,0,24,0,211,0,107,0,0,0,125,0,216,0,0,0,51,0,144,0,149,0,240,0,216,0,39,0,145,0,224,0,81,0,191,0,230,0,97,0,0,0,244,0,92,0,94,0,221,0,92,0,190,0,46,0);
signal scenario_full  : scenario_type := (0,0,13,31,185,31,12,31,78,31,237,31,175,31,126,31,87,31,87,30,186,31,80,31,80,30,225,31,139,31,14,31,17,31,227,31,124,31,35,31,7,31,7,30,197,31,197,30,11,31,170,31,170,30,213,31,213,30,67,31,59,31,92,31,200,31,138,31,4,31,4,30,111,31,121,31,28,31,28,30,28,29,28,28,134,31,100,31,249,31,46,31,48,31,152,31,118,31,60,31,43,31,81,31,81,30,111,31,189,31,2,31,43,31,147,31,93,31,250,31,250,30,99,31,10,31,161,31,220,31,134,31,76,31,27,31,27,30,106,31,7,31,90,31,242,31,230,31,128,31,62,31,11,31,235,31,194,31,238,31,14,31,176,31,176,30,69,31,161,31,161,30,72,31,119,31,119,30,239,31,219,31,22,31,22,30,115,31,115,30,203,31,247,31,171,31,151,31,151,30,151,29,46,31,197,31,117,31,168,31,168,30,168,29,60,31,77,31,29,31,85,31,87,31,210,31,27,31,27,30,230,31,127,31,100,31,49,31,49,30,241,31,54,31,54,30,166,31,166,30,83,31,205,31,69,31,164,31,115,31,166,31,14,31,210,31,210,30,119,31,157,31,237,31,85,31,166,31,75,31,75,30,75,29,163,31,132,31,132,30,96,31,56,31,54,31,94,31,11,31,44,31,44,30,132,31,52,31,28,31,28,30,235,31,235,30,249,31,147,31,112,31,190,31,190,30,254,31,103,31,12,31,114,31,7,31,7,31,78,31,114,31,114,30,75,31,75,30,99,31,99,30,142,31,23,31,134,31,134,30,15,31,15,30,220,31,234,31,194,31,205,31,101,31,108,31,134,31,127,31,51,31,170,31,42,31,78,31,60,31,60,30,165,31,165,30,237,31,82,31,237,31,34,31,171,31,102,31,143,31,143,30,175,31,128,31,113,31,113,30,207,31,116,31,243,31,41,31,94,31,94,30,214,31,197,31,104,31,37,31,163,31,162,31,99,31,79,31,197,31,218,31,22,31,229,31,220,31,238,31,201,31,201,30,201,29,201,28,180,31,219,31,219,30,219,29,219,28,200,31,129,31,24,31,240,31,210,31,112,31,6,31,112,31,127,31,71,31,140,31,198,31,14,31,87,31,238,31,91,31,113,31,148,31,22,31,126,31,26,31,190,31,218,31,14,31,24,31,88,31,137,31,67,31,58,31,212,31,214,31,188,31,219,31,219,30,197,31,143,31,5,31,23,31,116,31,128,31,253,31,123,31,224,31,159,31,93,31,113,31,40,31,40,30,147,31,20,31,207,31,187,31,201,31,217,31,1,31,107,31,199,31,107,31,30,31,30,30,106,31,106,30,249,31,1,31,115,31,238,31,48,31,5,31,136,31,115,31,13,31,93,31,93,30,160,31,172,31,51,31,63,31,192,31,51,31,92,31,209,31,26,31,159,31,159,30,116,31,155,31,155,30,215,31,213,31,198,31,253,31,125,31,200,31,211,31,20,31,30,31,233,31,86,31,143,31,116,31,116,30,242,31,3,31,3,30,154,31,228,31,58,31,58,30,250,31,163,31,45,31,45,30,68,31,246,31,246,30,49,31,233,31,59,31,59,30,215,31,129,31,247,31,247,30,80,31,55,31,97,31,153,31,140,31,159,31,159,30,47,31,225,31,201,31,105,31,105,30,13,31,150,31,52,31,215,31,16,31,239,31,135,31,199,31,156,31,140,31,140,30,196,31,220,31,153,31,104,31,46,31,115,31,115,30,115,29,5,31,86,31,163,31,218,31,16,31,16,30,16,29,227,31,108,31,19,31,41,31,41,30,129,31,19,31,19,30,27,31,191,31,70,31,215,31,81,31,96,31,86,31,21,31,10,31,90,31,56,31,88,31,59,31,100,31,100,30,247,31,103,31,103,30,205,31,205,30,80,31,35,31,201,31,201,30,32,31,38,31,103,31,103,30,171,31,171,30,164,31,18,31,250,31,236,31,100,31,151,31,46,31,233,31,206,31,206,30,81,31,81,30,175,31,175,30,251,31,251,30,177,31,227,31,227,30,25,31,25,30,25,31,174,31,193,31,209,31,133,31,109,31,185,31,185,30,246,31,229,31,159,31,200,31,200,30,49,31,49,30,251,31,251,30,3,31,44,31,96,31,15,31,139,31,120,31,173,31,83,31,83,30,49,31,131,31,207,31,207,30,61,31,61,30,252,31,147,31,183,31,13,31,215,31,215,30,215,29,3,31,115,31,56,31,243,31,61,31,61,31,61,30,244,31,190,31,206,31,150,31,150,30,96,31,85,31,137,31,137,30,189,31,189,30,84,31,214,31,124,31,106,31,211,31,76,31,23,31,117,31,190,31,190,30,46,31,156,31,41,31,78,31,78,30,235,31,235,30,67,31,208,31,109,31,38,31,160,31,242,31,237,31,237,30,153,31,222,31,222,30,19,31,57,31,115,31,212,31,31,31,196,31,55,31,85,31,237,31,240,31,62,31,191,31,29,31,29,30,49,31,247,31,101,31,66,31,27,31,65,31,130,31,183,31,186,31,186,30,232,31,199,31,241,31,215,31,42,31,141,31,65,31,63,31,183,31,122,31,28,31,43,31,196,31,132,31,28,31,155,31,53,31,15,31,15,30,133,31,133,30,133,29,25,31,25,30,59,31,250,31,237,31,237,30,190,31,190,30,96,31,216,31,129,31,129,30,129,29,79,31,52,31,136,31,244,31,103,31,150,31,221,31,221,30,48,31,238,31,144,31,58,31,71,31,128,31,126,31,218,31,244,31,23,31,230,31,18,31,2,31,148,31,148,30,148,29,176,31,19,31,198,31,198,30,133,31,23,31,174,31,248,31,142,31,107,31,36,31,32,31,5,31,5,30,111,31,111,30,216,31,244,31,244,30,244,29,139,31,203,31,37,31,195,31,120,31,68,31,13,31,254,31,28,31,141,31,155,31,155,30,10,31,226,31,226,30,70,31,70,30,70,29,70,28,21,31,75,31,75,30,75,29,114,31,133,31,74,31,190,31,224,31,118,31,6,31,89,31,225,31,67,31,80,31,80,30,121,31,121,30,178,31,60,31,186,31,254,31,38,31,38,30,204,31,160,31,171,31,66,31,31,31,4,31,179,31,180,31,126,31,34,31,165,31,165,30,180,31,180,30,191,31,249,31,157,31,191,31,191,30,64,31,159,31,145,31,145,30,129,31,209,31,252,31,32,31,32,30,79,31,103,31,102,31,174,31,151,31,151,30,155,31,155,30,111,31,150,31,77,31,220,31,155,31,155,30,95,31,83,31,240,31,60,31,60,30,128,31,117,31,123,31,123,30,58,31,58,30,211,31,214,31,18,31,18,30,210,31,147,31,165,31,105,31,105,30,101,31,127,31,26,31,17,31,237,31,170,31,254,31,24,31,44,31,198,31,13,31,106,31,80,31,188,31,127,31,151,31,218,31,234,31,218,31,246,31,253,31,65,31,189,31,189,30,19,31,74,31,186,31,186,30,166,31,166,30,166,29,141,31,216,31,216,30,216,29,80,31,84,31,244,31,13,31,82,31,82,30,40,31,40,30,248,31,217,31,51,31,151,31,151,30,151,29,171,31,171,30,46,31,171,31,94,31,226,31,177,31,123,31,87,31,166,31,9,31,17,31,37,31,37,30,151,31,147,31,60,31,61,31,61,30,12,31,12,30,12,29,190,31,226,31,226,30,93,31,162,31,58,31,105,31,57,31,120,31,154,31,179,31,50,31,45,31,45,30,240,31,177,31,174,31,26,31,189,31,216,31,249,31,247,31,76,31,32,31,93,31,125,31,50,31,209,31,143,31,109,31,18,31,199,31,1,31,89,31,194,31,194,30,218,31,189,31,96,31,96,30,139,31,16,31,63,31,33,31,214,31,28,31,28,30,158,31,158,30,50,31,240,31,205,31,103,31,172,31,230,31,254,31,110,31,213,31,29,31,180,31,176,31,177,31,228,31,109,31,200,31,133,31,84,31,254,31,254,30,254,29,33,31,14,31,16,31,16,30,151,31,132,31,55,31,89,31,7,31,223,31,223,30,130,31,130,30,156,31,225,31,24,31,24,31,211,31,107,31,107,30,125,31,216,31,216,30,51,31,144,31,149,31,240,31,216,31,39,31,145,31,224,31,81,31,191,31,230,31,97,31,97,30,244,31,92,31,94,31,221,31,92,31,190,31,46,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
