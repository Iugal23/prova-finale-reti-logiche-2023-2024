-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 178;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (103,0,0,0,25,0,0,0,38,0,0,0,49,0,34,0,0,0,10,0,31,0,204,0,58,0,73,0,249,0,217,0,96,0,140,0,72,0,0,0,234,0,241,0,56,0,232,0,94,0,69,0,0,0,247,0,0,0,17,0,136,0,32,0,111,0,0,0,242,0,157,0,150,0,111,0,88,0,202,0,80,0,0,0,0,0,189,0,113,0,0,0,113,0,199,0,143,0,109,0,98,0,70,0,195,0,1,0,99,0,45,0,0,0,81,0,8,0,108,0,84,0,208,0,31,0,151,0,161,0,0,0,156,0,104,0,183,0,143,0,172,0,232,0,110,0,212,0,0,0,0,0,163,0,228,0,121,0,208,0,136,0,2,0,26,0,35,0,138,0,39,0,224,0,159,0,115,0,111,0,93,0,0,0,0,0,135,0,48,0,146,0,218,0,248,0,0,0,84,0,19,0,0,0,3,0,160,0,0,0,0,0,68,0,0,0,201,0,79,0,218,0,0,0,116,0,109,0,54,0,94,0,24,0,136,0,103,0,216,0,0,0,125,0,89,0,206,0,0,0,91,0,54,0,90,0,17,0,87,0,32,0,105,0,141,0,139,0,90,0,234,0,50,0,62,0,180,0,248,0,0,0,246,0,0,0,243,0,13,0,19,0,103,0,159,0,0,0,107,0,0,0,126,0,122,0,172,0,13,0,50,0,116,0,0,0,109,0,29,0,65,0,177,0,95,0,235,0,118,0,0,0,0,0,71,0,183,0,61,0,206,0,191,0,31,0,129,0,120,0,0,0,116,0,0,0);
signal scenario_full  : scenario_type := (103,31,103,30,25,31,25,30,38,31,38,30,49,31,34,31,34,30,10,31,31,31,204,31,58,31,73,31,249,31,217,31,96,31,140,31,72,31,72,30,234,31,241,31,56,31,232,31,94,31,69,31,69,30,247,31,247,30,17,31,136,31,32,31,111,31,111,30,242,31,157,31,150,31,111,31,88,31,202,31,80,31,80,30,80,29,189,31,113,31,113,30,113,31,199,31,143,31,109,31,98,31,70,31,195,31,1,31,99,31,45,31,45,30,81,31,8,31,108,31,84,31,208,31,31,31,151,31,161,31,161,30,156,31,104,31,183,31,143,31,172,31,232,31,110,31,212,31,212,30,212,29,163,31,228,31,121,31,208,31,136,31,2,31,26,31,35,31,138,31,39,31,224,31,159,31,115,31,111,31,93,31,93,30,93,29,135,31,48,31,146,31,218,31,248,31,248,30,84,31,19,31,19,30,3,31,160,31,160,30,160,29,68,31,68,30,201,31,79,31,218,31,218,30,116,31,109,31,54,31,94,31,24,31,136,31,103,31,216,31,216,30,125,31,89,31,206,31,206,30,91,31,54,31,90,31,17,31,87,31,32,31,105,31,141,31,139,31,90,31,234,31,50,31,62,31,180,31,248,31,248,30,246,31,246,30,243,31,13,31,19,31,103,31,159,31,159,30,107,31,107,30,126,31,122,31,172,31,13,31,50,31,116,31,116,30,109,31,29,31,65,31,177,31,95,31,235,31,118,31,118,30,118,29,71,31,183,31,61,31,206,31,191,31,31,31,129,31,120,31,120,30,116,31,116,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
