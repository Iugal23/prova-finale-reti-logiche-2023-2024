-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_518 is
end project_tb_518;

architecture project_tb_arch_518 of project_tb_518 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 760;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (90,0,167,0,238,0,101,0,0,0,145,0,10,0,233,0,0,0,96,0,0,0,158,0,205,0,176,0,121,0,0,0,140,0,90,0,250,0,132,0,0,0,0,0,202,0,49,0,204,0,128,0,51,0,0,0,67,0,0,0,2,0,167,0,0,0,160,0,193,0,175,0,1,0,239,0,177,0,250,0,21,0,86,0,175,0,0,0,5,0,185,0,191,0,0,0,1,0,161,0,0,0,81,0,174,0,224,0,229,0,235,0,91,0,220,0,168,0,187,0,46,0,167,0,207,0,128,0,99,0,184,0,138,0,56,0,43,0,0,0,189,0,37,0,46,0,19,0,204,0,4,0,49,0,89,0,122,0,0,0,92,0,3,0,79,0,168,0,230,0,205,0,0,0,165,0,33,0,75,0,0,0,77,0,70,0,0,0,125,0,20,0,70,0,212,0,255,0,0,0,96,0,199,0,27,0,110,0,90,0,28,0,106,0,150,0,112,0,96,0,0,0,140,0,0,0,42,0,198,0,93,0,0,0,87,0,0,0,0,0,243,0,0,0,43,0,106,0,113,0,5,0,122,0,34,0,93,0,0,0,192,0,220,0,0,0,27,0,0,0,65,0,130,0,18,0,8,0,93,0,170,0,70,0,51,0,156,0,0,0,29,0,74,0,192,0,146,0,198,0,92,0,231,0,222,0,5,0,112,0,2,0,0,0,138,0,140,0,0,0,158,0,180,0,231,0,98,0,48,0,0,0,62,0,208,0,0,0,78,0,242,0,103,0,196,0,114,0,35,0,15,0,127,0,145,0,220,0,0,0,92,0,0,0,76,0,153,0,8,0,200,0,208,0,0,0,88,0,195,0,235,0,0,0,0,0,0,0,13,0,0,0,85,0,0,0,208,0,188,0,95,0,1,0,119,0,79,0,169,0,160,0,163,0,96,0,161,0,12,0,78,0,99,0,14,0,0,0,131,0,66,0,0,0,0,0,179,0,49,0,2,0,97,0,135,0,38,0,64,0,134,0,108,0,183,0,21,0,0,0,198,0,69,0,3,0,34,0,73,0,0,0,20,0,0,0,88,0,0,0,46,0,254,0,194,0,0,0,215,0,0,0,131,0,238,0,0,0,0,0,32,0,168,0,244,0,193,0,0,0,114,0,35,0,249,0,9,0,86,0,38,0,191,0,0,0,91,0,189,0,0,0,0,0,5,0,148,0,99,0,129,0,0,0,0,0,0,0,0,0,138,0,0,0,96,0,151,0,7,0,134,0,255,0,0,0,234,0,66,0,36,0,90,0,89,0,0,0,102,0,160,0,130,0,85,0,148,0,252,0,67,0,0,0,99,0,62,0,248,0,79,0,0,0,0,0,24,0,137,0,26,0,96,0,0,0,127,0,0,0,214,0,0,0,9,0,146,0,224,0,31,0,226,0,134,0,91,0,126,0,213,0,9,0,177,0,169,0,61,0,37,0,0,0,117,0,81,0,85,0,124,0,57,0,173,0,171,0,15,0,95,0,36,0,88,0,252,0,237,0,206,0,7,0,174,0,31,0,12,0,219,0,0,0,143,0,8,0,155,0,248,0,157,0,255,0,147,0,157,0,148,0,138,0,0,0,133,0,134,0,0,0,0,0,22,0,236,0,186,0,165,0,67,0,162,0,0,0,0,0,231,0,94,0,0,0,208,0,95,0,222,0,121,0,155,0,0,0,0,0,155,0,151,0,140,0,115,0,228,0,242,0,0,0,213,0,79,0,91,0,85,0,0,0,0,0,108,0,213,0,8,0,58,0,237,0,203,0,208,0,203,0,167,0,0,0,217,0,158,0,188,0,171,0,21,0,214,0,149,0,33,0,148,0,0,0,91,0,1,0,221,0,248,0,247,0,77,0,55,0,13,0,101,0,97,0,0,0,223,0,30,0,0,0,0,0,0,0,243,0,225,0,0,0,0,0,5,0,208,0,0,0,15,0,178,0,0,0,126,0,66,0,25,0,30,0,186,0,242,0,0,0,0,0,215,0,114,0,72,0,31,0,48,0,0,0,227,0,145,0,121,0,235,0,74,0,80,0,0,0,152,0,78,0,251,0,165,0,0,0,112,0,160,0,29,0,0,0,166,0,189,0,192,0,221,0,113,0,203,0,1,0,216,0,196,0,164,0,42,0,15,0,64,0,0,0,191,0,163,0,246,0,0,0,0,0,185,0,164,0,24,0,196,0,112,0,44,0,85,0,67,0,161,0,0,0,139,0,161,0,85,0,235,0,183,0,163,0,33,0,58,0,0,0,196,0,41,0,95,0,96,0,131,0,6,0,0,0,144,0,22,0,125,0,137,0,0,0,52,0,11,0,0,0,241,0,52,0,0,0,0,0,203,0,154,0,177,0,119,0,116,0,158,0,117,0,122,0,178,0,0,0,0,0,132,0,255,0,145,0,85,0,21,0,243,0,14,0,194,0,36,0,238,0,0,0,0,0,21,0,64,0,51,0,115,0,223,0,125,0,44,0,197,0,115,0,6,0,38,0,48,0,102,0,81,0,142,0,198,0,0,0,230,0,114,0,0,0,225,0,212,0,199,0,0,0,241,0,0,0,12,0,43,0,92,0,165,0,140,0,68,0,138,0,167,0,46,0,0,0,215,0,127,0,2,0,41,0,162,0,75,0,0,0,13,0,120,0,249,0,122,0,220,0,117,0,0,0,155,0,49,0,100,0,72,0,105,0,4,0,76,0,90,0,1,0,178,0,75,0,0,0,0,0,101,0,207,0,0,0,35,0,0,0,146,0,0,0,78,0,250,0,141,0,29,0,220,0,198,0,0,0,171,0,110,0,237,0,167,0,178,0,0,0,0,0,14,0,75,0,84,0,12,0,40,0,94,0,159,0,149,0,36,0,91,0,0,0,72,0,79,0,211,0,124,0,0,0,74,0,24,0,133,0,240,0,69,0,49,0,243,0,197,0,133,0,0,0,208,0,24,0,245,0,0,0,136,0,0,0,0,0,132,0,217,0,190,0,243,0,105,0,140,0,22,0,165,0,175,0,93,0,234,0,177,0,96,0,133,0,30,0,0,0,145,0,122,0,200,0,0,0,241,0,202,0,249,0,200,0,11,0,156,0,0,0,91,0,139,0,0,0,145,0,240,0,0,0,215,0,226,0,181,0,102,0,0,0,41,0,226,0,65,0,0,0,0,0,250,0,235,0,196,0,220,0,9,0,75,0,120,0,0,0,163,0,91,0,48,0,111,0,0,0,70,0,135,0,134,0,59,0,229,0,209,0,0,0,154,0,125,0,102,0,177,0,8,0,153,0,134,0,0,0,96,0,43,0,238,0,233,0,50,0,0,0,172,0,81,0,10,0,84,0,99,0,127,0,0,0,210,0,0,0,229,0,244,0,186,0,1,0,231,0,202,0,122,0,0,0);
signal scenario_full  : scenario_type := (90,31,167,31,238,31,101,31,101,30,145,31,10,31,233,31,233,30,96,31,96,30,158,31,205,31,176,31,121,31,121,30,140,31,90,31,250,31,132,31,132,30,132,29,202,31,49,31,204,31,128,31,51,31,51,30,67,31,67,30,2,31,167,31,167,30,160,31,193,31,175,31,1,31,239,31,177,31,250,31,21,31,86,31,175,31,175,30,5,31,185,31,191,31,191,30,1,31,161,31,161,30,81,31,174,31,224,31,229,31,235,31,91,31,220,31,168,31,187,31,46,31,167,31,207,31,128,31,99,31,184,31,138,31,56,31,43,31,43,30,189,31,37,31,46,31,19,31,204,31,4,31,49,31,89,31,122,31,122,30,92,31,3,31,79,31,168,31,230,31,205,31,205,30,165,31,33,31,75,31,75,30,77,31,70,31,70,30,125,31,20,31,70,31,212,31,255,31,255,30,96,31,199,31,27,31,110,31,90,31,28,31,106,31,150,31,112,31,96,31,96,30,140,31,140,30,42,31,198,31,93,31,93,30,87,31,87,30,87,29,243,31,243,30,43,31,106,31,113,31,5,31,122,31,34,31,93,31,93,30,192,31,220,31,220,30,27,31,27,30,65,31,130,31,18,31,8,31,93,31,170,31,70,31,51,31,156,31,156,30,29,31,74,31,192,31,146,31,198,31,92,31,231,31,222,31,5,31,112,31,2,31,2,30,138,31,140,31,140,30,158,31,180,31,231,31,98,31,48,31,48,30,62,31,208,31,208,30,78,31,242,31,103,31,196,31,114,31,35,31,15,31,127,31,145,31,220,31,220,30,92,31,92,30,76,31,153,31,8,31,200,31,208,31,208,30,88,31,195,31,235,31,235,30,235,29,235,28,13,31,13,30,85,31,85,30,208,31,188,31,95,31,1,31,119,31,79,31,169,31,160,31,163,31,96,31,161,31,12,31,78,31,99,31,14,31,14,30,131,31,66,31,66,30,66,29,179,31,49,31,2,31,97,31,135,31,38,31,64,31,134,31,108,31,183,31,21,31,21,30,198,31,69,31,3,31,34,31,73,31,73,30,20,31,20,30,88,31,88,30,46,31,254,31,194,31,194,30,215,31,215,30,131,31,238,31,238,30,238,29,32,31,168,31,244,31,193,31,193,30,114,31,35,31,249,31,9,31,86,31,38,31,191,31,191,30,91,31,189,31,189,30,189,29,5,31,148,31,99,31,129,31,129,30,129,29,129,28,129,27,138,31,138,30,96,31,151,31,7,31,134,31,255,31,255,30,234,31,66,31,36,31,90,31,89,31,89,30,102,31,160,31,130,31,85,31,148,31,252,31,67,31,67,30,99,31,62,31,248,31,79,31,79,30,79,29,24,31,137,31,26,31,96,31,96,30,127,31,127,30,214,31,214,30,9,31,146,31,224,31,31,31,226,31,134,31,91,31,126,31,213,31,9,31,177,31,169,31,61,31,37,31,37,30,117,31,81,31,85,31,124,31,57,31,173,31,171,31,15,31,95,31,36,31,88,31,252,31,237,31,206,31,7,31,174,31,31,31,12,31,219,31,219,30,143,31,8,31,155,31,248,31,157,31,255,31,147,31,157,31,148,31,138,31,138,30,133,31,134,31,134,30,134,29,22,31,236,31,186,31,165,31,67,31,162,31,162,30,162,29,231,31,94,31,94,30,208,31,95,31,222,31,121,31,155,31,155,30,155,29,155,31,151,31,140,31,115,31,228,31,242,31,242,30,213,31,79,31,91,31,85,31,85,30,85,29,108,31,213,31,8,31,58,31,237,31,203,31,208,31,203,31,167,31,167,30,217,31,158,31,188,31,171,31,21,31,214,31,149,31,33,31,148,31,148,30,91,31,1,31,221,31,248,31,247,31,77,31,55,31,13,31,101,31,97,31,97,30,223,31,30,31,30,30,30,29,30,28,243,31,225,31,225,30,225,29,5,31,208,31,208,30,15,31,178,31,178,30,126,31,66,31,25,31,30,31,186,31,242,31,242,30,242,29,215,31,114,31,72,31,31,31,48,31,48,30,227,31,145,31,121,31,235,31,74,31,80,31,80,30,152,31,78,31,251,31,165,31,165,30,112,31,160,31,29,31,29,30,166,31,189,31,192,31,221,31,113,31,203,31,1,31,216,31,196,31,164,31,42,31,15,31,64,31,64,30,191,31,163,31,246,31,246,30,246,29,185,31,164,31,24,31,196,31,112,31,44,31,85,31,67,31,161,31,161,30,139,31,161,31,85,31,235,31,183,31,163,31,33,31,58,31,58,30,196,31,41,31,95,31,96,31,131,31,6,31,6,30,144,31,22,31,125,31,137,31,137,30,52,31,11,31,11,30,241,31,52,31,52,30,52,29,203,31,154,31,177,31,119,31,116,31,158,31,117,31,122,31,178,31,178,30,178,29,132,31,255,31,145,31,85,31,21,31,243,31,14,31,194,31,36,31,238,31,238,30,238,29,21,31,64,31,51,31,115,31,223,31,125,31,44,31,197,31,115,31,6,31,38,31,48,31,102,31,81,31,142,31,198,31,198,30,230,31,114,31,114,30,225,31,212,31,199,31,199,30,241,31,241,30,12,31,43,31,92,31,165,31,140,31,68,31,138,31,167,31,46,31,46,30,215,31,127,31,2,31,41,31,162,31,75,31,75,30,13,31,120,31,249,31,122,31,220,31,117,31,117,30,155,31,49,31,100,31,72,31,105,31,4,31,76,31,90,31,1,31,178,31,75,31,75,30,75,29,101,31,207,31,207,30,35,31,35,30,146,31,146,30,78,31,250,31,141,31,29,31,220,31,198,31,198,30,171,31,110,31,237,31,167,31,178,31,178,30,178,29,14,31,75,31,84,31,12,31,40,31,94,31,159,31,149,31,36,31,91,31,91,30,72,31,79,31,211,31,124,31,124,30,74,31,24,31,133,31,240,31,69,31,49,31,243,31,197,31,133,31,133,30,208,31,24,31,245,31,245,30,136,31,136,30,136,29,132,31,217,31,190,31,243,31,105,31,140,31,22,31,165,31,175,31,93,31,234,31,177,31,96,31,133,31,30,31,30,30,145,31,122,31,200,31,200,30,241,31,202,31,249,31,200,31,11,31,156,31,156,30,91,31,139,31,139,30,145,31,240,31,240,30,215,31,226,31,181,31,102,31,102,30,41,31,226,31,65,31,65,30,65,29,250,31,235,31,196,31,220,31,9,31,75,31,120,31,120,30,163,31,91,31,48,31,111,31,111,30,70,31,135,31,134,31,59,31,229,31,209,31,209,30,154,31,125,31,102,31,177,31,8,31,153,31,134,31,134,30,96,31,43,31,238,31,233,31,50,31,50,30,172,31,81,31,10,31,84,31,99,31,127,31,127,30,210,31,210,30,229,31,244,31,186,31,1,31,231,31,202,31,122,31,122,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
