-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1020;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,85,0,83,0,160,0,194,0,77,0,0,0,0,0,1,0,0,0,0,0,67,0,73,0,26,0,106,0,0,0,0,0,0,0,243,0,97,0,248,0,0,0,198,0,12,0,233,0,15,0,65,0,226,0,23,0,0,0,129,0,59,0,174,0,0,0,130,0,54,0,217,0,195,0,110,0,117,0,5,0,99,0,153,0,67,0,226,0,134,0,43,0,106,0,114,0,205,0,0,0,1,0,0,0,212,0,0,0,205,0,93,0,0,0,231,0,37,0,19,0,23,0,131,0,181,0,0,0,0,0,89,0,4,0,0,0,142,0,99,0,0,0,69,0,23,0,243,0,252,0,253,0,64,0,29,0,228,0,79,0,0,0,166,0,12,0,10,0,0,0,44,0,130,0,232,0,134,0,0,0,34,0,103,0,117,0,254,0,44,0,28,0,71,0,170,0,0,0,145,0,0,0,0,0,90,0,226,0,132,0,175,0,0,0,198,0,192,0,198,0,252,0,168,0,111,0,253,0,0,0,0,0,255,0,105,0,241,0,224,0,84,0,79,0,0,0,69,0,26,0,54,0,218,0,0,0,65,0,164,0,165,0,108,0,107,0,186,0,72,0,0,0,14,0,155,0,216,0,0,0,0,0,0,0,0,0,112,0,0,0,0,0,116,0,84,0,152,0,0,0,0,0,114,0,0,0,138,0,218,0,0,0,122,0,49,0,0,0,175,0,0,0,106,0,226,0,44,0,139,0,101,0,171,0,159,0,0,0,25,0,43,0,249,0,244,0,232,0,0,0,0,0,148,0,194,0,255,0,252,0,0,0,163,0,237,0,4,0,0,0,0,0,185,0,89,0,253,0,158,0,233,0,12,0,4,0,0,0,231,0,170,0,0,0,169,0,151,0,0,0,198,0,119,0,138,0,137,0,224,0,50,0,0,0,70,0,78,0,17,0,28,0,205,0,12,0,0,0,120,0,0,0,24,0,129,0,224,0,0,0,0,0,145,0,167,0,170,0,0,0,9,0,147,0,0,0,116,0,88,0,0,0,242,0,145,0,128,0,100,0,1,0,110,0,239,0,0,0,218,0,197,0,55,0,233,0,147,0,145,0,163,0,58,0,213,0,123,0,0,0,82,0,158,0,0,0,160,0,184,0,16,0,105,0,51,0,217,0,0,0,113,0,184,0,189,0,251,0,0,0,133,0,92,0,127,0,165,0,0,0,147,0,168,0,0,0,0,0,162,0,59,0,93,0,245,0,0,0,168,0,167,0,0,0,140,0,59,0,184,0,0,0,2,0,203,0,0,0,226,0,0,0,65,0,198,0,245,0,174,0,33,0,125,0,0,0,46,0,165,0,148,0,110,0,3,0,242,0,0,0,151,0,65,0,0,0,154,0,64,0,119,0,0,0,229,0,31,0,98,0,0,0,102,0,233,0,0,0,87,0,155,0,171,0,144,0,229,0,208,0,83,0,253,0,0,0,11,0,233,0,70,0,0,0,2,0,103,0,87,0,246,0,106,0,255,0,39,0,176,0,75,0,210,0,68,0,12,0,130,0,186,0,125,0,0,0,121,0,240,0,202,0,164,0,213,0,0,0,161,0,158,0,164,0,35,0,0,0,0,0,3,0,0,0,43,0,0,0,0,0,135,0,98,0,0,0,235,0,228,0,111,0,28,0,0,0,0,0,112,0,0,0,118,0,195,0,123,0,84,0,0,0,32,0,194,0,51,0,121,0,23,0,4,0,67,0,23,0,0,0,156,0,0,0,146,0,196,0,4,0,199,0,16,0,72,0,0,0,4,0,112,0,58,0,136,0,203,0,52,0,193,0,0,0,0,0,105,0,154,0,116,0,20,0,202,0,34,0,7,0,56,0,61,0,228,0,173,0,160,0,0,0,0,0,0,0,145,0,36,0,125,0,213,0,21,0,216,0,82,0,67,0,0,0,53,0,64,0,223,0,78,0,125,0,0,0,167,0,227,0,89,0,182,0,166,0,167,0,188,0,118,0,69,0,223,0,0,0,109,0,56,0,102,0,0,0,83,0,109,0,0,0,160,0,183,0,59,0,43,0,87,0,187,0,94,0,32,0,0,0,149,0,252,0,180,0,16,0,0,0,142,0,103,0,35,0,213,0,219,0,9,0,126,0,236,0,207,0,90,0,0,0,119,0,0,0,244,0,36,0,245,0,114,0,0,0,167,0,0,0,250,0,147,0,97,0,184,0,210,0,44,0,234,0,34,0,0,0,87,0,94,0,159,0,123,0,231,0,156,0,151,0,80,0,24,0,78,0,71,0,0,0,159,0,109,0,179,0,209,0,0,0,0,0,4,0,193,0,209,0,194,0,21,0,0,0,9,0,11,0,228,0,195,0,206,0,0,0,154,0,242,0,7,0,195,0,75,0,191,0,98,0,79,0,82,0,165,0,119,0,79,0,79,0,0,0,0,0,240,0,4,0,172,0,144,0,148,0,249,0,0,0,112,0,196,0,172,0,155,0,5,0,73,0,157,0,121,0,223,0,70,0,246,0,0,0,159,0,138,0,31,0,41,0,194,0,217,0,1,0,93,0,176,0,133,0,28,0,0,0,0,0,113,0,9,0,0,0,0,0,250,0,87,0,153,0,213,0,11,0,0,0,254,0,226,0,0,0,0,0,0,0,80,0,252,0,0,0,0,0,0,0,7,0,0,0,0,0,229,0,0,0,0,0,66,0,17,0,0,0,176,0,0,0,150,0,85,0,181,0,164,0,183,0,5,0,161,0,147,0,209,0,50,0,91,0,156,0,0,0,24,0,200,0,0,0,145,0,250,0,0,0,0,0,0,0,100,0,223,0,77,0,222,0,9,0,135,0,55,0,246,0,116,0,181,0,122,0,88,0,244,0,0,0,190,0,0,0,150,0,19,0,0,0,126,0,152,0,0,0,207,0,138,0,240,0,233,0,67,0,105,0,211,0,248,0,206,0,231,0,0,0,210,0,0,0,0,0,252,0,82,0,93,0,124,0,0,0,236,0,104,0,0,0,0,0,63,0,20,0,100,0,36,0,190,0,161,0,0,0,168,0,209,0,114,0,117,0,100,0,0,0,14,0,0,0,41,0,0,0,72,0,0,0,95,0,16,0,210,0,67,0,143,0,204,0,35,0,61,0,0,0,0,0,222,0,132,0,216,0,76,0,0,0,179,0,186,0,84,0,232,0,0,0,4,0,112,0,105,0,0,0,0,0,25,0,0,0,157,0,20,0,188,0,0,0,65,0,191,0,188,0,92,0,0,0,40,0,174,0,56,0,97,0,183,0,16,0,0,0,33,0,72,0,148,0,54,0,212,0,91,0,212,0,65,0,48,0,188,0,245,0,0,0,45,0,195,0,234,0,175,0,121,0,0,0,197,0,166,0,78,0,112,0,38,0,70,0,245,0,181,0,6,0,225,0,35,0,246,0,12,0,119,0,62,0,37,0,126,0,186,0,4,0,0,0,9,0,200,0,0,0,98,0,255,0,181,0,217,0,242,0,34,0,240,0,49,0,0,0,104,0,0,0,0,0,198,0,4,0,23,0,180,0,109,0,180,0,44,0,50,0,0,0,0,0,0,0,110,0,208,0,0,0,36,0,188,0,1,0,0,0,140,0,202,0,54,0,0,0,8,0,65,0,0,0,102,0,0,0,80,0,70,0,213,0,155,0,210,0,195,0,129,0,212,0,139,0,0,0,190,0,59,0,219,0,112,0,128,0,192,0,86,0,170,0,61,0,0,0,235,0,205,0,77,0,121,0,246,0,0,0,90,0,0,0,0,0,5,0,68,0,239,0,0,0,0,0,191,0,173,0,173,0,208,0,67,0,213,0,59,0,112,0,121,0,217,0,0,0,148,0,41,0,143,0,44,0,227,0,24,0,241,0,253,0,32,0,91,0,157,0,121,0,20,0,37,0,169,0,0,0,96,0,0,0,0,0,142,0,57,0,0,0,151,0,153,0,207,0,21,0,52,0,206,0,129,0,221,0,168,0,0,0,7,0,18,0,16,0,240,0,120,0,0,0,186,0,101,0,70,0,0,0,72,0,162,0,246,0,0,0,238,0,53,0,61,0,58,0,162,0,31,0,238,0,0,0,5,0,62,0,52,0,169,0,200,0,141,0,47,0,0,0,1,0,55,0,151,0,18,0,91,0,109,0,198,0,176,0,162,0,81,0,9,0,200,0,38,0,82,0,151,0,0,0,0,0,0,0,103,0,107,0,2,0,0,0,0,0,138,0,236,0,188,0,0,0,0,0,203,0,60,0,173,0,64,0,0,0,0,0,0,0,236,0,221,0,62,0,246,0,253,0,163,0,79,0,37,0,87,0,82,0,181,0,160,0,204,0,214,0,3,0,147,0,100,0,0,0,100,0,149,0,211,0,107,0,86,0,211,0,83,0,0,0,168,0,60,0,0,0,117,0,124,0,1,0,212,0,108,0,78,0,108,0,116,0,103,0,0,0,71,0,0,0,95,0,0,0,0,0,0,0,10,0,235,0,67,0,0,0,0,0,153,0,0,0,0,0,0,0,0,0,228,0,19,0,0,0,239,0,217,0,6,0,0,0);
signal scenario_full  : scenario_type := (0,0,85,31,83,31,160,31,194,31,77,31,77,30,77,29,1,31,1,30,1,29,67,31,73,31,26,31,106,31,106,30,106,29,106,28,243,31,97,31,248,31,248,30,198,31,12,31,233,31,15,31,65,31,226,31,23,31,23,30,129,31,59,31,174,31,174,30,130,31,54,31,217,31,195,31,110,31,117,31,5,31,99,31,153,31,67,31,226,31,134,31,43,31,106,31,114,31,205,31,205,30,1,31,1,30,212,31,212,30,205,31,93,31,93,30,231,31,37,31,19,31,23,31,131,31,181,31,181,30,181,29,89,31,4,31,4,30,142,31,99,31,99,30,69,31,23,31,243,31,252,31,253,31,64,31,29,31,228,31,79,31,79,30,166,31,12,31,10,31,10,30,44,31,130,31,232,31,134,31,134,30,34,31,103,31,117,31,254,31,44,31,28,31,71,31,170,31,170,30,145,31,145,30,145,29,90,31,226,31,132,31,175,31,175,30,198,31,192,31,198,31,252,31,168,31,111,31,253,31,253,30,253,29,255,31,105,31,241,31,224,31,84,31,79,31,79,30,69,31,26,31,54,31,218,31,218,30,65,31,164,31,165,31,108,31,107,31,186,31,72,31,72,30,14,31,155,31,216,31,216,30,216,29,216,28,216,27,112,31,112,30,112,29,116,31,84,31,152,31,152,30,152,29,114,31,114,30,138,31,218,31,218,30,122,31,49,31,49,30,175,31,175,30,106,31,226,31,44,31,139,31,101,31,171,31,159,31,159,30,25,31,43,31,249,31,244,31,232,31,232,30,232,29,148,31,194,31,255,31,252,31,252,30,163,31,237,31,4,31,4,30,4,29,185,31,89,31,253,31,158,31,233,31,12,31,4,31,4,30,231,31,170,31,170,30,169,31,151,31,151,30,198,31,119,31,138,31,137,31,224,31,50,31,50,30,70,31,78,31,17,31,28,31,205,31,12,31,12,30,120,31,120,30,24,31,129,31,224,31,224,30,224,29,145,31,167,31,170,31,170,30,9,31,147,31,147,30,116,31,88,31,88,30,242,31,145,31,128,31,100,31,1,31,110,31,239,31,239,30,218,31,197,31,55,31,233,31,147,31,145,31,163,31,58,31,213,31,123,31,123,30,82,31,158,31,158,30,160,31,184,31,16,31,105,31,51,31,217,31,217,30,113,31,184,31,189,31,251,31,251,30,133,31,92,31,127,31,165,31,165,30,147,31,168,31,168,30,168,29,162,31,59,31,93,31,245,31,245,30,168,31,167,31,167,30,140,31,59,31,184,31,184,30,2,31,203,31,203,30,226,31,226,30,65,31,198,31,245,31,174,31,33,31,125,31,125,30,46,31,165,31,148,31,110,31,3,31,242,31,242,30,151,31,65,31,65,30,154,31,64,31,119,31,119,30,229,31,31,31,98,31,98,30,102,31,233,31,233,30,87,31,155,31,171,31,144,31,229,31,208,31,83,31,253,31,253,30,11,31,233,31,70,31,70,30,2,31,103,31,87,31,246,31,106,31,255,31,39,31,176,31,75,31,210,31,68,31,12,31,130,31,186,31,125,31,125,30,121,31,240,31,202,31,164,31,213,31,213,30,161,31,158,31,164,31,35,31,35,30,35,29,3,31,3,30,43,31,43,30,43,29,135,31,98,31,98,30,235,31,228,31,111,31,28,31,28,30,28,29,112,31,112,30,118,31,195,31,123,31,84,31,84,30,32,31,194,31,51,31,121,31,23,31,4,31,67,31,23,31,23,30,156,31,156,30,146,31,196,31,4,31,199,31,16,31,72,31,72,30,4,31,112,31,58,31,136,31,203,31,52,31,193,31,193,30,193,29,105,31,154,31,116,31,20,31,202,31,34,31,7,31,56,31,61,31,228,31,173,31,160,31,160,30,160,29,160,28,145,31,36,31,125,31,213,31,21,31,216,31,82,31,67,31,67,30,53,31,64,31,223,31,78,31,125,31,125,30,167,31,227,31,89,31,182,31,166,31,167,31,188,31,118,31,69,31,223,31,223,30,109,31,56,31,102,31,102,30,83,31,109,31,109,30,160,31,183,31,59,31,43,31,87,31,187,31,94,31,32,31,32,30,149,31,252,31,180,31,16,31,16,30,142,31,103,31,35,31,213,31,219,31,9,31,126,31,236,31,207,31,90,31,90,30,119,31,119,30,244,31,36,31,245,31,114,31,114,30,167,31,167,30,250,31,147,31,97,31,184,31,210,31,44,31,234,31,34,31,34,30,87,31,94,31,159,31,123,31,231,31,156,31,151,31,80,31,24,31,78,31,71,31,71,30,159,31,109,31,179,31,209,31,209,30,209,29,4,31,193,31,209,31,194,31,21,31,21,30,9,31,11,31,228,31,195,31,206,31,206,30,154,31,242,31,7,31,195,31,75,31,191,31,98,31,79,31,82,31,165,31,119,31,79,31,79,31,79,30,79,29,240,31,4,31,172,31,144,31,148,31,249,31,249,30,112,31,196,31,172,31,155,31,5,31,73,31,157,31,121,31,223,31,70,31,246,31,246,30,159,31,138,31,31,31,41,31,194,31,217,31,1,31,93,31,176,31,133,31,28,31,28,30,28,29,113,31,9,31,9,30,9,29,250,31,87,31,153,31,213,31,11,31,11,30,254,31,226,31,226,30,226,29,226,28,80,31,252,31,252,30,252,29,252,28,7,31,7,30,7,29,229,31,229,30,229,29,66,31,17,31,17,30,176,31,176,30,150,31,85,31,181,31,164,31,183,31,5,31,161,31,147,31,209,31,50,31,91,31,156,31,156,30,24,31,200,31,200,30,145,31,250,31,250,30,250,29,250,28,100,31,223,31,77,31,222,31,9,31,135,31,55,31,246,31,116,31,181,31,122,31,88,31,244,31,244,30,190,31,190,30,150,31,19,31,19,30,126,31,152,31,152,30,207,31,138,31,240,31,233,31,67,31,105,31,211,31,248,31,206,31,231,31,231,30,210,31,210,30,210,29,252,31,82,31,93,31,124,31,124,30,236,31,104,31,104,30,104,29,63,31,20,31,100,31,36,31,190,31,161,31,161,30,168,31,209,31,114,31,117,31,100,31,100,30,14,31,14,30,41,31,41,30,72,31,72,30,95,31,16,31,210,31,67,31,143,31,204,31,35,31,61,31,61,30,61,29,222,31,132,31,216,31,76,31,76,30,179,31,186,31,84,31,232,31,232,30,4,31,112,31,105,31,105,30,105,29,25,31,25,30,157,31,20,31,188,31,188,30,65,31,191,31,188,31,92,31,92,30,40,31,174,31,56,31,97,31,183,31,16,31,16,30,33,31,72,31,148,31,54,31,212,31,91,31,212,31,65,31,48,31,188,31,245,31,245,30,45,31,195,31,234,31,175,31,121,31,121,30,197,31,166,31,78,31,112,31,38,31,70,31,245,31,181,31,6,31,225,31,35,31,246,31,12,31,119,31,62,31,37,31,126,31,186,31,4,31,4,30,9,31,200,31,200,30,98,31,255,31,181,31,217,31,242,31,34,31,240,31,49,31,49,30,104,31,104,30,104,29,198,31,4,31,23,31,180,31,109,31,180,31,44,31,50,31,50,30,50,29,50,28,110,31,208,31,208,30,36,31,188,31,1,31,1,30,140,31,202,31,54,31,54,30,8,31,65,31,65,30,102,31,102,30,80,31,70,31,213,31,155,31,210,31,195,31,129,31,212,31,139,31,139,30,190,31,59,31,219,31,112,31,128,31,192,31,86,31,170,31,61,31,61,30,235,31,205,31,77,31,121,31,246,31,246,30,90,31,90,30,90,29,5,31,68,31,239,31,239,30,239,29,191,31,173,31,173,31,208,31,67,31,213,31,59,31,112,31,121,31,217,31,217,30,148,31,41,31,143,31,44,31,227,31,24,31,241,31,253,31,32,31,91,31,157,31,121,31,20,31,37,31,169,31,169,30,96,31,96,30,96,29,142,31,57,31,57,30,151,31,153,31,207,31,21,31,52,31,206,31,129,31,221,31,168,31,168,30,7,31,18,31,16,31,240,31,120,31,120,30,186,31,101,31,70,31,70,30,72,31,162,31,246,31,246,30,238,31,53,31,61,31,58,31,162,31,31,31,238,31,238,30,5,31,62,31,52,31,169,31,200,31,141,31,47,31,47,30,1,31,55,31,151,31,18,31,91,31,109,31,198,31,176,31,162,31,81,31,9,31,200,31,38,31,82,31,151,31,151,30,151,29,151,28,103,31,107,31,2,31,2,30,2,29,138,31,236,31,188,31,188,30,188,29,203,31,60,31,173,31,64,31,64,30,64,29,64,28,236,31,221,31,62,31,246,31,253,31,163,31,79,31,37,31,87,31,82,31,181,31,160,31,204,31,214,31,3,31,147,31,100,31,100,30,100,31,149,31,211,31,107,31,86,31,211,31,83,31,83,30,168,31,60,31,60,30,117,31,124,31,1,31,212,31,108,31,78,31,108,31,116,31,103,31,103,30,71,31,71,30,95,31,95,30,95,29,95,28,10,31,235,31,67,31,67,30,67,29,153,31,153,30,153,29,153,28,153,27,228,31,19,31,19,30,239,31,217,31,6,31,6,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
