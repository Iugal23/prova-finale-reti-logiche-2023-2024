-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_682 is
end project_tb_682;

architecture project_tb_arch_682 of project_tb_682 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 356;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,19,0,0,0,89,0,248,0,200,0,0,0,138,0,151,0,206,0,0,0,97,0,220,0,39,0,97,0,0,0,139,0,0,0,16,0,199,0,125,0,50,0,254,0,133,0,124,0,104,0,12,0,135,0,0,0,58,0,70,0,121,0,157,0,180,0,210,0,89,0,206,0,36,0,46,0,98,0,122,0,109,0,152,0,135,0,25,0,34,0,165,0,131,0,212,0,119,0,32,0,0,0,222,0,144,0,167,0,0,0,254,0,238,0,59,0,58,0,87,0,109,0,112,0,67,0,81,0,0,0,149,0,169,0,233,0,213,0,128,0,9,0,0,0,0,0,160,0,175,0,38,0,0,0,201,0,45,0,50,0,0,0,0,0,137,0,88,0,236,0,0,0,0,0,165,0,0,0,98,0,0,0,0,0,104,0,129,0,160,0,158,0,31,0,253,0,184,0,139,0,238,0,232,0,114,0,206,0,189,0,23,0,0,0,220,0,121,0,59,0,5,0,146,0,214,0,240,0,143,0,151,0,147,0,38,0,233,0,23,0,0,0,73,0,94,0,190,0,0,0,224,0,248,0,183,0,227,0,0,0,71,0,112,0,0,0,79,0,196,0,239,0,0,0,0,0,211,0,0,0,153,0,0,0,128,0,186,0,205,0,0,0,162,0,123,0,11,0,0,0,0,0,0,0,185,0,118,0,65,0,0,0,129,0,63,0,0,0,0,0,146,0,69,0,38,0,173,0,17,0,23,0,19,0,0,0,255,0,163,0,0,0,228,0,199,0,40,0,213,0,89,0,0,0,0,0,32,0,84,0,80,0,92,0,252,0,140,0,121,0,181,0,118,0,0,0,215,0,95,0,200,0,2,0,43,0,55,0,169,0,161,0,18,0,31,0,175,0,144,0,251,0,0,0,170,0,107,0,215,0,150,0,222,0,228,0,239,0,226,0,229,0,196,0,254,0,142,0,153,0,48,0,246,0,228,0,90,0,251,0,217,0,197,0,0,0,0,0,248,0,220,0,235,0,115,0,0,0,188,0,225,0,24,0,2,0,100,0,12,0,0,0,24,0,113,0,235,0,139,0,0,0,0,0,152,0,245,0,186,0,222,0,45,0,0,0,68,0,228,0,59,0,91,0,239,0,172,0,115,0,113,0,0,0,22,0,232,0,5,0,196,0,33,0,0,0,179,0,0,0,154,0,154,0,112,0,64,0,95,0,7,0,143,0,81,0,123,0,63,0,0,0,152,0,131,0,32,0,60,0,241,0,0,0,252,0,61,0,167,0,0,0,8,0,122,0,236,0,228,0,90,0,0,0,0,0,46,0,43,0,175,0,212,0,100,0,185,0,0,0,0,0,179,0,76,0,159,0,213,0,12,0,4,0,0,0,167,0,158,0,153,0,190,0,72,0,48,0,19,0,200,0,200,0,40,0,52,0,210,0,0,0,89,0,0,0,212,0,46,0,250,0,84,0,22,0,14,0,216,0,55,0,249,0,175,0,191,0,247,0,157,0,12,0,38,0,0,0,199,0,68,0,39,0,146,0,0,0,0,0,19,0,195,0,118,0,108,0,0,0,78,0,218,0,53,0,32,0,137,0);
signal scenario_full  : scenario_type := (0,0,19,31,19,30,89,31,248,31,200,31,200,30,138,31,151,31,206,31,206,30,97,31,220,31,39,31,97,31,97,30,139,31,139,30,16,31,199,31,125,31,50,31,254,31,133,31,124,31,104,31,12,31,135,31,135,30,58,31,70,31,121,31,157,31,180,31,210,31,89,31,206,31,36,31,46,31,98,31,122,31,109,31,152,31,135,31,25,31,34,31,165,31,131,31,212,31,119,31,32,31,32,30,222,31,144,31,167,31,167,30,254,31,238,31,59,31,58,31,87,31,109,31,112,31,67,31,81,31,81,30,149,31,169,31,233,31,213,31,128,31,9,31,9,30,9,29,160,31,175,31,38,31,38,30,201,31,45,31,50,31,50,30,50,29,137,31,88,31,236,31,236,30,236,29,165,31,165,30,98,31,98,30,98,29,104,31,129,31,160,31,158,31,31,31,253,31,184,31,139,31,238,31,232,31,114,31,206,31,189,31,23,31,23,30,220,31,121,31,59,31,5,31,146,31,214,31,240,31,143,31,151,31,147,31,38,31,233,31,23,31,23,30,73,31,94,31,190,31,190,30,224,31,248,31,183,31,227,31,227,30,71,31,112,31,112,30,79,31,196,31,239,31,239,30,239,29,211,31,211,30,153,31,153,30,128,31,186,31,205,31,205,30,162,31,123,31,11,31,11,30,11,29,11,28,185,31,118,31,65,31,65,30,129,31,63,31,63,30,63,29,146,31,69,31,38,31,173,31,17,31,23,31,19,31,19,30,255,31,163,31,163,30,228,31,199,31,40,31,213,31,89,31,89,30,89,29,32,31,84,31,80,31,92,31,252,31,140,31,121,31,181,31,118,31,118,30,215,31,95,31,200,31,2,31,43,31,55,31,169,31,161,31,18,31,31,31,175,31,144,31,251,31,251,30,170,31,107,31,215,31,150,31,222,31,228,31,239,31,226,31,229,31,196,31,254,31,142,31,153,31,48,31,246,31,228,31,90,31,251,31,217,31,197,31,197,30,197,29,248,31,220,31,235,31,115,31,115,30,188,31,225,31,24,31,2,31,100,31,12,31,12,30,24,31,113,31,235,31,139,31,139,30,139,29,152,31,245,31,186,31,222,31,45,31,45,30,68,31,228,31,59,31,91,31,239,31,172,31,115,31,113,31,113,30,22,31,232,31,5,31,196,31,33,31,33,30,179,31,179,30,154,31,154,31,112,31,64,31,95,31,7,31,143,31,81,31,123,31,63,31,63,30,152,31,131,31,32,31,60,31,241,31,241,30,252,31,61,31,167,31,167,30,8,31,122,31,236,31,228,31,90,31,90,30,90,29,46,31,43,31,175,31,212,31,100,31,185,31,185,30,185,29,179,31,76,31,159,31,213,31,12,31,4,31,4,30,167,31,158,31,153,31,190,31,72,31,48,31,19,31,200,31,200,31,40,31,52,31,210,31,210,30,89,31,89,30,212,31,46,31,250,31,84,31,22,31,14,31,216,31,55,31,249,31,175,31,191,31,247,31,157,31,12,31,38,31,38,30,199,31,68,31,39,31,146,31,146,30,146,29,19,31,195,31,118,31,108,31,108,30,78,31,218,31,53,31,32,31,137,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
