-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 396;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,138,0,86,0,137,0,143,0,38,0,168,0,195,0,182,0,51,0,182,0,121,0,156,0,218,0,198,0,242,0,86,0,156,0,0,0,104,0,0,0,197,0,0,0,0,0,0,0,32,0,234,0,5,0,20,0,0,0,0,0,0,0,67,0,232,0,0,0,80,0,198,0,52,0,204,0,119,0,92,0,12,0,0,0,198,0,7,0,188,0,109,0,0,0,156,0,13,0,215,0,0,0,217,0,196,0,252,0,60,0,207,0,0,0,0,0,74,0,151,0,0,0,166,0,28,0,44,0,0,0,137,0,78,0,175,0,0,0,169,0,59,0,40,0,72,0,0,0,0,0,184,0,0,0,0,0,111,0,0,0,141,0,138,0,97,0,0,0,76,0,19,0,154,0,45,0,95,0,210,0,252,0,79,0,16,0,50,0,94,0,230,0,4,0,32,0,133,0,69,0,247,0,0,0,29,0,84,0,124,0,236,0,232,0,0,0,148,0,194,0,141,0,75,0,0,0,46,0,211,0,201,0,218,0,0,0,87,0,212,0,111,0,0,0,69,0,0,0,13,0,69,0,235,0,7,0,222,0,28,0,130,0,124,0,181,0,71,0,175,0,59,0,191,0,139,0,0,0,128,0,5,0,60,0,0,0,2,0,0,0,200,0,0,0,124,0,28,0,64,0,112,0,224,0,241,0,158,0,22,0,0,0,240,0,0,0,0,0,132,0,231,0,102,0,24,0,35,0,75,0,15,0,77,0,75,0,101,0,113,0,22,0,75,0,24,0,0,0,109,0,230,0,32,0,0,0,202,0,0,0,53,0,152,0,0,0,252,0,151,0,0,0,65,0,145,0,9,0,123,0,0,0,97,0,144,0,175,0,0,0,177,0,183,0,0,0,33,0,0,0,16,0,172,0,78,0,60,0,128,0,245,0,171,0,172,0,146,0,74,0,227,0,117,0,178,0,215,0,83,0,0,0,0,0,60,0,131,0,74,0,31,0,210,0,0,0,90,0,36,0,226,0,93,0,89,0,0,0,195,0,0,0,154,0,93,0,254,0,0,0,26,0,0,0,117,0,76,0,120,0,107,0,191,0,241,0,148,0,251,0,217,0,15,0,0,0,250,0,207,0,240,0,108,0,255,0,179,0,10,0,52,0,158,0,206,0,94,0,35,0,0,0,132,0,183,0,103,0,0,0,0,0,220,0,130,0,157,0,0,0,77,0,199,0,158,0,90,0,195,0,202,0,225,0,0,0,217,0,168,0,0,0,36,0,114,0,219,0,0,0,0,0,213,0,43,0,52,0,159,0,153,0,214,0,210,0,123,0,128,0,15,0,200,0,102,0,136,0,82,0,232,0,225,0,191,0,219,0,0,0,146,0,239,0,128,0,94,0,0,0,38,0,125,0,71,0,84,0,212,0,137,0,64,0,78,0,3,0,55,0,226,0,40,0,57,0,238,0,64,0,215,0,9,0,190,0,193,0,106,0,230,0,154,0,15,0,38,0,0,0,167,0,236,0,73,0,105,0,135,0,165,0,185,0,42,0,0,0,122,0,203,0,138,0,0,0,250,0,8,0,102,0,31,0,228,0,226,0,212,0,226,0,140,0,173,0,214,0,244,0,52,0,0,0,0,0,233,0,187,0,13,0,4,0,82,0,68,0,0,0,106,0,202,0,0,0,95,0,187,0,134,0,104,0,14,0,171,0,206,0,161,0,60,0,0,0,215,0,64,0,145,0,130,0,161,0,235,0,196,0,39,0,250,0,198,0,212,0,227,0);
signal scenario_full  : scenario_type := (0,0,138,31,86,31,137,31,143,31,38,31,168,31,195,31,182,31,51,31,182,31,121,31,156,31,218,31,198,31,242,31,86,31,156,31,156,30,104,31,104,30,197,31,197,30,197,29,197,28,32,31,234,31,5,31,20,31,20,30,20,29,20,28,67,31,232,31,232,30,80,31,198,31,52,31,204,31,119,31,92,31,12,31,12,30,198,31,7,31,188,31,109,31,109,30,156,31,13,31,215,31,215,30,217,31,196,31,252,31,60,31,207,31,207,30,207,29,74,31,151,31,151,30,166,31,28,31,44,31,44,30,137,31,78,31,175,31,175,30,169,31,59,31,40,31,72,31,72,30,72,29,184,31,184,30,184,29,111,31,111,30,141,31,138,31,97,31,97,30,76,31,19,31,154,31,45,31,95,31,210,31,252,31,79,31,16,31,50,31,94,31,230,31,4,31,32,31,133,31,69,31,247,31,247,30,29,31,84,31,124,31,236,31,232,31,232,30,148,31,194,31,141,31,75,31,75,30,46,31,211,31,201,31,218,31,218,30,87,31,212,31,111,31,111,30,69,31,69,30,13,31,69,31,235,31,7,31,222,31,28,31,130,31,124,31,181,31,71,31,175,31,59,31,191,31,139,31,139,30,128,31,5,31,60,31,60,30,2,31,2,30,200,31,200,30,124,31,28,31,64,31,112,31,224,31,241,31,158,31,22,31,22,30,240,31,240,30,240,29,132,31,231,31,102,31,24,31,35,31,75,31,15,31,77,31,75,31,101,31,113,31,22,31,75,31,24,31,24,30,109,31,230,31,32,31,32,30,202,31,202,30,53,31,152,31,152,30,252,31,151,31,151,30,65,31,145,31,9,31,123,31,123,30,97,31,144,31,175,31,175,30,177,31,183,31,183,30,33,31,33,30,16,31,172,31,78,31,60,31,128,31,245,31,171,31,172,31,146,31,74,31,227,31,117,31,178,31,215,31,83,31,83,30,83,29,60,31,131,31,74,31,31,31,210,31,210,30,90,31,36,31,226,31,93,31,89,31,89,30,195,31,195,30,154,31,93,31,254,31,254,30,26,31,26,30,117,31,76,31,120,31,107,31,191,31,241,31,148,31,251,31,217,31,15,31,15,30,250,31,207,31,240,31,108,31,255,31,179,31,10,31,52,31,158,31,206,31,94,31,35,31,35,30,132,31,183,31,103,31,103,30,103,29,220,31,130,31,157,31,157,30,77,31,199,31,158,31,90,31,195,31,202,31,225,31,225,30,217,31,168,31,168,30,36,31,114,31,219,31,219,30,219,29,213,31,43,31,52,31,159,31,153,31,214,31,210,31,123,31,128,31,15,31,200,31,102,31,136,31,82,31,232,31,225,31,191,31,219,31,219,30,146,31,239,31,128,31,94,31,94,30,38,31,125,31,71,31,84,31,212,31,137,31,64,31,78,31,3,31,55,31,226,31,40,31,57,31,238,31,64,31,215,31,9,31,190,31,193,31,106,31,230,31,154,31,15,31,38,31,38,30,167,31,236,31,73,31,105,31,135,31,165,31,185,31,42,31,42,30,122,31,203,31,138,31,138,30,250,31,8,31,102,31,31,31,228,31,226,31,212,31,226,31,140,31,173,31,214,31,244,31,52,31,52,30,52,29,233,31,187,31,13,31,4,31,82,31,68,31,68,30,106,31,202,31,202,30,95,31,187,31,134,31,104,31,14,31,171,31,206,31,161,31,60,31,60,30,215,31,64,31,145,31,130,31,161,31,235,31,196,31,39,31,250,31,198,31,212,31,227,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
