-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_545 is
end project_tb_545;

architecture project_tb_arch_545 of project_tb_545 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 692;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (121,0,0,0,0,0,227,0,226,0,243,0,251,0,0,0,94,0,177,0,152,0,56,0,237,0,78,0,0,0,0,0,4,0,102,0,178,0,0,0,0,0,114,0,194,0,0,0,118,0,0,0,253,0,0,0,189,0,158,0,210,0,29,0,0,0,0,0,247,0,0,0,114,0,45,0,0,0,61,0,0,0,0,0,0,0,89,0,227,0,94,0,0,0,71,0,199,0,93,0,174,0,86,0,236,0,0,0,0,0,26,0,165,0,0,0,125,0,177,0,0,0,0,0,0,0,170,0,181,0,0,0,226,0,148,0,62,0,52,0,146,0,116,0,0,0,202,0,72,0,0,0,26,0,88,0,5,0,173,0,86,0,86,0,180,0,125,0,133,0,176,0,195,0,23,0,41,0,227,0,176,0,48,0,96,0,185,0,19,0,125,0,45,0,242,0,185,0,66,0,4,0,91,0,45,0,0,0,164,0,0,0,140,0,116,0,111,0,47,0,43,0,0,0,109,0,0,0,124,0,0,0,104,0,154,0,140,0,132,0,107,0,9,0,76,0,125,0,93,0,32,0,0,0,178,0,108,0,0,0,176,0,108,0,47,0,0,0,87,0,152,0,233,0,43,0,123,0,17,0,52,0,59,0,0,0,246,0,87,0,44,0,112,0,184,0,0,0,0,0,87,0,141,0,72,0,229,0,0,0,34,0,17,0,128,0,9,0,227,0,0,0,220,0,175,0,0,0,0,0,177,0,125,0,223,0,0,0,115,0,195,0,131,0,0,0,29,0,59,0,235,0,155,0,124,0,30,0,69,0,200,0,174,0,135,0,226,0,53,0,69,0,119,0,92,0,190,0,0,0,154,0,46,0,0,0,131,0,11,0,17,0,0,0,220,0,32,0,144,0,0,0,0,0,179,0,0,0,254,0,83,0,117,0,5,0,63,0,127,0,0,0,193,0,216,0,15,0,0,0,0,0,78,0,223,0,42,0,38,0,59,0,0,0,0,0,236,0,134,0,72,0,0,0,164,0,47,0,236,0,122,0,27,0,112,0,45,0,70,0,0,0,204,0,71,0,45,0,88,0,0,0,0,0,0,0,189,0,226,0,61,0,172,0,0,0,47,0,100,0,130,0,100,0,0,0,195,0,84,0,0,0,3,0,128,0,0,0,205,0,230,0,143,0,0,0,219,0,74,0,21,0,0,0,3,0,247,0,103,0,202,0,238,0,93,0,114,0,192,0,139,0,0,0,86,0,135,0,0,0,137,0,0,0,64,0,203,0,143,0,74,0,97,0,0,0,206,0,109,0,97,0,209,0,0,0,255,0,0,0,0,0,0,0,34,0,225,0,0,0,252,0,0,0,0,0,196,0,0,0,212,0,0,0,158,0,10,0,47,0,161,0,28,0,34,0,11,0,3,0,205,0,96,0,159,0,74,0,214,0,193,0,66,0,206,0,184,0,0,0,218,0,84,0,141,0,239,0,107,0,27,0,110,0,46,0,217,0,16,0,12,0,200,0,51,0,212,0,0,0,153,0,0,0,38,0,91,0,150,0,5,0,174,0,0,0,121,0,0,0,250,0,0,0,53,0,71,0,135,0,156,0,114,0,142,0,193,0,0,0,39,0,0,0,149,0,210,0,222,0,0,0,241,0,242,0,194,0,0,0,66,0,0,0,184,0,0,0,1,0,0,0,178,0,0,0,150,0,199,0,0,0,201,0,94,0,141,0,208,0,176,0,4,0,254,0,137,0,13,0,19,0,177,0,195,0,93,0,208,0,158,0,160,0,29,0,58,0,140,0,54,0,186,0,79,0,93,0,60,0,216,0,248,0,36,0,64,0,48,0,0,0,170,0,0,0,95,0,15,0,155,0,131,0,50,0,12,0,0,0,154,0,0,0,0,0,69,0,0,0,50,0,189,0,102,0,82,0,0,0,188,0,246,0,234,0,103,0,193,0,137,0,0,0,0,0,216,0,248,0,110,0,172,0,130,0,150,0,114,0,0,0,21,0,172,0,199,0,15,0,207,0,51,0,80,0,0,0,0,0,35,0,126,0,245,0,53,0,222,0,0,0,117,0,0,0,9,0,89,0,97,0,108,0,131,0,0,0,0,0,117,0,61,0,207,0,0,0,5,0,0,0,236,0,81,0,223,0,65,0,174,0,16,0,95,0,206,0,166,0,109,0,0,0,5,0,0,0,182,0,221,0,84,0,85,0,254,0,186,0,0,0,178,0,167,0,195,0,218,0,0,0,0,0,0,0,79,0,0,0,50,0,197,0,177,0,0,0,0,0,193,0,165,0,0,0,227,0,191,0,203,0,238,0,0,0,26,0,0,0,132,0,184,0,84,0,52,0,0,0,204,0,147,0,203,0,42,0,0,0,176,0,153,0,0,0,214,0,56,0,25,0,38,0,222,0,24,0,236,0,0,0,163,0,11,0,18,0,229,0,70,0,68,0,185,0,0,0,0,0,31,0,179,0,198,0,55,0,87,0,76,0,0,0,37,0,113,0,228,0,94,0,0,0,199,0,73,0,210,0,0,0,60,0,68,0,75,0,171,0,170,0,10,0,0,0,127,0,0,0,221,0,44,0,0,0,0,0,120,0,238,0,190,0,17,0,177,0,219,0,185,0,16,0,72,0,14,0,28,0,230,0,0,0,157,0,38,0,235,0,88,0,248,0,153,0,0,0,0,0,195,0,57,0,176,0,224,0,24,0,12,0,0,0,166,0,23,0,13,0,30,0,0,0,13,0,9,0,0,0,82,0,252,0,6,0,63,0,127,0,45,0,197,0,76,0,21,0,191,0,106,0,0,0,165,0,186,0,213,0,87,0,0,0,199,0,0,0,184,0,10,0,243,0,0,0,0,0,29,0,78,0,129,0,0,0,0,0,92,0,176,0,86,0,121,0,214,0,203,0,136,0,111,0,53,0,255,0,111,0,158,0,44,0,112,0,212,0,175,0,0,0,93,0,0,0,212,0,126,0,162,0,52,0,137,0,76,0,178,0,0,0,52,0,0,0,215,0,0,0,136,0,183,0,93,0,219,0,171,0,179,0,78,0,129,0,65,0,75,0,0,0,174,0,0,0,189,0,205,0,177,0,0,0);
signal scenario_full  : scenario_type := (121,31,121,30,121,29,227,31,226,31,243,31,251,31,251,30,94,31,177,31,152,31,56,31,237,31,78,31,78,30,78,29,4,31,102,31,178,31,178,30,178,29,114,31,194,31,194,30,118,31,118,30,253,31,253,30,189,31,158,31,210,31,29,31,29,30,29,29,247,31,247,30,114,31,45,31,45,30,61,31,61,30,61,29,61,28,89,31,227,31,94,31,94,30,71,31,199,31,93,31,174,31,86,31,236,31,236,30,236,29,26,31,165,31,165,30,125,31,177,31,177,30,177,29,177,28,170,31,181,31,181,30,226,31,148,31,62,31,52,31,146,31,116,31,116,30,202,31,72,31,72,30,26,31,88,31,5,31,173,31,86,31,86,31,180,31,125,31,133,31,176,31,195,31,23,31,41,31,227,31,176,31,48,31,96,31,185,31,19,31,125,31,45,31,242,31,185,31,66,31,4,31,91,31,45,31,45,30,164,31,164,30,140,31,116,31,111,31,47,31,43,31,43,30,109,31,109,30,124,31,124,30,104,31,154,31,140,31,132,31,107,31,9,31,76,31,125,31,93,31,32,31,32,30,178,31,108,31,108,30,176,31,108,31,47,31,47,30,87,31,152,31,233,31,43,31,123,31,17,31,52,31,59,31,59,30,246,31,87,31,44,31,112,31,184,31,184,30,184,29,87,31,141,31,72,31,229,31,229,30,34,31,17,31,128,31,9,31,227,31,227,30,220,31,175,31,175,30,175,29,177,31,125,31,223,31,223,30,115,31,195,31,131,31,131,30,29,31,59,31,235,31,155,31,124,31,30,31,69,31,200,31,174,31,135,31,226,31,53,31,69,31,119,31,92,31,190,31,190,30,154,31,46,31,46,30,131,31,11,31,17,31,17,30,220,31,32,31,144,31,144,30,144,29,179,31,179,30,254,31,83,31,117,31,5,31,63,31,127,31,127,30,193,31,216,31,15,31,15,30,15,29,78,31,223,31,42,31,38,31,59,31,59,30,59,29,236,31,134,31,72,31,72,30,164,31,47,31,236,31,122,31,27,31,112,31,45,31,70,31,70,30,204,31,71,31,45,31,88,31,88,30,88,29,88,28,189,31,226,31,61,31,172,31,172,30,47,31,100,31,130,31,100,31,100,30,195,31,84,31,84,30,3,31,128,31,128,30,205,31,230,31,143,31,143,30,219,31,74,31,21,31,21,30,3,31,247,31,103,31,202,31,238,31,93,31,114,31,192,31,139,31,139,30,86,31,135,31,135,30,137,31,137,30,64,31,203,31,143,31,74,31,97,31,97,30,206,31,109,31,97,31,209,31,209,30,255,31,255,30,255,29,255,28,34,31,225,31,225,30,252,31,252,30,252,29,196,31,196,30,212,31,212,30,158,31,10,31,47,31,161,31,28,31,34,31,11,31,3,31,205,31,96,31,159,31,74,31,214,31,193,31,66,31,206,31,184,31,184,30,218,31,84,31,141,31,239,31,107,31,27,31,110,31,46,31,217,31,16,31,12,31,200,31,51,31,212,31,212,30,153,31,153,30,38,31,91,31,150,31,5,31,174,31,174,30,121,31,121,30,250,31,250,30,53,31,71,31,135,31,156,31,114,31,142,31,193,31,193,30,39,31,39,30,149,31,210,31,222,31,222,30,241,31,242,31,194,31,194,30,66,31,66,30,184,31,184,30,1,31,1,30,178,31,178,30,150,31,199,31,199,30,201,31,94,31,141,31,208,31,176,31,4,31,254,31,137,31,13,31,19,31,177,31,195,31,93,31,208,31,158,31,160,31,29,31,58,31,140,31,54,31,186,31,79,31,93,31,60,31,216,31,248,31,36,31,64,31,48,31,48,30,170,31,170,30,95,31,15,31,155,31,131,31,50,31,12,31,12,30,154,31,154,30,154,29,69,31,69,30,50,31,189,31,102,31,82,31,82,30,188,31,246,31,234,31,103,31,193,31,137,31,137,30,137,29,216,31,248,31,110,31,172,31,130,31,150,31,114,31,114,30,21,31,172,31,199,31,15,31,207,31,51,31,80,31,80,30,80,29,35,31,126,31,245,31,53,31,222,31,222,30,117,31,117,30,9,31,89,31,97,31,108,31,131,31,131,30,131,29,117,31,61,31,207,31,207,30,5,31,5,30,236,31,81,31,223,31,65,31,174,31,16,31,95,31,206,31,166,31,109,31,109,30,5,31,5,30,182,31,221,31,84,31,85,31,254,31,186,31,186,30,178,31,167,31,195,31,218,31,218,30,218,29,218,28,79,31,79,30,50,31,197,31,177,31,177,30,177,29,193,31,165,31,165,30,227,31,191,31,203,31,238,31,238,30,26,31,26,30,132,31,184,31,84,31,52,31,52,30,204,31,147,31,203,31,42,31,42,30,176,31,153,31,153,30,214,31,56,31,25,31,38,31,222,31,24,31,236,31,236,30,163,31,11,31,18,31,229,31,70,31,68,31,185,31,185,30,185,29,31,31,179,31,198,31,55,31,87,31,76,31,76,30,37,31,113,31,228,31,94,31,94,30,199,31,73,31,210,31,210,30,60,31,68,31,75,31,171,31,170,31,10,31,10,30,127,31,127,30,221,31,44,31,44,30,44,29,120,31,238,31,190,31,17,31,177,31,219,31,185,31,16,31,72,31,14,31,28,31,230,31,230,30,157,31,38,31,235,31,88,31,248,31,153,31,153,30,153,29,195,31,57,31,176,31,224,31,24,31,12,31,12,30,166,31,23,31,13,31,30,31,30,30,13,31,9,31,9,30,82,31,252,31,6,31,63,31,127,31,45,31,197,31,76,31,21,31,191,31,106,31,106,30,165,31,186,31,213,31,87,31,87,30,199,31,199,30,184,31,10,31,243,31,243,30,243,29,29,31,78,31,129,31,129,30,129,29,92,31,176,31,86,31,121,31,214,31,203,31,136,31,111,31,53,31,255,31,111,31,158,31,44,31,112,31,212,31,175,31,175,30,93,31,93,30,212,31,126,31,162,31,52,31,137,31,76,31,178,31,178,30,52,31,52,30,215,31,215,30,136,31,183,31,93,31,219,31,171,31,179,31,78,31,129,31,65,31,75,31,75,30,174,31,174,30,189,31,205,31,177,31,177,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
