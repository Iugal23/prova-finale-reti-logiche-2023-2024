-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 956;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,160,0,0,0,50,0,133,0,102,0,0,0,125,0,158,0,26,0,80,0,0,0,61,0,133,0,243,0,102,0,77,0,220,0,21,0,176,0,186,0,77,0,86,0,101,0,183,0,97,0,143,0,250,0,33,0,0,0,12,0,81,0,23,0,183,0,194,0,183,0,0,0,152,0,233,0,139,0,243,0,0,0,0,0,164,0,63,0,152,0,0,0,101,0,46,0,142,0,0,0,0,0,189,0,0,0,0,0,144,0,244,0,134,0,204,0,235,0,220,0,153,0,234,0,157,0,30,0,0,0,220,0,137,0,68,0,246,0,195,0,139,0,240,0,243,0,0,0,211,0,13,0,25,0,79,0,209,0,121,0,172,0,59,0,205,0,91,0,211,0,35,0,127,0,97,0,97,0,157,0,22,0,231,0,230,0,229,0,9,0,0,0,128,0,53,0,166,0,0,0,217,0,0,0,0,0,0,0,71,0,117,0,0,0,39,0,204,0,46,0,0,0,95,0,0,0,197,0,0,0,151,0,61,0,142,0,44,0,164,0,55,0,59,0,32,0,215,0,93,0,91,0,93,0,0,0,207,0,22,0,198,0,77,0,123,0,79,0,69,0,55,0,202,0,81,0,0,0,231,0,17,0,185,0,0,0,181,0,180,0,233,0,143,0,139,0,0,0,122,0,0,0,0,0,0,0,103,0,33,0,0,0,166,0,97,0,0,0,0,0,67,0,0,0,0,0,84,0,0,0,0,0,49,0,213,0,13,0,0,0,151,0,133,0,0,0,150,0,0,0,0,0,191,0,0,0,148,0,212,0,128,0,152,0,0,0,132,0,219,0,89,0,16,0,237,0,0,0,94,0,0,0,6,0,95,0,249,0,173,0,47,0,118,0,242,0,25,0,226,0,29,0,169,0,122,0,0,0,222,0,0,0,212,0,23,0,0,0,77,0,140,0,199,0,56,0,80,0,172,0,10,0,0,0,170,0,147,0,0,0,156,0,123,0,176,0,58,0,0,0,82,0,223,0,56,0,221,0,112,0,179,0,210,0,184,0,98,0,0,0,237,0,119,0,99,0,254,0,165,0,0,0,203,0,228,0,120,0,141,0,0,0,0,0,221,0,27,0,101,0,0,0,38,0,218,0,0,0,47,0,32,0,35,0,136,0,42,0,241,0,214,0,0,0,176,0,208,0,176,0,108,0,153,0,2,0,6,0,0,0,142,0,152,0,105,0,0,0,199,0,199,0,0,0,211,0,74,0,0,0,39,0,188,0,0,0,16,0,224,0,127,0,249,0,140,0,133,0,59,0,240,0,155,0,150,0,241,0,16,0,254,0,101,0,42,0,68,0,143,0,59,0,196,0,6,0,0,0,42,0,129,0,44,0,49,0,0,0,233,0,83,0,229,0,0,0,235,0,31,0,210,0,187,0,76,0,124,0,91,0,228,0,6,0,0,0,23,0,91,0,184,0,0,0,121,0,0,0,203,0,3,0,0,0,239,0,0,0,147,0,185,0,0,0,43,0,17,0,0,0,231,0,197,0,14,0,198,0,145,0,0,0,148,0,0,0,224,0,58,0,146,0,126,0,75,0,154,0,34,0,218,0,189,0,104,0,0,0,93,0,0,0,81,0,0,0,130,0,10,0,156,0,14,0,144,0,0,0,122,0,250,0,229,0,163,0,165,0,85,0,39,0,0,0,12,0,0,0,16,0,181,0,0,0,167,0,0,0,63,0,140,0,159,0,63,0,232,0,0,0,233,0,34,0,202,0,180,0,228,0,4,0,33,0,41,0,130,0,164,0,177,0,0,0,241,0,245,0,43,0,192,0,30,0,196,0,142,0,127,0,87,0,208,0,56,0,51,0,11,0,205,0,240,0,251,0,254,0,192,0,103,0,5,0,202,0,144,0,212,0,0,0,154,0,3,0,221,0,0,0,141,0,46,0,209,0,147,0,250,0,111,0,46,0,173,0,103,0,196,0,61,0,0,0,16,0,38,0,205,0,158,0,81,0,38,0,0,0,124,0,14,0,199,0,53,0,53,0,0,0,164,0,0,0,0,0,85,0,224,0,93,0,78,0,101,0,196,0,0,0,0,0,96,0,58,0,0,0,21,0,42,0,199,0,158,0,157,0,197,0,0,0,0,0,0,0,112,0,199,0,188,0,24,0,252,0,0,0,241,0,185,0,158,0,159,0,0,0,151,0,0,0,0,0,134,0,28,0,63,0,67,0,159,0,231,0,200,0,45,0,13,0,0,0,0,0,67,0,69,0,0,0,128,0,83,0,199,0,122,0,0,0,0,0,159,0,223,0,0,0,90,0,127,0,182,0,0,0,128,0,105,0,162,0,134,0,7,0,21,0,0,0,253,0,0,0,60,0,165,0,74,0,0,0,189,0,112,0,120,0,13,0,0,0,208,0,124,0,249,0,35,0,165,0,28,0,151,0,99,0,120,0,0,0,90,0,247,0,219,0,48,0,149,0,0,0,0,0,75,0,0,0,171,0,0,0,0,0,47,0,182,0,0,0,243,0,75,0,138,0,247,0,9,0,189,0,43,0,255,0,0,0,137,0,0,0,0,0,18,0,0,0,206,0,232,0,14,0,41,0,174,0,122,0,104,0,151,0,247,0,110,0,32,0,120,0,155,0,0,0,146,0,251,0,197,0,0,0,182,0,0,0,14,0,58,0,94,0,88,0,207,0,220,0,187,0,190,0,199,0,60,0,0,0,147,0,1,0,72,0,0,0,162,0,125,0,50,0,0,0,69,0,165,0,191,0,244,0,0,0,160,0,214,0,0,0,13,0,250,0,205,0,36,0,227,0,154,0,100,0,77,0,39,0,0,0,105,0,2,0,109,0,75,0,151,0,160,0,35,0,0,0,77,0,0,0,0,0,0,0,90,0,0,0,55,0,209,0,235,0,153,0,198,0,13,0,241,0,232,0,0,0,82,0,0,0,93,0,0,0,178,0,211,0,195,0,0,0,0,0,0,0,218,0,130,0,73,0,173,0,200,0,146,0,225,0,83,0,124,0,67,0,174,0,119,0,248,0,19,0,127,0,14,0,205,0,39,0,234,0,151,0,118,0,250,0,84,0,5,0,251,0,157,0,104,0,229,0,48,0,0,0,57,0,206,0,0,0,200,0,126,0,64,0,0,0,31,0,197,0,0,0,223,0,226,0,113,0,81,0,0,0,66,0,62,0,153,0,0,0,248,0,189,0,0,0,60,0,201,0,219,0,0,0,255,0,59,0,74,0,187,0,70,0,53,0,0,0,200,0,204,0,158,0,193,0,114,0,0,0,0,0,192,0,163,0,53,0,130,0,237,0,41,0,140,0,0,0,178,0,0,0,248,0,243,0,73,0,0,0,139,0,35,0,0,0,148,0,248,0,149,0,172,0,100,0,105,0,101,0,83,0,242,0,200,0,99,0,203,0,111,0,210,0,138,0,0,0,0,0,0,0,93,0,195,0,100,0,82,0,93,0,103,0,185,0,174,0,24,0,117,0,36,0,91,0,140,0,236,0,75,0,26,0,174,0,0,0,21,0,211,0,0,0,164,0,136,0,45,0,0,0,0,0,0,0,123,0,198,0,0,0,90,0,0,0,0,0,230,0,203,0,192,0,189,0,70,0,192,0,4,0,245,0,198,0,12,0,202,0,102,0,7,0,152,0,187,0,123,0,247,0,0,0,237,0,193,0,86,0,182,0,61,0,248,0,0,0,23,0,156,0,93,0,159,0,243,0,0,0,16,0,60,0,0,0,180,0,212,0,83,0,104,0,89,0,0,0,144,0,10,0,4,0,86,0,191,0,224,0,207,0,0,0,0,0,0,0,157,0,196,0,168,0,193,0,0,0,79,0,0,0,60,0,0,0,103,0,228,0,222,0,72,0,34,0,46,0,0,0,182,0,14,0,18,0,240,0,232,0,59,0,184,0,0,0,19,0,146,0,167,0,209,0,115,0,67,0,63,0,148,0,90,0,68,0,0,0,63,0,42,0,239,0,92,0,0,0,209,0,30,0,198,0,240,0,141,0,180,0,213,0,178,0,83,0,55,0,240,0,0,0,146,0,0,0,0,0,73,0,224,0,220,0,101,0,141,0,149,0,214,0,85,0,225,0,201,0,160,0,0,0,0,0,0,0,0,0,235,0,121,0,250,0,247,0,181,0,254,0,0,0,38,0,6,0,111,0,160,0,237,0,218,0,0,0,242,0,222,0,124,0,149,0,171,0,24,0,73,0,61,0,0,0,122,0,36,0,0,0,147,0,148,0,154,0,241,0,0,0);
signal scenario_full  : scenario_type := (232,31,160,31,160,30,50,31,133,31,102,31,102,30,125,31,158,31,26,31,80,31,80,30,61,31,133,31,243,31,102,31,77,31,220,31,21,31,176,31,186,31,77,31,86,31,101,31,183,31,97,31,143,31,250,31,33,31,33,30,12,31,81,31,23,31,183,31,194,31,183,31,183,30,152,31,233,31,139,31,243,31,243,30,243,29,164,31,63,31,152,31,152,30,101,31,46,31,142,31,142,30,142,29,189,31,189,30,189,29,144,31,244,31,134,31,204,31,235,31,220,31,153,31,234,31,157,31,30,31,30,30,220,31,137,31,68,31,246,31,195,31,139,31,240,31,243,31,243,30,211,31,13,31,25,31,79,31,209,31,121,31,172,31,59,31,205,31,91,31,211,31,35,31,127,31,97,31,97,31,157,31,22,31,231,31,230,31,229,31,9,31,9,30,128,31,53,31,166,31,166,30,217,31,217,30,217,29,217,28,71,31,117,31,117,30,39,31,204,31,46,31,46,30,95,31,95,30,197,31,197,30,151,31,61,31,142,31,44,31,164,31,55,31,59,31,32,31,215,31,93,31,91,31,93,31,93,30,207,31,22,31,198,31,77,31,123,31,79,31,69,31,55,31,202,31,81,31,81,30,231,31,17,31,185,31,185,30,181,31,180,31,233,31,143,31,139,31,139,30,122,31,122,30,122,29,122,28,103,31,33,31,33,30,166,31,97,31,97,30,97,29,67,31,67,30,67,29,84,31,84,30,84,29,49,31,213,31,13,31,13,30,151,31,133,31,133,30,150,31,150,30,150,29,191,31,191,30,148,31,212,31,128,31,152,31,152,30,132,31,219,31,89,31,16,31,237,31,237,30,94,31,94,30,6,31,95,31,249,31,173,31,47,31,118,31,242,31,25,31,226,31,29,31,169,31,122,31,122,30,222,31,222,30,212,31,23,31,23,30,77,31,140,31,199,31,56,31,80,31,172,31,10,31,10,30,170,31,147,31,147,30,156,31,123,31,176,31,58,31,58,30,82,31,223,31,56,31,221,31,112,31,179,31,210,31,184,31,98,31,98,30,237,31,119,31,99,31,254,31,165,31,165,30,203,31,228,31,120,31,141,31,141,30,141,29,221,31,27,31,101,31,101,30,38,31,218,31,218,30,47,31,32,31,35,31,136,31,42,31,241,31,214,31,214,30,176,31,208,31,176,31,108,31,153,31,2,31,6,31,6,30,142,31,152,31,105,31,105,30,199,31,199,31,199,30,211,31,74,31,74,30,39,31,188,31,188,30,16,31,224,31,127,31,249,31,140,31,133,31,59,31,240,31,155,31,150,31,241,31,16,31,254,31,101,31,42,31,68,31,143,31,59,31,196,31,6,31,6,30,42,31,129,31,44,31,49,31,49,30,233,31,83,31,229,31,229,30,235,31,31,31,210,31,187,31,76,31,124,31,91,31,228,31,6,31,6,30,23,31,91,31,184,31,184,30,121,31,121,30,203,31,3,31,3,30,239,31,239,30,147,31,185,31,185,30,43,31,17,31,17,30,231,31,197,31,14,31,198,31,145,31,145,30,148,31,148,30,224,31,58,31,146,31,126,31,75,31,154,31,34,31,218,31,189,31,104,31,104,30,93,31,93,30,81,31,81,30,130,31,10,31,156,31,14,31,144,31,144,30,122,31,250,31,229,31,163,31,165,31,85,31,39,31,39,30,12,31,12,30,16,31,181,31,181,30,167,31,167,30,63,31,140,31,159,31,63,31,232,31,232,30,233,31,34,31,202,31,180,31,228,31,4,31,33,31,41,31,130,31,164,31,177,31,177,30,241,31,245,31,43,31,192,31,30,31,196,31,142,31,127,31,87,31,208,31,56,31,51,31,11,31,205,31,240,31,251,31,254,31,192,31,103,31,5,31,202,31,144,31,212,31,212,30,154,31,3,31,221,31,221,30,141,31,46,31,209,31,147,31,250,31,111,31,46,31,173,31,103,31,196,31,61,31,61,30,16,31,38,31,205,31,158,31,81,31,38,31,38,30,124,31,14,31,199,31,53,31,53,31,53,30,164,31,164,30,164,29,85,31,224,31,93,31,78,31,101,31,196,31,196,30,196,29,96,31,58,31,58,30,21,31,42,31,199,31,158,31,157,31,197,31,197,30,197,29,197,28,112,31,199,31,188,31,24,31,252,31,252,30,241,31,185,31,158,31,159,31,159,30,151,31,151,30,151,29,134,31,28,31,63,31,67,31,159,31,231,31,200,31,45,31,13,31,13,30,13,29,67,31,69,31,69,30,128,31,83,31,199,31,122,31,122,30,122,29,159,31,223,31,223,30,90,31,127,31,182,31,182,30,128,31,105,31,162,31,134,31,7,31,21,31,21,30,253,31,253,30,60,31,165,31,74,31,74,30,189,31,112,31,120,31,13,31,13,30,208,31,124,31,249,31,35,31,165,31,28,31,151,31,99,31,120,31,120,30,90,31,247,31,219,31,48,31,149,31,149,30,149,29,75,31,75,30,171,31,171,30,171,29,47,31,182,31,182,30,243,31,75,31,138,31,247,31,9,31,189,31,43,31,255,31,255,30,137,31,137,30,137,29,18,31,18,30,206,31,232,31,14,31,41,31,174,31,122,31,104,31,151,31,247,31,110,31,32,31,120,31,155,31,155,30,146,31,251,31,197,31,197,30,182,31,182,30,14,31,58,31,94,31,88,31,207,31,220,31,187,31,190,31,199,31,60,31,60,30,147,31,1,31,72,31,72,30,162,31,125,31,50,31,50,30,69,31,165,31,191,31,244,31,244,30,160,31,214,31,214,30,13,31,250,31,205,31,36,31,227,31,154,31,100,31,77,31,39,31,39,30,105,31,2,31,109,31,75,31,151,31,160,31,35,31,35,30,77,31,77,30,77,29,77,28,90,31,90,30,55,31,209,31,235,31,153,31,198,31,13,31,241,31,232,31,232,30,82,31,82,30,93,31,93,30,178,31,211,31,195,31,195,30,195,29,195,28,218,31,130,31,73,31,173,31,200,31,146,31,225,31,83,31,124,31,67,31,174,31,119,31,248,31,19,31,127,31,14,31,205,31,39,31,234,31,151,31,118,31,250,31,84,31,5,31,251,31,157,31,104,31,229,31,48,31,48,30,57,31,206,31,206,30,200,31,126,31,64,31,64,30,31,31,197,31,197,30,223,31,226,31,113,31,81,31,81,30,66,31,62,31,153,31,153,30,248,31,189,31,189,30,60,31,201,31,219,31,219,30,255,31,59,31,74,31,187,31,70,31,53,31,53,30,200,31,204,31,158,31,193,31,114,31,114,30,114,29,192,31,163,31,53,31,130,31,237,31,41,31,140,31,140,30,178,31,178,30,248,31,243,31,73,31,73,30,139,31,35,31,35,30,148,31,248,31,149,31,172,31,100,31,105,31,101,31,83,31,242,31,200,31,99,31,203,31,111,31,210,31,138,31,138,30,138,29,138,28,93,31,195,31,100,31,82,31,93,31,103,31,185,31,174,31,24,31,117,31,36,31,91,31,140,31,236,31,75,31,26,31,174,31,174,30,21,31,211,31,211,30,164,31,136,31,45,31,45,30,45,29,45,28,123,31,198,31,198,30,90,31,90,30,90,29,230,31,203,31,192,31,189,31,70,31,192,31,4,31,245,31,198,31,12,31,202,31,102,31,7,31,152,31,187,31,123,31,247,31,247,30,237,31,193,31,86,31,182,31,61,31,248,31,248,30,23,31,156,31,93,31,159,31,243,31,243,30,16,31,60,31,60,30,180,31,212,31,83,31,104,31,89,31,89,30,144,31,10,31,4,31,86,31,191,31,224,31,207,31,207,30,207,29,207,28,157,31,196,31,168,31,193,31,193,30,79,31,79,30,60,31,60,30,103,31,228,31,222,31,72,31,34,31,46,31,46,30,182,31,14,31,18,31,240,31,232,31,59,31,184,31,184,30,19,31,146,31,167,31,209,31,115,31,67,31,63,31,148,31,90,31,68,31,68,30,63,31,42,31,239,31,92,31,92,30,209,31,30,31,198,31,240,31,141,31,180,31,213,31,178,31,83,31,55,31,240,31,240,30,146,31,146,30,146,29,73,31,224,31,220,31,101,31,141,31,149,31,214,31,85,31,225,31,201,31,160,31,160,30,160,29,160,28,160,27,235,31,121,31,250,31,247,31,181,31,254,31,254,30,38,31,6,31,111,31,160,31,237,31,218,31,218,30,242,31,222,31,124,31,149,31,171,31,24,31,73,31,61,31,61,30,122,31,36,31,36,30,147,31,148,31,154,31,241,31,241,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
