-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 982;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,252,0,0,0,34,0,35,0,84,0,103,0,246,0,0,0,0,0,0,0,50,0,169,0,0,0,0,0,176,0,187,0,1,0,168,0,212,0,14,0,0,0,102,0,231,0,220,0,100,0,172,0,33,0,18,0,24,0,0,0,0,0,217,0,0,0,130,0,22,0,222,0,164,0,75,0,60,0,160,0,201,0,253,0,74,0,255,0,150,0,3,0,0,0,191,0,25,0,122,0,205,0,217,0,26,0,253,0,190,0,207,0,0,0,220,0,67,0,14,0,171,0,0,0,0,0,92,0,129,0,80,0,187,0,37,0,93,0,0,0,75,0,191,0,0,0,9,0,105,0,189,0,0,0,91,0,224,0,38,0,139,0,0,0,0,0,234,0,6,0,98,0,138,0,184,0,108,0,0,0,101,0,0,0,176,0,234,0,98,0,109,0,198,0,109,0,76,0,27,0,0,0,146,0,249,0,229,0,189,0,74,0,89,0,234,0,0,0,214,0,0,0,0,0,47,0,72,0,170,0,16,0,129,0,98,0,0,0,23,0,48,0,0,0,246,0,203,0,149,0,213,0,222,0,218,0,0,0,246,0,96,0,163,0,19,0,14,0,0,0,135,0,0,0,2,0,148,0,98,0,0,0,157,0,203,0,117,0,0,0,86,0,240,0,0,0,0,0,163,0,79,0,0,0,100,0,69,0,208,0,190,0,0,0,197,0,189,0,63,0,0,0,71,0,168,0,110,0,141,0,150,0,170,0,237,0,0,0,192,0,212,0,219,0,157,0,55,0,141,0,167,0,0,0,145,0,0,0,122,0,229,0,0,0,24,0,159,0,0,0,0,0,0,0,105,0,37,0,0,0,207,0,255,0,24,0,82,0,80,0,220,0,0,0,140,0,113,0,40,0,20,0,170,0,53,0,94,0,7,0,0,0,76,0,206,0,179,0,40,0,144,0,12,0,12,0,0,0,134,0,187,0,15,0,121,0,24,0,44,0,6,0,76,0,0,0,45,0,233,0,41,0,43,0,163,0,171,0,242,0,139,0,177,0,119,0,173,0,0,0,16,0,193,0,228,0,214,0,191,0,71,0,0,0,3,0,93,0,174,0,250,0,41,0,140,0,250,0,104,0,0,0,112,0,241,0,124,0,140,0,118,0,176,0,100,0,167,0,116,0,0,0,75,0,129,0,29,0,213,0,163,0,100,0,226,0,61,0,186,0,68,0,14,0,169,0,0,0,204,0,0,0,75,0,45,0,0,0,0,0,223,0,220,0,165,0,117,0,97,0,5,0,92,0,157,0,77,0,58,0,158,0,26,0,223,0,193,0,0,0,115,0,174,0,200,0,161,0,67,0,0,0,0,0,221,0,57,0,188,0,78,0,90,0,217,0,165,0,250,0,0,0,166,0,0,0,208,0,0,0,78,0,70,0,49,0,231,0,148,0,113,0,250,0,152,0,180,0,0,0,0,0,138,0,92,0,200,0,244,0,33,0,0,0,152,0,73,0,0,0,84,0,242,0,149,0,166,0,155,0,248,0,98,0,0,0,26,0,191,0,0,0,14,0,152,0,16,0,165,0,225,0,199,0,119,0,57,0,25,0,188,0,174,0,106,0,123,0,232,0,124,0,85,0,78,0,33,0,73,0,0,0,151,0,56,0,0,0,72,0,202,0,0,0,144,0,213,0,0,0,200,0,72,0,0,0,43,0,0,0,6,0,0,0,74,0,181,0,35,0,128,0,157,0,104,0,35,0,219,0,43,0,138,0,126,0,113,0,124,0,60,0,160,0,138,0,0,0,0,0,0,0,192,0,125,0,0,0,0,0,252,0,69,0,178,0,208,0,109,0,238,0,34,0,179,0,54,0,94,0,239,0,7,0,206,0,94,0,135,0,8,0,0,0,97,0,26,0,20,0,221,0,205,0,96,0,92,0,14,0,70,0,0,0,0,0,119,0,10,0,97,0,220,0,0,0,56,0,26,0,0,0,213,0,228,0,223,0,168,0,0,0,0,0,77,0,163,0,24,0,253,0,224,0,40,0,51,0,0,0,239,0,252,0,0,0,154,0,0,0,0,0,102,0,179,0,135,0,119,0,223,0,175,0,0,0,78,0,160,0,0,0,0,0,147,0,230,0,243,0,0,0,226,0,134,0,177,0,79,0,63,0,205,0,74,0,43,0,9,0,97,0,217,0,19,0,193,0,82,0,202,0,53,0,195,0,79,0,85,0,194,0,73,0,188,0,190,0,253,0,96,0,219,0,0,0,0,0,115,0,0,0,70,0,61,0,65,0,0,0,0,0,166,0,0,0,250,0,217,0,136,0,159,0,154,0,220,0,21,0,17,0,0,0,0,0,71,0,193,0,20,0,0,0,69,0,88,0,107,0,43,0,91,0,75,0,96,0,210,0,76,0,158,0,249,0,85,0,31,0,189,0,239,0,120,0,152,0,34,0,20,0,78,0,2,0,72,0,56,0,76,0,134,0,199,0,0,0,214,0,26,0,212,0,0,0,32,0,239,0,15,0,237,0,206,0,136,0,0,0,0,0,48,0,218,0,199,0,202,0,52,0,57,0,245,0,120,0,141,0,3,0,101,0,121,0,13,0,33,0,216,0,0,0,177,0,55,0,0,0,131,0,154,0,219,0,156,0,178,0,173,0,143,0,68,0,32,0,174,0,135,0,70,0,149,0,9,0,179,0,14,0,140,0,156,0,160,0,0,0,33,0,79,0,0,0,0,0,16,0,110,0,145,0,113,0,241,0,57,0,110,0,143,0,6,0,110,0,243,0,152,0,101,0,165,0,216,0,25,0,157,0,0,0,113,0,53,0,0,0,200,0,232,0,89,0,111,0,232,0,0,0,169,0,170,0,32,0,53,0,225,0,48,0,0,0,30,0,6,0,43,0,100,0,41,0,145,0,172,0,8,0,167,0,10,0,147,0,237,0,0,0,222,0,14,0,201,0,40,0,7,0,169,0,92,0,0,0,99,0,0,0,131,0,216,0,0,0,247,0,37,0,77,0,106,0,95,0,0,0,123,0,0,0,5,0,173,0,255,0,0,0,229,0,169,0,169,0,6,0,0,0,248,0,138,0,174,0,0,0,233,0,0,0,17,0,0,0,57,0,252,0,137,0,104,0,209,0,172,0,237,0,224,0,212,0,207,0,133,0,130,0,63,0,199,0,59,0,13,0,236,0,202,0,112,0,197,0,198,0,253,0,198,0,0,0,208,0,46,0,15,0,78,0,0,0,108,0,0,0,167,0,66,0,52,0,188,0,0,0,157,0,191,0,228,0,0,0,183,0,214,0,18,0,232,0,159,0,214,0,177,0,0,0,239,0,197,0,173,0,28,0,77,0,0,0,163,0,167,0,0,0,0,0,0,0,14,0,247,0,0,0,216,0,3,0,0,0,193,0,141,0,57,0,43,0,254,0,17,0,201,0,63,0,175,0,181,0,117,0,166,0,250,0,239,0,194,0,4,0,13,0,139,0,124,0,0,0,145,0,133,0,239,0,183,0,173,0,132,0,102,0,237,0,0,0,0,0,109,0,100,0,0,0,122,0,225,0,237,0,243,0,251,0,0,0,124,0,0,0,0,0,105,0,0,0,72,0,30,0,116,0,181,0,33,0,220,0,68,0,95,0,213,0,77,0,117,0,0,0,75,0,70,0,0,0,116,0,169,0,0,0,0,0,65,0,238,0,63,0,24,0,112,0,64,0,0,0,52,0,184,0,15,0,0,0,142,0,143,0,31,0,129,0,2,0,141,0,0,0,220,0,14,0,196,0,141,0,100,0,57,0,229,0,114,0,80,0,193,0,72,0,22,0,0,0,110,0,164,0,185,0,0,0,39,0,137,0,242,0,0,0,218,0,223,0,195,0,30,0,244,0,46,0,65,0,0,0,66,0,96,0,68,0,240,0,92,0,0,0,93,0,1,0,155,0,232,0,89,0,55,0,165,0,177,0,80,0,43,0,128,0,0,0,102,0,65,0,123,0,158,0,0,0,103,0,158,0,0,0,0,0,205,0,193,0,103,0,0,0,149,0,7,0,26,0,0,0,158,0,148,0,132,0,0,0,68,0,173,0,97,0,0,0,141,0,253,0,205,0,126,0,230,0,0,0,205,0,0,0,168,0,61,0,89,0,53,0,151,0,42,0,0,0,201,0,186,0,0,0,55,0,229,0,226,0,219,0,239,0,0,0,0,0,183,0,64,0,147,0,0,0,225,0,42,0,139,0,231,0,92,0,255,0,0,0,0,0,68,0,5,0,112,0,0,0,149,0,183,0,181,0,231,0,176,0,0,0,48,0,0,0,228,0,206,0,0,0,179,0,218,0,154,0,134,0,139,0,0,0,247,0,149,0,48,0,147,0,88,0,251,0,130,0,53,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,252,31,252,30,34,31,35,31,84,31,103,31,246,31,246,30,246,29,246,28,50,31,169,31,169,30,169,29,176,31,187,31,1,31,168,31,212,31,14,31,14,30,102,31,231,31,220,31,100,31,172,31,33,31,18,31,24,31,24,30,24,29,217,31,217,30,130,31,22,31,222,31,164,31,75,31,60,31,160,31,201,31,253,31,74,31,255,31,150,31,3,31,3,30,191,31,25,31,122,31,205,31,217,31,26,31,253,31,190,31,207,31,207,30,220,31,67,31,14,31,171,31,171,30,171,29,92,31,129,31,80,31,187,31,37,31,93,31,93,30,75,31,191,31,191,30,9,31,105,31,189,31,189,30,91,31,224,31,38,31,139,31,139,30,139,29,234,31,6,31,98,31,138,31,184,31,108,31,108,30,101,31,101,30,176,31,234,31,98,31,109,31,198,31,109,31,76,31,27,31,27,30,146,31,249,31,229,31,189,31,74,31,89,31,234,31,234,30,214,31,214,30,214,29,47,31,72,31,170,31,16,31,129,31,98,31,98,30,23,31,48,31,48,30,246,31,203,31,149,31,213,31,222,31,218,31,218,30,246,31,96,31,163,31,19,31,14,31,14,30,135,31,135,30,2,31,148,31,98,31,98,30,157,31,203,31,117,31,117,30,86,31,240,31,240,30,240,29,163,31,79,31,79,30,100,31,69,31,208,31,190,31,190,30,197,31,189,31,63,31,63,30,71,31,168,31,110,31,141,31,150,31,170,31,237,31,237,30,192,31,212,31,219,31,157,31,55,31,141,31,167,31,167,30,145,31,145,30,122,31,229,31,229,30,24,31,159,31,159,30,159,29,159,28,105,31,37,31,37,30,207,31,255,31,24,31,82,31,80,31,220,31,220,30,140,31,113,31,40,31,20,31,170,31,53,31,94,31,7,31,7,30,76,31,206,31,179,31,40,31,144,31,12,31,12,31,12,30,134,31,187,31,15,31,121,31,24,31,44,31,6,31,76,31,76,30,45,31,233,31,41,31,43,31,163,31,171,31,242,31,139,31,177,31,119,31,173,31,173,30,16,31,193,31,228,31,214,31,191,31,71,31,71,30,3,31,93,31,174,31,250,31,41,31,140,31,250,31,104,31,104,30,112,31,241,31,124,31,140,31,118,31,176,31,100,31,167,31,116,31,116,30,75,31,129,31,29,31,213,31,163,31,100,31,226,31,61,31,186,31,68,31,14,31,169,31,169,30,204,31,204,30,75,31,45,31,45,30,45,29,223,31,220,31,165,31,117,31,97,31,5,31,92,31,157,31,77,31,58,31,158,31,26,31,223,31,193,31,193,30,115,31,174,31,200,31,161,31,67,31,67,30,67,29,221,31,57,31,188,31,78,31,90,31,217,31,165,31,250,31,250,30,166,31,166,30,208,31,208,30,78,31,70,31,49,31,231,31,148,31,113,31,250,31,152,31,180,31,180,30,180,29,138,31,92,31,200,31,244,31,33,31,33,30,152,31,73,31,73,30,84,31,242,31,149,31,166,31,155,31,248,31,98,31,98,30,26,31,191,31,191,30,14,31,152,31,16,31,165,31,225,31,199,31,119,31,57,31,25,31,188,31,174,31,106,31,123,31,232,31,124,31,85,31,78,31,33,31,73,31,73,30,151,31,56,31,56,30,72,31,202,31,202,30,144,31,213,31,213,30,200,31,72,31,72,30,43,31,43,30,6,31,6,30,74,31,181,31,35,31,128,31,157,31,104,31,35,31,219,31,43,31,138,31,126,31,113,31,124,31,60,31,160,31,138,31,138,30,138,29,138,28,192,31,125,31,125,30,125,29,252,31,69,31,178,31,208,31,109,31,238,31,34,31,179,31,54,31,94,31,239,31,7,31,206,31,94,31,135,31,8,31,8,30,97,31,26,31,20,31,221,31,205,31,96,31,92,31,14,31,70,31,70,30,70,29,119,31,10,31,97,31,220,31,220,30,56,31,26,31,26,30,213,31,228,31,223,31,168,31,168,30,168,29,77,31,163,31,24,31,253,31,224,31,40,31,51,31,51,30,239,31,252,31,252,30,154,31,154,30,154,29,102,31,179,31,135,31,119,31,223,31,175,31,175,30,78,31,160,31,160,30,160,29,147,31,230,31,243,31,243,30,226,31,134,31,177,31,79,31,63,31,205,31,74,31,43,31,9,31,97,31,217,31,19,31,193,31,82,31,202,31,53,31,195,31,79,31,85,31,194,31,73,31,188,31,190,31,253,31,96,31,219,31,219,30,219,29,115,31,115,30,70,31,61,31,65,31,65,30,65,29,166,31,166,30,250,31,217,31,136,31,159,31,154,31,220,31,21,31,17,31,17,30,17,29,71,31,193,31,20,31,20,30,69,31,88,31,107,31,43,31,91,31,75,31,96,31,210,31,76,31,158,31,249,31,85,31,31,31,189,31,239,31,120,31,152,31,34,31,20,31,78,31,2,31,72,31,56,31,76,31,134,31,199,31,199,30,214,31,26,31,212,31,212,30,32,31,239,31,15,31,237,31,206,31,136,31,136,30,136,29,48,31,218,31,199,31,202,31,52,31,57,31,245,31,120,31,141,31,3,31,101,31,121,31,13,31,33,31,216,31,216,30,177,31,55,31,55,30,131,31,154,31,219,31,156,31,178,31,173,31,143,31,68,31,32,31,174,31,135,31,70,31,149,31,9,31,179,31,14,31,140,31,156,31,160,31,160,30,33,31,79,31,79,30,79,29,16,31,110,31,145,31,113,31,241,31,57,31,110,31,143,31,6,31,110,31,243,31,152,31,101,31,165,31,216,31,25,31,157,31,157,30,113,31,53,31,53,30,200,31,232,31,89,31,111,31,232,31,232,30,169,31,170,31,32,31,53,31,225,31,48,31,48,30,30,31,6,31,43,31,100,31,41,31,145,31,172,31,8,31,167,31,10,31,147,31,237,31,237,30,222,31,14,31,201,31,40,31,7,31,169,31,92,31,92,30,99,31,99,30,131,31,216,31,216,30,247,31,37,31,77,31,106,31,95,31,95,30,123,31,123,30,5,31,173,31,255,31,255,30,229,31,169,31,169,31,6,31,6,30,248,31,138,31,174,31,174,30,233,31,233,30,17,31,17,30,57,31,252,31,137,31,104,31,209,31,172,31,237,31,224,31,212,31,207,31,133,31,130,31,63,31,199,31,59,31,13,31,236,31,202,31,112,31,197,31,198,31,253,31,198,31,198,30,208,31,46,31,15,31,78,31,78,30,108,31,108,30,167,31,66,31,52,31,188,31,188,30,157,31,191,31,228,31,228,30,183,31,214,31,18,31,232,31,159,31,214,31,177,31,177,30,239,31,197,31,173,31,28,31,77,31,77,30,163,31,167,31,167,30,167,29,167,28,14,31,247,31,247,30,216,31,3,31,3,30,193,31,141,31,57,31,43,31,254,31,17,31,201,31,63,31,175,31,181,31,117,31,166,31,250,31,239,31,194,31,4,31,13,31,139,31,124,31,124,30,145,31,133,31,239,31,183,31,173,31,132,31,102,31,237,31,237,30,237,29,109,31,100,31,100,30,122,31,225,31,237,31,243,31,251,31,251,30,124,31,124,30,124,29,105,31,105,30,72,31,30,31,116,31,181,31,33,31,220,31,68,31,95,31,213,31,77,31,117,31,117,30,75,31,70,31,70,30,116,31,169,31,169,30,169,29,65,31,238,31,63,31,24,31,112,31,64,31,64,30,52,31,184,31,15,31,15,30,142,31,143,31,31,31,129,31,2,31,141,31,141,30,220,31,14,31,196,31,141,31,100,31,57,31,229,31,114,31,80,31,193,31,72,31,22,31,22,30,110,31,164,31,185,31,185,30,39,31,137,31,242,31,242,30,218,31,223,31,195,31,30,31,244,31,46,31,65,31,65,30,66,31,96,31,68,31,240,31,92,31,92,30,93,31,1,31,155,31,232,31,89,31,55,31,165,31,177,31,80,31,43,31,128,31,128,30,102,31,65,31,123,31,158,31,158,30,103,31,158,31,158,30,158,29,205,31,193,31,103,31,103,30,149,31,7,31,26,31,26,30,158,31,148,31,132,31,132,30,68,31,173,31,97,31,97,30,141,31,253,31,205,31,126,31,230,31,230,30,205,31,205,30,168,31,61,31,89,31,53,31,151,31,42,31,42,30,201,31,186,31,186,30,55,31,229,31,226,31,219,31,239,31,239,30,239,29,183,31,64,31,147,31,147,30,225,31,42,31,139,31,231,31,92,31,255,31,255,30,255,29,68,31,5,31,112,31,112,30,149,31,183,31,181,31,231,31,176,31,176,30,48,31,48,30,228,31,206,31,206,30,179,31,218,31,154,31,134,31,139,31,139,30,247,31,149,31,48,31,147,31,88,31,251,31,130,31,53,31,53,30,53,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
