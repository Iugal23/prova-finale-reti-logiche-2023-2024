-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 292;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,0,0,13,0,200,0,37,0,85,0,10,0,242,0,115,0,252,0,172,0,60,0,236,0,16,0,134,0,44,0,116,0,164,0,0,0,73,0,0,0,95,0,0,0,0,0,25,0,79,0,217,0,8,0,114,0,0,0,0,0,133,0,218,0,62,0,176,0,117,0,0,0,0,0,49,0,66,0,91,0,0,0,44,0,20,0,244,0,187,0,26,0,189,0,70,0,174,0,198,0,201,0,214,0,71,0,119,0,72,0,0,0,244,0,13,0,232,0,6,0,100,0,162,0,206,0,45,0,114,0,0,0,87,0,225,0,103,0,161,0,114,0,142,0,92,0,219,0,80,0,221,0,157,0,0,0,199,0,0,0,0,0,54,0,156,0,0,0,0,0,0,0,202,0,102,0,0,0,0,0,0,0,30,0,189,0,98,0,0,0,118,0,216,0,0,0,241,0,131,0,165,0,156,0,5,0,0,0,31,0,210,0,255,0,132,0,107,0,63,0,244,0,1,0,13,0,229,0,221,0,115,0,202,0,201,0,206,0,122,0,93,0,120,0,0,0,113,0,1,0,0,0,219,0,43,0,184,0,86,0,234,0,110,0,50,0,0,0,252,0,245,0,195,0,177,0,0,0,96,0,156,0,0,0,132,0,183,0,0,0,11,0,24,0,5,0,67,0,44,0,90,0,254,0,0,0,179,0,205,0,253,0,180,0,0,0,223,0,0,0,158,0,0,0,67,0,0,0,0,0,0,0,13,0,70,0,65,0,230,0,100,0,61,0,36,0,0,0,188,0,0,0,0,0,134,0,1,0,0,0,104,0,161,0,0,0,93,0,6,0,0,0,37,0,159,0,0,0,0,0,89,0,104,0,59,0,116,0,185,0,161,0,60,0,14,0,0,0,102,0,215,0,184,0,198,0,30,0,92,0,142,0,187,0,35,0,116,0,178,0,164,0,5,0,236,0,144,0,219,0,0,0,26,0,200,0,100,0,47,0,133,0,94,0,0,0,0,0,149,0,79,0,95,0,0,0,192,0,0,0,206,0,108,0,187,0,237,0,34,0,167,0,45,0,115,0,205,0,0,0,101,0,64,0,17,0,185,0,197,0,150,0,0,0,7,0,63,0,156,0,0,0,89,0,245,0,168,0,37,0,62,0,76,0,35,0,160,0,0,0,0,0,246,0,89,0,215,0,3,0,200,0,0,0,170,0,0,0,0,0,93,0,122,0,53,0,118,0,6,0,73,0,130,0,219,0,94,0,0,0,144,0,240,0,0,0,196,0,103,0,0,0,101,0,145,0,127,0,57,0,223,0);
signal scenario_full  : scenario_type := (128,31,128,30,13,31,200,31,37,31,85,31,10,31,242,31,115,31,252,31,172,31,60,31,236,31,16,31,134,31,44,31,116,31,164,31,164,30,73,31,73,30,95,31,95,30,95,29,25,31,79,31,217,31,8,31,114,31,114,30,114,29,133,31,218,31,62,31,176,31,117,31,117,30,117,29,49,31,66,31,91,31,91,30,44,31,20,31,244,31,187,31,26,31,189,31,70,31,174,31,198,31,201,31,214,31,71,31,119,31,72,31,72,30,244,31,13,31,232,31,6,31,100,31,162,31,206,31,45,31,114,31,114,30,87,31,225,31,103,31,161,31,114,31,142,31,92,31,219,31,80,31,221,31,157,31,157,30,199,31,199,30,199,29,54,31,156,31,156,30,156,29,156,28,202,31,102,31,102,30,102,29,102,28,30,31,189,31,98,31,98,30,118,31,216,31,216,30,241,31,131,31,165,31,156,31,5,31,5,30,31,31,210,31,255,31,132,31,107,31,63,31,244,31,1,31,13,31,229,31,221,31,115,31,202,31,201,31,206,31,122,31,93,31,120,31,120,30,113,31,1,31,1,30,219,31,43,31,184,31,86,31,234,31,110,31,50,31,50,30,252,31,245,31,195,31,177,31,177,30,96,31,156,31,156,30,132,31,183,31,183,30,11,31,24,31,5,31,67,31,44,31,90,31,254,31,254,30,179,31,205,31,253,31,180,31,180,30,223,31,223,30,158,31,158,30,67,31,67,30,67,29,67,28,13,31,70,31,65,31,230,31,100,31,61,31,36,31,36,30,188,31,188,30,188,29,134,31,1,31,1,30,104,31,161,31,161,30,93,31,6,31,6,30,37,31,159,31,159,30,159,29,89,31,104,31,59,31,116,31,185,31,161,31,60,31,14,31,14,30,102,31,215,31,184,31,198,31,30,31,92,31,142,31,187,31,35,31,116,31,178,31,164,31,5,31,236,31,144,31,219,31,219,30,26,31,200,31,100,31,47,31,133,31,94,31,94,30,94,29,149,31,79,31,95,31,95,30,192,31,192,30,206,31,108,31,187,31,237,31,34,31,167,31,45,31,115,31,205,31,205,30,101,31,64,31,17,31,185,31,197,31,150,31,150,30,7,31,63,31,156,31,156,30,89,31,245,31,168,31,37,31,62,31,76,31,35,31,160,31,160,30,160,29,246,31,89,31,215,31,3,31,200,31,200,30,170,31,170,30,170,29,93,31,122,31,53,31,118,31,6,31,73,31,130,31,219,31,94,31,94,30,144,31,240,31,240,30,196,31,103,31,103,30,101,31,145,31,127,31,57,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
