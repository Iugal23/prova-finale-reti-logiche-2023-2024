-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 305;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,168,0,0,0,92,0,58,0,172,0,110,0,13,0,158,0,0,0,198,0,170,0,0,0,127,0,82,0,0,0,214,0,0,0,120,0,114,0,225,0,0,0,0,0,0,0,49,0,181,0,72,0,11,0,81,0,179,0,29,0,0,0,0,0,242,0,144,0,195,0,36,0,196,0,83,0,0,0,175,0,82,0,0,0,0,0,244,0,211,0,102,0,247,0,121,0,61,0,174,0,50,0,144,0,18,0,0,0,58,0,122,0,0,0,176,0,0,0,55,0,0,0,17,0,0,0,0,0,173,0,192,0,17,0,77,0,2,0,235,0,91,0,161,0,138,0,193,0,88,0,136,0,89,0,119,0,205,0,125,0,191,0,171,0,243,0,80,0,98,0,40,0,62,0,149,0,238,0,0,0,0,0,12,0,105,0,250,0,209,0,0,0,255,0,0,0,26,0,176,0,254,0,199,0,116,0,39,0,0,0,107,0,42,0,37,0,181,0,0,0,231,0,0,0,133,0,136,0,208,0,3,0,119,0,21,0,58,0,131,0,229,0,138,0,0,0,148,0,248,0,200,0,0,0,0,0,0,0,0,0,228,0,125,0,23,0,72,0,0,0,104,0,150,0,0,0,172,0,44,0,0,0,78,0,0,0,237,0,137,0,66,0,73,0,85,0,211,0,119,0,208,0,30,0,0,0,114,0,0,0,0,0,0,0,89,0,42,0,0,0,0,0,109,0,50,0,46,0,0,0,187,0,166,0,34,0,171,0,130,0,0,0,0,0,0,0,162,0,0,0,0,0,160,0,0,0,2,0,237,0,176,0,0,0,27,0,232,0,0,0,133,0,213,0,217,0,85,0,199,0,156,0,108,0,38,0,235,0,181,0,220,0,157,0,185,0,117,0,67,0,0,0,140,0,66,0,133,0,0,0,168,0,14,0,68,0,222,0,159,0,78,0,0,0,109,0,23,0,0,0,16,0,0,0,24,0,207,0,5,0,217,0,117,0,251,0,122,0,199,0,36,0,0,0,28,0,47,0,0,0,0,0,164,0,0,0,0,0,218,0,157,0,135,0,0,0,24,0,45,0,0,0,238,0,0,0,0,0,0,0,0,0,97,0,106,0,111,0,89,0,103,0,19,0,121,0,0,0,92,0,68,0,81,0,143,0,113,0,159,0,133,0,0,0,214,0,0,0,169,0,0,0,187,0,128,0,200,0,24,0,121,0,134,0,129,0,8,0,0,0,150,0,15,0,0,0,154,0,0,0,22,0,116,0,170,0,178,0,104,0,0,0,0,0,80,0,0,0,153,0,78,0,158,0,206,0,12,0,130,0,188,0,0,0,0,0,3,0,182,0,147,0,36,0,225,0,153,0);
signal scenario_full  : scenario_type := (189,31,168,31,168,30,92,31,58,31,172,31,110,31,13,31,158,31,158,30,198,31,170,31,170,30,127,31,82,31,82,30,214,31,214,30,120,31,114,31,225,31,225,30,225,29,225,28,49,31,181,31,72,31,11,31,81,31,179,31,29,31,29,30,29,29,242,31,144,31,195,31,36,31,196,31,83,31,83,30,175,31,82,31,82,30,82,29,244,31,211,31,102,31,247,31,121,31,61,31,174,31,50,31,144,31,18,31,18,30,58,31,122,31,122,30,176,31,176,30,55,31,55,30,17,31,17,30,17,29,173,31,192,31,17,31,77,31,2,31,235,31,91,31,161,31,138,31,193,31,88,31,136,31,89,31,119,31,205,31,125,31,191,31,171,31,243,31,80,31,98,31,40,31,62,31,149,31,238,31,238,30,238,29,12,31,105,31,250,31,209,31,209,30,255,31,255,30,26,31,176,31,254,31,199,31,116,31,39,31,39,30,107,31,42,31,37,31,181,31,181,30,231,31,231,30,133,31,136,31,208,31,3,31,119,31,21,31,58,31,131,31,229,31,138,31,138,30,148,31,248,31,200,31,200,30,200,29,200,28,200,27,228,31,125,31,23,31,72,31,72,30,104,31,150,31,150,30,172,31,44,31,44,30,78,31,78,30,237,31,137,31,66,31,73,31,85,31,211,31,119,31,208,31,30,31,30,30,114,31,114,30,114,29,114,28,89,31,42,31,42,30,42,29,109,31,50,31,46,31,46,30,187,31,166,31,34,31,171,31,130,31,130,30,130,29,130,28,162,31,162,30,162,29,160,31,160,30,2,31,237,31,176,31,176,30,27,31,232,31,232,30,133,31,213,31,217,31,85,31,199,31,156,31,108,31,38,31,235,31,181,31,220,31,157,31,185,31,117,31,67,31,67,30,140,31,66,31,133,31,133,30,168,31,14,31,68,31,222,31,159,31,78,31,78,30,109,31,23,31,23,30,16,31,16,30,24,31,207,31,5,31,217,31,117,31,251,31,122,31,199,31,36,31,36,30,28,31,47,31,47,30,47,29,164,31,164,30,164,29,218,31,157,31,135,31,135,30,24,31,45,31,45,30,238,31,238,30,238,29,238,28,238,27,97,31,106,31,111,31,89,31,103,31,19,31,121,31,121,30,92,31,68,31,81,31,143,31,113,31,159,31,133,31,133,30,214,31,214,30,169,31,169,30,187,31,128,31,200,31,24,31,121,31,134,31,129,31,8,31,8,30,150,31,15,31,15,30,154,31,154,30,22,31,116,31,170,31,178,31,104,31,104,30,104,29,80,31,80,30,153,31,78,31,158,31,206,31,12,31,130,31,188,31,188,30,188,29,3,31,182,31,147,31,36,31,225,31,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
