-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 778;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,12,0,0,0,168,0,166,0,0,0,0,0,56,0,201,0,110,0,159,0,8,0,119,0,236,0,103,0,255,0,75,0,132,0,61,0,65,0,219,0,194,0,85,0,0,0,3,0,30,0,0,0,1,0,94,0,42,0,104,0,241,0,78,0,0,0,92,0,222,0,61,0,220,0,20,0,218,0,104,0,0,0,0,0,157,0,100,0,251,0,128,0,0,0,241,0,59,0,148,0,1,0,112,0,113,0,192,0,203,0,65,0,4,0,83,0,127,0,133,0,177,0,8,0,0,0,172,0,0,0,109,0,219,0,94,0,77,0,220,0,40,0,82,0,156,0,93,0,95,0,221,0,239,0,30,0,0,0,112,0,34,0,94,0,5,0,191,0,0,0,143,0,195,0,138,0,0,0,41,0,171,0,240,0,132,0,0,0,224,0,149,0,154,0,218,0,90,0,0,0,72,0,0,0,152,0,114,0,147,0,39,0,141,0,86,0,67,0,7,0,36,0,203,0,55,0,116,0,3,0,216,0,72,0,187,0,110,0,0,0,182,0,0,0,19,0,167,0,26,0,132,0,119,0,123,0,12,0,0,0,11,0,0,0,104,0,61,0,242,0,40,0,30,0,244,0,0,0,204,0,170,0,236,0,128,0,29,0,162,0,179,0,244,0,49,0,0,0,17,0,206,0,61,0,118,0,192,0,53,0,232,0,253,0,117,0,216,0,188,0,114,0,0,0,116,0,0,0,185,0,77,0,221,0,0,0,101,0,144,0,0,0,50,0,192,0,199,0,0,0,43,0,217,0,242,0,167,0,96,0,11,0,0,0,0,0,242,0,0,0,146,0,44,0,105,0,85,0,137,0,167,0,110,0,146,0,227,0,43,0,104,0,224,0,43,0,87,0,187,0,235,0,131,0,186,0,108,0,220,0,97,0,0,0,0,0,0,0,137,0,26,0,0,0,115,0,239,0,109,0,15,0,195,0,109,0,0,0,219,0,68,0,103,0,184,0,83,0,176,0,128,0,33,0,0,0,208,0,235,0,186,0,100,0,246,0,88,0,88,0,165,0,19,0,47,0,8,0,154,0,162,0,169,0,0,0,206,0,112,0,195,0,153,0,168,0,185,0,138,0,0,0,120,0,246,0,0,0,0,0,157,0,107,0,209,0,174,0,148,0,0,0,143,0,173,0,0,0,107,0,233,0,89,0,122,0,64,0,104,0,186,0,0,0,14,0,185,0,170,0,0,0,32,0,197,0,123,0,127,0,59,0,228,0,90,0,155,0,227,0,213,0,12,0,159,0,148,0,0,0,64,0,106,0,79,0,128,0,0,0,1,0,128,0,233,0,95,0,122,0,178,0,27,0,10,0,164,0,76,0,0,0,158,0,0,0,0,0,129,0,42,0,121,0,244,0,149,0,164,0,0,0,225,0,246,0,0,0,158,0,0,0,89,0,22,0,158,0,19,0,232,0,36,0,29,0,46,0,187,0,171,0,55,0,59,0,0,0,40,0,124,0,83,0,88,0,6,0,0,0,138,0,0,0,165,0,181,0,177,0,65,0,57,0,60,0,24,0,209,0,248,0,176,0,40,0,53,0,40,0,154,0,65,0,164,0,27,0,118,0,175,0,51,0,0,0,248,0,170,0,208,0,188,0,122,0,0,0,167,0,147,0,103,0,5,0,77,0,240,0,96,0,0,0,204,0,140,0,63,0,58,0,76,0,219,0,0,0,79,0,233,0,35,0,86,0,0,0,247,0,154,0,239,0,0,0,221,0,253,0,0,0,128,0,169,0,0,0,107,0,215,0,0,0,159,0,0,0,0,0,254,0,202,0,0,0,206,0,141,0,132,0,75,0,95,0,233,0,83,0,223,0,0,0,198,0,241,0,25,0,0,0,142,0,148,0,0,0,0,0,32,0,238,0,90,0,74,0,0,0,8,0,185,0,0,0,145,0,228,0,157,0,78,0,12,0,196,0,138,0,231,0,0,0,223,0,153,0,0,0,218,0,156,0,0,0,246,0,0,0,0,0,13,0,0,0,28,0,166,0,245,0,6,0,13,0,193,0,14,0,64,0,0,0,0,0,214,0,170,0,56,0,104,0,245,0,203,0,0,0,0,0,133,0,187,0,120,0,0,0,68,0,106,0,150,0,115,0,0,0,0,0,0,0,68,0,179,0,252,0,140,0,99,0,251,0,20,0,251,0,0,0,0,0,95,0,158,0,232,0,180,0,90,0,176,0,0,0,0,0,202,0,242,0,243,0,118,0,81,0,141,0,62,0,146,0,33,0,0,0,191,0,195,0,0,0,9,0,147,0,0,0,100,0,169,0,214,0,17,0,183,0,0,0,243,0,251,0,0,0,243,0,65,0,148,0,37,0,46,0,3,0,0,0,190,0,35,0,125,0,51,0,215,0,35,0,0,0,0,0,205,0,81,0,23,0,42,0,71,0,148,0,74,0,117,0,230,0,249,0,55,0,23,0,159,0,72,0,195,0,167,0,159,0,0,0,0,0,4,0,164,0,17,0,192,0,44,0,0,0,162,0,200,0,4,0,91,0,0,0,0,0,38,0,224,0,82,0,145,0,249,0,82,0,144,0,206,0,129,0,23,0,48,0,62,0,99,0,97,0,54,0,0,0,246,0,20,0,0,0,41,0,93,0,0,0,36,0,208,0,121,0,0,0,164,0,0,0,61,0,219,0,0,0,53,0,169,0,0,0,66,0,103,0,17,0,0,0,138,0,156,0,237,0,1,0,104,0,186,0,0,0,138,0,71,0,85,0,241,0,160,0,252,0,103,0,245,0,179,0,46,0,186,0,170,0,165,0,46,0,158,0,135,0,23,0,97,0,53,0,170,0,90,0,48,0,192,0,0,0,219,0,0,0,4,0,0,0,0,0,80,0,66,0,116,0,201,0,136,0,176,0,187,0,125,0,63,0,7,0,74,0,222,0,0,0,190,0,175,0,231,0,208,0,21,0,215,0,0,0,100,0,36,0,117,0,188,0,60,0,123,0,77,0,145,0,0,0,32,0,101,0,68,0,116,0,0,0,63,0,126,0,163,0,134,0,0,0,120,0,104,0,14,0,105,0,246,0,83,0,200,0,58,0,224,0,0,0,187,0,170,0,172,0,111,0,208,0,156,0,10,0,0,0,143,0,89,0,0,0,65,0,0,0,124,0,6,0,211,0,168,0,20,0,77,0,92,0,174,0,105,0,38,0,85,0,13,0,0,0,84,0,131,0,52,0,0,0,164,0,36,0,150,0,162,0,14,0,0,0,233,0,231,0,213,0,0,0,115,0,0,0,54,0,231,0,38,0,0,0,92,0,139,0,155,0,17,0,36,0,101,0,102,0,147,0,29,0,0,0,115,0,247,0,136,0,0,0,20,0,31,0,100,0,0,0,222,0,121,0,25,0,138,0,83,0,44,0,193,0,209,0,108,0,187,0,43,0,94,0,205,0,6,0,104,0,0,0,116,0,230,0,201,0);
signal scenario_full  : scenario_type := (136,31,12,31,12,30,168,31,166,31,166,30,166,29,56,31,201,31,110,31,159,31,8,31,119,31,236,31,103,31,255,31,75,31,132,31,61,31,65,31,219,31,194,31,85,31,85,30,3,31,30,31,30,30,1,31,94,31,42,31,104,31,241,31,78,31,78,30,92,31,222,31,61,31,220,31,20,31,218,31,104,31,104,30,104,29,157,31,100,31,251,31,128,31,128,30,241,31,59,31,148,31,1,31,112,31,113,31,192,31,203,31,65,31,4,31,83,31,127,31,133,31,177,31,8,31,8,30,172,31,172,30,109,31,219,31,94,31,77,31,220,31,40,31,82,31,156,31,93,31,95,31,221,31,239,31,30,31,30,30,112,31,34,31,94,31,5,31,191,31,191,30,143,31,195,31,138,31,138,30,41,31,171,31,240,31,132,31,132,30,224,31,149,31,154,31,218,31,90,31,90,30,72,31,72,30,152,31,114,31,147,31,39,31,141,31,86,31,67,31,7,31,36,31,203,31,55,31,116,31,3,31,216,31,72,31,187,31,110,31,110,30,182,31,182,30,19,31,167,31,26,31,132,31,119,31,123,31,12,31,12,30,11,31,11,30,104,31,61,31,242,31,40,31,30,31,244,31,244,30,204,31,170,31,236,31,128,31,29,31,162,31,179,31,244,31,49,31,49,30,17,31,206,31,61,31,118,31,192,31,53,31,232,31,253,31,117,31,216,31,188,31,114,31,114,30,116,31,116,30,185,31,77,31,221,31,221,30,101,31,144,31,144,30,50,31,192,31,199,31,199,30,43,31,217,31,242,31,167,31,96,31,11,31,11,30,11,29,242,31,242,30,146,31,44,31,105,31,85,31,137,31,167,31,110,31,146,31,227,31,43,31,104,31,224,31,43,31,87,31,187,31,235,31,131,31,186,31,108,31,220,31,97,31,97,30,97,29,97,28,137,31,26,31,26,30,115,31,239,31,109,31,15,31,195,31,109,31,109,30,219,31,68,31,103,31,184,31,83,31,176,31,128,31,33,31,33,30,208,31,235,31,186,31,100,31,246,31,88,31,88,31,165,31,19,31,47,31,8,31,154,31,162,31,169,31,169,30,206,31,112,31,195,31,153,31,168,31,185,31,138,31,138,30,120,31,246,31,246,30,246,29,157,31,107,31,209,31,174,31,148,31,148,30,143,31,173,31,173,30,107,31,233,31,89,31,122,31,64,31,104,31,186,31,186,30,14,31,185,31,170,31,170,30,32,31,197,31,123,31,127,31,59,31,228,31,90,31,155,31,227,31,213,31,12,31,159,31,148,31,148,30,64,31,106,31,79,31,128,31,128,30,1,31,128,31,233,31,95,31,122,31,178,31,27,31,10,31,164,31,76,31,76,30,158,31,158,30,158,29,129,31,42,31,121,31,244,31,149,31,164,31,164,30,225,31,246,31,246,30,158,31,158,30,89,31,22,31,158,31,19,31,232,31,36,31,29,31,46,31,187,31,171,31,55,31,59,31,59,30,40,31,124,31,83,31,88,31,6,31,6,30,138,31,138,30,165,31,181,31,177,31,65,31,57,31,60,31,24,31,209,31,248,31,176,31,40,31,53,31,40,31,154,31,65,31,164,31,27,31,118,31,175,31,51,31,51,30,248,31,170,31,208,31,188,31,122,31,122,30,167,31,147,31,103,31,5,31,77,31,240,31,96,31,96,30,204,31,140,31,63,31,58,31,76,31,219,31,219,30,79,31,233,31,35,31,86,31,86,30,247,31,154,31,239,31,239,30,221,31,253,31,253,30,128,31,169,31,169,30,107,31,215,31,215,30,159,31,159,30,159,29,254,31,202,31,202,30,206,31,141,31,132,31,75,31,95,31,233,31,83,31,223,31,223,30,198,31,241,31,25,31,25,30,142,31,148,31,148,30,148,29,32,31,238,31,90,31,74,31,74,30,8,31,185,31,185,30,145,31,228,31,157,31,78,31,12,31,196,31,138,31,231,31,231,30,223,31,153,31,153,30,218,31,156,31,156,30,246,31,246,30,246,29,13,31,13,30,28,31,166,31,245,31,6,31,13,31,193,31,14,31,64,31,64,30,64,29,214,31,170,31,56,31,104,31,245,31,203,31,203,30,203,29,133,31,187,31,120,31,120,30,68,31,106,31,150,31,115,31,115,30,115,29,115,28,68,31,179,31,252,31,140,31,99,31,251,31,20,31,251,31,251,30,251,29,95,31,158,31,232,31,180,31,90,31,176,31,176,30,176,29,202,31,242,31,243,31,118,31,81,31,141,31,62,31,146,31,33,31,33,30,191,31,195,31,195,30,9,31,147,31,147,30,100,31,169,31,214,31,17,31,183,31,183,30,243,31,251,31,251,30,243,31,65,31,148,31,37,31,46,31,3,31,3,30,190,31,35,31,125,31,51,31,215,31,35,31,35,30,35,29,205,31,81,31,23,31,42,31,71,31,148,31,74,31,117,31,230,31,249,31,55,31,23,31,159,31,72,31,195,31,167,31,159,31,159,30,159,29,4,31,164,31,17,31,192,31,44,31,44,30,162,31,200,31,4,31,91,31,91,30,91,29,38,31,224,31,82,31,145,31,249,31,82,31,144,31,206,31,129,31,23,31,48,31,62,31,99,31,97,31,54,31,54,30,246,31,20,31,20,30,41,31,93,31,93,30,36,31,208,31,121,31,121,30,164,31,164,30,61,31,219,31,219,30,53,31,169,31,169,30,66,31,103,31,17,31,17,30,138,31,156,31,237,31,1,31,104,31,186,31,186,30,138,31,71,31,85,31,241,31,160,31,252,31,103,31,245,31,179,31,46,31,186,31,170,31,165,31,46,31,158,31,135,31,23,31,97,31,53,31,170,31,90,31,48,31,192,31,192,30,219,31,219,30,4,31,4,30,4,29,80,31,66,31,116,31,201,31,136,31,176,31,187,31,125,31,63,31,7,31,74,31,222,31,222,30,190,31,175,31,231,31,208,31,21,31,215,31,215,30,100,31,36,31,117,31,188,31,60,31,123,31,77,31,145,31,145,30,32,31,101,31,68,31,116,31,116,30,63,31,126,31,163,31,134,31,134,30,120,31,104,31,14,31,105,31,246,31,83,31,200,31,58,31,224,31,224,30,187,31,170,31,172,31,111,31,208,31,156,31,10,31,10,30,143,31,89,31,89,30,65,31,65,30,124,31,6,31,211,31,168,31,20,31,77,31,92,31,174,31,105,31,38,31,85,31,13,31,13,30,84,31,131,31,52,31,52,30,164,31,36,31,150,31,162,31,14,31,14,30,233,31,231,31,213,31,213,30,115,31,115,30,54,31,231,31,38,31,38,30,92,31,139,31,155,31,17,31,36,31,101,31,102,31,147,31,29,31,29,30,115,31,247,31,136,31,136,30,20,31,31,31,100,31,100,30,222,31,121,31,25,31,138,31,83,31,44,31,193,31,209,31,108,31,187,31,43,31,94,31,205,31,6,31,104,31,104,30,116,31,230,31,201,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
