-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 707;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (8,0,249,0,0,0,0,0,53,0,172,0,0,0,187,0,234,0,0,0,221,0,250,0,0,0,192,0,0,0,72,0,0,0,34,0,190,0,79,0,247,0,147,0,130,0,0,0,37,0,0,0,37,0,0,0,0,0,3,0,98,0,0,0,0,0,128,0,110,0,199,0,0,0,0,0,64,0,0,0,0,0,0,0,0,0,29,0,192,0,81,0,202,0,40,0,200,0,237,0,142,0,75,0,160,0,85,0,0,0,214,0,234,0,87,0,158,0,93,0,78,0,47,0,176,0,179,0,3,0,198,0,0,0,117,0,168,0,162,0,120,0,234,0,60,0,0,0,44,0,83,0,219,0,0,0,220,0,186,0,0,0,240,0,0,0,174,0,129,0,230,0,153,0,142,0,169,0,0,0,185,0,235,0,203,0,231,0,17,0,37,0,153,0,177,0,207,0,195,0,122,0,218,0,0,0,82,0,7,0,0,0,93,0,0,0,254,0,156,0,6,0,25,0,125,0,197,0,0,0,0,0,70,0,18,0,0,0,140,0,0,0,112,0,116,0,180,0,54,0,0,0,54,0,239,0,156,0,169,0,177,0,102,0,243,0,91,0,248,0,0,0,0,0,0,0,132,0,183,0,0,0,0,0,75,0,186,0,6,0,57,0,253,0,156,0,126,0,64,0,77,0,59,0,70,0,170,0,0,0,0,0,70,0,67,0,95,0,31,0,53,0,165,0,41,0,149,0,98,0,158,0,68,0,248,0,0,0,96,0,2,0,10,0,155,0,223,0,93,0,32,0,154,0,121,0,98,0,138,0,26,0,207,0,237,0,119,0,0,0,0,0,193,0,0,0,161,0,163,0,211,0,72,0,170,0,0,0,0,0,6,0,0,0,169,0,5,0,0,0,215,0,115,0,210,0,73,0,147,0,67,0,177,0,20,0,7,0,28,0,0,0,145,0,245,0,118,0,46,0,0,0,247,0,101,0,232,0,0,0,18,0,247,0,229,0,35,0,100,0,75,0,131,0,91,0,33,0,167,0,110,0,124,0,198,0,141,0,133,0,186,0,175,0,255,0,126,0,154,0,4,0,12,0,33,0,131,0,159,0,165,0,97,0,115,0,55,0,93,0,30,0,79,0,15,0,104,0,228,0,194,0,111,0,40,0,103,0,85,0,88,0,18,0,0,0,0,0,54,0,93,0,37,0,194,0,0,0,54,0,58,0,247,0,196,0,0,0,0,0,238,0,141,0,244,0,139,0,191,0,69,0,207,0,201,0,0,0,165,0,231,0,0,0,191,0,82,0,24,0,15,0,86,0,87,0,25,0,252,0,113,0,36,0,105,0,38,0,52,0,215,0,0,0,0,0,189,0,72,0,205,0,100,0,148,0,146,0,87,0,62,0,7,0,254,0,9,0,0,0,167,0,240,0,218,0,0,0,168,0,193,0,0,0,108,0,218,0,236,0,0,0,0,0,123,0,50,0,48,0,8,0,71,0,110,0,47,0,78,0,203,0,89,0,188,0,0,0,43,0,0,0,36,0,254,0,102,0,151,0,215,0,165,0,204,0,146,0,131,0,90,0,181,0,140,0,200,0,112,0,211,0,70,0,163,0,114,0,44,0,0,0,6,0,59,0,196,0,67,0,143,0,27,0,48,0,28,0,255,0,202,0,224,0,237,0,0,0,118,0,174,0,83,0,89,0,0,0,56,0,213,0,0,0,222,0,110,0,91,0,59,0,179,0,224,0,110,0,108,0,45,0,0,0,71,0,100,0,83,0,0,0,0,0,194,0,110,0,81,0,174,0,254,0,156,0,230,0,182,0,66,0,141,0,0,0,251,0,0,0,75,0,235,0,63,0,46,0,0,0,186,0,238,0,0,0,248,0,0,0,249,0,62,0,226,0,170,0,130,0,0,0,247,0,77,0,156,0,0,0,233,0,230,0,0,0,0,0,0,0,47,0,104,0,166,0,117,0,227,0,0,0,179,0,67,0,127,0,13,0,0,0,70,0,0,0,0,0,80,0,142,0,0,0,3,0,223,0,84,0,229,0,0,0,94,0,199,0,15,0,39,0,42,0,77,0,217,0,0,0,45,0,8,0,94,0,0,0,227,0,17,0,88,0,103,0,4,0,149,0,205,0,0,0,214,0,141,0,255,0,129,0,248,0,0,0,59,0,0,0,189,0,0,0,31,0,47,0,91,0,87,0,132,0,173,0,0,0,214,0,97,0,160,0,0,0,73,0,168,0,216,0,209,0,67,0,18,0,120,0,232,0,0,0,91,0,228,0,46,0,42,0,241,0,73,0,183,0,208,0,40,0,127,0,76,0,149,0,176,0,73,0,122,0,0,0,112,0,253,0,0,0,220,0,183,0,108,0,0,0,246,0,205,0,152,0,0,0,95,0,71,0,225,0,109,0,55,0,229,0,33,0,0,0,0,0,0,0,0,0,0,0,105,0,0,0,69,0,73,0,218,0,30,0,247,0,135,0,193,0,0,0,211,0,56,0,41,0,0,0,124,0,124,0,249,0,38,0,101,0,124,0,237,0,208,0,141,0,212,0,18,0,111,0,0,0,98,0,160,0,240,0,0,0,0,0,81,0,24,0,254,0,186,0,14,0,0,0,202,0,4,0,21,0,181,0,0,0,10,0,98,0,199,0,166,0,246,0,158,0,147,0,0,0,90,0,243,0,4,0,0,0,78,0,158,0,176,0,197,0,163,0,66,0,5,0,150,0,0,0,0,0,0,0,199,0,0,0,148,0,210,0,0,0,115,0,0,0,57,0,39,0,228,0,165,0,118,0,61,0,156,0,159,0,140,0,227,0,5,0,14,0,33,0,131,0,240,0,0,0,238,0,166,0,238,0,48,0,29,0,0,0,144,0,70,0,0,0,109,0,0,0,0,0,0,0,13,0,0,0,0,0,0,0,0,0,118,0,0,0,231,0,240,0,139,0,79,0,191,0,0,0,177,0,0,0,44,0,30,0,91,0,250,0,248,0,0,0,0,0,235,0,181,0,216,0,110,0,179,0,125,0,49,0,27,0,136,0,252,0,175,0,28,0,80,0,181,0,126,0,0,0,249,0,189,0,107,0,0,0,79,0,143,0,163,0,0,0,86,0,35,0,0,0,45,0,173,0,199,0,241,0,236,0,191,0,0,0,174,0,106,0,52,0);
signal scenario_full  : scenario_type := (8,31,249,31,249,30,249,29,53,31,172,31,172,30,187,31,234,31,234,30,221,31,250,31,250,30,192,31,192,30,72,31,72,30,34,31,190,31,79,31,247,31,147,31,130,31,130,30,37,31,37,30,37,31,37,30,37,29,3,31,98,31,98,30,98,29,128,31,110,31,199,31,199,30,199,29,64,31,64,30,64,29,64,28,64,27,29,31,192,31,81,31,202,31,40,31,200,31,237,31,142,31,75,31,160,31,85,31,85,30,214,31,234,31,87,31,158,31,93,31,78,31,47,31,176,31,179,31,3,31,198,31,198,30,117,31,168,31,162,31,120,31,234,31,60,31,60,30,44,31,83,31,219,31,219,30,220,31,186,31,186,30,240,31,240,30,174,31,129,31,230,31,153,31,142,31,169,31,169,30,185,31,235,31,203,31,231,31,17,31,37,31,153,31,177,31,207,31,195,31,122,31,218,31,218,30,82,31,7,31,7,30,93,31,93,30,254,31,156,31,6,31,25,31,125,31,197,31,197,30,197,29,70,31,18,31,18,30,140,31,140,30,112,31,116,31,180,31,54,31,54,30,54,31,239,31,156,31,169,31,177,31,102,31,243,31,91,31,248,31,248,30,248,29,248,28,132,31,183,31,183,30,183,29,75,31,186,31,6,31,57,31,253,31,156,31,126,31,64,31,77,31,59,31,70,31,170,31,170,30,170,29,70,31,67,31,95,31,31,31,53,31,165,31,41,31,149,31,98,31,158,31,68,31,248,31,248,30,96,31,2,31,10,31,155,31,223,31,93,31,32,31,154,31,121,31,98,31,138,31,26,31,207,31,237,31,119,31,119,30,119,29,193,31,193,30,161,31,163,31,211,31,72,31,170,31,170,30,170,29,6,31,6,30,169,31,5,31,5,30,215,31,115,31,210,31,73,31,147,31,67,31,177,31,20,31,7,31,28,31,28,30,145,31,245,31,118,31,46,31,46,30,247,31,101,31,232,31,232,30,18,31,247,31,229,31,35,31,100,31,75,31,131,31,91,31,33,31,167,31,110,31,124,31,198,31,141,31,133,31,186,31,175,31,255,31,126,31,154,31,4,31,12,31,33,31,131,31,159,31,165,31,97,31,115,31,55,31,93,31,30,31,79,31,15,31,104,31,228,31,194,31,111,31,40,31,103,31,85,31,88,31,18,31,18,30,18,29,54,31,93,31,37,31,194,31,194,30,54,31,58,31,247,31,196,31,196,30,196,29,238,31,141,31,244,31,139,31,191,31,69,31,207,31,201,31,201,30,165,31,231,31,231,30,191,31,82,31,24,31,15,31,86,31,87,31,25,31,252,31,113,31,36,31,105,31,38,31,52,31,215,31,215,30,215,29,189,31,72,31,205,31,100,31,148,31,146,31,87,31,62,31,7,31,254,31,9,31,9,30,167,31,240,31,218,31,218,30,168,31,193,31,193,30,108,31,218,31,236,31,236,30,236,29,123,31,50,31,48,31,8,31,71,31,110,31,47,31,78,31,203,31,89,31,188,31,188,30,43,31,43,30,36,31,254,31,102,31,151,31,215,31,165,31,204,31,146,31,131,31,90,31,181,31,140,31,200,31,112,31,211,31,70,31,163,31,114,31,44,31,44,30,6,31,59,31,196,31,67,31,143,31,27,31,48,31,28,31,255,31,202,31,224,31,237,31,237,30,118,31,174,31,83,31,89,31,89,30,56,31,213,31,213,30,222,31,110,31,91,31,59,31,179,31,224,31,110,31,108,31,45,31,45,30,71,31,100,31,83,31,83,30,83,29,194,31,110,31,81,31,174,31,254,31,156,31,230,31,182,31,66,31,141,31,141,30,251,31,251,30,75,31,235,31,63,31,46,31,46,30,186,31,238,31,238,30,248,31,248,30,249,31,62,31,226,31,170,31,130,31,130,30,247,31,77,31,156,31,156,30,233,31,230,31,230,30,230,29,230,28,47,31,104,31,166,31,117,31,227,31,227,30,179,31,67,31,127,31,13,31,13,30,70,31,70,30,70,29,80,31,142,31,142,30,3,31,223,31,84,31,229,31,229,30,94,31,199,31,15,31,39,31,42,31,77,31,217,31,217,30,45,31,8,31,94,31,94,30,227,31,17,31,88,31,103,31,4,31,149,31,205,31,205,30,214,31,141,31,255,31,129,31,248,31,248,30,59,31,59,30,189,31,189,30,31,31,47,31,91,31,87,31,132,31,173,31,173,30,214,31,97,31,160,31,160,30,73,31,168,31,216,31,209,31,67,31,18,31,120,31,232,31,232,30,91,31,228,31,46,31,42,31,241,31,73,31,183,31,208,31,40,31,127,31,76,31,149,31,176,31,73,31,122,31,122,30,112,31,253,31,253,30,220,31,183,31,108,31,108,30,246,31,205,31,152,31,152,30,95,31,71,31,225,31,109,31,55,31,229,31,33,31,33,30,33,29,33,28,33,27,33,26,105,31,105,30,69,31,73,31,218,31,30,31,247,31,135,31,193,31,193,30,211,31,56,31,41,31,41,30,124,31,124,31,249,31,38,31,101,31,124,31,237,31,208,31,141,31,212,31,18,31,111,31,111,30,98,31,160,31,240,31,240,30,240,29,81,31,24,31,254,31,186,31,14,31,14,30,202,31,4,31,21,31,181,31,181,30,10,31,98,31,199,31,166,31,246,31,158,31,147,31,147,30,90,31,243,31,4,31,4,30,78,31,158,31,176,31,197,31,163,31,66,31,5,31,150,31,150,30,150,29,150,28,199,31,199,30,148,31,210,31,210,30,115,31,115,30,57,31,39,31,228,31,165,31,118,31,61,31,156,31,159,31,140,31,227,31,5,31,14,31,33,31,131,31,240,31,240,30,238,31,166,31,238,31,48,31,29,31,29,30,144,31,70,31,70,30,109,31,109,30,109,29,109,28,13,31,13,30,13,29,13,28,13,27,118,31,118,30,231,31,240,31,139,31,79,31,191,31,191,30,177,31,177,30,44,31,30,31,91,31,250,31,248,31,248,30,248,29,235,31,181,31,216,31,110,31,179,31,125,31,49,31,27,31,136,31,252,31,175,31,28,31,80,31,181,31,126,31,126,30,249,31,189,31,107,31,107,30,79,31,143,31,163,31,163,30,86,31,35,31,35,30,45,31,173,31,199,31,241,31,236,31,191,31,191,30,174,31,106,31,52,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
