-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_111 is
end project_tb_111;

architecture project_tb_arch_111 of project_tb_111 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 664;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (217,0,0,0,0,0,47,0,169,0,116,0,113,0,185,0,0,0,219,0,3,0,0,0,1,0,185,0,254,0,191,0,100,0,22,0,105,0,165,0,136,0,96,0,0,0,0,0,242,0,0,0,0,0,0,0,238,0,0,0,173,0,11,0,226,0,167,0,192,0,134,0,42,0,92,0,219,0,0,0,154,0,97,0,136,0,56,0,154,0,230,0,160,0,86,0,29,0,179,0,85,0,153,0,58,0,56,0,163,0,0,0,223,0,91,0,198,0,159,0,85,0,0,0,49,0,255,0,165,0,73,0,0,0,0,0,2,0,124,0,0,0,0,0,0,0,116,0,48,0,93,0,0,0,211,0,130,0,118,0,0,0,0,0,209,0,228,0,248,0,178,0,223,0,20,0,5,0,34,0,151,0,189,0,162,0,145,0,239,0,0,0,26,0,229,0,3,0,82,0,40,0,249,0,193,0,0,0,103,0,221,0,38,0,46,0,234,0,157,0,241,0,92,0,0,0,94,0,0,0,210,0,0,0,59,0,187,0,17,0,214,0,187,0,197,0,150,0,161,0,63,0,0,0,0,0,197,0,0,0,138,0,0,0,0,0,0,0,139,0,192,0,175,0,60,0,61,0,0,0,136,0,172,0,0,0,167,0,59,0,147,0,0,0,0,0,43,0,161,0,49,0,206,0,171,0,158,0,72,0,3,0,159,0,200,0,207,0,144,0,0,0,0,0,64,0,170,0,60,0,144,0,0,0,184,0,0,0,18,0,0,0,219,0,166,0,244,0,0,0,219,0,0,0,0,0,222,0,86,0,192,0,39,0,183,0,237,0,25,0,118,0,0,0,53,0,199,0,249,0,219,0,195,0,137,0,185,0,147,0,228,0,66,0,52,0,195,0,24,0,140,0,106,0,0,0,59,0,35,0,34,0,146,0,0,0,182,0,0,0,207,0,30,0,176,0,178,0,41,0,0,0,103,0,179,0,128,0,47,0,189,0,8,0,203,0,170,0,0,0,165,0,24,0,98,0,0,0,102,0,149,0,209,0,92,0,196,0,157,0,125,0,4,0,191,0,85,0,250,0,10,0,66,0,0,0,225,0,26,0,0,0,159,0,0,0,233,0,189,0,73,0,0,0,216,0,56,0,163,0,197,0,234,0,237,0,85,0,174,0,0,0,105,0,72,0,72,0,96,0,19,0,119,0,192,0,84,0,141,0,223,0,218,0,167,0,85,0,152,0,103,0,239,0,0,0,0,0,44,0,160,0,39,0,178,0,55,0,178,0,21,0,32,0,0,0,0,0,168,0,220,0,76,0,185,0,89,0,136,0,211,0,0,0,195,0,67,0,189,0,245,0,0,0,0,0,86,0,0,0,248,0,246,0,60,0,0,0,183,0,0,0,0,0,177,0,26,0,199,0,67,0,50,0,219,0,174,0,114,0,133,0,59,0,142,0,68,0,7,0,89,0,52,0,107,0,0,0,0,0,179,0,170,0,128,0,61,0,195,0,155,0,196,0,2,0,112,0,0,0,161,0,89,0,90,0,193,0,0,0,30,0,130,0,104,0,180,0,102,0,35,0,255,0,144,0,221,0,174,0,136,0,90,0,200,0,176,0,211,0,84,0,19,0,215,0,245,0,222,0,224,0,40,0,174,0,106,0,195,0,0,0,53,0,13,0,155,0,158,0,68,0,189,0,204,0,0,0,189,0,184,0,0,0,227,0,131,0,243,0,130,0,1,0,38,0,0,0,83,0,113,0,28,0,212,0,170,0,147,0,125,0,0,0,208,0,146,0,214,0,43,0,248,0,0,0,182,0,0,0,0,0,117,0,209,0,234,0,57,0,221,0,0,0,231,0,245,0,146,0,0,0,0,0,5,0,121,0,61,0,148,0,147,0,154,0,2,0,225,0,153,0,0,0,26,0,40,0,141,0,190,0,25,0,33,0,9,0,215,0,0,0,249,0,89,0,88,0,246,0,70,0,72,0,225,0,181,0,200,0,0,0,14,0,0,0,78,0,47,0,94,0,209,0,59,0,185,0,12,0,63,0,218,0,78,0,253,0,39,0,103,0,191,0,0,0,0,0,0,0,0,0,108,0,15,0,128,0,81,0,113,0,80,0,26,0,37,0,184,0,0,0,96,0,0,0,221,0,78,0,107,0,48,0,0,0,0,0,0,0,0,0,24,0,165,0,219,0,203,0,0,0,26,0,0,0,0,0,228,0,145,0,175,0,0,0,94,0,244,0,148,0,184,0,144,0,72,0,255,0,59,0,0,0,0,0,0,0,235,0,0,0,234,0,3,0,0,0,64,0,252,0,0,0,63,0,216,0,143,0,0,0,240,0,88,0,181,0,198,0,134,0,69,0,185,0,186,0,192,0,143,0,0,0,255,0,76,0,0,0,24,0,60,0,208,0,96,0,0,0,63,0,199,0,188,0,0,0,143,0,242,0,124,0,224,0,49,0,12,0,0,0,195,0,226,0,0,0,0,0,117,0,157,0,248,0,44,0,252,0,0,0,0,0,195,0,63,0,72,0,29,0,48,0,135,0,0,0,0,0,111,0,140,0,122,0,0,0,80,0,70,0,249,0,232,0,0,0,219,0,0,0,183,0,29,0,217,0,132,0,180,0,193,0,0,0,248,0,168,0,28,0,13,0,11,0,113,0,111,0,0,0,131,0,13,0,17,0,0,0,65,0,91,0,227,0,117,0,181,0,39,0,2,0,246,0,73,0,28,0,109,0,148,0,0,0,61,0,0,0,35,0,15,0,13,0,0,0,82,0,193,0,78,0,49,0,150,0,61,0,0,0,0,0,143,0,229,0,29,0,0,0,0,0,13,0,0,0,253,0,122,0,29,0,210,0,21,0,156,0,170,0,216,0,69,0,133,0,9,0,0,0,228,0,49,0,25,0,0,0,172,0,4,0,163,0,15,0,102,0,108,0,0,0,0,0,209,0,134,0,3,0,228,0,0,0,134,0);
signal scenario_full  : scenario_type := (217,31,217,30,217,29,47,31,169,31,116,31,113,31,185,31,185,30,219,31,3,31,3,30,1,31,185,31,254,31,191,31,100,31,22,31,105,31,165,31,136,31,96,31,96,30,96,29,242,31,242,30,242,29,242,28,238,31,238,30,173,31,11,31,226,31,167,31,192,31,134,31,42,31,92,31,219,31,219,30,154,31,97,31,136,31,56,31,154,31,230,31,160,31,86,31,29,31,179,31,85,31,153,31,58,31,56,31,163,31,163,30,223,31,91,31,198,31,159,31,85,31,85,30,49,31,255,31,165,31,73,31,73,30,73,29,2,31,124,31,124,30,124,29,124,28,116,31,48,31,93,31,93,30,211,31,130,31,118,31,118,30,118,29,209,31,228,31,248,31,178,31,223,31,20,31,5,31,34,31,151,31,189,31,162,31,145,31,239,31,239,30,26,31,229,31,3,31,82,31,40,31,249,31,193,31,193,30,103,31,221,31,38,31,46,31,234,31,157,31,241,31,92,31,92,30,94,31,94,30,210,31,210,30,59,31,187,31,17,31,214,31,187,31,197,31,150,31,161,31,63,31,63,30,63,29,197,31,197,30,138,31,138,30,138,29,138,28,139,31,192,31,175,31,60,31,61,31,61,30,136,31,172,31,172,30,167,31,59,31,147,31,147,30,147,29,43,31,161,31,49,31,206,31,171,31,158,31,72,31,3,31,159,31,200,31,207,31,144,31,144,30,144,29,64,31,170,31,60,31,144,31,144,30,184,31,184,30,18,31,18,30,219,31,166,31,244,31,244,30,219,31,219,30,219,29,222,31,86,31,192,31,39,31,183,31,237,31,25,31,118,31,118,30,53,31,199,31,249,31,219,31,195,31,137,31,185,31,147,31,228,31,66,31,52,31,195,31,24,31,140,31,106,31,106,30,59,31,35,31,34,31,146,31,146,30,182,31,182,30,207,31,30,31,176,31,178,31,41,31,41,30,103,31,179,31,128,31,47,31,189,31,8,31,203,31,170,31,170,30,165,31,24,31,98,31,98,30,102,31,149,31,209,31,92,31,196,31,157,31,125,31,4,31,191,31,85,31,250,31,10,31,66,31,66,30,225,31,26,31,26,30,159,31,159,30,233,31,189,31,73,31,73,30,216,31,56,31,163,31,197,31,234,31,237,31,85,31,174,31,174,30,105,31,72,31,72,31,96,31,19,31,119,31,192,31,84,31,141,31,223,31,218,31,167,31,85,31,152,31,103,31,239,31,239,30,239,29,44,31,160,31,39,31,178,31,55,31,178,31,21,31,32,31,32,30,32,29,168,31,220,31,76,31,185,31,89,31,136,31,211,31,211,30,195,31,67,31,189,31,245,31,245,30,245,29,86,31,86,30,248,31,246,31,60,31,60,30,183,31,183,30,183,29,177,31,26,31,199,31,67,31,50,31,219,31,174,31,114,31,133,31,59,31,142,31,68,31,7,31,89,31,52,31,107,31,107,30,107,29,179,31,170,31,128,31,61,31,195,31,155,31,196,31,2,31,112,31,112,30,161,31,89,31,90,31,193,31,193,30,30,31,130,31,104,31,180,31,102,31,35,31,255,31,144,31,221,31,174,31,136,31,90,31,200,31,176,31,211,31,84,31,19,31,215,31,245,31,222,31,224,31,40,31,174,31,106,31,195,31,195,30,53,31,13,31,155,31,158,31,68,31,189,31,204,31,204,30,189,31,184,31,184,30,227,31,131,31,243,31,130,31,1,31,38,31,38,30,83,31,113,31,28,31,212,31,170,31,147,31,125,31,125,30,208,31,146,31,214,31,43,31,248,31,248,30,182,31,182,30,182,29,117,31,209,31,234,31,57,31,221,31,221,30,231,31,245,31,146,31,146,30,146,29,5,31,121,31,61,31,148,31,147,31,154,31,2,31,225,31,153,31,153,30,26,31,40,31,141,31,190,31,25,31,33,31,9,31,215,31,215,30,249,31,89,31,88,31,246,31,70,31,72,31,225,31,181,31,200,31,200,30,14,31,14,30,78,31,47,31,94,31,209,31,59,31,185,31,12,31,63,31,218,31,78,31,253,31,39,31,103,31,191,31,191,30,191,29,191,28,191,27,108,31,15,31,128,31,81,31,113,31,80,31,26,31,37,31,184,31,184,30,96,31,96,30,221,31,78,31,107,31,48,31,48,30,48,29,48,28,48,27,24,31,165,31,219,31,203,31,203,30,26,31,26,30,26,29,228,31,145,31,175,31,175,30,94,31,244,31,148,31,184,31,144,31,72,31,255,31,59,31,59,30,59,29,59,28,235,31,235,30,234,31,3,31,3,30,64,31,252,31,252,30,63,31,216,31,143,31,143,30,240,31,88,31,181,31,198,31,134,31,69,31,185,31,186,31,192,31,143,31,143,30,255,31,76,31,76,30,24,31,60,31,208,31,96,31,96,30,63,31,199,31,188,31,188,30,143,31,242,31,124,31,224,31,49,31,12,31,12,30,195,31,226,31,226,30,226,29,117,31,157,31,248,31,44,31,252,31,252,30,252,29,195,31,63,31,72,31,29,31,48,31,135,31,135,30,135,29,111,31,140,31,122,31,122,30,80,31,70,31,249,31,232,31,232,30,219,31,219,30,183,31,29,31,217,31,132,31,180,31,193,31,193,30,248,31,168,31,28,31,13,31,11,31,113,31,111,31,111,30,131,31,13,31,17,31,17,30,65,31,91,31,227,31,117,31,181,31,39,31,2,31,246,31,73,31,28,31,109,31,148,31,148,30,61,31,61,30,35,31,15,31,13,31,13,30,82,31,193,31,78,31,49,31,150,31,61,31,61,30,61,29,143,31,229,31,29,31,29,30,29,29,13,31,13,30,253,31,122,31,29,31,210,31,21,31,156,31,170,31,216,31,69,31,133,31,9,31,9,30,228,31,49,31,25,31,25,30,172,31,4,31,163,31,15,31,102,31,108,31,108,30,108,29,209,31,134,31,3,31,228,31,228,30,134,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
