-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 779;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,104,0,251,0,0,0,240,0,0,0,242,0,56,0,48,0,170,0,175,0,181,0,195,0,36,0,211,0,159,0,218,0,147,0,0,0,0,0,0,0,131,0,147,0,189,0,0,0,232,0,178,0,41,0,34,0,32,0,116,0,0,0,203,0,84,0,0,0,0,0,122,0,97,0,47,0,0,0,0,0,0,0,25,0,224,0,204,0,0,0,151,0,90,0,225,0,187,0,90,0,33,0,163,0,16,0,95,0,246,0,20,0,0,0,139,0,174,0,133,0,154,0,0,0,240,0,247,0,0,0,130,0,187,0,173,0,0,0,130,0,0,0,125,0,8,0,241,0,185,0,210,0,5,0,150,0,201,0,164,0,41,0,139,0,95,0,102,0,136,0,0,0,1,0,132,0,183,0,0,0,52,0,250,0,254,0,3,0,0,0,73,0,0,0,251,0,157,0,143,0,234,0,124,0,164,0,5,0,206,0,154,0,43,0,121,0,80,0,176,0,134,0,78,0,181,0,148,0,248,0,172,0,136,0,215,0,7,0,134,0,113,0,15,0,70,0,211,0,150,0,57,0,65,0,0,0,0,0,0,0,0,0,34,0,0,0,34,0,154,0,57,0,156,0,85,0,18,0,100,0,199,0,116,0,186,0,160,0,57,0,129,0,104,0,75,0,120,0,0,0,0,0,168,0,209,0,0,0,168,0,161,0,242,0,179,0,48,0,222,0,224,0,252,0,0,0,228,0,66,0,177,0,253,0,0,0,89,0,89,0,0,0,79,0,9,0,94,0,0,0,44,0,36,0,173,0,114,0,113,0,0,0,74,0,0,0,174,0,125,0,45,0,141,0,98,0,21,0,135,0,37,0,0,0,138,0,209,0,33,0,47,0,182,0,177,0,154,0,97,0,69,0,125,0,0,0,0,0,253,0,2,0,58,0,4,0,17,0,52,0,12,0,238,0,0,0,24,0,235,0,123,0,148,0,162,0,0,0,114,0,0,0,0,0,122,0,85,0,100,0,13,0,139,0,245,0,175,0,253,0,200,0,250,0,47,0,8,0,37,0,223,0,133,0,42,0,0,0,203,0,156,0,174,0,127,0,249,0,20,0,237,0,0,0,22,0,239,0,22,0,8,0,1,0,0,0,165,0,20,0,0,0,0,0,166,0,0,0,0,0,82,0,229,0,201,0,0,0,184,0,0,0,20,0,81,0,32,0,0,0,202,0,219,0,196,0,12,0,112,0,81,0,226,0,0,0,68,0,172,0,120,0,149,0,0,0,57,0,134,0,108,0,0,0,112,0,161,0,18,0,0,0,201,0,36,0,194,0,90,0,21,0,16,0,0,0,82,0,162,0,49,0,174,0,30,0,142,0,98,0,109,0,92,0,202,0,223,0,244,0,80,0,36,0,207,0,154,0,0,0,27,0,16,0,24,0,170,0,0,0,54,0,0,0,157,0,37,0,245,0,254,0,0,0,248,0,17,0,0,0,230,0,182,0,173,0,237,0,42,0,203,0,104,0,253,0,184,0,107,0,0,0,181,0,59,0,140,0,251,0,137,0,84,0,39,0,90,0,222,0,199,0,182,0,64,0,0,0,118,0,166,0,105,0,129,0,182,0,233,0,229,0,155,0,90,0,77,0,0,0,79,0,58,0,176,0,226,0,67,0,0,0,0,0,149,0,0,0,0,0,59,0,72,0,201,0,219,0,0,0,42,0,234,0,0,0,212,0,174,0,60,0,215,0,181,0,0,0,0,0,156,0,0,0,230,0,196,0,212,0,135,0,61,0,78,0,0,0,29,0,127,0,0,0,120,0,12,0,235,0,168,0,146,0,216,0,51,0,44,0,21,0,0,0,212,0,106,0,122,0,0,0,186,0,0,0,0,0,91,0,46,0,186,0,182,0,27,0,65,0,0,0,104,0,0,0,127,0,51,0,222,0,0,0,64,0,0,0,124,0,0,0,144,0,0,0,208,0,81,0,110,0,234,0,218,0,154,0,87,0,249,0,145,0,43,0,182,0,64,0,219,0,218,0,244,0,0,0,129,0,166,0,199,0,175,0,65,0,0,0,112,0,183,0,0,0,254,0,7,0,220,0,0,0,82,0,68,0,242,0,0,0,188,0,157,0,0,0,0,0,213,0,0,0,0,0,210,0,215,0,177,0,118,0,178,0,245,0,146,0,230,0,19,0,228,0,215,0,55,0,95,0,95,0,69,0,192,0,31,0,0,0,214,0,247,0,38,0,141,0,103,0,105,0,165,0,53,0,125,0,120,0,28,0,5,0,70,0,105,0,221,0,120,0,149,0,209,0,5,0,168,0,214,0,77,0,0,0,200,0,0,0,66,0,108,0,40,0,170,0,0,0,179,0,3,0,155,0,10,0,247,0,78,0,72,0,44,0,0,0,0,0,173,0,61,0,191,0,0,0,188,0,0,0,171,0,13,0,0,0,237,0,0,0,42,0,188,0,18,0,145,0,202,0,192,0,98,0,54,0,0,0,5,0,233,0,0,0,0,0,136,0,0,0,159,0,0,0,201,0,37,0,82,0,144,0,13,0,198,0,0,0,178,0,31,0,13,0,0,0,240,0,187,0,240,0,27,0,24,0,48,0,227,0,148,0,0,0,113,0,242,0,208,0,179,0,0,0,48,0,212,0,92,0,139,0,24,0,12,0,51,0,232,0,95,0,114,0,57,0,48,0,0,0,231,0,150,0,42,0,81,0,116,0,119,0,0,0,71,0,0,0,0,0,39,0,67,0,83,0,138,0,20,0,46,0,188,0,0,0,204,0,0,0,0,0,185,0,208,0,209,0,217,0,55,0,29,0,43,0,124,0,166,0,32,0,0,0,36,0,62,0,0,0,147,0,45,0,149,0,4,0,10,0,234,0,0,0,0,0,199,0,195,0,17,0,0,0,204,0,59,0,0,0,137,0,242,0,4,0,162,0,0,0,245,0,125,0,254,0,164,0,0,0,0,0,0,0,87,0,212,0,16,0,111,0,4,0,0,0,168,0,0,0,10,0,121,0,166,0,0,0,151,0,229,0,103,0,212,0,247,0,162,0,153,0,249,0,199,0,0,0,37,0,207,0,168,0,113,0,16,0,92,0,0,0,255,0,0,0,245,0,55,0,0,0,140,0,85,0,0,0,238,0,158,0,76,0,205,0,195,0,38,0,116,0,211,0,236,0,69,0,86,0,37,0,97,0,142,0,155,0,170,0,130,0,49,0,0,0,0,0,0,0,0,0,195,0,114,0,0,0,14,0,0,0,47,0,10,0,0,0,224,0,44,0,25,0,17,0,95,0,0,0,206,0,45,0,131,0,40,0,188,0,182,0,93,0,65,0,105,0,152,0,0,0,133,0,0,0,254,0,0,0,57,0,62,0,204,0,162,0,0,0,221,0,69,0,7,0,0,0,215,0,109,0,0,0,171,0,144,0,77,0,68,0,34,0,189,0,0,0,12,0,249,0,0,0,95,0,27,0,80,0,131,0);
signal scenario_full  : scenario_type := (0,0,104,31,251,31,251,30,240,31,240,30,242,31,56,31,48,31,170,31,175,31,181,31,195,31,36,31,211,31,159,31,218,31,147,31,147,30,147,29,147,28,131,31,147,31,189,31,189,30,232,31,178,31,41,31,34,31,32,31,116,31,116,30,203,31,84,31,84,30,84,29,122,31,97,31,47,31,47,30,47,29,47,28,25,31,224,31,204,31,204,30,151,31,90,31,225,31,187,31,90,31,33,31,163,31,16,31,95,31,246,31,20,31,20,30,139,31,174,31,133,31,154,31,154,30,240,31,247,31,247,30,130,31,187,31,173,31,173,30,130,31,130,30,125,31,8,31,241,31,185,31,210,31,5,31,150,31,201,31,164,31,41,31,139,31,95,31,102,31,136,31,136,30,1,31,132,31,183,31,183,30,52,31,250,31,254,31,3,31,3,30,73,31,73,30,251,31,157,31,143,31,234,31,124,31,164,31,5,31,206,31,154,31,43,31,121,31,80,31,176,31,134,31,78,31,181,31,148,31,248,31,172,31,136,31,215,31,7,31,134,31,113,31,15,31,70,31,211,31,150,31,57,31,65,31,65,30,65,29,65,28,65,27,34,31,34,30,34,31,154,31,57,31,156,31,85,31,18,31,100,31,199,31,116,31,186,31,160,31,57,31,129,31,104,31,75,31,120,31,120,30,120,29,168,31,209,31,209,30,168,31,161,31,242,31,179,31,48,31,222,31,224,31,252,31,252,30,228,31,66,31,177,31,253,31,253,30,89,31,89,31,89,30,79,31,9,31,94,31,94,30,44,31,36,31,173,31,114,31,113,31,113,30,74,31,74,30,174,31,125,31,45,31,141,31,98,31,21,31,135,31,37,31,37,30,138,31,209,31,33,31,47,31,182,31,177,31,154,31,97,31,69,31,125,31,125,30,125,29,253,31,2,31,58,31,4,31,17,31,52,31,12,31,238,31,238,30,24,31,235,31,123,31,148,31,162,31,162,30,114,31,114,30,114,29,122,31,85,31,100,31,13,31,139,31,245,31,175,31,253,31,200,31,250,31,47,31,8,31,37,31,223,31,133,31,42,31,42,30,203,31,156,31,174,31,127,31,249,31,20,31,237,31,237,30,22,31,239,31,22,31,8,31,1,31,1,30,165,31,20,31,20,30,20,29,166,31,166,30,166,29,82,31,229,31,201,31,201,30,184,31,184,30,20,31,81,31,32,31,32,30,202,31,219,31,196,31,12,31,112,31,81,31,226,31,226,30,68,31,172,31,120,31,149,31,149,30,57,31,134,31,108,31,108,30,112,31,161,31,18,31,18,30,201,31,36,31,194,31,90,31,21,31,16,31,16,30,82,31,162,31,49,31,174,31,30,31,142,31,98,31,109,31,92,31,202,31,223,31,244,31,80,31,36,31,207,31,154,31,154,30,27,31,16,31,24,31,170,31,170,30,54,31,54,30,157,31,37,31,245,31,254,31,254,30,248,31,17,31,17,30,230,31,182,31,173,31,237,31,42,31,203,31,104,31,253,31,184,31,107,31,107,30,181,31,59,31,140,31,251,31,137,31,84,31,39,31,90,31,222,31,199,31,182,31,64,31,64,30,118,31,166,31,105,31,129,31,182,31,233,31,229,31,155,31,90,31,77,31,77,30,79,31,58,31,176,31,226,31,67,31,67,30,67,29,149,31,149,30,149,29,59,31,72,31,201,31,219,31,219,30,42,31,234,31,234,30,212,31,174,31,60,31,215,31,181,31,181,30,181,29,156,31,156,30,230,31,196,31,212,31,135,31,61,31,78,31,78,30,29,31,127,31,127,30,120,31,12,31,235,31,168,31,146,31,216,31,51,31,44,31,21,31,21,30,212,31,106,31,122,31,122,30,186,31,186,30,186,29,91,31,46,31,186,31,182,31,27,31,65,31,65,30,104,31,104,30,127,31,51,31,222,31,222,30,64,31,64,30,124,31,124,30,144,31,144,30,208,31,81,31,110,31,234,31,218,31,154,31,87,31,249,31,145,31,43,31,182,31,64,31,219,31,218,31,244,31,244,30,129,31,166,31,199,31,175,31,65,31,65,30,112,31,183,31,183,30,254,31,7,31,220,31,220,30,82,31,68,31,242,31,242,30,188,31,157,31,157,30,157,29,213,31,213,30,213,29,210,31,215,31,177,31,118,31,178,31,245,31,146,31,230,31,19,31,228,31,215,31,55,31,95,31,95,31,69,31,192,31,31,31,31,30,214,31,247,31,38,31,141,31,103,31,105,31,165,31,53,31,125,31,120,31,28,31,5,31,70,31,105,31,221,31,120,31,149,31,209,31,5,31,168,31,214,31,77,31,77,30,200,31,200,30,66,31,108,31,40,31,170,31,170,30,179,31,3,31,155,31,10,31,247,31,78,31,72,31,44,31,44,30,44,29,173,31,61,31,191,31,191,30,188,31,188,30,171,31,13,31,13,30,237,31,237,30,42,31,188,31,18,31,145,31,202,31,192,31,98,31,54,31,54,30,5,31,233,31,233,30,233,29,136,31,136,30,159,31,159,30,201,31,37,31,82,31,144,31,13,31,198,31,198,30,178,31,31,31,13,31,13,30,240,31,187,31,240,31,27,31,24,31,48,31,227,31,148,31,148,30,113,31,242,31,208,31,179,31,179,30,48,31,212,31,92,31,139,31,24,31,12,31,51,31,232,31,95,31,114,31,57,31,48,31,48,30,231,31,150,31,42,31,81,31,116,31,119,31,119,30,71,31,71,30,71,29,39,31,67,31,83,31,138,31,20,31,46,31,188,31,188,30,204,31,204,30,204,29,185,31,208,31,209,31,217,31,55,31,29,31,43,31,124,31,166,31,32,31,32,30,36,31,62,31,62,30,147,31,45,31,149,31,4,31,10,31,234,31,234,30,234,29,199,31,195,31,17,31,17,30,204,31,59,31,59,30,137,31,242,31,4,31,162,31,162,30,245,31,125,31,254,31,164,31,164,30,164,29,164,28,87,31,212,31,16,31,111,31,4,31,4,30,168,31,168,30,10,31,121,31,166,31,166,30,151,31,229,31,103,31,212,31,247,31,162,31,153,31,249,31,199,31,199,30,37,31,207,31,168,31,113,31,16,31,92,31,92,30,255,31,255,30,245,31,55,31,55,30,140,31,85,31,85,30,238,31,158,31,76,31,205,31,195,31,38,31,116,31,211,31,236,31,69,31,86,31,37,31,97,31,142,31,155,31,170,31,130,31,49,31,49,30,49,29,49,28,49,27,195,31,114,31,114,30,14,31,14,30,47,31,10,31,10,30,224,31,44,31,25,31,17,31,95,31,95,30,206,31,45,31,131,31,40,31,188,31,182,31,93,31,65,31,105,31,152,31,152,30,133,31,133,30,254,31,254,30,57,31,62,31,204,31,162,31,162,30,221,31,69,31,7,31,7,30,215,31,109,31,109,30,171,31,144,31,77,31,68,31,34,31,189,31,189,30,12,31,249,31,249,30,95,31,27,31,80,31,131,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
