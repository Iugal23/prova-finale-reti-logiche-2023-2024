-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_888 is
end project_tb_888;

architecture project_tb_arch_888 of project_tb_888 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 275;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (226,0,236,0,209,0,182,0,58,0,143,0,103,0,81,0,93,0,121,0,96,0,218,0,7,0,0,0,81,0,245,0,197,0,192,0,76,0,95,0,0,0,176,0,0,0,205,0,28,0,64,0,173,0,226,0,0,0,64,0,53,0,0,0,237,0,90,0,168,0,0,0,60,0,189,0,211,0,0,0,237,0,85,0,208,0,157,0,43,0,0,0,0,0,199,0,119,0,146,0,0,0,130,0,0,0,216,0,104,0,65,0,233,0,103,0,71,0,9,0,233,0,116,0,140,0,175,0,143,0,248,0,0,0,140,0,100,0,101,0,0,0,51,0,6,0,90,0,0,0,196,0,76,0,34,0,52,0,0,0,0,0,232,0,46,0,0,0,118,0,0,0,0,0,197,0,121,0,0,0,10,0,0,0,88,0,0,0,0,0,132,0,88,0,248,0,156,0,43,0,110,0,0,0,89,0,144,0,134,0,0,0,178,0,148,0,136,0,0,0,159,0,210,0,122,0,0,0,0,0,189,0,81,0,39,0,28,0,222,0,0,0,177,0,246,0,146,0,81,0,243,0,200,0,186,0,23,0,24,0,0,0,63,0,0,0,239,0,0,0,108,0,0,0,218,0,54,0,248,0,81,0,135,0,218,0,213,0,0,0,129,0,0,0,167,0,0,0,145,0,171,0,114,0,233,0,137,0,61,0,35,0,0,0,108,0,0,0,4,0,15,0,204,0,162,0,221,0,0,0,231,0,8,0,159,0,148,0,0,0,0,0,126,0,133,0,0,0,48,0,254,0,177,0,70,0,12,0,0,0,11,0,42,0,14,0,250,0,0,0,0,0,78,0,35,0,0,0,234,0,76,0,0,0,59,0,62,0,0,0,112,0,0,0,237,0,147,0,0,0,131,0,210,0,111,0,0,0,16,0,85,0,0,0,97,0,56,0,0,0,79,0,0,0,110,0,104,0,23,0,8,0,90,0,217,0,226,0,143,0,0,0,159,0,45,0,161,0,0,0,243,0,184,0,231,0,254,0,116,0,3,0,0,0,126,0,128,0,138,0,24,0,0,0,204,0,158,0,210,0,47,0,145,0,204,0,247,0,59,0,60,0,103,0,234,0,0,0,127,0,206,0,121,0,0,0,93,0,215,0,74,0,0,0,19,0,51,0,248,0,86,0,182,0,233,0,0,0,208,0,0,0,248,0,19,0,239,0,132,0,168,0,0,0,0,0,155,0,252,0);
signal scenario_full  : scenario_type := (226,31,236,31,209,31,182,31,58,31,143,31,103,31,81,31,93,31,121,31,96,31,218,31,7,31,7,30,81,31,245,31,197,31,192,31,76,31,95,31,95,30,176,31,176,30,205,31,28,31,64,31,173,31,226,31,226,30,64,31,53,31,53,30,237,31,90,31,168,31,168,30,60,31,189,31,211,31,211,30,237,31,85,31,208,31,157,31,43,31,43,30,43,29,199,31,119,31,146,31,146,30,130,31,130,30,216,31,104,31,65,31,233,31,103,31,71,31,9,31,233,31,116,31,140,31,175,31,143,31,248,31,248,30,140,31,100,31,101,31,101,30,51,31,6,31,90,31,90,30,196,31,76,31,34,31,52,31,52,30,52,29,232,31,46,31,46,30,118,31,118,30,118,29,197,31,121,31,121,30,10,31,10,30,88,31,88,30,88,29,132,31,88,31,248,31,156,31,43,31,110,31,110,30,89,31,144,31,134,31,134,30,178,31,148,31,136,31,136,30,159,31,210,31,122,31,122,30,122,29,189,31,81,31,39,31,28,31,222,31,222,30,177,31,246,31,146,31,81,31,243,31,200,31,186,31,23,31,24,31,24,30,63,31,63,30,239,31,239,30,108,31,108,30,218,31,54,31,248,31,81,31,135,31,218,31,213,31,213,30,129,31,129,30,167,31,167,30,145,31,171,31,114,31,233,31,137,31,61,31,35,31,35,30,108,31,108,30,4,31,15,31,204,31,162,31,221,31,221,30,231,31,8,31,159,31,148,31,148,30,148,29,126,31,133,31,133,30,48,31,254,31,177,31,70,31,12,31,12,30,11,31,42,31,14,31,250,31,250,30,250,29,78,31,35,31,35,30,234,31,76,31,76,30,59,31,62,31,62,30,112,31,112,30,237,31,147,31,147,30,131,31,210,31,111,31,111,30,16,31,85,31,85,30,97,31,56,31,56,30,79,31,79,30,110,31,104,31,23,31,8,31,90,31,217,31,226,31,143,31,143,30,159,31,45,31,161,31,161,30,243,31,184,31,231,31,254,31,116,31,3,31,3,30,126,31,128,31,138,31,24,31,24,30,204,31,158,31,210,31,47,31,145,31,204,31,247,31,59,31,60,31,103,31,234,31,234,30,127,31,206,31,121,31,121,30,93,31,215,31,74,31,74,30,19,31,51,31,248,31,86,31,182,31,233,31,233,30,208,31,208,30,248,31,19,31,239,31,132,31,168,31,168,30,168,29,155,31,252,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
