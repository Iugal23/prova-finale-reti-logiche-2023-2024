-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_180 is
end project_tb_180;

architecture project_tb_arch_180 of project_tb_180 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 981;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (107,0,0,0,25,0,202,0,21,0,117,0,77,0,28,0,9,0,89,0,225,0,112,0,117,0,0,0,58,0,136,0,69,0,204,0,142,0,217,0,255,0,88,0,152,0,0,0,27,0,0,0,243,0,148,0,29,0,77,0,7,0,2,0,101,0,0,0,95,0,0,0,50,0,97,0,58,0,210,0,142,0,0,0,0,0,0,0,59,0,82,0,116,0,40,0,248,0,0,0,204,0,0,0,0,0,47,0,35,0,0,0,182,0,226,0,0,0,43,0,252,0,0,0,93,0,234,0,183,0,0,0,53,0,30,0,0,0,0,0,128,0,171,0,62,0,177,0,0,0,53,0,79,0,165,0,62,0,13,0,0,0,126,0,47,0,123,0,248,0,139,0,149,0,56,0,91,0,0,0,46,0,0,0,83,0,186,0,242,0,0,0,0,0,212,0,38,0,0,0,95,0,43,0,0,0,245,0,51,0,143,0,112,0,71,0,35,0,116,0,0,0,149,0,14,0,102,0,208,0,10,0,157,0,0,0,192,0,0,0,0,0,165,0,199,0,80,0,0,0,124,0,40,0,54,0,244,0,90,0,0,0,0,0,97,0,134,0,107,0,0,0,61,0,246,0,0,0,87,0,0,0,237,0,135,0,115,0,130,0,204,0,158,0,226,0,253,0,0,0,224,0,76,0,75,0,0,0,142,0,242,0,80,0,207,0,0,0,221,0,0,0,0,0,18,0,198,0,46,0,124,0,0,0,195,0,0,0,137,0,167,0,0,0,208,0,21,0,200,0,0,0,100,0,252,0,110,0,0,0,117,0,210,0,65,0,57,0,4,0,100,0,100,0,219,0,5,0,110,0,74,0,4,0,52,0,59,0,224,0,117,0,70,0,76,0,33,0,0,0,0,0,254,0,60,0,177,0,0,0,101,0,181,0,215,0,105,0,4,0,34,0,0,0,82,0,14,0,12,0,212,0,0,0,0,0,56,0,137,0,55,0,0,0,35,0,88,0,182,0,86,0,0,0,171,0,0,0,0,0,74,0,252,0,0,0,157,0,36,0,0,0,139,0,166,0,100,0,140,0,0,0,0,0,0,0,0,0,114,0,48,0,255,0,47,0,111,0,124,0,177,0,169,0,232,0,184,0,0,0,0,0,27,0,0,0,0,0,0,0,0,0,0,0,162,0,0,0,136,0,48,0,119,0,0,0,44,0,46,0,230,0,197,0,98,0,117,0,147,0,167,0,186,0,0,0,134,0,237,0,91,0,119,0,81,0,144,0,4,0,199,0,190,0,20,0,108,0,0,0,0,0,74,0,0,0,30,0,0,0,61,0,175,0,110,0,23,0,0,0,0,0,219,0,108,0,28,0,250,0,88,0,0,0,237,0,167,0,54,0,243,0,67,0,94,0,0,0,57,0,5,0,115,0,91,0,110,0,128,0,252,0,255,0,0,0,46,0,83,0,23,0,33,0,237,0,0,0,0,0,0,0,0,0,0,0,242,0,0,0,73,0,0,0,89,0,0,0,167,0,239,0,0,0,70,0,43,0,235,0,48,0,0,0,6,0,0,0,150,0,0,0,141,0,136,0,25,0,198,0,0,0,0,0,251,0,76,0,29,0,236,0,113,0,38,0,166,0,49,0,233,0,100,0,78,0,0,0,216,0,33,0,176,0,120,0,130,0,254,0,164,0,113,0,0,0,100,0,91,0,0,0,0,0,50,0,151,0,238,0,124,0,49,0,22,0,133,0,235,0,0,0,109,0,216,0,248,0,67,0,0,0,192,0,219,0,63,0,158,0,78,0,241,0,49,0,225,0,213,0,224,0,106,0,250,0,183,0,22,0,43,0,227,0,189,0,35,0,239,0,155,0,28,0,156,0,124,0,45,0,63,0,0,0,0,0,114,0,185,0,133,0,0,0,0,0,50,0,11,0,166,0,93,0,99,0,28,0,109,0,58,0,0,0,130,0,61,0,197,0,229,0,52,0,130,0,122,0,237,0,0,0,122,0,143,0,90,0,0,0,240,0,0,0,171,0,192,0,49,0,0,0,183,0,0,0,225,0,52,0,92,0,88,0,143,0,180,0,115,0,0,0,103,0,0,0,174,0,0,0,0,0,5,0,63,0,119,0,0,0,35,0,0,0,56,0,237,0,250,0,246,0,255,0,18,0,0,0,0,0,9,0,106,0,167,0,64,0,131,0,185,0,0,0,184,0,0,0,191,0,252,0,0,0,127,0,13,0,106,0,114,0,0,0,170,0,14,0,149,0,241,0,222,0,231,0,0,0,55,0,239,0,61,0,0,0,184,0,112,0,96,0,2,0,41,0,188,0,157,0,4,0,172,0,83,0,0,0,21,0,139,0,253,0,13,0,98,0,200,0,29,0,37,0,0,0,93,0,28,0,0,0,0,0,56,0,12,0,219,0,243,0,18,0,252,0,145,0,0,0,218,0,148,0,97,0,245,0,46,0,0,0,0,0,60,0,5,0,235,0,0,0,235,0,98,0,248,0,0,0,3,0,138,0,129,0,0,0,49,0,0,0,31,0,6,0,159,0,158,0,165,0,128,0,167,0,188,0,51,0,81,0,240,0,13,0,163,0,243,0,0,0,83,0,133,0,236,0,3,0,220,0,187,0,165,0,3,0,13,0,218,0,0,0,242,0,7,0,217,0,0,0,111,0,149,0,0,0,182,0,0,0,41,0,32,0,7,0,14,0,67,0,0,0,74,0,186,0,180,0,0,0,89,0,143,0,238,0,143,0,0,0,0,0,48,0,50,0,187,0,89,0,114,0,77,0,247,0,91,0,68,0,191,0,80,0,155,0,43,0,220,0,201,0,74,0,173,0,161,0,23,0,10,0,56,0,139,0,222,0,0,0,108,0,163,0,0,0,68,0,202,0,200,0,108,0,174,0,0,0,41,0,108,0,46,0,73,0,105,0,71,0,0,0,177,0,17,0,0,0,23,0,14,0,143,0,121,0,49,0,209,0,179,0,63,0,13,0,2,0,0,0,104,0,13,0,0,0,155,0,0,0,110,0,37,0,0,0,127,0,0,0,0,0,241,0,255,0,0,0,158,0,30,0,115,0,130,0,34,0,231,0,228,0,161,0,0,0,125,0,182,0,247,0,208,0,0,0,253,0,0,0,38,0,21,0,181,0,55,0,22,0,25,0,214,0,74,0,10,0,115,0,217,0,195,0,203,0,184,0,0,0,28,0,96,0,0,0,41,0,216,0,107,0,0,0,192,0,31,0,0,0,232,0,0,0,199,0,23,0,49,0,49,0,206,0,187,0,102,0,70,0,0,0,240,0,163,0,0,0,0,0,0,0,62,0,24,0,141,0,33,0,199,0,46,0,233,0,75,0,83,0,0,0,36,0,0,0,158,0,0,0,3,0,0,0,211,0,119,0,224,0,0,0,109,0,114,0,97,0,0,0,0,0,0,0,46,0,16,0,93,0,55,0,216,0,131,0,189,0,86,0,186,0,0,0,229,0,132,0,181,0,229,0,116,0,251,0,24,0,81,0,150,0,190,0,176,0,145,0,171,0,130,0,135,0,222,0,206,0,248,0,72,0,112,0,177,0,243,0,7,0,192,0,66,0,0,0,168,0,171,0,43,0,0,0,242,0,237,0,65,0,57,0,0,0,136,0,120,0,171,0,0,0,249,0,42,0,47,0,240,0,235,0,169,0,6,0,25,0,255,0,66,0,69,0,214,0,60,0,58,0,167,0,20,0,0,0,95,0,136,0,106,0,174,0,255,0,90,0,109,0,132,0,207,0,20,0,104,0,0,0,193,0,68,0,0,0,239,0,199,0,215,0,214,0,149,0,26,0,30,0,0,0,52,0,199,0,215,0,243,0,23,0,203,0,57,0,0,0,26,0,186,0,83,0,91,0,13,0,5,0,176,0,5,0,0,0,116,0,104,0,38,0,61,0,134,0,94,0,123,0,14,0,102,0,61,0,61,0,54,0,0,0,143,0,105,0,224,0,235,0,158,0,26,0,0,0,174,0,0,0,21,0,53,0,246,0,6,0,49,0,90,0,194,0,156,0,43,0,0,0,211,0,137,0,71,0,147,0,53,0,0,0,64,0,50,0,0,0,0,0,31,0,254,0,0,0,43,0,131,0,18,0,130,0,54,0,0,0,0,0,124,0,183,0,165,0,59,0,141,0,0,0,0,0,0,0,0,0,166,0,17,0,47,0,170,0,136,0,40,0,150,0,119,0,192,0,218,0,135,0,254,0,0,0,81,0,0,0,157,0,207,0,144,0,0,0,0,0,0,0,160,0,0,0,207,0,0,0,0,0,166,0,68,0,0,0,100,0,23,0,81,0,236,0,183,0,0,0,164,0,0,0,96,0,234,0,200,0,19,0,253,0,155,0,215,0,207,0,206,0);
signal scenario_full  : scenario_type := (107,31,107,30,25,31,202,31,21,31,117,31,77,31,28,31,9,31,89,31,225,31,112,31,117,31,117,30,58,31,136,31,69,31,204,31,142,31,217,31,255,31,88,31,152,31,152,30,27,31,27,30,243,31,148,31,29,31,77,31,7,31,2,31,101,31,101,30,95,31,95,30,50,31,97,31,58,31,210,31,142,31,142,30,142,29,142,28,59,31,82,31,116,31,40,31,248,31,248,30,204,31,204,30,204,29,47,31,35,31,35,30,182,31,226,31,226,30,43,31,252,31,252,30,93,31,234,31,183,31,183,30,53,31,30,31,30,30,30,29,128,31,171,31,62,31,177,31,177,30,53,31,79,31,165,31,62,31,13,31,13,30,126,31,47,31,123,31,248,31,139,31,149,31,56,31,91,31,91,30,46,31,46,30,83,31,186,31,242,31,242,30,242,29,212,31,38,31,38,30,95,31,43,31,43,30,245,31,51,31,143,31,112,31,71,31,35,31,116,31,116,30,149,31,14,31,102,31,208,31,10,31,157,31,157,30,192,31,192,30,192,29,165,31,199,31,80,31,80,30,124,31,40,31,54,31,244,31,90,31,90,30,90,29,97,31,134,31,107,31,107,30,61,31,246,31,246,30,87,31,87,30,237,31,135,31,115,31,130,31,204,31,158,31,226,31,253,31,253,30,224,31,76,31,75,31,75,30,142,31,242,31,80,31,207,31,207,30,221,31,221,30,221,29,18,31,198,31,46,31,124,31,124,30,195,31,195,30,137,31,167,31,167,30,208,31,21,31,200,31,200,30,100,31,252,31,110,31,110,30,117,31,210,31,65,31,57,31,4,31,100,31,100,31,219,31,5,31,110,31,74,31,4,31,52,31,59,31,224,31,117,31,70,31,76,31,33,31,33,30,33,29,254,31,60,31,177,31,177,30,101,31,181,31,215,31,105,31,4,31,34,31,34,30,82,31,14,31,12,31,212,31,212,30,212,29,56,31,137,31,55,31,55,30,35,31,88,31,182,31,86,31,86,30,171,31,171,30,171,29,74,31,252,31,252,30,157,31,36,31,36,30,139,31,166,31,100,31,140,31,140,30,140,29,140,28,140,27,114,31,48,31,255,31,47,31,111,31,124,31,177,31,169,31,232,31,184,31,184,30,184,29,27,31,27,30,27,29,27,28,27,27,27,26,162,31,162,30,136,31,48,31,119,31,119,30,44,31,46,31,230,31,197,31,98,31,117,31,147,31,167,31,186,31,186,30,134,31,237,31,91,31,119,31,81,31,144,31,4,31,199,31,190,31,20,31,108,31,108,30,108,29,74,31,74,30,30,31,30,30,61,31,175,31,110,31,23,31,23,30,23,29,219,31,108,31,28,31,250,31,88,31,88,30,237,31,167,31,54,31,243,31,67,31,94,31,94,30,57,31,5,31,115,31,91,31,110,31,128,31,252,31,255,31,255,30,46,31,83,31,23,31,33,31,237,31,237,30,237,29,237,28,237,27,237,26,242,31,242,30,73,31,73,30,89,31,89,30,167,31,239,31,239,30,70,31,43,31,235,31,48,31,48,30,6,31,6,30,150,31,150,30,141,31,136,31,25,31,198,31,198,30,198,29,251,31,76,31,29,31,236,31,113,31,38,31,166,31,49,31,233,31,100,31,78,31,78,30,216,31,33,31,176,31,120,31,130,31,254,31,164,31,113,31,113,30,100,31,91,31,91,30,91,29,50,31,151,31,238,31,124,31,49,31,22,31,133,31,235,31,235,30,109,31,216,31,248,31,67,31,67,30,192,31,219,31,63,31,158,31,78,31,241,31,49,31,225,31,213,31,224,31,106,31,250,31,183,31,22,31,43,31,227,31,189,31,35,31,239,31,155,31,28,31,156,31,124,31,45,31,63,31,63,30,63,29,114,31,185,31,133,31,133,30,133,29,50,31,11,31,166,31,93,31,99,31,28,31,109,31,58,31,58,30,130,31,61,31,197,31,229,31,52,31,130,31,122,31,237,31,237,30,122,31,143,31,90,31,90,30,240,31,240,30,171,31,192,31,49,31,49,30,183,31,183,30,225,31,52,31,92,31,88,31,143,31,180,31,115,31,115,30,103,31,103,30,174,31,174,30,174,29,5,31,63,31,119,31,119,30,35,31,35,30,56,31,237,31,250,31,246,31,255,31,18,31,18,30,18,29,9,31,106,31,167,31,64,31,131,31,185,31,185,30,184,31,184,30,191,31,252,31,252,30,127,31,13,31,106,31,114,31,114,30,170,31,14,31,149,31,241,31,222,31,231,31,231,30,55,31,239,31,61,31,61,30,184,31,112,31,96,31,2,31,41,31,188,31,157,31,4,31,172,31,83,31,83,30,21,31,139,31,253,31,13,31,98,31,200,31,29,31,37,31,37,30,93,31,28,31,28,30,28,29,56,31,12,31,219,31,243,31,18,31,252,31,145,31,145,30,218,31,148,31,97,31,245,31,46,31,46,30,46,29,60,31,5,31,235,31,235,30,235,31,98,31,248,31,248,30,3,31,138,31,129,31,129,30,49,31,49,30,31,31,6,31,159,31,158,31,165,31,128,31,167,31,188,31,51,31,81,31,240,31,13,31,163,31,243,31,243,30,83,31,133,31,236,31,3,31,220,31,187,31,165,31,3,31,13,31,218,31,218,30,242,31,7,31,217,31,217,30,111,31,149,31,149,30,182,31,182,30,41,31,32,31,7,31,14,31,67,31,67,30,74,31,186,31,180,31,180,30,89,31,143,31,238,31,143,31,143,30,143,29,48,31,50,31,187,31,89,31,114,31,77,31,247,31,91,31,68,31,191,31,80,31,155,31,43,31,220,31,201,31,74,31,173,31,161,31,23,31,10,31,56,31,139,31,222,31,222,30,108,31,163,31,163,30,68,31,202,31,200,31,108,31,174,31,174,30,41,31,108,31,46,31,73,31,105,31,71,31,71,30,177,31,17,31,17,30,23,31,14,31,143,31,121,31,49,31,209,31,179,31,63,31,13,31,2,31,2,30,104,31,13,31,13,30,155,31,155,30,110,31,37,31,37,30,127,31,127,30,127,29,241,31,255,31,255,30,158,31,30,31,115,31,130,31,34,31,231,31,228,31,161,31,161,30,125,31,182,31,247,31,208,31,208,30,253,31,253,30,38,31,21,31,181,31,55,31,22,31,25,31,214,31,74,31,10,31,115,31,217,31,195,31,203,31,184,31,184,30,28,31,96,31,96,30,41,31,216,31,107,31,107,30,192,31,31,31,31,30,232,31,232,30,199,31,23,31,49,31,49,31,206,31,187,31,102,31,70,31,70,30,240,31,163,31,163,30,163,29,163,28,62,31,24,31,141,31,33,31,199,31,46,31,233,31,75,31,83,31,83,30,36,31,36,30,158,31,158,30,3,31,3,30,211,31,119,31,224,31,224,30,109,31,114,31,97,31,97,30,97,29,97,28,46,31,16,31,93,31,55,31,216,31,131,31,189,31,86,31,186,31,186,30,229,31,132,31,181,31,229,31,116,31,251,31,24,31,81,31,150,31,190,31,176,31,145,31,171,31,130,31,135,31,222,31,206,31,248,31,72,31,112,31,177,31,243,31,7,31,192,31,66,31,66,30,168,31,171,31,43,31,43,30,242,31,237,31,65,31,57,31,57,30,136,31,120,31,171,31,171,30,249,31,42,31,47,31,240,31,235,31,169,31,6,31,25,31,255,31,66,31,69,31,214,31,60,31,58,31,167,31,20,31,20,30,95,31,136,31,106,31,174,31,255,31,90,31,109,31,132,31,207,31,20,31,104,31,104,30,193,31,68,31,68,30,239,31,199,31,215,31,214,31,149,31,26,31,30,31,30,30,52,31,199,31,215,31,243,31,23,31,203,31,57,31,57,30,26,31,186,31,83,31,91,31,13,31,5,31,176,31,5,31,5,30,116,31,104,31,38,31,61,31,134,31,94,31,123,31,14,31,102,31,61,31,61,31,54,31,54,30,143,31,105,31,224,31,235,31,158,31,26,31,26,30,174,31,174,30,21,31,53,31,246,31,6,31,49,31,90,31,194,31,156,31,43,31,43,30,211,31,137,31,71,31,147,31,53,31,53,30,64,31,50,31,50,30,50,29,31,31,254,31,254,30,43,31,131,31,18,31,130,31,54,31,54,30,54,29,124,31,183,31,165,31,59,31,141,31,141,30,141,29,141,28,141,27,166,31,17,31,47,31,170,31,136,31,40,31,150,31,119,31,192,31,218,31,135,31,254,31,254,30,81,31,81,30,157,31,207,31,144,31,144,30,144,29,144,28,160,31,160,30,207,31,207,30,207,29,166,31,68,31,68,30,100,31,23,31,81,31,236,31,183,31,183,30,164,31,164,30,96,31,234,31,200,31,19,31,253,31,155,31,215,31,207,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
