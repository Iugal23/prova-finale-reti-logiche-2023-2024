-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_692 is
end project_tb_692;

architecture project_tb_arch_692 of project_tb_692 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 274;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (121,0,0,0,223,0,154,0,0,0,103,0,185,0,0,0,38,0,110,0,95,0,216,0,48,0,32,0,175,0,44,0,0,0,0,0,0,0,112,0,0,0,42,0,151,0,181,0,0,0,0,0,64,0,79,0,167,0,56,0,0,0,76,0,0,0,68,0,48,0,121,0,33,0,154,0,30,0,222,0,247,0,129,0,196,0,0,0,191,0,40,0,80,0,57,0,220,0,50,0,166,0,109,0,0,0,234,0,18,0,0,0,71,0,30,0,152,0,0,0,85,0,0,0,198,0,0,0,223,0,0,0,0,0,158,0,5,0,164,0,74,0,0,0,72,0,150,0,214,0,137,0,235,0,0,0,167,0,56,0,0,0,0,0,5,0,0,0,68,0,149,0,0,0,19,0,0,0,211,0,58,0,222,0,177,0,0,0,61,0,19,0,179,0,108,0,70,0,33,0,146,0,100,0,240,0,0,0,11,0,120,0,0,0,114,0,197,0,226,0,39,0,91,0,0,0,182,0,0,0,19,0,70,0,121,0,174,0,125,0,0,0,228,0,117,0,0,0,0,0,94,0,0,0,160,0,56,0,90,0,0,0,20,0,160,0,210,0,0,0,58,0,81,0,130,0,192,0,32,0,11,0,137,0,237,0,115,0,228,0,157,0,125,0,146,0,193,0,183,0,206,0,151,0,124,0,0,0,0,0,151,0,0,0,51,0,0,0,183,0,145,0,161,0,0,0,188,0,87,0,170,0,27,0,0,0,52,0,110,0,91,0,0,0,147,0,16,0,218,0,210,0,24,0,10,0,11,0,174,0,92,0,248,0,21,0,31,0,0,0,237,0,17,0,0,0,79,0,0,0,168,0,239,0,87,0,0,0,255,0,240,0,56,0,105,0,9,0,163,0,219,0,174,0,137,0,0,0,114,0,0,0,229,0,146,0,189,0,74,0,0,0,253,0,53,0,94,0,8,0,63,0,12,0,247,0,79,0,119,0,210,0,70,0,95,0,32,0,174,0,166,0,181,0,49,0,82,0,247,0,49,0,254,0,137,0,21,0,173,0,0,0,0,0,0,0,108,0,0,0,243,0,231,0,172,0,248,0,225,0,3,0,98,0,206,0,0,0,5,0,55,0,84,0,169,0,0,0,196,0,190,0,217,0,158,0,123,0,0,0,2,0,236,0,52,0,217,0,237,0,170,0,0,0,68,0,44,0,2,0,105,0,117,0,147,0,182,0);
signal scenario_full  : scenario_type := (121,31,121,30,223,31,154,31,154,30,103,31,185,31,185,30,38,31,110,31,95,31,216,31,48,31,32,31,175,31,44,31,44,30,44,29,44,28,112,31,112,30,42,31,151,31,181,31,181,30,181,29,64,31,79,31,167,31,56,31,56,30,76,31,76,30,68,31,48,31,121,31,33,31,154,31,30,31,222,31,247,31,129,31,196,31,196,30,191,31,40,31,80,31,57,31,220,31,50,31,166,31,109,31,109,30,234,31,18,31,18,30,71,31,30,31,152,31,152,30,85,31,85,30,198,31,198,30,223,31,223,30,223,29,158,31,5,31,164,31,74,31,74,30,72,31,150,31,214,31,137,31,235,31,235,30,167,31,56,31,56,30,56,29,5,31,5,30,68,31,149,31,149,30,19,31,19,30,211,31,58,31,222,31,177,31,177,30,61,31,19,31,179,31,108,31,70,31,33,31,146,31,100,31,240,31,240,30,11,31,120,31,120,30,114,31,197,31,226,31,39,31,91,31,91,30,182,31,182,30,19,31,70,31,121,31,174,31,125,31,125,30,228,31,117,31,117,30,117,29,94,31,94,30,160,31,56,31,90,31,90,30,20,31,160,31,210,31,210,30,58,31,81,31,130,31,192,31,32,31,11,31,137,31,237,31,115,31,228,31,157,31,125,31,146,31,193,31,183,31,206,31,151,31,124,31,124,30,124,29,151,31,151,30,51,31,51,30,183,31,145,31,161,31,161,30,188,31,87,31,170,31,27,31,27,30,52,31,110,31,91,31,91,30,147,31,16,31,218,31,210,31,24,31,10,31,11,31,174,31,92,31,248,31,21,31,31,31,31,30,237,31,17,31,17,30,79,31,79,30,168,31,239,31,87,31,87,30,255,31,240,31,56,31,105,31,9,31,163,31,219,31,174,31,137,31,137,30,114,31,114,30,229,31,146,31,189,31,74,31,74,30,253,31,53,31,94,31,8,31,63,31,12,31,247,31,79,31,119,31,210,31,70,31,95,31,32,31,174,31,166,31,181,31,49,31,82,31,247,31,49,31,254,31,137,31,21,31,173,31,173,30,173,29,173,28,108,31,108,30,243,31,231,31,172,31,248,31,225,31,3,31,98,31,206,31,206,30,5,31,55,31,84,31,169,31,169,30,196,31,190,31,217,31,158,31,123,31,123,30,2,31,236,31,52,31,217,31,237,31,170,31,170,30,68,31,44,31,2,31,105,31,117,31,147,31,182,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
