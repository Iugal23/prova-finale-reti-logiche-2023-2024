-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 726;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,147,0,115,0,211,0,134,0,155,0,195,0,0,0,0,0,237,0,199,0,8,0,255,0,96,0,59,0,179,0,72,0,0,0,238,0,254,0,62,0,34,0,92,0,112,0,39,0,238,0,0,0,0,0,0,0,9,0,164,0,0,0,49,0,10,0,174,0,44,0,231,0,59,0,60,0,3,0,32,0,139,0,183,0,78,0,247,0,0,0,148,0,107,0,182,0,38,0,183,0,58,0,0,0,0,0,159,0,0,0,10,0,97,0,117,0,167,0,0,0,104,0,104,0,220,0,182,0,111,0,83,0,122,0,4,0,150,0,245,0,0,0,146,0,83,0,119,0,67,0,200,0,36,0,15,0,72,0,137,0,0,0,213,0,49,0,132,0,5,0,224,0,0,0,200,0,3,0,187,0,10,0,163,0,66,0,148,0,218,0,55,0,62,0,158,0,161,0,40,0,128,0,122,0,191,0,96,0,124,0,0,0,63,0,103,0,71,0,33,0,12,0,36,0,17,0,0,0,17,0,0,0,114,0,121,0,0,0,245,0,225,0,0,0,107,0,214,0,0,0,39,0,0,0,0,0,246,0,0,0,110,0,1,0,116,0,0,0,253,0,206,0,87,0,195,0,173,0,83,0,233,0,160,0,0,0,98,0,0,0,198,0,0,0,92,0,0,0,78,0,212,0,0,0,118,0,0,0,246,0,62,0,34,0,34,0,136,0,133,0,0,0,186,0,250,0,214,0,24,0,245,0,0,0,148,0,120,0,0,0,65,0,0,0,253,0,0,0,159,0,103,0,200,0,166,0,187,0,0,0,236,0,0,0,179,0,0,0,194,0,42,0,56,0,181,0,247,0,0,0,46,0,194,0,149,0,108,0,95,0,202,0,255,0,239,0,64,0,190,0,149,0,69,0,99,0,0,0,99,0,185,0,53,0,35,0,139,0,124,0,243,0,0,0,5,0,131,0,242,0,17,0,139,0,193,0,11,0,58,0,87,0,137,0,36,0,222,0,104,0,46,0,185,0,107,0,0,0,252,0,92,0,241,0,45,0,48,0,115,0,229,0,12,0,85,0,6,0,157,0,20,0,37,0,140,0,0,0,185,0,209,0,0,0,0,0,190,0,145,0,41,0,135,0,244,0,155,0,242,0,141,0,221,0,0,0,195,0,235,0,0,0,92,0,0,0,248,0,135,0,239,0,0,0,179,0,186,0,43,0,72,0,16,0,0,0,92,0,47,0,57,0,240,0,16,0,135,0,133,0,0,0,0,0,203,0,212,0,62,0,0,0,156,0,192,0,218,0,180,0,171,0,5,0,143,0,0,0,185,0,74,0,0,0,124,0,183,0,0,0,36,0,75,0,146,0,219,0,88,0,137,0,2,0,172,0,250,0,236,0,226,0,52,0,89,0,88,0,110,0,105,0,221,0,249,0,202,0,170,0,0,0,2,0,225,0,0,0,181,0,74,0,86,0,145,0,232,0,154,0,186,0,132,0,93,0,194,0,34,0,19,0,212,0,0,0,13,0,0,0,213,0,62,0,0,0,122,0,158,0,194,0,186,0,104,0,214,0,199,0,65,0,229,0,225,0,243,0,0,0,162,0,175,0,230,0,122,0,50,0,0,0,0,0,238,0,51,0,0,0,0,0,192,0,52,0,123,0,0,0,243,0,218,0,98,0,0,0,81,0,36,0,156,0,218,0,82,0,214,0,203,0,160,0,222,0,79,0,182,0,112,0,65,0,40,0,138,0,0,0,68,0,119,0,177,0,197,0,156,0,1,0,168,0,103,0,0,0,0,0,126,0,0,0,200,0,101,0,95,0,118,0,119,0,133,0,0,0,200,0,22,0,0,0,199,0,0,0,125,0,0,0,0,0,146,0,133,0,55,0,161,0,213,0,0,0,64,0,0,0,0,0,0,0,41,0,43,0,0,0,111,0,144,0,13,0,243,0,219,0,68,0,117,0,56,0,53,0,123,0,143,0,0,0,0,0,0,0,182,0,108,0,7,0,29,0,65,0,0,0,32,0,80,0,0,0,88,0,0,0,93,0,0,0,50,0,103,0,243,0,162,0,193,0,0,0,3,0,0,0,59,0,212,0,145,0,0,0,226,0,173,0,182,0,0,0,0,0,12,0,0,0,127,0,215,0,69,0,18,0,183,0,19,0,225,0,0,0,93,0,227,0,79,0,159,0,6,0,135,0,107,0,89,0,190,0,242,0,0,0,200,0,198,0,177,0,245,0,20,0,41,0,174,0,0,0,198,0,0,0,106,0,250,0,161,0,199,0,176,0,0,0,0,0,80,0,74,0,31,0,123,0,111,0,160,0,10,0,139,0,0,0,217,0,137,0,43,0,139,0,108,0,97,0,36,0,220,0,134,0,79,0,91,0,92,0,145,0,128,0,58,0,0,0,128,0,0,0,27,0,38,0,243,0,37,0,78,0,88,0,188,0,205,0,150,0,220,0,9,0,162,0,20,0,65,0,105,0,203,0,0,0,172,0,0,0,81,0,117,0,47,0,160,0,223,0,211,0,213,0,100,0,207,0,0,0,202,0,204,0,216,0,195,0,243,0,157,0,0,0,137,0,237,0,10,0,220,0,10,0,176,0,81,0,0,0,61,0,180,0,33,0,43,0,99,0,74,0,226,0,112,0,154,0,221,0,118,0,21,0,167,0,46,0,121,0,46,0,133,0,14,0,0,0,86,0,0,0,121,0,100,0,60,0,0,0,120,0,63,0,27,0,0,0,252,0,190,0,86,0,99,0,191,0,20,0,0,0,2,0,92,0,0,0,234,0,179,0,177,0,127,0,11,0,230,0,166,0,70,0,244,0,240,0,146,0,26,0,86,0,174,0,0,0,81,0,122,0,20,0,0,0,44,0,71,0,241,0,164,0,128,0,158,0,176,0,0,0,117,0,110,0,186,0,66,0,0,0,253,0,223,0,54,0,122,0,13,0,0,0,252,0,32,0,4,0,13,0,127,0,0,0,0,0,0,0,86,0,93,0,0,0,225,0,0,0,0,0,19,0,136,0,13,0,203,0,0,0,0,0,4,0,0,0,0,0,0,0,115,0,248,0,0,0,199,0,30,0,65,0,185,0,18,0,0,0,218,0,111,0,113,0,0,0,178,0,107,0,236,0,122,0,126,0,35,0,43,0,178,0,0,0,94,0,172,0,21,0,196,0,243,0,58,0,126,0,52,0,232,0,0,0,72,0,0,0,120,0,148,0,37,0,210,0,59,0,105,0,241,0);
signal scenario_full  : scenario_type := (6,31,147,31,115,31,211,31,134,31,155,31,195,31,195,30,195,29,237,31,199,31,8,31,255,31,96,31,59,31,179,31,72,31,72,30,238,31,254,31,62,31,34,31,92,31,112,31,39,31,238,31,238,30,238,29,238,28,9,31,164,31,164,30,49,31,10,31,174,31,44,31,231,31,59,31,60,31,3,31,32,31,139,31,183,31,78,31,247,31,247,30,148,31,107,31,182,31,38,31,183,31,58,31,58,30,58,29,159,31,159,30,10,31,97,31,117,31,167,31,167,30,104,31,104,31,220,31,182,31,111,31,83,31,122,31,4,31,150,31,245,31,245,30,146,31,83,31,119,31,67,31,200,31,36,31,15,31,72,31,137,31,137,30,213,31,49,31,132,31,5,31,224,31,224,30,200,31,3,31,187,31,10,31,163,31,66,31,148,31,218,31,55,31,62,31,158,31,161,31,40,31,128,31,122,31,191,31,96,31,124,31,124,30,63,31,103,31,71,31,33,31,12,31,36,31,17,31,17,30,17,31,17,30,114,31,121,31,121,30,245,31,225,31,225,30,107,31,214,31,214,30,39,31,39,30,39,29,246,31,246,30,110,31,1,31,116,31,116,30,253,31,206,31,87,31,195,31,173,31,83,31,233,31,160,31,160,30,98,31,98,30,198,31,198,30,92,31,92,30,78,31,212,31,212,30,118,31,118,30,246,31,62,31,34,31,34,31,136,31,133,31,133,30,186,31,250,31,214,31,24,31,245,31,245,30,148,31,120,31,120,30,65,31,65,30,253,31,253,30,159,31,103,31,200,31,166,31,187,31,187,30,236,31,236,30,179,31,179,30,194,31,42,31,56,31,181,31,247,31,247,30,46,31,194,31,149,31,108,31,95,31,202,31,255,31,239,31,64,31,190,31,149,31,69,31,99,31,99,30,99,31,185,31,53,31,35,31,139,31,124,31,243,31,243,30,5,31,131,31,242,31,17,31,139,31,193,31,11,31,58,31,87,31,137,31,36,31,222,31,104,31,46,31,185,31,107,31,107,30,252,31,92,31,241,31,45,31,48,31,115,31,229,31,12,31,85,31,6,31,157,31,20,31,37,31,140,31,140,30,185,31,209,31,209,30,209,29,190,31,145,31,41,31,135,31,244,31,155,31,242,31,141,31,221,31,221,30,195,31,235,31,235,30,92,31,92,30,248,31,135,31,239,31,239,30,179,31,186,31,43,31,72,31,16,31,16,30,92,31,47,31,57,31,240,31,16,31,135,31,133,31,133,30,133,29,203,31,212,31,62,31,62,30,156,31,192,31,218,31,180,31,171,31,5,31,143,31,143,30,185,31,74,31,74,30,124,31,183,31,183,30,36,31,75,31,146,31,219,31,88,31,137,31,2,31,172,31,250,31,236,31,226,31,52,31,89,31,88,31,110,31,105,31,221,31,249,31,202,31,170,31,170,30,2,31,225,31,225,30,181,31,74,31,86,31,145,31,232,31,154,31,186,31,132,31,93,31,194,31,34,31,19,31,212,31,212,30,13,31,13,30,213,31,62,31,62,30,122,31,158,31,194,31,186,31,104,31,214,31,199,31,65,31,229,31,225,31,243,31,243,30,162,31,175,31,230,31,122,31,50,31,50,30,50,29,238,31,51,31,51,30,51,29,192,31,52,31,123,31,123,30,243,31,218,31,98,31,98,30,81,31,36,31,156,31,218,31,82,31,214,31,203,31,160,31,222,31,79,31,182,31,112,31,65,31,40,31,138,31,138,30,68,31,119,31,177,31,197,31,156,31,1,31,168,31,103,31,103,30,103,29,126,31,126,30,200,31,101,31,95,31,118,31,119,31,133,31,133,30,200,31,22,31,22,30,199,31,199,30,125,31,125,30,125,29,146,31,133,31,55,31,161,31,213,31,213,30,64,31,64,30,64,29,64,28,41,31,43,31,43,30,111,31,144,31,13,31,243,31,219,31,68,31,117,31,56,31,53,31,123,31,143,31,143,30,143,29,143,28,182,31,108,31,7,31,29,31,65,31,65,30,32,31,80,31,80,30,88,31,88,30,93,31,93,30,50,31,103,31,243,31,162,31,193,31,193,30,3,31,3,30,59,31,212,31,145,31,145,30,226,31,173,31,182,31,182,30,182,29,12,31,12,30,127,31,215,31,69,31,18,31,183,31,19,31,225,31,225,30,93,31,227,31,79,31,159,31,6,31,135,31,107,31,89,31,190,31,242,31,242,30,200,31,198,31,177,31,245,31,20,31,41,31,174,31,174,30,198,31,198,30,106,31,250,31,161,31,199,31,176,31,176,30,176,29,80,31,74,31,31,31,123,31,111,31,160,31,10,31,139,31,139,30,217,31,137,31,43,31,139,31,108,31,97,31,36,31,220,31,134,31,79,31,91,31,92,31,145,31,128,31,58,31,58,30,128,31,128,30,27,31,38,31,243,31,37,31,78,31,88,31,188,31,205,31,150,31,220,31,9,31,162,31,20,31,65,31,105,31,203,31,203,30,172,31,172,30,81,31,117,31,47,31,160,31,223,31,211,31,213,31,100,31,207,31,207,30,202,31,204,31,216,31,195,31,243,31,157,31,157,30,137,31,237,31,10,31,220,31,10,31,176,31,81,31,81,30,61,31,180,31,33,31,43,31,99,31,74,31,226,31,112,31,154,31,221,31,118,31,21,31,167,31,46,31,121,31,46,31,133,31,14,31,14,30,86,31,86,30,121,31,100,31,60,31,60,30,120,31,63,31,27,31,27,30,252,31,190,31,86,31,99,31,191,31,20,31,20,30,2,31,92,31,92,30,234,31,179,31,177,31,127,31,11,31,230,31,166,31,70,31,244,31,240,31,146,31,26,31,86,31,174,31,174,30,81,31,122,31,20,31,20,30,44,31,71,31,241,31,164,31,128,31,158,31,176,31,176,30,117,31,110,31,186,31,66,31,66,30,253,31,223,31,54,31,122,31,13,31,13,30,252,31,32,31,4,31,13,31,127,31,127,30,127,29,127,28,86,31,93,31,93,30,225,31,225,30,225,29,19,31,136,31,13,31,203,31,203,30,203,29,4,31,4,30,4,29,4,28,115,31,248,31,248,30,199,31,30,31,65,31,185,31,18,31,18,30,218,31,111,31,113,31,113,30,178,31,107,31,236,31,122,31,126,31,35,31,43,31,178,31,178,30,94,31,172,31,21,31,196,31,243,31,58,31,126,31,52,31,232,31,232,30,72,31,72,30,120,31,148,31,37,31,210,31,59,31,105,31,241,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
