-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 896;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (215,0,0,0,205,0,79,0,130,0,83,0,45,0,248,0,30,0,0,0,175,0,69,0,107,0,234,0,128,0,22,0,0,0,0,0,6,0,133,0,213,0,7,0,222,0,91,0,231,0,62,0,32,0,143,0,0,0,0,0,28,0,60,0,0,0,13,0,121,0,255,0,208,0,240,0,69,0,123,0,184,0,85,0,0,0,58,0,170,0,117,0,28,0,220,0,10,0,183,0,66,0,236,0,101,0,6,0,234,0,166,0,21,0,0,0,165,0,3,0,199,0,158,0,78,0,84,0,160,0,217,0,0,0,180,0,53,0,12,0,89,0,247,0,90,0,109,0,231,0,0,0,226,0,184,0,53,0,7,0,0,0,0,0,212,0,135,0,21,0,243,0,150,0,232,0,20,0,215,0,209,0,207,0,59,0,32,0,206,0,0,0,200,0,224,0,163,0,54,0,92,0,39,0,102,0,40,0,27,0,130,0,96,0,71,0,180,0,92,0,0,0,154,0,0,0,82,0,171,0,175,0,195,0,125,0,56,0,116,0,0,0,116,0,22,0,50,0,0,0,144,0,0,0,49,0,238,0,63,0,0,0,25,0,184,0,209,0,8,0,0,0,69,0,11,0,131,0,0,0,68,0,0,0,234,0,0,0,168,0,15,0,29,0,248,0,238,0,135,0,0,0,221,0,129,0,70,0,134,0,0,0,0,0,197,0,186,0,15,0,9,0,34,0,0,0,44,0,189,0,126,0,0,0,136,0,115,0,0,0,159,0,208,0,64,0,0,0,137,0,235,0,21,0,0,0,93,0,0,0,223,0,0,0,190,0,0,0,170,0,239,0,168,0,0,0,89,0,111,0,235,0,14,0,0,0,13,0,242,0,246,0,0,0,186,0,241,0,235,0,110,0,206,0,38,0,183,0,108,0,103,0,7,0,108,0,243,0,92,0,249,0,238,0,0,0,181,0,220,0,0,0,129,0,85,0,77,0,173,0,0,0,228,0,149,0,66,0,13,0,213,0,200,0,35,0,0,0,0,0,92,0,156,0,113,0,245,0,41,0,199,0,23,0,13,0,109,0,147,0,117,0,0,0,253,0,170,0,63,0,76,0,0,0,125,0,0,0,56,0,0,0,226,0,90,0,250,0,169,0,253,0,13,0,248,0,0,0,85,0,71,0,156,0,205,0,152,0,148,0,76,0,0,0,131,0,253,0,182,0,69,0,0,0,251,0,29,0,0,0,47,0,240,0,166,0,219,0,123,0,217,0,92,0,52,0,171,0,153,0,0,0,49,0,211,0,27,0,196,0,0,0,110,0,148,0,98,0,128,0,126,0,130,0,214,0,203,0,121,0,189,0,140,0,234,0,227,0,0,0,199,0,12,0,32,0,226,0,66,0,176,0,134,0,162,0,168,0,120,0,251,0,186,0,170,0,246,0,65,0,85,0,119,0,0,0,24,0,134,0,200,0,224,0,166,0,18,0,52,0,140,0,87,0,0,0,0,0,91,0,44,0,0,0,0,0,57,0,64,0,77,0,0,0,253,0,116,0,255,0,41,0,108,0,117,0,0,0,92,0,11,0,172,0,119,0,27,0,111,0,17,0,2,0,159,0,226,0,71,0,119,0,13,0,0,0,0,0,151,0,129,0,24,0,174,0,158,0,105,0,220,0,0,0,170,0,85,0,170,0,0,0,212,0,0,0,188,0,202,0,106,0,44,0,120,0,129,0,0,0,5,0,126,0,245,0,17,0,0,0,246,0,181,0,0,0,0,0,6,0,45,0,131,0,114,0,116,0,0,0,216,0,52,0,0,0,24,0,43,0,7,0,83,0,0,0,71,0,124,0,3,0,36,0,128,0,234,0,235,0,188,0,9,0,234,0,93,0,222,0,0,0,203,0,216,0,62,0,106,0,165,0,134,0,227,0,0,0,30,0,25,0,49,0,221,0,44,0,0,0,0,0,135,0,121,0,137,0,0,0,130,0,219,0,169,0,0,0,247,0,193,0,97,0,111,0,70,0,96,0,179,0,97,0,23,0,206,0,253,0,153,0,43,0,144,0,0,0,255,0,247,0,253,0,65,0,0,0,210,0,249,0,152,0,178,0,0,0,126,0,58,0,212,0,43,0,204,0,235,0,149,0,83,0,0,0,189,0,0,0,151,0,116,0,112,0,214,0,162,0,105,0,144,0,139,0,26,0,0,0,103,0,143,0,0,0,229,0,231,0,250,0,205,0,34,0,59,0,174,0,245,0,0,0,102,0,115,0,92,0,169,0,134,0,60,0,143,0,56,0,236,0,103,0,122,0,160,0,218,0,167,0,37,0,230,0,0,0,26,0,0,0,165,0,232,0,144,0,218,0,0,0,122,0,0,0,234,0,84,0,219,0,160,0,200,0,206,0,37,0,33,0,8,0,148,0,53,0,118,0,162,0,55,0,167,0,185,0,9,0,253,0,166,0,0,0,25,0,121,0,135,0,41,0,0,0,173,0,17,0,229,0,224,0,184,0,29,0,175,0,0,0,74,0,8,0,229,0,179,0,255,0,69,0,255,0,206,0,10,0,97,0,236,0,0,0,142,0,118,0,165,0,70,0,63,0,171,0,34,0,48,0,18,0,250,0,137,0,216,0,0,0,8,0,88,0,147,0,8,0,148,0,0,0,0,0,0,0,187,0,31,0,255,0,114,0,15,0,181,0,220,0,129,0,138,0,103,0,38,0,119,0,85,0,205,0,152,0,186,0,94,0,9,0,0,0,45,0,129,0,132,0,0,0,130,0,84,0,22,0,232,0,26,0,244,0,0,0,74,0,241,0,20,0,228,0,65,0,0,0,238,0,44,0,61,0,151,0,0,0,31,0,196,0,138,0,59,0,241,0,202,0,113,0,216,0,247,0,69,0,72,0,0,0,105,0,0,0,0,0,46,0,0,0,121,0,238,0,188,0,85,0,0,0,106,0,51,0,0,0,188,0,153,0,75,0,179,0,84,0,222,0,58,0,0,0,44,0,101,0,23,0,0,0,135,0,0,0,84,0,101,0,184,0,132,0,0,0,148,0,65,0,170,0,204,0,29,0,71,0,0,0,228,0,165,0,67,0,128,0,238,0,186,0,162,0,182,0,30,0,161,0,183,0,180,0,161,0,162,0,72,0,93,0,0,0,87,0,0,0,108,0,0,0,0,0,50,0,109,0,34,0,165,0,177,0,240,0,0,0,251,0,49,0,207,0,194,0,160,0,32,0,104,0,137,0,76,0,142,0,46,0,52,0,244,0,0,0,161,0,0,0,210,0,0,0,56,0,137,0,57,0,126,0,28,0,0,0,125,0,0,0,198,0,250,0,0,0,47,0,0,0,0,0,184,0,0,0,59,0,214,0,157,0,0,0,75,0,38,0,52,0,0,0,217,0,250,0,2,0,7,0,22,0,11,0,59,0,0,0,158,0,180,0,110,0,37,0,0,0,41,0,209,0,133,0,197,0,0,0,20,0,21,0,199,0,40,0,0,0,119,0,213,0,86,0,219,0,0,0,151,0,198,0,213,0,232,0,157,0,0,0,181,0,52,0,35,0,188,0,196,0,71,0,102,0,0,0,69,0,40,0,99,0,244,0,32,0,40,0,89,0,49,0,0,0,222,0,138,0,189,0,0,0,148,0,116,0,132,0,145,0,86,0,0,0,213,0,62,0,118,0,51,0,128,0,9,0,154,0,27,0,0,0,21,0,0,0,89,0,0,0,187,0,193,0,186,0,223,0,186,0,134,0,58,0,101,0,0,0,115,0,154,0,242,0,138,0,185,0,46,0,7,0,173,0,120,0,241,0,116,0,0,0,153,0,199,0,29,0,217,0,116,0,0,0,0,0,223,0,34,0,129,0,152,0,0,0,0,0,194,0,220,0,0,0,203,0,161,0,145,0,20,0,0,0,26,0,180,0,225,0,198,0,112,0,227,0,0,0,51,0,213,0,0,0,42,0,78,0,229,0,0,0,0,0,106,0,212,0,135,0,179,0,109,0,136,0,0,0,43,0);
signal scenario_full  : scenario_type := (215,31,215,30,205,31,79,31,130,31,83,31,45,31,248,31,30,31,30,30,175,31,69,31,107,31,234,31,128,31,22,31,22,30,22,29,6,31,133,31,213,31,7,31,222,31,91,31,231,31,62,31,32,31,143,31,143,30,143,29,28,31,60,31,60,30,13,31,121,31,255,31,208,31,240,31,69,31,123,31,184,31,85,31,85,30,58,31,170,31,117,31,28,31,220,31,10,31,183,31,66,31,236,31,101,31,6,31,234,31,166,31,21,31,21,30,165,31,3,31,199,31,158,31,78,31,84,31,160,31,217,31,217,30,180,31,53,31,12,31,89,31,247,31,90,31,109,31,231,31,231,30,226,31,184,31,53,31,7,31,7,30,7,29,212,31,135,31,21,31,243,31,150,31,232,31,20,31,215,31,209,31,207,31,59,31,32,31,206,31,206,30,200,31,224,31,163,31,54,31,92,31,39,31,102,31,40,31,27,31,130,31,96,31,71,31,180,31,92,31,92,30,154,31,154,30,82,31,171,31,175,31,195,31,125,31,56,31,116,31,116,30,116,31,22,31,50,31,50,30,144,31,144,30,49,31,238,31,63,31,63,30,25,31,184,31,209,31,8,31,8,30,69,31,11,31,131,31,131,30,68,31,68,30,234,31,234,30,168,31,15,31,29,31,248,31,238,31,135,31,135,30,221,31,129,31,70,31,134,31,134,30,134,29,197,31,186,31,15,31,9,31,34,31,34,30,44,31,189,31,126,31,126,30,136,31,115,31,115,30,159,31,208,31,64,31,64,30,137,31,235,31,21,31,21,30,93,31,93,30,223,31,223,30,190,31,190,30,170,31,239,31,168,31,168,30,89,31,111,31,235,31,14,31,14,30,13,31,242,31,246,31,246,30,186,31,241,31,235,31,110,31,206,31,38,31,183,31,108,31,103,31,7,31,108,31,243,31,92,31,249,31,238,31,238,30,181,31,220,31,220,30,129,31,85,31,77,31,173,31,173,30,228,31,149,31,66,31,13,31,213,31,200,31,35,31,35,30,35,29,92,31,156,31,113,31,245,31,41,31,199,31,23,31,13,31,109,31,147,31,117,31,117,30,253,31,170,31,63,31,76,31,76,30,125,31,125,30,56,31,56,30,226,31,90,31,250,31,169,31,253,31,13,31,248,31,248,30,85,31,71,31,156,31,205,31,152,31,148,31,76,31,76,30,131,31,253,31,182,31,69,31,69,30,251,31,29,31,29,30,47,31,240,31,166,31,219,31,123,31,217,31,92,31,52,31,171,31,153,31,153,30,49,31,211,31,27,31,196,31,196,30,110,31,148,31,98,31,128,31,126,31,130,31,214,31,203,31,121,31,189,31,140,31,234,31,227,31,227,30,199,31,12,31,32,31,226,31,66,31,176,31,134,31,162,31,168,31,120,31,251,31,186,31,170,31,246,31,65,31,85,31,119,31,119,30,24,31,134,31,200,31,224,31,166,31,18,31,52,31,140,31,87,31,87,30,87,29,91,31,44,31,44,30,44,29,57,31,64,31,77,31,77,30,253,31,116,31,255,31,41,31,108,31,117,31,117,30,92,31,11,31,172,31,119,31,27,31,111,31,17,31,2,31,159,31,226,31,71,31,119,31,13,31,13,30,13,29,151,31,129,31,24,31,174,31,158,31,105,31,220,31,220,30,170,31,85,31,170,31,170,30,212,31,212,30,188,31,202,31,106,31,44,31,120,31,129,31,129,30,5,31,126,31,245,31,17,31,17,30,246,31,181,31,181,30,181,29,6,31,45,31,131,31,114,31,116,31,116,30,216,31,52,31,52,30,24,31,43,31,7,31,83,31,83,30,71,31,124,31,3,31,36,31,128,31,234,31,235,31,188,31,9,31,234,31,93,31,222,31,222,30,203,31,216,31,62,31,106,31,165,31,134,31,227,31,227,30,30,31,25,31,49,31,221,31,44,31,44,30,44,29,135,31,121,31,137,31,137,30,130,31,219,31,169,31,169,30,247,31,193,31,97,31,111,31,70,31,96,31,179,31,97,31,23,31,206,31,253,31,153,31,43,31,144,31,144,30,255,31,247,31,253,31,65,31,65,30,210,31,249,31,152,31,178,31,178,30,126,31,58,31,212,31,43,31,204,31,235,31,149,31,83,31,83,30,189,31,189,30,151,31,116,31,112,31,214,31,162,31,105,31,144,31,139,31,26,31,26,30,103,31,143,31,143,30,229,31,231,31,250,31,205,31,34,31,59,31,174,31,245,31,245,30,102,31,115,31,92,31,169,31,134,31,60,31,143,31,56,31,236,31,103,31,122,31,160,31,218,31,167,31,37,31,230,31,230,30,26,31,26,30,165,31,232,31,144,31,218,31,218,30,122,31,122,30,234,31,84,31,219,31,160,31,200,31,206,31,37,31,33,31,8,31,148,31,53,31,118,31,162,31,55,31,167,31,185,31,9,31,253,31,166,31,166,30,25,31,121,31,135,31,41,31,41,30,173,31,17,31,229,31,224,31,184,31,29,31,175,31,175,30,74,31,8,31,229,31,179,31,255,31,69,31,255,31,206,31,10,31,97,31,236,31,236,30,142,31,118,31,165,31,70,31,63,31,171,31,34,31,48,31,18,31,250,31,137,31,216,31,216,30,8,31,88,31,147,31,8,31,148,31,148,30,148,29,148,28,187,31,31,31,255,31,114,31,15,31,181,31,220,31,129,31,138,31,103,31,38,31,119,31,85,31,205,31,152,31,186,31,94,31,9,31,9,30,45,31,129,31,132,31,132,30,130,31,84,31,22,31,232,31,26,31,244,31,244,30,74,31,241,31,20,31,228,31,65,31,65,30,238,31,44,31,61,31,151,31,151,30,31,31,196,31,138,31,59,31,241,31,202,31,113,31,216,31,247,31,69,31,72,31,72,30,105,31,105,30,105,29,46,31,46,30,121,31,238,31,188,31,85,31,85,30,106,31,51,31,51,30,188,31,153,31,75,31,179,31,84,31,222,31,58,31,58,30,44,31,101,31,23,31,23,30,135,31,135,30,84,31,101,31,184,31,132,31,132,30,148,31,65,31,170,31,204,31,29,31,71,31,71,30,228,31,165,31,67,31,128,31,238,31,186,31,162,31,182,31,30,31,161,31,183,31,180,31,161,31,162,31,72,31,93,31,93,30,87,31,87,30,108,31,108,30,108,29,50,31,109,31,34,31,165,31,177,31,240,31,240,30,251,31,49,31,207,31,194,31,160,31,32,31,104,31,137,31,76,31,142,31,46,31,52,31,244,31,244,30,161,31,161,30,210,31,210,30,56,31,137,31,57,31,126,31,28,31,28,30,125,31,125,30,198,31,250,31,250,30,47,31,47,30,47,29,184,31,184,30,59,31,214,31,157,31,157,30,75,31,38,31,52,31,52,30,217,31,250,31,2,31,7,31,22,31,11,31,59,31,59,30,158,31,180,31,110,31,37,31,37,30,41,31,209,31,133,31,197,31,197,30,20,31,21,31,199,31,40,31,40,30,119,31,213,31,86,31,219,31,219,30,151,31,198,31,213,31,232,31,157,31,157,30,181,31,52,31,35,31,188,31,196,31,71,31,102,31,102,30,69,31,40,31,99,31,244,31,32,31,40,31,89,31,49,31,49,30,222,31,138,31,189,31,189,30,148,31,116,31,132,31,145,31,86,31,86,30,213,31,62,31,118,31,51,31,128,31,9,31,154,31,27,31,27,30,21,31,21,30,89,31,89,30,187,31,193,31,186,31,223,31,186,31,134,31,58,31,101,31,101,30,115,31,154,31,242,31,138,31,185,31,46,31,7,31,173,31,120,31,241,31,116,31,116,30,153,31,199,31,29,31,217,31,116,31,116,30,116,29,223,31,34,31,129,31,152,31,152,30,152,29,194,31,220,31,220,30,203,31,161,31,145,31,20,31,20,30,26,31,180,31,225,31,198,31,112,31,227,31,227,30,51,31,213,31,213,30,42,31,78,31,229,31,229,30,229,29,106,31,212,31,135,31,179,31,109,31,136,31,136,30,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
