-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_789 is
end project_tb_789;

architecture project_tb_arch_789 of project_tb_789 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 986;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (47,0,0,0,46,0,198,0,47,0,84,0,165,0,194,0,157,0,57,0,208,0,81,0,253,0,68,0,50,0,110,0,45,0,88,0,155,0,216,0,48,0,19,0,223,0,107,0,193,0,242,0,22,0,0,0,0,0,0,0,229,0,0,0,171,0,0,0,0,0,0,0,77,0,19,0,90,0,186,0,29,0,49,0,0,0,212,0,100,0,225,0,251,0,106,0,237,0,0,0,237,0,188,0,220,0,54,0,133,0,239,0,186,0,0,0,247,0,183,0,117,0,82,0,0,0,0,0,242,0,74,0,0,0,45,0,43,0,149,0,186,0,217,0,198,0,113,0,88,0,25,0,169,0,182,0,0,0,172,0,0,0,93,0,91,0,0,0,116,0,125,0,131,0,190,0,85,0,70,0,31,0,214,0,113,0,0,0,47,0,79,0,229,0,0,0,143,0,160,0,0,0,62,0,149,0,78,0,236,0,221,0,100,0,167,0,0,0,0,0,146,0,49,0,0,0,0,0,54,0,47,0,0,0,34,0,66,0,0,0,79,0,254,0,112,0,231,0,110,0,20,0,224,0,243,0,70,0,83,0,117,0,10,0,163,0,0,0,0,0,184,0,238,0,249,0,95,0,32,0,27,0,208,0,208,0,213,0,205,0,247,0,0,0,36,0,9,0,149,0,105,0,189,0,0,0,55,0,204,0,0,0,247,0,170,0,0,0,205,0,184,0,67,0,205,0,198,0,0,0,43,0,105,0,249,0,225,0,243,0,201,0,0,0,62,0,49,0,123,0,65,0,233,0,108,0,15,0,224,0,186,0,193,0,2,0,134,0,62,0,221,0,52,0,0,0,249,0,80,0,0,0,7,0,162,0,0,0,164,0,244,0,123,0,139,0,12,0,111,0,0,0,176,0,0,0,31,0,179,0,46,0,7,0,0,0,98,0,155,0,141,0,131,0,147,0,195,0,135,0,231,0,198,0,0,0,241,0,0,0,0,0,0,0,140,0,97,0,220,0,71,0,181,0,234,0,156,0,0,0,158,0,213,0,78,0,0,0,196,0,0,0,153,0,0,0,0,0,25,0,119,0,130,0,144,0,203,0,0,0,145,0,133,0,170,0,95,0,254,0,0,0,77,0,36,0,71,0,214,0,0,0,0,0,76,0,78,0,62,0,218,0,40,0,0,0,101,0,220,0,152,0,125,0,136,0,229,0,101,0,0,0,0,0,69,0,0,0,59,0,63,0,253,0,9,0,236,0,252,0,235,0,0,0,245,0,0,0,203,0,9,0,199,0,59,0,0,0,0,0,236,0,21,0,0,0,163,0,244,0,182,0,207,0,0,0,41,0,0,0,152,0,116,0,0,0,193,0,83,0,108,0,174,0,109,0,25,0,38,0,203,0,98,0,0,0,219,0,134,0,0,0,0,0,87,0,25,0,93,0,0,0,152,0,230,0,252,0,182,0,243,0,207,0,193,0,0,0,70,0,83,0,0,0,73,0,0,0,195,0,72,0,138,0,151,0,111,0,43,0,12,0,0,0,101,0,251,0,27,0,253,0,140,0,111,0,207,0,0,0,227,0,22,0,39,0,254,0,39,0,206,0,0,0,65,0,190,0,221,0,184,0,0,0,0,0,123,0,95,0,171,0,0,0,134,0,87,0,0,0,0,0,176,0,0,0,39,0,142,0,249,0,0,0,79,0,94,0,59,0,102,0,143,0,68,0,157,0,134,0,218,0,140,0,111,0,4,0,37,0,211,0,191,0,87,0,19,0,154,0,148,0,193,0,43,0,104,0,204,0,133,0,136,0,0,0,198,0,0,0,54,0,207,0,109,0,0,0,0,0,0,0,13,0,191,0,29,0,118,0,0,0,240,0,138,0,120,0,206,0,7,0,0,0,231,0,79,0,76,0,58,0,13,0,0,0,97,0,170,0,135,0,0,0,6,0,0,0,208,0,242,0,238,0,0,0,163,0,48,0,150,0,0,0,61,0,85,0,36,0,0,0,218,0,145,0,184,0,0,0,11,0,51,0,94,0,132,0,59,0,219,0,237,0,156,0,87,0,238,0,199,0,0,0,213,0,130,0,0,0,54,0,147,0,200,0,213,0,0,0,203,0,0,0,138,0,19,0,206,0,200,0,155,0,0,0,188,0,97,0,128,0,136,0,44,0,70,0,172,0,88,0,224,0,156,0,43,0,146,0,229,0,0,0,103,0,0,0,27,0,161,0,61,0,0,0,89,0,187,0,0,0,50,0,143,0,4,0,68,0,47,0,155,0,32,0,0,0,125,0,67,0,0,0,213,0,0,0,170,0,190,0,0,0,242,0,229,0,138,0,21,0,245,0,158,0,11,0,10,0,106,0,252,0,125,0,0,0,34,0,80,0,0,0,203,0,0,0,89,0,0,0,62,0,0,0,171,0,211,0,117,0,204,0,185,0,0,0,46,0,0,0,0,0,2,0,233,0,0,0,87,0,62,0,176,0,31,0,0,0,0,0,73,0,68,0,30,0,72,0,3,0,22,0,172,0,33,0,0,0,177,0,203,0,33,0,118,0,140,0,164,0,1,0,104,0,119,0,177,0,153,0,0,0,244,0,176,0,145,0,40,0,0,0,170,0,181,0,247,0,0,0,0,0,0,0,112,0,32,0,217,0,161,0,0,0,0,0,0,0,92,0,26,0,0,0,127,0,232,0,1,0,0,0,0,0,158,0,43,0,59,0,184,0,14,0,77,0,76,0,12,0,0,0,181,0,236,0,0,0,20,0,241,0,87,0,123,0,229,0,151,0,217,0,182,0,0,0,187,0,2,0,0,0,164,0,0,0,49,0,79,0,199,0,111,0,0,0,0,0,252,0,20,0,0,0,112,0,246,0,0,0,94,0,12,0,89,0,215,0,0,0,148,0,193,0,6,0,39,0,209,0,18,0,236,0,200,0,147,0,14,0,166,0,183,0,210,0,23,0,0,0,198,0,232,0,140,0,238,0,175,0,11,0,81,0,39,0,197,0,161,0,186,0,165,0,47,0,165,0,0,0,7,0,136,0,108,0,29,0,98,0,63,0,110,0,192,0,100,0,139,0,124,0,13,0,244,0,89,0,251,0,0,0,0,0,27,0,35,0,225,0,80,0,221,0,22,0,177,0,38,0,203,0,0,0,152,0,4,0,0,0,252,0,0,0,28,0,195,0,203,0,112,0,0,0,202,0,0,0,144,0,226,0,173,0,43,0,186,0,0,0,35,0,0,0,127,0,247,0,155,0,175,0,27,0,0,0,30,0,115,0,39,0,0,0,67,0,60,0,0,0,192,0,50,0,141,0,235,0,90,0,202,0,237,0,69,0,247,0,161,0,203,0,25,0,76,0,129,0,73,0,100,0,202,0,49,0,81,0,207,0,95,0,196,0,0,0,0,0,20,0,0,0,185,0,255,0,80,0,0,0,131,0,0,0,201,0,68,0,105,0,144,0,97,0,8,0,102,0,71,0,218,0,0,0,215,0,126,0,110,0,114,0,156,0,6,0,140,0,102,0,108,0,91,0,0,0,185,0,157,0,128,0,0,0,144,0,195,0,190,0,0,0,179,0,110,0,0,0,19,0,0,0,0,0,105,0,217,0,7,0,173,0,131,0,73,0,174,0,218,0,37,0,218,0,161,0,41,0,30,0,0,0,77,0,1,0,37,0,45,0,110,0,164,0,30,0,33,0,225,0,0,0,197,0,216,0,0,0,100,0,99,0,108,0,230,0,0,0,26,0,33,0,5,0,0,0,111,0,50,0,93,0,14,0,219,0,53,0,137,0,20,0,94,0,0,0,0,0,184,0,0,0,0,0,145,0,245,0,246,0,21,0,0,0,198,0,68,0,0,0,234,0,143,0,245,0,202,0,54,0,164,0,110,0,53,0,30,0,41,0,78,0,154,0,0,0,249,0,40,0,0,0,78,0,0,0,140,0,156,0,161,0,20,0,102,0,183,0,107,0,100,0,250,0,0,0,144,0,180,0,230,0,220,0,31,0,43,0,155,0,0,0,55,0,246,0,90,0,0,0,0,0,0,0,225,0,13,0,129,0,248,0,66,0,23,0,108,0,9,0,0,0,232,0,0,0,41,0,241,0,248,0,126,0,238,0,248,0,224,0,101,0,196,0,42,0,16,0,0,0,0,0,182,0,1,0,122,0,69,0,0,0,0,0,209,0,31,0,18,0,45,0,3,0,28,0,233,0,0,0,137,0,210,0,0,0,0,0,175,0,13,0,241,0,176,0,57,0,76,0,0,0,177,0,189,0,0,0,60,0,141,0,0,0,170,0,0,0,0,0,114,0,134,0,0,0,20,0,68,0,142,0,200,0,129,0,148,0,168,0,48,0,141,0,2,0,189,0,61,0,188,0,109,0,187,0,111,0,179,0,82,0,109,0,8,0,193,0,0,0);
signal scenario_full  : scenario_type := (47,31,47,30,46,31,198,31,47,31,84,31,165,31,194,31,157,31,57,31,208,31,81,31,253,31,68,31,50,31,110,31,45,31,88,31,155,31,216,31,48,31,19,31,223,31,107,31,193,31,242,31,22,31,22,30,22,29,22,28,229,31,229,30,171,31,171,30,171,29,171,28,77,31,19,31,90,31,186,31,29,31,49,31,49,30,212,31,100,31,225,31,251,31,106,31,237,31,237,30,237,31,188,31,220,31,54,31,133,31,239,31,186,31,186,30,247,31,183,31,117,31,82,31,82,30,82,29,242,31,74,31,74,30,45,31,43,31,149,31,186,31,217,31,198,31,113,31,88,31,25,31,169,31,182,31,182,30,172,31,172,30,93,31,91,31,91,30,116,31,125,31,131,31,190,31,85,31,70,31,31,31,214,31,113,31,113,30,47,31,79,31,229,31,229,30,143,31,160,31,160,30,62,31,149,31,78,31,236,31,221,31,100,31,167,31,167,30,167,29,146,31,49,31,49,30,49,29,54,31,47,31,47,30,34,31,66,31,66,30,79,31,254,31,112,31,231,31,110,31,20,31,224,31,243,31,70,31,83,31,117,31,10,31,163,31,163,30,163,29,184,31,238,31,249,31,95,31,32,31,27,31,208,31,208,31,213,31,205,31,247,31,247,30,36,31,9,31,149,31,105,31,189,31,189,30,55,31,204,31,204,30,247,31,170,31,170,30,205,31,184,31,67,31,205,31,198,31,198,30,43,31,105,31,249,31,225,31,243,31,201,31,201,30,62,31,49,31,123,31,65,31,233,31,108,31,15,31,224,31,186,31,193,31,2,31,134,31,62,31,221,31,52,31,52,30,249,31,80,31,80,30,7,31,162,31,162,30,164,31,244,31,123,31,139,31,12,31,111,31,111,30,176,31,176,30,31,31,179,31,46,31,7,31,7,30,98,31,155,31,141,31,131,31,147,31,195,31,135,31,231,31,198,31,198,30,241,31,241,30,241,29,241,28,140,31,97,31,220,31,71,31,181,31,234,31,156,31,156,30,158,31,213,31,78,31,78,30,196,31,196,30,153,31,153,30,153,29,25,31,119,31,130,31,144,31,203,31,203,30,145,31,133,31,170,31,95,31,254,31,254,30,77,31,36,31,71,31,214,31,214,30,214,29,76,31,78,31,62,31,218,31,40,31,40,30,101,31,220,31,152,31,125,31,136,31,229,31,101,31,101,30,101,29,69,31,69,30,59,31,63,31,253,31,9,31,236,31,252,31,235,31,235,30,245,31,245,30,203,31,9,31,199,31,59,31,59,30,59,29,236,31,21,31,21,30,163,31,244,31,182,31,207,31,207,30,41,31,41,30,152,31,116,31,116,30,193,31,83,31,108,31,174,31,109,31,25,31,38,31,203,31,98,31,98,30,219,31,134,31,134,30,134,29,87,31,25,31,93,31,93,30,152,31,230,31,252,31,182,31,243,31,207,31,193,31,193,30,70,31,83,31,83,30,73,31,73,30,195,31,72,31,138,31,151,31,111,31,43,31,12,31,12,30,101,31,251,31,27,31,253,31,140,31,111,31,207,31,207,30,227,31,22,31,39,31,254,31,39,31,206,31,206,30,65,31,190,31,221,31,184,31,184,30,184,29,123,31,95,31,171,31,171,30,134,31,87,31,87,30,87,29,176,31,176,30,39,31,142,31,249,31,249,30,79,31,94,31,59,31,102,31,143,31,68,31,157,31,134,31,218,31,140,31,111,31,4,31,37,31,211,31,191,31,87,31,19,31,154,31,148,31,193,31,43,31,104,31,204,31,133,31,136,31,136,30,198,31,198,30,54,31,207,31,109,31,109,30,109,29,109,28,13,31,191,31,29,31,118,31,118,30,240,31,138,31,120,31,206,31,7,31,7,30,231,31,79,31,76,31,58,31,13,31,13,30,97,31,170,31,135,31,135,30,6,31,6,30,208,31,242,31,238,31,238,30,163,31,48,31,150,31,150,30,61,31,85,31,36,31,36,30,218,31,145,31,184,31,184,30,11,31,51,31,94,31,132,31,59,31,219,31,237,31,156,31,87,31,238,31,199,31,199,30,213,31,130,31,130,30,54,31,147,31,200,31,213,31,213,30,203,31,203,30,138,31,19,31,206,31,200,31,155,31,155,30,188,31,97,31,128,31,136,31,44,31,70,31,172,31,88,31,224,31,156,31,43,31,146,31,229,31,229,30,103,31,103,30,27,31,161,31,61,31,61,30,89,31,187,31,187,30,50,31,143,31,4,31,68,31,47,31,155,31,32,31,32,30,125,31,67,31,67,30,213,31,213,30,170,31,190,31,190,30,242,31,229,31,138,31,21,31,245,31,158,31,11,31,10,31,106,31,252,31,125,31,125,30,34,31,80,31,80,30,203,31,203,30,89,31,89,30,62,31,62,30,171,31,211,31,117,31,204,31,185,31,185,30,46,31,46,30,46,29,2,31,233,31,233,30,87,31,62,31,176,31,31,31,31,30,31,29,73,31,68,31,30,31,72,31,3,31,22,31,172,31,33,31,33,30,177,31,203,31,33,31,118,31,140,31,164,31,1,31,104,31,119,31,177,31,153,31,153,30,244,31,176,31,145,31,40,31,40,30,170,31,181,31,247,31,247,30,247,29,247,28,112,31,32,31,217,31,161,31,161,30,161,29,161,28,92,31,26,31,26,30,127,31,232,31,1,31,1,30,1,29,158,31,43,31,59,31,184,31,14,31,77,31,76,31,12,31,12,30,181,31,236,31,236,30,20,31,241,31,87,31,123,31,229,31,151,31,217,31,182,31,182,30,187,31,2,31,2,30,164,31,164,30,49,31,79,31,199,31,111,31,111,30,111,29,252,31,20,31,20,30,112,31,246,31,246,30,94,31,12,31,89,31,215,31,215,30,148,31,193,31,6,31,39,31,209,31,18,31,236,31,200,31,147,31,14,31,166,31,183,31,210,31,23,31,23,30,198,31,232,31,140,31,238,31,175,31,11,31,81,31,39,31,197,31,161,31,186,31,165,31,47,31,165,31,165,30,7,31,136,31,108,31,29,31,98,31,63,31,110,31,192,31,100,31,139,31,124,31,13,31,244,31,89,31,251,31,251,30,251,29,27,31,35,31,225,31,80,31,221,31,22,31,177,31,38,31,203,31,203,30,152,31,4,31,4,30,252,31,252,30,28,31,195,31,203,31,112,31,112,30,202,31,202,30,144,31,226,31,173,31,43,31,186,31,186,30,35,31,35,30,127,31,247,31,155,31,175,31,27,31,27,30,30,31,115,31,39,31,39,30,67,31,60,31,60,30,192,31,50,31,141,31,235,31,90,31,202,31,237,31,69,31,247,31,161,31,203,31,25,31,76,31,129,31,73,31,100,31,202,31,49,31,81,31,207,31,95,31,196,31,196,30,196,29,20,31,20,30,185,31,255,31,80,31,80,30,131,31,131,30,201,31,68,31,105,31,144,31,97,31,8,31,102,31,71,31,218,31,218,30,215,31,126,31,110,31,114,31,156,31,6,31,140,31,102,31,108,31,91,31,91,30,185,31,157,31,128,31,128,30,144,31,195,31,190,31,190,30,179,31,110,31,110,30,19,31,19,30,19,29,105,31,217,31,7,31,173,31,131,31,73,31,174,31,218,31,37,31,218,31,161,31,41,31,30,31,30,30,77,31,1,31,37,31,45,31,110,31,164,31,30,31,33,31,225,31,225,30,197,31,216,31,216,30,100,31,99,31,108,31,230,31,230,30,26,31,33,31,5,31,5,30,111,31,50,31,93,31,14,31,219,31,53,31,137,31,20,31,94,31,94,30,94,29,184,31,184,30,184,29,145,31,245,31,246,31,21,31,21,30,198,31,68,31,68,30,234,31,143,31,245,31,202,31,54,31,164,31,110,31,53,31,30,31,41,31,78,31,154,31,154,30,249,31,40,31,40,30,78,31,78,30,140,31,156,31,161,31,20,31,102,31,183,31,107,31,100,31,250,31,250,30,144,31,180,31,230,31,220,31,31,31,43,31,155,31,155,30,55,31,246,31,90,31,90,30,90,29,90,28,225,31,13,31,129,31,248,31,66,31,23,31,108,31,9,31,9,30,232,31,232,30,41,31,241,31,248,31,126,31,238,31,248,31,224,31,101,31,196,31,42,31,16,31,16,30,16,29,182,31,1,31,122,31,69,31,69,30,69,29,209,31,31,31,18,31,45,31,3,31,28,31,233,31,233,30,137,31,210,31,210,30,210,29,175,31,13,31,241,31,176,31,57,31,76,31,76,30,177,31,189,31,189,30,60,31,141,31,141,30,170,31,170,30,170,29,114,31,134,31,134,30,20,31,68,31,142,31,200,31,129,31,148,31,168,31,48,31,141,31,2,31,189,31,61,31,188,31,109,31,187,31,111,31,179,31,82,31,109,31,8,31,193,31,193,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
