-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 400;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (58,0,180,0,210,0,64,0,0,0,0,0,139,0,160,0,0,0,59,0,154,0,131,0,76,0,0,0,2,0,120,0,98,0,225,0,60,0,0,0,175,0,0,0,250,0,173,0,116,0,4,0,170,0,122,0,0,0,197,0,206,0,184,0,126,0,63,0,76,0,130,0,55,0,57,0,0,0,135,0,108,0,54,0,130,0,184,0,69,0,199,0,11,0,215,0,67,0,31,0,43,0,0,0,137,0,0,0,198,0,69,0,133,0,186,0,0,0,10,0,192,0,17,0,27,0,57,0,7,0,211,0,3,0,115,0,187,0,111,0,0,0,117,0,109,0,176,0,226,0,20,0,0,0,0,0,156,0,206,0,20,0,158,0,21,0,235,0,0,0,0,0,124,0,9,0,55,0,87,0,1,0,187,0,28,0,0,0,163,0,154,0,0,0,28,0,227,0,0,0,85,0,243,0,107,0,128,0,0,0,2,0,205,0,0,0,0,0,70,0,97,0,143,0,194,0,162,0,74,0,19,0,0,0,27,0,114,0,155,0,212,0,109,0,39,0,245,0,95,0,47,0,249,0,79,0,89,0,82,0,154,0,150,0,92,0,165,0,0,0,56,0,34,0,131,0,78,0,90,0,243,0,12,0,94,0,0,0,247,0,0,0,0,0,134,0,178,0,30,0,14,0,0,0,0,0,82,0,158,0,0,0,71,0,55,0,82,0,0,0,11,0,130,0,51,0,38,0,124,0,46,0,160,0,225,0,168,0,183,0,196,0,48,0,146,0,145,0,207,0,148,0,161,0,56,0,237,0,190,0,96,0,0,0,0,0,218,0,142,0,0,0,0,0,0,0,184,0,0,0,135,0,22,0,206,0,161,0,0,0,229,0,221,0,174,0,0,0,0,0,38,0,51,0,139,0,188,0,0,0,203,0,113,0,78,0,0,0,134,0,0,0,0,0,0,0,67,0,116,0,27,0,185,0,39,0,10,0,248,0,18,0,177,0,187,0,0,0,51,0,117,0,63,0,100,0,0,0,249,0,59,0,73,0,11,0,0,0,5,0,229,0,0,0,201,0,87,0,119,0,213,0,173,0,79,0,253,0,84,0,0,0,116,0,250,0,25,0,0,0,204,0,26,0,70,0,67,0,63,0,5,0,249,0,222,0,103,0,0,0,30,0,183,0,48,0,113,0,97,0,234,0,17,0,247,0,170,0,252,0,217,0,0,0,100,0,0,0,99,0,52,0,27,0,0,0,153,0,147,0,233,0,167,0,154,0,139,0,230,0,0,0,61,0,19,0,79,0,171,0,0,0,25,0,125,0,108,0,238,0,48,0,4,0,0,0,205,0,217,0,0,0,141,0,64,0,5,0,0,0,0,0,0,0,225,0,120,0,148,0,199,0,0,0,24,0,92,0,151,0,68,0,64,0,1,0,171,0,253,0,59,0,38,0,142,0,15,0,170,0,34,0,96,0,117,0,146,0,58,0,184,0,151,0,41,0,24,0,252,0,0,0,144,0,132,0,153,0,0,0,252,0,9,0,196,0,57,0,45,0,0,0,37,0,159,0,0,0,237,0,0,0,134,0,108,0,0,0,118,0,0,0,221,0,76,0,170,0,15,0,169,0,98,0,51,0,0,0,0,0,210,0,129,0,7,0,229,0,0,0,154,0,0,0,177,0,109,0,132,0,13,0,103,0,25,0,0,0,0,0,188,0,159,0,0,0,132,0,23,0,148,0,151,0,125,0,0,0,0,0,140,0,230,0,0,0,164,0,0,0,51,0,0,0,101,0,0,0,50,0);
signal scenario_full  : scenario_type := (58,31,180,31,210,31,64,31,64,30,64,29,139,31,160,31,160,30,59,31,154,31,131,31,76,31,76,30,2,31,120,31,98,31,225,31,60,31,60,30,175,31,175,30,250,31,173,31,116,31,4,31,170,31,122,31,122,30,197,31,206,31,184,31,126,31,63,31,76,31,130,31,55,31,57,31,57,30,135,31,108,31,54,31,130,31,184,31,69,31,199,31,11,31,215,31,67,31,31,31,43,31,43,30,137,31,137,30,198,31,69,31,133,31,186,31,186,30,10,31,192,31,17,31,27,31,57,31,7,31,211,31,3,31,115,31,187,31,111,31,111,30,117,31,109,31,176,31,226,31,20,31,20,30,20,29,156,31,206,31,20,31,158,31,21,31,235,31,235,30,235,29,124,31,9,31,55,31,87,31,1,31,187,31,28,31,28,30,163,31,154,31,154,30,28,31,227,31,227,30,85,31,243,31,107,31,128,31,128,30,2,31,205,31,205,30,205,29,70,31,97,31,143,31,194,31,162,31,74,31,19,31,19,30,27,31,114,31,155,31,212,31,109,31,39,31,245,31,95,31,47,31,249,31,79,31,89,31,82,31,154,31,150,31,92,31,165,31,165,30,56,31,34,31,131,31,78,31,90,31,243,31,12,31,94,31,94,30,247,31,247,30,247,29,134,31,178,31,30,31,14,31,14,30,14,29,82,31,158,31,158,30,71,31,55,31,82,31,82,30,11,31,130,31,51,31,38,31,124,31,46,31,160,31,225,31,168,31,183,31,196,31,48,31,146,31,145,31,207,31,148,31,161,31,56,31,237,31,190,31,96,31,96,30,96,29,218,31,142,31,142,30,142,29,142,28,184,31,184,30,135,31,22,31,206,31,161,31,161,30,229,31,221,31,174,31,174,30,174,29,38,31,51,31,139,31,188,31,188,30,203,31,113,31,78,31,78,30,134,31,134,30,134,29,134,28,67,31,116,31,27,31,185,31,39,31,10,31,248,31,18,31,177,31,187,31,187,30,51,31,117,31,63,31,100,31,100,30,249,31,59,31,73,31,11,31,11,30,5,31,229,31,229,30,201,31,87,31,119,31,213,31,173,31,79,31,253,31,84,31,84,30,116,31,250,31,25,31,25,30,204,31,26,31,70,31,67,31,63,31,5,31,249,31,222,31,103,31,103,30,30,31,183,31,48,31,113,31,97,31,234,31,17,31,247,31,170,31,252,31,217,31,217,30,100,31,100,30,99,31,52,31,27,31,27,30,153,31,147,31,233,31,167,31,154,31,139,31,230,31,230,30,61,31,19,31,79,31,171,31,171,30,25,31,125,31,108,31,238,31,48,31,4,31,4,30,205,31,217,31,217,30,141,31,64,31,5,31,5,30,5,29,5,28,225,31,120,31,148,31,199,31,199,30,24,31,92,31,151,31,68,31,64,31,1,31,171,31,253,31,59,31,38,31,142,31,15,31,170,31,34,31,96,31,117,31,146,31,58,31,184,31,151,31,41,31,24,31,252,31,252,30,144,31,132,31,153,31,153,30,252,31,9,31,196,31,57,31,45,31,45,30,37,31,159,31,159,30,237,31,237,30,134,31,108,31,108,30,118,31,118,30,221,31,76,31,170,31,15,31,169,31,98,31,51,31,51,30,51,29,210,31,129,31,7,31,229,31,229,30,154,31,154,30,177,31,109,31,132,31,13,31,103,31,25,31,25,30,25,29,188,31,159,31,159,30,132,31,23,31,148,31,151,31,125,31,125,30,125,29,140,31,230,31,230,30,164,31,164,30,51,31,51,30,101,31,101,30,50,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
