-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_189 is
end project_tb_189;

architecture project_tb_arch_189 of project_tb_189 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 686;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (58,0,121,0,182,0,133,0,159,0,144,0,179,0,15,0,184,0,9,0,0,0,4,0,208,0,24,0,216,0,208,0,34,0,6,0,128,0,40,0,30,0,0,0,30,0,168,0,112,0,50,0,64,0,98,0,43,0,0,0,0,0,130,0,30,0,168,0,212,0,195,0,0,0,5,0,199,0,245,0,217,0,27,0,27,0,160,0,9,0,146,0,238,0,238,0,0,0,152,0,241,0,228,0,81,0,0,0,157,0,9,0,0,0,217,0,245,0,0,0,18,0,108,0,23,0,31,0,113,0,4,0,0,0,20,0,249,0,159,0,54,0,43,0,180,0,82,0,225,0,165,0,211,0,133,0,5,0,0,0,148,0,51,0,192,0,0,0,13,0,0,0,181,0,250,0,0,0,0,0,187,0,175,0,18,0,28,0,238,0,0,0,255,0,141,0,138,0,187,0,126,0,159,0,7,0,83,0,211,0,0,0,0,0,0,0,82,0,14,0,69,0,168,0,140,0,243,0,156,0,38,0,54,0,157,0,0,0,73,0,226,0,0,0,0,0,105,0,79,0,0,0,0,0,0,0,233,0,0,0,192,0,23,0,62,0,0,0,95,0,51,0,166,0,137,0,237,0,155,0,255,0,149,0,106,0,0,0,150,0,0,0,231,0,0,0,17,0,1,0,110,0,115,0,156,0,222,0,253,0,154,0,156,0,0,0,119,0,166,0,3,0,221,0,0,0,29,0,43,0,0,0,225,0,180,0,0,0,151,0,235,0,23,0,62,0,53,0,0,0,102,0,5,0,162,0,195,0,0,0,0,0,104,0,0,0,110,0,143,0,31,0,248,0,231,0,187,0,217,0,13,0,253,0,115,0,142,0,87,0,11,0,180,0,167,0,0,0,180,0,0,0,0,0,74,0,164,0,137,0,12,0,157,0,0,0,131,0,200,0,102,0,226,0,0,0,56,0,91,0,246,0,114,0,125,0,255,0,0,0,144,0,224,0,147,0,36,0,96,0,94,0,104,0,93,0,147,0,29,0,223,0,174,0,183,0,181,0,231,0,56,0,122,0,184,0,146,0,29,0,155,0,223,0,49,0,234,0,73,0,127,0,226,0,161,0,130,0,204,0,192,0,0,0,72,0,0,0,32,0,191,0,214,0,14,0,104,0,94,0,103,0,38,0,252,0,173,0,147,0,0,0,98,0,20,0,131,0,7,0,160,0,237,0,198,0,109,0,33,0,0,0,169,0,169,0,204,0,73,0,229,0,0,0,45,0,167,0,208,0,42,0,0,0,71,0,0,0,233,0,33,0,252,0,52,0,81,0,0,0,193,0,0,0,50,0,217,0,0,0,54,0,182,0,231,0,0,0,0,0,0,0,225,0,0,0,62,0,0,0,26,0,84,0,180,0,148,0,213,0,193,0,0,0,51,0,215,0,0,0,152,0,190,0,0,0,3,0,0,0,129,0,0,0,53,0,150,0,0,0,104,0,132,0,14,0,0,0,111,0,142,0,192,0,170,0,41,0,237,0,0,0,139,0,66,0,63,0,242,0,107,0,0,0,251,0,253,0,160,0,253,0,164,0,153,0,0,0,167,0,0,0,0,0,16,0,78,0,251,0,134,0,162,0,70,0,124,0,156,0,35,0,0,0,0,0,26,0,0,0,137,0,0,0,43,0,0,0,184,0,0,0,145,0,92,0,75,0,104,0,40,0,10,0,148,0,221,0,238,0,98,0,220,0,158,0,64,0,109,0,222,0,224,0,29,0,0,0,0,0,0,0,185,0,122,0,157,0,0,0,247,0,0,0,0,0,49,0,63,0,226,0,104,0,0,0,174,0,0,0,0,0,84,0,0,0,67,0,43,0,166,0,0,0,45,0,0,0,71,0,186,0,181,0,136,0,0,0,229,0,148,0,23,0,180,0,64,0,0,0,0,0,0,0,242,0,201,0,0,0,202,0,66,0,114,0,100,0,99,0,218,0,198,0,60,0,0,0,146,0,51,0,196,0,21,0,97,0,161,0,0,0,113,0,0,0,57,0,199,0,214,0,141,0,188,0,109,0,96,0,0,0,236,0,233,0,0,0,71,0,255,0,165,0,0,0,168,0,0,0,140,0,176,0,228,0,0,0,95,0,80,0,206,0,134,0,0,0,214,0,125,0,119,0,8,0,233,0,219,0,0,0,109,0,189,0,0,0,3,0,221,0,196,0,216,0,82,0,230,0,71,0,179,0,60,0,231,0,205,0,0,0,0,0,0,0,240,0,181,0,255,0,30,0,0,0,84,0,88,0,248,0,151,0,198,0,170,0,251,0,169,0,162,0,193,0,0,0,14,0,38,0,45,0,30,0,5,0,0,0,200,0,198,0,236,0,98,0,117,0,0,0,214,0,176,0,0,0,254,0,60,0,247,0,242,0,35,0,129,0,214,0,0,0,28,0,45,0,78,0,231,0,129,0,0,0,39,0,149,0,0,0,199,0,26,0,139,0,2,0,108,0,201,0,43,0,83,0,3,0,157,0,201,0,29,0,93,0,156,0,114,0,131,0,50,0,216,0,192,0,147,0,229,0,117,0,119,0,0,0,131,0,25,0,176,0,0,0,17,0,43,0,66,0,189,0,79,0,74,0,37,0,180,0,72,0,189,0,0,0,40,0,157,0,0,0,47,0,134,0,250,0,0,0,81,0,139,0,188,0,0,0,0,0,85,0,33,0,0,0,254,0,71,0,117,0,57,0,116,0,80,0,72,0,83,0,0,0,0,0,14,0,92,0,44,0,18,0,103,0,134,0,169,0,214,0,214,0,173,0,63,0,0,0,251,0,174,0,185,0,152,0,247,0,0,0,174,0,0,0,243,0,0,0,0,0,125,0,163,0,66,0,37,0,240,0,220,0,0,0,0,0,214,0,90,0,61,0,214,0,215,0,0,0,89,0,203,0,8,0,253,0,0,0,136,0,10,0,78,0,39,0,0,0,162,0,180,0,57,0,0,0,132,0,201,0,140,0,229,0,189,0,56,0,30,0,1,0,159,0,23,0,145,0,216,0,85,0,0,0,44,0,0,0,203,0,21,0,23,0,121,0);
signal scenario_full  : scenario_type := (58,31,121,31,182,31,133,31,159,31,144,31,179,31,15,31,184,31,9,31,9,30,4,31,208,31,24,31,216,31,208,31,34,31,6,31,128,31,40,31,30,31,30,30,30,31,168,31,112,31,50,31,64,31,98,31,43,31,43,30,43,29,130,31,30,31,168,31,212,31,195,31,195,30,5,31,199,31,245,31,217,31,27,31,27,31,160,31,9,31,146,31,238,31,238,31,238,30,152,31,241,31,228,31,81,31,81,30,157,31,9,31,9,30,217,31,245,31,245,30,18,31,108,31,23,31,31,31,113,31,4,31,4,30,20,31,249,31,159,31,54,31,43,31,180,31,82,31,225,31,165,31,211,31,133,31,5,31,5,30,148,31,51,31,192,31,192,30,13,31,13,30,181,31,250,31,250,30,250,29,187,31,175,31,18,31,28,31,238,31,238,30,255,31,141,31,138,31,187,31,126,31,159,31,7,31,83,31,211,31,211,30,211,29,211,28,82,31,14,31,69,31,168,31,140,31,243,31,156,31,38,31,54,31,157,31,157,30,73,31,226,31,226,30,226,29,105,31,79,31,79,30,79,29,79,28,233,31,233,30,192,31,23,31,62,31,62,30,95,31,51,31,166,31,137,31,237,31,155,31,255,31,149,31,106,31,106,30,150,31,150,30,231,31,231,30,17,31,1,31,110,31,115,31,156,31,222,31,253,31,154,31,156,31,156,30,119,31,166,31,3,31,221,31,221,30,29,31,43,31,43,30,225,31,180,31,180,30,151,31,235,31,23,31,62,31,53,31,53,30,102,31,5,31,162,31,195,31,195,30,195,29,104,31,104,30,110,31,143,31,31,31,248,31,231,31,187,31,217,31,13,31,253,31,115,31,142,31,87,31,11,31,180,31,167,31,167,30,180,31,180,30,180,29,74,31,164,31,137,31,12,31,157,31,157,30,131,31,200,31,102,31,226,31,226,30,56,31,91,31,246,31,114,31,125,31,255,31,255,30,144,31,224,31,147,31,36,31,96,31,94,31,104,31,93,31,147,31,29,31,223,31,174,31,183,31,181,31,231,31,56,31,122,31,184,31,146,31,29,31,155,31,223,31,49,31,234,31,73,31,127,31,226,31,161,31,130,31,204,31,192,31,192,30,72,31,72,30,32,31,191,31,214,31,14,31,104,31,94,31,103,31,38,31,252,31,173,31,147,31,147,30,98,31,20,31,131,31,7,31,160,31,237,31,198,31,109,31,33,31,33,30,169,31,169,31,204,31,73,31,229,31,229,30,45,31,167,31,208,31,42,31,42,30,71,31,71,30,233,31,33,31,252,31,52,31,81,31,81,30,193,31,193,30,50,31,217,31,217,30,54,31,182,31,231,31,231,30,231,29,231,28,225,31,225,30,62,31,62,30,26,31,84,31,180,31,148,31,213,31,193,31,193,30,51,31,215,31,215,30,152,31,190,31,190,30,3,31,3,30,129,31,129,30,53,31,150,31,150,30,104,31,132,31,14,31,14,30,111,31,142,31,192,31,170,31,41,31,237,31,237,30,139,31,66,31,63,31,242,31,107,31,107,30,251,31,253,31,160,31,253,31,164,31,153,31,153,30,167,31,167,30,167,29,16,31,78,31,251,31,134,31,162,31,70,31,124,31,156,31,35,31,35,30,35,29,26,31,26,30,137,31,137,30,43,31,43,30,184,31,184,30,145,31,92,31,75,31,104,31,40,31,10,31,148,31,221,31,238,31,98,31,220,31,158,31,64,31,109,31,222,31,224,31,29,31,29,30,29,29,29,28,185,31,122,31,157,31,157,30,247,31,247,30,247,29,49,31,63,31,226,31,104,31,104,30,174,31,174,30,174,29,84,31,84,30,67,31,43,31,166,31,166,30,45,31,45,30,71,31,186,31,181,31,136,31,136,30,229,31,148,31,23,31,180,31,64,31,64,30,64,29,64,28,242,31,201,31,201,30,202,31,66,31,114,31,100,31,99,31,218,31,198,31,60,31,60,30,146,31,51,31,196,31,21,31,97,31,161,31,161,30,113,31,113,30,57,31,199,31,214,31,141,31,188,31,109,31,96,31,96,30,236,31,233,31,233,30,71,31,255,31,165,31,165,30,168,31,168,30,140,31,176,31,228,31,228,30,95,31,80,31,206,31,134,31,134,30,214,31,125,31,119,31,8,31,233,31,219,31,219,30,109,31,189,31,189,30,3,31,221,31,196,31,216,31,82,31,230,31,71,31,179,31,60,31,231,31,205,31,205,30,205,29,205,28,240,31,181,31,255,31,30,31,30,30,84,31,88,31,248,31,151,31,198,31,170,31,251,31,169,31,162,31,193,31,193,30,14,31,38,31,45,31,30,31,5,31,5,30,200,31,198,31,236,31,98,31,117,31,117,30,214,31,176,31,176,30,254,31,60,31,247,31,242,31,35,31,129,31,214,31,214,30,28,31,45,31,78,31,231,31,129,31,129,30,39,31,149,31,149,30,199,31,26,31,139,31,2,31,108,31,201,31,43,31,83,31,3,31,157,31,201,31,29,31,93,31,156,31,114,31,131,31,50,31,216,31,192,31,147,31,229,31,117,31,119,31,119,30,131,31,25,31,176,31,176,30,17,31,43,31,66,31,189,31,79,31,74,31,37,31,180,31,72,31,189,31,189,30,40,31,157,31,157,30,47,31,134,31,250,31,250,30,81,31,139,31,188,31,188,30,188,29,85,31,33,31,33,30,254,31,71,31,117,31,57,31,116,31,80,31,72,31,83,31,83,30,83,29,14,31,92,31,44,31,18,31,103,31,134,31,169,31,214,31,214,31,173,31,63,31,63,30,251,31,174,31,185,31,152,31,247,31,247,30,174,31,174,30,243,31,243,30,243,29,125,31,163,31,66,31,37,31,240,31,220,31,220,30,220,29,214,31,90,31,61,31,214,31,215,31,215,30,89,31,203,31,8,31,253,31,253,30,136,31,10,31,78,31,39,31,39,30,162,31,180,31,57,31,57,30,132,31,201,31,140,31,229,31,189,31,56,31,30,31,1,31,159,31,23,31,145,31,216,31,85,31,85,30,44,31,44,30,203,31,21,31,23,31,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
