-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 723;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (130,0,0,0,16,0,89,0,0,0,209,0,0,0,77,0,155,0,192,0,126,0,0,0,0,0,103,0,114,0,65,0,220,0,154,0,0,0,164,0,102,0,194,0,67,0,246,0,47,0,0,0,108,0,0,0,0,0,27,0,87,0,11,0,50,0,0,0,233,0,153,0,94,0,67,0,146,0,139,0,206,0,24,0,0,0,125,0,48,0,0,0,198,0,0,0,213,0,1,0,114,0,0,0,0,0,209,0,43,0,114,0,70,0,134,0,173,0,0,0,175,0,0,0,11,0,0,0,164,0,0,0,0,0,36,0,72,0,0,0,50,0,115,0,214,0,33,0,199,0,68,0,57,0,139,0,196,0,167,0,189,0,75,0,0,0,235,0,77,0,160,0,0,0,0,0,51,0,37,0,41,0,146,0,73,0,195,0,82,0,56,0,72,0,28,0,215,0,234,0,0,0,149,0,0,0,0,0,0,0,69,0,0,0,215,0,82,0,162,0,133,0,139,0,253,0,38,0,173,0,184,0,191,0,0,0,90,0,175,0,222,0,251,0,250,0,97,0,0,0,0,0,0,0,54,0,115,0,227,0,36,0,9,0,141,0,148,0,0,0,242,0,213,0,195,0,128,0,144,0,66,0,67,0,0,0,79,0,134,0,0,0,0,0,130,0,0,0,210,0,130,0,135,0,0,0,0,0,0,0,168,0,151,0,0,0,84,0,131,0,0,0,1,0,154,0,34,0,0,0,58,0,50,0,105,0,139,0,238,0,9,0,0,0,0,0,194,0,156,0,0,0,0,0,110,0,98,0,148,0,24,0,0,0,143,0,103,0,0,0,147,0,202,0,190,0,0,0,0,0,113,0,172,0,0,0,1,0,120,0,0,0,222,0,0,0,251,0,169,0,72,0,0,0,127,0,15,0,83,0,81,0,0,0,213,0,115,0,0,0,0,0,0,0,219,0,0,0,61,0,160,0,0,0,66,0,48,0,70,0,111,0,169,0,0,0,211,0,214,0,135,0,0,0,183,0,241,0,113,0,83,0,122,0,12,0,9,0,45,0,195,0,0,0,247,0,23,0,208,0,189,0,32,0,47,0,16,0,249,0,193,0,216,0,0,0,31,0,158,0,99,0,201,0,56,0,0,0,175,0,202,0,0,0,134,0,0,0,107,0,79,0,65,0,245,0,164,0,186,0,133,0,26,0,111,0,18,0,0,0,218,0,160,0,0,0,217,0,30,0,102,0,0,0,150,0,217,0,237,0,8,0,150,0,233,0,73,0,0,0,150,0,0,0,0,0,47,0,129,0,38,0,240,0,0,0,253,0,112,0,250,0,119,0,120,0,0,0,133,0,238,0,0,0,0,0,0,0,51,0,6,0,109,0,28,0,29,0,40,0,119,0,15,0,74,0,0,0,14,0,47,0,132,0,91,0,0,0,29,0,69,0,124,0,193,0,184,0,0,0,81,0,139,0,245,0,142,0,224,0,205,0,0,0,217,0,0,0,138,0,208,0,41,0,105,0,198,0,163,0,229,0,0,0,0,0,153,0,0,0,5,0,136,0,36,0,165,0,55,0,224,0,94,0,89,0,63,0,103,0,138,0,51,0,136,0,31,0,40,0,192,0,146,0,152,0,204,0,88,0,173,0,0,0,200,0,0,0,6,0,178,0,231,0,48,0,226,0,148,0,53,0,19,0,232,0,0,0,0,0,49,0,156,0,169,0,142,0,117,0,109,0,49,0,98,0,81,0,202,0,214,0,0,0,199,0,0,0,0,0,233,0,207,0,193,0,0,0,207,0,4,0,215,0,0,0,0,0,175,0,29,0,236,0,126,0,34,0,66,0,145,0,236,0,232,0,80,0,51,0,171,0,237,0,252,0,146,0,49,0,25,0,146,0,0,0,252,0,106,0,226,0,64,0,87,0,0,0,0,0,0,0,38,0,0,0,62,0,25,0,74,0,12,0,124,0,137,0,224,0,120,0,183,0,103,0,238,0,238,0,35,0,141,0,54,0,0,0,37,0,176,0,223,0,171,0,2,0,148,0,147,0,243,0,151,0,0,0,238,0,70,0,206,0,94,0,57,0,58,0,146,0,65,0,0,0,184,0,95,0,153,0,35,0,20,0,19,0,165,0,138,0,9,0,56,0,21,0,129,0,0,0,137,0,0,0,65,0,237,0,85,0,159,0,153,0,59,0,82,0,38,0,237,0,251,0,174,0,0,0,227,0,0,0,207,0,241,0,51,0,9,0,114,0,0,0,70,0,232,0,219,0,125,0,242,0,255,0,248,0,82,0,105,0,0,0,42,0,214,0,214,0,124,0,143,0,252,0,135,0,0,0,224,0,88,0,179,0,229,0,0,0,160,0,143,0,28,0,214,0,120,0,12,0,113,0,43,0,47,0,39,0,80,0,127,0,243,0,168,0,79,0,50,0,80,0,219,0,0,0,0,0,93,0,235,0,178,0,113,0,236,0,187,0,16,0,0,0,97,0,218,0,253,0,126,0,203,0,189,0,231,0,0,0,231,0,0,0,0,0,43,0,8,0,130,0,85,0,54,0,139,0,167,0,63,0,0,0,70,0,65,0,65,0,54,0,186,0,81,0,235,0,0,0,44,0,0,0,170,0,108,0,153,0,50,0,0,0,247,0,0,0,254,0,229,0,150,0,246,0,91,0,0,0,0,0,200,0,184,0,196,0,140,0,30,0,0,0,149,0,247,0,54,0,30,0,145,0,168,0,151,0,215,0,98,0,0,0,0,0,182,0,11,0,41,0,88,0,213,0,0,0,159,0,113,0,176,0,125,0,32,0,104,0,112,0,228,0,93,0,123,0,50,0,182,0,49,0,113,0,220,0,204,0,207,0,44,0,0,0,0,0,170,0,22,0,219,0,138,0,239,0,173,0,0,0,0,0,41,0,25,0,0,0,112,0,0,0,21,0,86,0,117,0,176,0,140,0,0,0,243,0,115,0,236,0,49,0,209,0,222,0,0,0,0,0,0,0,0,0,161,0,59,0,102,0,48,0,76,0,116,0,0,0,0,0,0,0,0,0,211,0,97,0,0,0,96,0,80,0,112,0,47,0,52,0,248,0,165,0,0,0,43,0,0,0,68,0,17,0,149,0,33,0,0,0,247,0,7,0,55,0,151,0,181,0,59,0,0,0,0,0,137,0,0,0,187,0,135,0,125,0,24,0,82,0,0,0,111,0,199,0,109,0,0,0,66,0,83,0,42,0,77,0,251,0);
signal scenario_full  : scenario_type := (130,31,130,30,16,31,89,31,89,30,209,31,209,30,77,31,155,31,192,31,126,31,126,30,126,29,103,31,114,31,65,31,220,31,154,31,154,30,164,31,102,31,194,31,67,31,246,31,47,31,47,30,108,31,108,30,108,29,27,31,87,31,11,31,50,31,50,30,233,31,153,31,94,31,67,31,146,31,139,31,206,31,24,31,24,30,125,31,48,31,48,30,198,31,198,30,213,31,1,31,114,31,114,30,114,29,209,31,43,31,114,31,70,31,134,31,173,31,173,30,175,31,175,30,11,31,11,30,164,31,164,30,164,29,36,31,72,31,72,30,50,31,115,31,214,31,33,31,199,31,68,31,57,31,139,31,196,31,167,31,189,31,75,31,75,30,235,31,77,31,160,31,160,30,160,29,51,31,37,31,41,31,146,31,73,31,195,31,82,31,56,31,72,31,28,31,215,31,234,31,234,30,149,31,149,30,149,29,149,28,69,31,69,30,215,31,82,31,162,31,133,31,139,31,253,31,38,31,173,31,184,31,191,31,191,30,90,31,175,31,222,31,251,31,250,31,97,31,97,30,97,29,97,28,54,31,115,31,227,31,36,31,9,31,141,31,148,31,148,30,242,31,213,31,195,31,128,31,144,31,66,31,67,31,67,30,79,31,134,31,134,30,134,29,130,31,130,30,210,31,130,31,135,31,135,30,135,29,135,28,168,31,151,31,151,30,84,31,131,31,131,30,1,31,154,31,34,31,34,30,58,31,50,31,105,31,139,31,238,31,9,31,9,30,9,29,194,31,156,31,156,30,156,29,110,31,98,31,148,31,24,31,24,30,143,31,103,31,103,30,147,31,202,31,190,31,190,30,190,29,113,31,172,31,172,30,1,31,120,31,120,30,222,31,222,30,251,31,169,31,72,31,72,30,127,31,15,31,83,31,81,31,81,30,213,31,115,31,115,30,115,29,115,28,219,31,219,30,61,31,160,31,160,30,66,31,48,31,70,31,111,31,169,31,169,30,211,31,214,31,135,31,135,30,183,31,241,31,113,31,83,31,122,31,12,31,9,31,45,31,195,31,195,30,247,31,23,31,208,31,189,31,32,31,47,31,16,31,249,31,193,31,216,31,216,30,31,31,158,31,99,31,201,31,56,31,56,30,175,31,202,31,202,30,134,31,134,30,107,31,79,31,65,31,245,31,164,31,186,31,133,31,26,31,111,31,18,31,18,30,218,31,160,31,160,30,217,31,30,31,102,31,102,30,150,31,217,31,237,31,8,31,150,31,233,31,73,31,73,30,150,31,150,30,150,29,47,31,129,31,38,31,240,31,240,30,253,31,112,31,250,31,119,31,120,31,120,30,133,31,238,31,238,30,238,29,238,28,51,31,6,31,109,31,28,31,29,31,40,31,119,31,15,31,74,31,74,30,14,31,47,31,132,31,91,31,91,30,29,31,69,31,124,31,193,31,184,31,184,30,81,31,139,31,245,31,142,31,224,31,205,31,205,30,217,31,217,30,138,31,208,31,41,31,105,31,198,31,163,31,229,31,229,30,229,29,153,31,153,30,5,31,136,31,36,31,165,31,55,31,224,31,94,31,89,31,63,31,103,31,138,31,51,31,136,31,31,31,40,31,192,31,146,31,152,31,204,31,88,31,173,31,173,30,200,31,200,30,6,31,178,31,231,31,48,31,226,31,148,31,53,31,19,31,232,31,232,30,232,29,49,31,156,31,169,31,142,31,117,31,109,31,49,31,98,31,81,31,202,31,214,31,214,30,199,31,199,30,199,29,233,31,207,31,193,31,193,30,207,31,4,31,215,31,215,30,215,29,175,31,29,31,236,31,126,31,34,31,66,31,145,31,236,31,232,31,80,31,51,31,171,31,237,31,252,31,146,31,49,31,25,31,146,31,146,30,252,31,106,31,226,31,64,31,87,31,87,30,87,29,87,28,38,31,38,30,62,31,25,31,74,31,12,31,124,31,137,31,224,31,120,31,183,31,103,31,238,31,238,31,35,31,141,31,54,31,54,30,37,31,176,31,223,31,171,31,2,31,148,31,147,31,243,31,151,31,151,30,238,31,70,31,206,31,94,31,57,31,58,31,146,31,65,31,65,30,184,31,95,31,153,31,35,31,20,31,19,31,165,31,138,31,9,31,56,31,21,31,129,31,129,30,137,31,137,30,65,31,237,31,85,31,159,31,153,31,59,31,82,31,38,31,237,31,251,31,174,31,174,30,227,31,227,30,207,31,241,31,51,31,9,31,114,31,114,30,70,31,232,31,219,31,125,31,242,31,255,31,248,31,82,31,105,31,105,30,42,31,214,31,214,31,124,31,143,31,252,31,135,31,135,30,224,31,88,31,179,31,229,31,229,30,160,31,143,31,28,31,214,31,120,31,12,31,113,31,43,31,47,31,39,31,80,31,127,31,243,31,168,31,79,31,50,31,80,31,219,31,219,30,219,29,93,31,235,31,178,31,113,31,236,31,187,31,16,31,16,30,97,31,218,31,253,31,126,31,203,31,189,31,231,31,231,30,231,31,231,30,231,29,43,31,8,31,130,31,85,31,54,31,139,31,167,31,63,31,63,30,70,31,65,31,65,31,54,31,186,31,81,31,235,31,235,30,44,31,44,30,170,31,108,31,153,31,50,31,50,30,247,31,247,30,254,31,229,31,150,31,246,31,91,31,91,30,91,29,200,31,184,31,196,31,140,31,30,31,30,30,149,31,247,31,54,31,30,31,145,31,168,31,151,31,215,31,98,31,98,30,98,29,182,31,11,31,41,31,88,31,213,31,213,30,159,31,113,31,176,31,125,31,32,31,104,31,112,31,228,31,93,31,123,31,50,31,182,31,49,31,113,31,220,31,204,31,207,31,44,31,44,30,44,29,170,31,22,31,219,31,138,31,239,31,173,31,173,30,173,29,41,31,25,31,25,30,112,31,112,30,21,31,86,31,117,31,176,31,140,31,140,30,243,31,115,31,236,31,49,31,209,31,222,31,222,30,222,29,222,28,222,27,161,31,59,31,102,31,48,31,76,31,116,31,116,30,116,29,116,28,116,27,211,31,97,31,97,30,96,31,80,31,112,31,47,31,52,31,248,31,165,31,165,30,43,31,43,30,68,31,17,31,149,31,33,31,33,30,247,31,7,31,55,31,151,31,181,31,59,31,59,30,59,29,137,31,137,30,187,31,135,31,125,31,24,31,82,31,82,30,111,31,199,31,109,31,109,30,66,31,83,31,42,31,77,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
