-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_864 is
end project_tb_864;

architecture project_tb_arch_864 of project_tb_864 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 719;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (84,0,232,0,91,0,225,0,97,0,179,0,31,0,38,0,73,0,0,0,0,0,220,0,58,0,144,0,185,0,219,0,0,0,27,0,0,0,174,0,97,0,250,0,198,0,121,0,225,0,0,0,0,0,199,0,0,0,15,0,7,0,0,0,0,0,214,0,223,0,0,0,185,0,1,0,111,0,140,0,6,0,0,0,87,0,0,0,0,0,173,0,0,0,0,0,106,0,175,0,78,0,132,0,85,0,85,0,194,0,121,0,0,0,88,0,246,0,241,0,50,0,91,0,55,0,0,0,29,0,85,0,142,0,201,0,0,0,149,0,117,0,0,0,152,0,109,0,172,0,170,0,16,0,0,0,177,0,44,0,101,0,92,0,182,0,0,0,0,0,63,0,232,0,68,0,208,0,110,0,118,0,152,0,237,0,0,0,168,0,202,0,96,0,212,0,0,0,112,0,160,0,0,0,0,0,201,0,0,0,148,0,78,0,108,0,136,0,85,0,0,0,0,0,0,0,0,0,203,0,0,0,113,0,45,0,95,0,176,0,227,0,142,0,185,0,0,0,0,0,108,0,138,0,74,0,76,0,80,0,102,0,0,0,39,0,105,0,148,0,173,0,0,0,0,0,125,0,0,0,177,0,98,0,121,0,0,0,194,0,11,0,209,0,37,0,58,0,166,0,52,0,18,0,19,0,67,0,34,0,0,0,125,0,36,0,55,0,35,0,0,0,70,0,8,0,7,0,8,0,47,0,171,0,122,0,227,0,76,0,222,0,0,0,0,0,72,0,163,0,0,0,0,0,202,0,9,0,18,0,95,0,0,0,0,0,205,0,14,0,112,0,1,0,138,0,177,0,48,0,149,0,241,0,210,0,0,0,49,0,246,0,150,0,206,0,222,0,80,0,0,0,229,0,1,0,71,0,199,0,120,0,222,0,123,0,39,0,159,0,206,0,248,0,150,0,93,0,125,0,93,0,146,0,58,0,134,0,190,0,212,0,74,0,0,0,97,0,85,0,15,0,62,0,217,0,236,0,142,0,111,0,16,0,232,0,235,0,0,0,254,0,0,0,61,0,0,0,84,0,112,0,8,0,0,0,0,0,70,0,144,0,184,0,244,0,105,0,156,0,220,0,82,0,71,0,241,0,88,0,0,0,152,0,229,0,109,0,0,0,218,0,235,0,24,0,225,0,187,0,230,0,41,0,0,0,204,0,143,0,17,0,71,0,122,0,133,0,177,0,216,0,252,0,103,0,153,0,162,0,50,0,94,0,89,0,225,0,112,0,0,0,184,0,0,0,0,0,0,0,0,0,60,0,31,0,0,0,136,0,218,0,49,0,143,0,145,0,220,0,0,0,103,0,198,0,49,0,225,0,35,0,224,0,140,0,168,0,127,0,95,0,104,0,244,0,130,0,30,0,224,0,221,0,80,0,35,0,177,0,233,0,94,0,110,0,144,0,63,0,215,0,205,0,80,0,113,0,132,0,241,0,182,0,183,0,42,0,221,0,116,0,251,0,106,0,4,0,220,0,226,0,0,0,65,0,224,0,8,0,252,0,110,0,228,0,0,0,157,0,245,0,103,0,224,0,163,0,0,0,0,0,0,0,239,0,0,0,226,0,230,0,185,0,201,0,79,0,150,0,46,0,249,0,115,0,0,0,56,0,81,0,62,0,97,0,118,0,139,0,82,0,60,0,30,0,0,0,152,0,0,0,233,0,0,0,249,0,0,0,190,0,87,0,120,0,31,0,150,0,112,0,211,0,151,0,221,0,0,0,59,0,201,0,189,0,24,0,62,0,75,0,178,0,47,0,0,0,168,0,0,0,232,0,4,0,72,0,162,0,67,0,232,0,39,0,16,0,133,0,0,0,3,0,90,0,162,0,0,0,0,0,140,0,102,0,255,0,200,0,218,0,122,0,0,0,24,0,147,0,0,0,125,0,208,0,161,0,0,0,0,0,31,0,20,0,159,0,154,0,101,0,85,0,221,0,27,0,62,0,13,0,237,0,174,0,195,0,10,0,105,0,206,0,0,0,0,0,78,0,195,0,189,0,43,0,0,0,85,0,0,0,181,0,141,0,0,0,135,0,111,0,46,0,39,0,172,0,5,0,220,0,36,0,88,0,250,0,0,0,127,0,64,0,76,0,0,0,6,0,60,0,253,0,0,0,88,0,206,0,154,0,177,0,27,0,132,0,142,0,255,0,82,0,98,0,0,0,229,0,240,0,0,0,0,0,180,0,81,0,103,0,44,0,120,0,184,0,0,0,91,0,0,0,214,0,31,0,137,0,40,0,0,0,0,0,0,0,127,0,137,0,241,0,159,0,220,0,0,0,227,0,247,0,166,0,22,0,0,0,0,0,152,0,242,0,241,0,240,0,9,0,0,0,204,0,145,0,160,0,175,0,115,0,16,0,202,0,205,0,0,0,65,0,168,0,214,0,20,0,0,0,253,0,0,0,0,0,89,0,159,0,5,0,113,0,13,0,0,0,0,0,132,0,180,0,146,0,0,0,4,0,249,0,111,0,0,0,136,0,167,0,109,0,225,0,4,0,186,0,151,0,28,0,0,0,42,0,105,0,38,0,162,0,40,0,129,0,141,0,135,0,22,0,140,0,68,0,129,0,157,0,53,0,0,0,162,0,143,0,57,0,41,0,125,0,217,0,221,0,248,0,248,0,0,0,0,0,63,0,197,0,157,0,43,0,79,0,0,0,97,0,186,0,0,0,152,0,123,0,0,0,0,0,0,0,179,0,41,0,0,0,230,0,0,0,43,0,10,0,107,0,131,0,65,0,0,0,114,0,130,0,13,0,65,0,50,0,185,0,57,0,211,0,239,0,207,0,0,0,0,0,98,0,79,0,106,0,155,0,0,0,0,0,245,0,206,0,0,0,239,0,0,0,243,0,68,0,48,0,196,0,222,0,196,0,254,0,102,0,0,0,58,0,0,0,118,0,148,0,0,0,64,0,0,0,124,0,116,0,47,0,225,0,170,0,103,0,27,0,15,0,60,0,36,0,183,0,224,0,160,0,107,0,86,0,241,0,0,0,82,0,177,0,126,0,8,0,8,0,0,0,111,0,40,0,134,0,177,0,0,0,0,0,148,0,92,0,212,0,153,0,0,0,183,0,39,0,212,0,91,0,0,0,14,0,7,0,207,0,0,0,63,0,125,0,66,0,221,0,0,0,230,0,49,0,31,0,128,0,128,0,28,0,0,0,154,0);
signal scenario_full  : scenario_type := (84,31,232,31,91,31,225,31,97,31,179,31,31,31,38,31,73,31,73,30,73,29,220,31,58,31,144,31,185,31,219,31,219,30,27,31,27,30,174,31,97,31,250,31,198,31,121,31,225,31,225,30,225,29,199,31,199,30,15,31,7,31,7,30,7,29,214,31,223,31,223,30,185,31,1,31,111,31,140,31,6,31,6,30,87,31,87,30,87,29,173,31,173,30,173,29,106,31,175,31,78,31,132,31,85,31,85,31,194,31,121,31,121,30,88,31,246,31,241,31,50,31,91,31,55,31,55,30,29,31,85,31,142,31,201,31,201,30,149,31,117,31,117,30,152,31,109,31,172,31,170,31,16,31,16,30,177,31,44,31,101,31,92,31,182,31,182,30,182,29,63,31,232,31,68,31,208,31,110,31,118,31,152,31,237,31,237,30,168,31,202,31,96,31,212,31,212,30,112,31,160,31,160,30,160,29,201,31,201,30,148,31,78,31,108,31,136,31,85,31,85,30,85,29,85,28,85,27,203,31,203,30,113,31,45,31,95,31,176,31,227,31,142,31,185,31,185,30,185,29,108,31,138,31,74,31,76,31,80,31,102,31,102,30,39,31,105,31,148,31,173,31,173,30,173,29,125,31,125,30,177,31,98,31,121,31,121,30,194,31,11,31,209,31,37,31,58,31,166,31,52,31,18,31,19,31,67,31,34,31,34,30,125,31,36,31,55,31,35,31,35,30,70,31,8,31,7,31,8,31,47,31,171,31,122,31,227,31,76,31,222,31,222,30,222,29,72,31,163,31,163,30,163,29,202,31,9,31,18,31,95,31,95,30,95,29,205,31,14,31,112,31,1,31,138,31,177,31,48,31,149,31,241,31,210,31,210,30,49,31,246,31,150,31,206,31,222,31,80,31,80,30,229,31,1,31,71,31,199,31,120,31,222,31,123,31,39,31,159,31,206,31,248,31,150,31,93,31,125,31,93,31,146,31,58,31,134,31,190,31,212,31,74,31,74,30,97,31,85,31,15,31,62,31,217,31,236,31,142,31,111,31,16,31,232,31,235,31,235,30,254,31,254,30,61,31,61,30,84,31,112,31,8,31,8,30,8,29,70,31,144,31,184,31,244,31,105,31,156,31,220,31,82,31,71,31,241,31,88,31,88,30,152,31,229,31,109,31,109,30,218,31,235,31,24,31,225,31,187,31,230,31,41,31,41,30,204,31,143,31,17,31,71,31,122,31,133,31,177,31,216,31,252,31,103,31,153,31,162,31,50,31,94,31,89,31,225,31,112,31,112,30,184,31,184,30,184,29,184,28,184,27,60,31,31,31,31,30,136,31,218,31,49,31,143,31,145,31,220,31,220,30,103,31,198,31,49,31,225,31,35,31,224,31,140,31,168,31,127,31,95,31,104,31,244,31,130,31,30,31,224,31,221,31,80,31,35,31,177,31,233,31,94,31,110,31,144,31,63,31,215,31,205,31,80,31,113,31,132,31,241,31,182,31,183,31,42,31,221,31,116,31,251,31,106,31,4,31,220,31,226,31,226,30,65,31,224,31,8,31,252,31,110,31,228,31,228,30,157,31,245,31,103,31,224,31,163,31,163,30,163,29,163,28,239,31,239,30,226,31,230,31,185,31,201,31,79,31,150,31,46,31,249,31,115,31,115,30,56,31,81,31,62,31,97,31,118,31,139,31,82,31,60,31,30,31,30,30,152,31,152,30,233,31,233,30,249,31,249,30,190,31,87,31,120,31,31,31,150,31,112,31,211,31,151,31,221,31,221,30,59,31,201,31,189,31,24,31,62,31,75,31,178,31,47,31,47,30,168,31,168,30,232,31,4,31,72,31,162,31,67,31,232,31,39,31,16,31,133,31,133,30,3,31,90,31,162,31,162,30,162,29,140,31,102,31,255,31,200,31,218,31,122,31,122,30,24,31,147,31,147,30,125,31,208,31,161,31,161,30,161,29,31,31,20,31,159,31,154,31,101,31,85,31,221,31,27,31,62,31,13,31,237,31,174,31,195,31,10,31,105,31,206,31,206,30,206,29,78,31,195,31,189,31,43,31,43,30,85,31,85,30,181,31,141,31,141,30,135,31,111,31,46,31,39,31,172,31,5,31,220,31,36,31,88,31,250,31,250,30,127,31,64,31,76,31,76,30,6,31,60,31,253,31,253,30,88,31,206,31,154,31,177,31,27,31,132,31,142,31,255,31,82,31,98,31,98,30,229,31,240,31,240,30,240,29,180,31,81,31,103,31,44,31,120,31,184,31,184,30,91,31,91,30,214,31,31,31,137,31,40,31,40,30,40,29,40,28,127,31,137,31,241,31,159,31,220,31,220,30,227,31,247,31,166,31,22,31,22,30,22,29,152,31,242,31,241,31,240,31,9,31,9,30,204,31,145,31,160,31,175,31,115,31,16,31,202,31,205,31,205,30,65,31,168,31,214,31,20,31,20,30,253,31,253,30,253,29,89,31,159,31,5,31,113,31,13,31,13,30,13,29,132,31,180,31,146,31,146,30,4,31,249,31,111,31,111,30,136,31,167,31,109,31,225,31,4,31,186,31,151,31,28,31,28,30,42,31,105,31,38,31,162,31,40,31,129,31,141,31,135,31,22,31,140,31,68,31,129,31,157,31,53,31,53,30,162,31,143,31,57,31,41,31,125,31,217,31,221,31,248,31,248,31,248,30,248,29,63,31,197,31,157,31,43,31,79,31,79,30,97,31,186,31,186,30,152,31,123,31,123,30,123,29,123,28,179,31,41,31,41,30,230,31,230,30,43,31,10,31,107,31,131,31,65,31,65,30,114,31,130,31,13,31,65,31,50,31,185,31,57,31,211,31,239,31,207,31,207,30,207,29,98,31,79,31,106,31,155,31,155,30,155,29,245,31,206,31,206,30,239,31,239,30,243,31,68,31,48,31,196,31,222,31,196,31,254,31,102,31,102,30,58,31,58,30,118,31,148,31,148,30,64,31,64,30,124,31,116,31,47,31,225,31,170,31,103,31,27,31,15,31,60,31,36,31,183,31,224,31,160,31,107,31,86,31,241,31,241,30,82,31,177,31,126,31,8,31,8,31,8,30,111,31,40,31,134,31,177,31,177,30,177,29,148,31,92,31,212,31,153,31,153,30,183,31,39,31,212,31,91,31,91,30,14,31,7,31,207,31,207,30,63,31,125,31,66,31,221,31,221,30,230,31,49,31,31,31,128,31,128,31,28,31,28,30,154,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
