-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_795 is
end project_tb_795;

architecture project_tb_arch_795 of project_tb_795 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 452;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (230,0,33,0,0,0,138,0,100,0,15,0,135,0,18,0,148,0,0,0,0,0,0,0,32,0,180,0,217,0,119,0,192,0,227,0,0,0,0,0,230,0,182,0,77,0,6,0,15,0,213,0,109,0,93,0,242,0,165,0,173,0,45,0,205,0,82,0,55,0,198,0,161,0,227,0,30,0,6,0,160,0,33,0,53,0,12,0,113,0,0,0,194,0,0,0,140,0,0,0,86,0,0,0,189,0,16,0,0,0,0,0,90,0,2,0,202,0,0,0,129,0,176,0,89,0,36,0,61,0,238,0,195,0,165,0,237,0,65,0,70,0,174,0,187,0,147,0,0,0,243,0,245,0,29,0,0,0,0,0,236,0,9,0,36,0,0,0,0,0,151,0,0,0,90,0,0,0,221,0,0,0,13,0,134,0,0,0,35,0,0,0,0,0,231,0,163,0,145,0,79,0,28,0,0,0,68,0,207,0,159,0,204,0,141,0,123,0,130,0,0,0,0,0,0,0,83,0,247,0,0,0,196,0,149,0,104,0,197,0,150,0,112,0,210,0,16,0,5,0,10,0,117,0,8,0,121,0,179,0,235,0,112,0,0,0,79,0,79,0,0,0,198,0,74,0,202,0,133,0,19,0,224,0,93,0,18,0,243,0,90,0,80,0,0,0,2,0,0,0,212,0,219,0,111,0,240,0,0,0,110,0,102,0,185,0,39,0,0,0,0,0,126,0,0,0,39,0,99,0,81,0,205,0,0,0,153,0,0,0,110,0,205,0,7,0,228,0,0,0,25,0,68,0,0,0,126,0,137,0,0,0,0,0,79,0,0,0,46,0,158,0,60,0,57,0,112,0,148,0,177,0,230,0,210,0,136,0,36,0,200,0,201,0,29,0,176,0,203,0,240,0,210,0,0,0,14,0,46,0,63,0,214,0,155,0,15,0,0,0,80,0,171,0,130,0,216,0,12,0,147,0,64,0,154,0,253,0,99,0,7,0,113,0,67,0,64,0,120,0,149,0,96,0,210,0,113,0,252,0,8,0,0,0,0,0,23,0,202,0,120,0,157,0,239,0,0,0,65,0,104,0,181,0,71,0,102,0,249,0,0,0,185,0,104,0,248,0,146,0,105,0,0,0,177,0,177,0,49,0,130,0,186,0,62,0,7,0,224,0,88,0,208,0,101,0,3,0,86,0,56,0,132,0,25,0,0,0,232,0,0,0,38,0,0,0,40,0,240,0,173,0,246,0,31,0,126,0,62,0,0,0,215,0,78,0,241,0,39,0,0,0,53,0,226,0,146,0,0,0,238,0,131,0,0,0,233,0,153,0,224,0,246,0,122,0,180,0,125,0,70,0,0,0,176,0,155,0,80,0,31,0,122,0,169,0,1,0,50,0,28,0,153,0,71,0,0,0,218,0,139,0,189,0,18,0,151,0,54,0,113,0,17,0,246,0,0,0,139,0,85,0,228,0,0,0,0,0,145,0,55,0,84,0,96,0,238,0,0,0,237,0,126,0,146,0,194,0,93,0,32,0,110,0,88,0,184,0,0,0,145,0,0,0,227,0,210,0,127,0,221,0,54,0,190,0,204,0,109,0,217,0,24,0,13,0,0,0,108,0,172,0,0,0,75,0,55,0,0,0,108,0,242,0,0,0,0,0,145,0,64,0,0,0,238,0,0,0,176,0,88,0,193,0,0,0,0,0,119,0,0,0,73,0,10,0,0,0,14,0,60,0,62,0,62,0,180,0,0,0,86,0,190,0,235,0,43,0,236,0,19,0,195,0,162,0,56,0,38,0,200,0,142,0,235,0,0,0,65,0,181,0,0,0,8,0,20,0,103,0,194,0,0,0,187,0,26,0,66,0,29,0,0,0,74,0,139,0,106,0,133,0,0,0,113,0,48,0,228,0,53,0,199,0,0,0,31,0,197,0,219,0,30,0,9,0,0,0,203,0,29,0,226,0,117,0,208,0,236,0,0,0,174,0,0,0,15,0,151,0,203,0,40,0,10,0,48,0,0,0,244,0,129,0);
signal scenario_full  : scenario_type := (230,31,33,31,33,30,138,31,100,31,15,31,135,31,18,31,148,31,148,30,148,29,148,28,32,31,180,31,217,31,119,31,192,31,227,31,227,30,227,29,230,31,182,31,77,31,6,31,15,31,213,31,109,31,93,31,242,31,165,31,173,31,45,31,205,31,82,31,55,31,198,31,161,31,227,31,30,31,6,31,160,31,33,31,53,31,12,31,113,31,113,30,194,31,194,30,140,31,140,30,86,31,86,30,189,31,16,31,16,30,16,29,90,31,2,31,202,31,202,30,129,31,176,31,89,31,36,31,61,31,238,31,195,31,165,31,237,31,65,31,70,31,174,31,187,31,147,31,147,30,243,31,245,31,29,31,29,30,29,29,236,31,9,31,36,31,36,30,36,29,151,31,151,30,90,31,90,30,221,31,221,30,13,31,134,31,134,30,35,31,35,30,35,29,231,31,163,31,145,31,79,31,28,31,28,30,68,31,207,31,159,31,204,31,141,31,123,31,130,31,130,30,130,29,130,28,83,31,247,31,247,30,196,31,149,31,104,31,197,31,150,31,112,31,210,31,16,31,5,31,10,31,117,31,8,31,121,31,179,31,235,31,112,31,112,30,79,31,79,31,79,30,198,31,74,31,202,31,133,31,19,31,224,31,93,31,18,31,243,31,90,31,80,31,80,30,2,31,2,30,212,31,219,31,111,31,240,31,240,30,110,31,102,31,185,31,39,31,39,30,39,29,126,31,126,30,39,31,99,31,81,31,205,31,205,30,153,31,153,30,110,31,205,31,7,31,228,31,228,30,25,31,68,31,68,30,126,31,137,31,137,30,137,29,79,31,79,30,46,31,158,31,60,31,57,31,112,31,148,31,177,31,230,31,210,31,136,31,36,31,200,31,201,31,29,31,176,31,203,31,240,31,210,31,210,30,14,31,46,31,63,31,214,31,155,31,15,31,15,30,80,31,171,31,130,31,216,31,12,31,147,31,64,31,154,31,253,31,99,31,7,31,113,31,67,31,64,31,120,31,149,31,96,31,210,31,113,31,252,31,8,31,8,30,8,29,23,31,202,31,120,31,157,31,239,31,239,30,65,31,104,31,181,31,71,31,102,31,249,31,249,30,185,31,104,31,248,31,146,31,105,31,105,30,177,31,177,31,49,31,130,31,186,31,62,31,7,31,224,31,88,31,208,31,101,31,3,31,86,31,56,31,132,31,25,31,25,30,232,31,232,30,38,31,38,30,40,31,240,31,173,31,246,31,31,31,126,31,62,31,62,30,215,31,78,31,241,31,39,31,39,30,53,31,226,31,146,31,146,30,238,31,131,31,131,30,233,31,153,31,224,31,246,31,122,31,180,31,125,31,70,31,70,30,176,31,155,31,80,31,31,31,122,31,169,31,1,31,50,31,28,31,153,31,71,31,71,30,218,31,139,31,189,31,18,31,151,31,54,31,113,31,17,31,246,31,246,30,139,31,85,31,228,31,228,30,228,29,145,31,55,31,84,31,96,31,238,31,238,30,237,31,126,31,146,31,194,31,93,31,32,31,110,31,88,31,184,31,184,30,145,31,145,30,227,31,210,31,127,31,221,31,54,31,190,31,204,31,109,31,217,31,24,31,13,31,13,30,108,31,172,31,172,30,75,31,55,31,55,30,108,31,242,31,242,30,242,29,145,31,64,31,64,30,238,31,238,30,176,31,88,31,193,31,193,30,193,29,119,31,119,30,73,31,10,31,10,30,14,31,60,31,62,31,62,31,180,31,180,30,86,31,190,31,235,31,43,31,236,31,19,31,195,31,162,31,56,31,38,31,200,31,142,31,235,31,235,30,65,31,181,31,181,30,8,31,20,31,103,31,194,31,194,30,187,31,26,31,66,31,29,31,29,30,74,31,139,31,106,31,133,31,133,30,113,31,48,31,228,31,53,31,199,31,199,30,31,31,197,31,219,31,30,31,9,31,9,30,203,31,29,31,226,31,117,31,208,31,236,31,236,30,174,31,174,30,15,31,151,31,203,31,40,31,10,31,48,31,48,30,244,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
