-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 759;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,14,0,101,0,0,0,132,0,209,0,0,0,227,0,156,0,182,0,153,0,20,0,0,0,176,0,183,0,63,0,71,0,242,0,220,0,87,0,229,0,8,0,160,0,32,0,84,0,58,0,208,0,112,0,0,0,241,0,49,0,0,0,29,0,238,0,72,0,19,0,59,0,117,0,235,0,182,0,147,0,102,0,88,0,0,0,0,0,213,0,68,0,210,0,241,0,137,0,67,0,86,0,179,0,79,0,104,0,139,0,210,0,166,0,0,0,68,0,172,0,0,0,95,0,209,0,140,0,55,0,164,0,0,0,252,0,99,0,0,0,251,0,244,0,135,0,45,0,217,0,0,0,46,0,244,0,127,0,0,0,103,0,0,0,165,0,28,0,135,0,140,0,2,0,179,0,115,0,0,0,198,0,244,0,194,0,46,0,254,0,216,0,102,0,88,0,204,0,177,0,243,0,0,0,46,0,0,0,157,0,1,0,74,0,45,0,148,0,0,0,153,0,63,0,126,0,87,0,227,0,199,0,59,0,0,0,242,0,240,0,102,0,145,0,97,0,106,0,184,0,120,0,133,0,161,0,53,0,205,0,176,0,0,0,108,0,219,0,232,0,252,0,174,0,27,0,238,0,68,0,38,0,252,0,66,0,236,0,152,0,132,0,0,0,0,0,172,0,128,0,0,0,183,0,206,0,240,0,94,0,188,0,4,0,47,0,38,0,0,0,238,0,101,0,255,0,241,0,240,0,158,0,3,0,149,0,101,0,76,0,49,0,220,0,174,0,174,0,0,0,217,0,11,0,94,0,239,0,9,0,0,0,182,0,254,0,208,0,255,0,47,0,14,0,97,0,207,0,196,0,224,0,51,0,69,0,3,0,20,0,103,0,161,0,85,0,149,0,0,0,174,0,198,0,170,0,185,0,88,0,9,0,139,0,186,0,114,0,40,0,0,0,83,0,214,0,0,0,213,0,49,0,120,0,202,0,195,0,165,0,157,0,145,0,0,0,244,0,0,0,241,0,132,0,89,0,221,0,110,0,173,0,246,0,242,0,125,0,85,0,180,0,152,0,0,0,191,0,98,0,251,0,0,0,45,0,164,0,221,0,210,0,0,0,89,0,38,0,117,0,63,0,0,0,253,0,169,0,116,0,0,0,80,0,55,0,253,0,166,0,208,0,179,0,217,0,123,0,245,0,207,0,200,0,239,0,200,0,129,0,104,0,243,0,171,0,160,0,192,0,176,0,0,0,65,0,166,0,225,0,145,0,103,0,14,0,25,0,34,0,125,0,43,0,235,0,38,0,201,0,170,0,61,0,0,0,210,0,245,0,63,0,0,0,0,0,117,0,63,0,208,0,204,0,0,0,131,0,163,0,146,0,0,0,18,0,193,0,179,0,171,0,135,0,104,0,0,0,59,0,5,0,7,0,87,0,171,0,205,0,72,0,0,0,34,0,18,0,69,0,181,0,140,0,68,0,165,0,0,0,213,0,0,0,0,0,253,0,1,0,33,0,249,0,0,0,83,0,245,0,23,0,147,0,0,0,123,0,225,0,0,0,84,0,5,0,216,0,154,0,50,0,83,0,85,0,117,0,119,0,191,0,202,0,31,0,31,0,32,0,229,0,78,0,56,0,0,0,251,0,0,0,0,0,248,0,20,0,53,0,208,0,0,0,0,0,146,0,220,0,208,0,106,0,216,0,245,0,0,0,16,0,34,0,97,0,235,0,84,0,113,0,91,0,132,0,113,0,159,0,156,0,207,0,95,0,45,0,164,0,29,0,58,0,236,0,2,0,201,0,0,0,0,0,176,0,28,0,53,0,168,0,0,0,171,0,181,0,146,0,235,0,67,0,231,0,0,0,64,0,147,0,111,0,237,0,10,0,133,0,229,0,41,0,0,0,0,0,131,0,36,0,223,0,9,0,40,0,184,0,17,0,61,0,205,0,170,0,64,0,212,0,26,0,81,0,58,0,247,0,20,0,0,0,150,0,38,0,153,0,109,0,73,0,22,0,0,0,0,0,73,0,203,0,26,0,208,0,149,0,0,0,140,0,43,0,247,0,0,0,200,0,0,0,249,0,52,0,64,0,32,0,247,0,50,0,0,0,236,0,99,0,128,0,144,0,106,0,0,0,154,0,138,0,0,0,207,0,89,0,254,0,11,0,0,0,13,0,24,0,157,0,133,0,41,0,59,0,106,0,31,0,66,0,151,0,48,0,62,0,165,0,220,0,77,0,210,0,209,0,113,0,95,0,161,0,0,0,33,0,41,0,0,0,49,0,237,0,0,0,132,0,154,0,209,0,168,0,20,0,0,0,201,0,112,0,218,0,242,0,0,0,153,0,75,0,53,0,182,0,63,0,181,0,138,0,5,0,214,0,107,0,65,0,94,0,39,0,211,0,98,0,0,0,23,0,94,0,113,0,200,0,219,0,64,0,38,0,62,0,247,0,178,0,0,0,13,0,71,0,26,0,33,0,236,0,226,0,176,0,171,0,77,0,7,0,227,0,0,0,221,0,71,0,112,0,73,0,220,0,238,0,188,0,175,0,232,0,85,0,136,0,0,0,0,0,123,0,45,0,0,0,245,0,15,0,0,0,13,0,187,0,170,0,132,0,22,0,5,0,238,0,39,0,237,0,215,0,127,0,137,0,14,0,176,0,41,0,0,0,47,0,83,0,0,0,168,0,81,0,134,0,0,0,202,0,207,0,83,0,87,0,0,0,242,0,77,0,248,0,54,0,168,0,116,0,0,0,0,0,82,0,100,0,0,0,173,0,162,0,0,0,213,0,214,0,139,0,3,0,72,0,235,0,0,0,170,0,99,0,0,0,241,0,113,0,0,0,0,0,64,0,203,0,0,0,0,0,0,0,32,0,0,0,0,0,234,0,150,0,151,0,23,0,0,0,194,0,97,0,0,0,240,0,199,0,192,0,197,0,50,0,207,0,232,0,126,0,254,0,0,0,133,0,177,0,159,0,85,0,78,0,78,0,80,0,113,0,50,0,178,0,118,0,118,0,115,0,239,0,48,0,228,0,73,0,180,0,50,0,145,0,123,0,166,0,128,0,0,0,205,0,22,0,150,0,90,0,219,0,48,0,237,0,134,0,143,0,143,0,28,0,0,0,42,0,0,0,60,0,39,0,52,0,0,0,247,0,20,0,179,0,181,0,42,0,174,0,126,0,126,0,143,0,22,0,175,0,147,0,0,0,83,0,237,0,101,0,253,0,0,0,33,0,45,0,0,0,74,0,221,0,6,0,55,0,151,0,36,0,0,0,68,0,0,0,0,0,0,0,56,0,239,0,213,0,26,0,3,0,41,0,27,0,188,0,27,0,235,0,226,0,254,0,174,0,96,0,87,0,169,0,145,0,222,0,179,0,91,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,14,31,101,31,101,30,132,31,209,31,209,30,227,31,156,31,182,31,153,31,20,31,20,30,176,31,183,31,63,31,71,31,242,31,220,31,87,31,229,31,8,31,160,31,32,31,84,31,58,31,208,31,112,31,112,30,241,31,49,31,49,30,29,31,238,31,72,31,19,31,59,31,117,31,235,31,182,31,147,31,102,31,88,31,88,30,88,29,213,31,68,31,210,31,241,31,137,31,67,31,86,31,179,31,79,31,104,31,139,31,210,31,166,31,166,30,68,31,172,31,172,30,95,31,209,31,140,31,55,31,164,31,164,30,252,31,99,31,99,30,251,31,244,31,135,31,45,31,217,31,217,30,46,31,244,31,127,31,127,30,103,31,103,30,165,31,28,31,135,31,140,31,2,31,179,31,115,31,115,30,198,31,244,31,194,31,46,31,254,31,216,31,102,31,88,31,204,31,177,31,243,31,243,30,46,31,46,30,157,31,1,31,74,31,45,31,148,31,148,30,153,31,63,31,126,31,87,31,227,31,199,31,59,31,59,30,242,31,240,31,102,31,145,31,97,31,106,31,184,31,120,31,133,31,161,31,53,31,205,31,176,31,176,30,108,31,219,31,232,31,252,31,174,31,27,31,238,31,68,31,38,31,252,31,66,31,236,31,152,31,132,31,132,30,132,29,172,31,128,31,128,30,183,31,206,31,240,31,94,31,188,31,4,31,47,31,38,31,38,30,238,31,101,31,255,31,241,31,240,31,158,31,3,31,149,31,101,31,76,31,49,31,220,31,174,31,174,31,174,30,217,31,11,31,94,31,239,31,9,31,9,30,182,31,254,31,208,31,255,31,47,31,14,31,97,31,207,31,196,31,224,31,51,31,69,31,3,31,20,31,103,31,161,31,85,31,149,31,149,30,174,31,198,31,170,31,185,31,88,31,9,31,139,31,186,31,114,31,40,31,40,30,83,31,214,31,214,30,213,31,49,31,120,31,202,31,195,31,165,31,157,31,145,31,145,30,244,31,244,30,241,31,132,31,89,31,221,31,110,31,173,31,246,31,242,31,125,31,85,31,180,31,152,31,152,30,191,31,98,31,251,31,251,30,45,31,164,31,221,31,210,31,210,30,89,31,38,31,117,31,63,31,63,30,253,31,169,31,116,31,116,30,80,31,55,31,253,31,166,31,208,31,179,31,217,31,123,31,245,31,207,31,200,31,239,31,200,31,129,31,104,31,243,31,171,31,160,31,192,31,176,31,176,30,65,31,166,31,225,31,145,31,103,31,14,31,25,31,34,31,125,31,43,31,235,31,38,31,201,31,170,31,61,31,61,30,210,31,245,31,63,31,63,30,63,29,117,31,63,31,208,31,204,31,204,30,131,31,163,31,146,31,146,30,18,31,193,31,179,31,171,31,135,31,104,31,104,30,59,31,5,31,7,31,87,31,171,31,205,31,72,31,72,30,34,31,18,31,69,31,181,31,140,31,68,31,165,31,165,30,213,31,213,30,213,29,253,31,1,31,33,31,249,31,249,30,83,31,245,31,23,31,147,31,147,30,123,31,225,31,225,30,84,31,5,31,216,31,154,31,50,31,83,31,85,31,117,31,119,31,191,31,202,31,31,31,31,31,32,31,229,31,78,31,56,31,56,30,251,31,251,30,251,29,248,31,20,31,53,31,208,31,208,30,208,29,146,31,220,31,208,31,106,31,216,31,245,31,245,30,16,31,34,31,97,31,235,31,84,31,113,31,91,31,132,31,113,31,159,31,156,31,207,31,95,31,45,31,164,31,29,31,58,31,236,31,2,31,201,31,201,30,201,29,176,31,28,31,53,31,168,31,168,30,171,31,181,31,146,31,235,31,67,31,231,31,231,30,64,31,147,31,111,31,237,31,10,31,133,31,229,31,41,31,41,30,41,29,131,31,36,31,223,31,9,31,40,31,184,31,17,31,61,31,205,31,170,31,64,31,212,31,26,31,81,31,58,31,247,31,20,31,20,30,150,31,38,31,153,31,109,31,73,31,22,31,22,30,22,29,73,31,203,31,26,31,208,31,149,31,149,30,140,31,43,31,247,31,247,30,200,31,200,30,249,31,52,31,64,31,32,31,247,31,50,31,50,30,236,31,99,31,128,31,144,31,106,31,106,30,154,31,138,31,138,30,207,31,89,31,254,31,11,31,11,30,13,31,24,31,157,31,133,31,41,31,59,31,106,31,31,31,66,31,151,31,48,31,62,31,165,31,220,31,77,31,210,31,209,31,113,31,95,31,161,31,161,30,33,31,41,31,41,30,49,31,237,31,237,30,132,31,154,31,209,31,168,31,20,31,20,30,201,31,112,31,218,31,242,31,242,30,153,31,75,31,53,31,182,31,63,31,181,31,138,31,5,31,214,31,107,31,65,31,94,31,39,31,211,31,98,31,98,30,23,31,94,31,113,31,200,31,219,31,64,31,38,31,62,31,247,31,178,31,178,30,13,31,71,31,26,31,33,31,236,31,226,31,176,31,171,31,77,31,7,31,227,31,227,30,221,31,71,31,112,31,73,31,220,31,238,31,188,31,175,31,232,31,85,31,136,31,136,30,136,29,123,31,45,31,45,30,245,31,15,31,15,30,13,31,187,31,170,31,132,31,22,31,5,31,238,31,39,31,237,31,215,31,127,31,137,31,14,31,176,31,41,31,41,30,47,31,83,31,83,30,168,31,81,31,134,31,134,30,202,31,207,31,83,31,87,31,87,30,242,31,77,31,248,31,54,31,168,31,116,31,116,30,116,29,82,31,100,31,100,30,173,31,162,31,162,30,213,31,214,31,139,31,3,31,72,31,235,31,235,30,170,31,99,31,99,30,241,31,113,31,113,30,113,29,64,31,203,31,203,30,203,29,203,28,32,31,32,30,32,29,234,31,150,31,151,31,23,31,23,30,194,31,97,31,97,30,240,31,199,31,192,31,197,31,50,31,207,31,232,31,126,31,254,31,254,30,133,31,177,31,159,31,85,31,78,31,78,31,80,31,113,31,50,31,178,31,118,31,118,31,115,31,239,31,48,31,228,31,73,31,180,31,50,31,145,31,123,31,166,31,128,31,128,30,205,31,22,31,150,31,90,31,219,31,48,31,237,31,134,31,143,31,143,31,28,31,28,30,42,31,42,30,60,31,39,31,52,31,52,30,247,31,20,31,179,31,181,31,42,31,174,31,126,31,126,31,143,31,22,31,175,31,147,31,147,30,83,31,237,31,101,31,253,31,253,30,33,31,45,31,45,30,74,31,221,31,6,31,55,31,151,31,36,31,36,30,68,31,68,30,68,29,68,28,56,31,239,31,213,31,26,31,3,31,41,31,27,31,188,31,27,31,235,31,226,31,254,31,174,31,96,31,87,31,169,31,145,31,222,31,179,31,91,31,91,30,91,29,91,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
