-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 835;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (226,0,78,0,146,0,10,0,140,0,0,0,80,0,195,0,0,0,17,0,47,0,187,0,174,0,0,0,214,0,225,0,31,0,79,0,189,0,141,0,239,0,33,0,197,0,0,0,152,0,146,0,189,0,242,0,244,0,221,0,188,0,119,0,207,0,188,0,248,0,107,0,32,0,42,0,158,0,0,0,54,0,65,0,0,0,141,0,0,0,0,0,237,0,88,0,0,0,87,0,171,0,0,0,128,0,99,0,16,0,49,0,169,0,58,0,244,0,0,0,78,0,144,0,7,0,171,0,0,0,184,0,67,0,137,0,51,0,0,0,22,0,149,0,0,0,22,0,17,0,29,0,250,0,76,0,168,0,192,0,0,0,107,0,0,0,177,0,219,0,6,0,141,0,21,0,183,0,0,0,246,0,28,0,85,0,0,0,185,0,235,0,108,0,0,0,145,0,52,0,255,0,54,0,212,0,101,0,160,0,83,0,213,0,30,0,68,0,113,0,0,0,233,0,205,0,190,0,0,0,206,0,229,0,18,0,173,0,163,0,49,0,232,0,82,0,214,0,0,0,218,0,45,0,7,0,0,0,155,0,0,0,0,0,153,0,0,0,112,0,0,0,70,0,74,0,0,0,99,0,171,0,198,0,0,0,26,0,0,0,0,0,156,0,192,0,214,0,169,0,0,0,0,0,39,0,115,0,226,0,15,0,28,0,242,0,84,0,2,0,163,0,0,0,99,0,91,0,241,0,44,0,182,0,0,0,136,0,53,0,9,0,103,0,46,0,0,0,0,0,9,0,177,0,34,0,177,0,73,0,121,0,184,0,105,0,0,0,53,0,230,0,0,0,161,0,0,0,75,0,136,0,133,0,101,0,211,0,98,0,108,0,197,0,237,0,141,0,42,0,191,0,84,0,9,0,149,0,82,0,0,0,240,0,3,0,219,0,163,0,51,0,0,0,0,0,0,0,48,0,69,0,106,0,26,0,253,0,0,0,234,0,33,0,29,0,91,0,0,0,63,0,207,0,5,0,91,0,241,0,125,0,31,0,31,0,90,0,170,0,11,0,0,0,67,0,0,0,71,0,223,0,151,0,138,0,172,0,229,0,38,0,0,0,58,0,25,0,0,0,105,0,63,0,182,0,54,0,159,0,167,0,0,0,189,0,171,0,0,0,18,0,181,0,191,0,178,0,132,0,237,0,30,0,139,0,130,0,0,0,0,0,57,0,0,0,204,0,217,0,229,0,167,0,59,0,42,0,235,0,0,0,0,0,191,0,0,0,0,0,209,0,0,0,0,0,41,0,109,0,12,0,179,0,99,0,192,0,176,0,23,0,127,0,0,0,0,0,5,0,223,0,0,0,147,0,24,0,96,0,113,0,97,0,0,0,87,0,230,0,127,0,66,0,252,0,74,0,94,0,221,0,64,0,158,0,0,0,0,0,233,0,203,0,51,0,75,0,40,0,24,0,0,0,62,0,18,0,113,0,159,0,0,0,166,0,0,0,154,0,23,0,0,0,0,0,166,0,188,0,0,0,254,0,144,0,68,0,0,0,149,0,118,0,59,0,130,0,0,0,172,0,205,0,157,0,93,0,0,0,10,0,0,0,0,0,109,0,31,0,0,0,89,0,50,0,187,0,113,0,0,0,71,0,34,0,235,0,194,0,247,0,177,0,67,0,107,0,137,0,39,0,244,0,163,0,26,0,229,0,252,0,16,0,61,0,0,0,195,0,0,0,99,0,74,0,240,0,79,0,230,0,66,0,178,0,252,0,31,0,83,0,27,0,0,0,0,0,20,0,241,0,28,0,195,0,165,0,104,0,245,0,64,0,83,0,174,0,32,0,158,0,131,0,219,0,69,0,6,0,180,0,108,0,144,0,0,0,0,0,83,0,0,0,219,0,237,0,0,0,0,0,0,0,172,0,114,0,200,0,129,0,213,0,34,0,210,0,175,0,157,0,114,0,24,0,124,0,0,0,143,0,250,0,209,0,50,0,234,0,63,0,0,0,91,0,48,0,116,0,191,0,209,0,172,0,253,0,176,0,79,0,180,0,101,0,190,0,0,0,46,0,0,0,81,0,43,0,43,0,0,0,1,0,54,0,0,0,0,0,140,0,42,0,75,0,77,0,54,0,44,0,176,0,79,0,58,0,49,0,137,0,82,0,1,0,79,0,131,0,3,0,94,0,130,0,117,0,24,0,149,0,45,0,146,0,141,0,249,0,8,0,168,0,73,0,25,0,0,0,78,0,66,0,166,0,241,0,117,0,160,0,133,0,172,0,238,0,205,0,211,0,0,0,217,0,167,0,94,0,24,0,34,0,0,0,2,0,90,0,251,0,179,0,30,0,0,0,55,0,0,0,120,0,139,0,0,0,35,0,17,0,176,0,0,0,0,0,159,0,139,0,0,0,158,0,106,0,138,0,211,0,82,0,110,0,145,0,209,0,219,0,189,0,199,0,26,0,85,0,11,0,2,0,84,0,0,0,168,0,190,0,167,0,0,0,0,0,211,0,0,0,6,0,237,0,0,0,174,0,118,0,206,0,1,0,0,0,0,0,0,0,113,0,131,0,73,0,69,0,0,0,0,0,182,0,203,0,20,0,0,0,219,0,0,0,83,0,22,0,142,0,138,0,114,0,3,0,243,0,0,0,0,0,155,0,68,0,20,0,129,0,70,0,0,0,135,0,0,0,101,0,159,0,30,0,0,0,192,0,95,0,0,0,205,0,47,0,91,0,0,0,55,0,251,0,237,0,16,0,50,0,99,0,171,0,52,0,87,0,118,0,247,0,249,0,93,0,0,0,155,0,1,0,236,0,245,0,204,0,0,0,52,0,0,0,199,0,235,0,80,0,145,0,66,0,169,0,128,0,21,0,125,0,8,0,88,0,76,0,3,0,57,0,133,0,85,0,211,0,0,0,75,0,129,0,0,0,115,0,153,0,152,0,193,0,173,0,92,0,40,0,46,0,21,0,155,0,224,0,110,0,186,0,215,0,61,0,131,0,207,0,0,0,193,0,18,0,38,0,253,0,168,0,172,0,235,0,0,0,102,0,0,0,189,0,208,0,164,0,0,0,0,0,0,0,61,0,6,0,0,0,61,0,175,0,46,0,0,0,57,0,0,0,180,0,103,0,24,0,239,0,242,0,206,0,252,0,71,0,149,0,240,0,81,0,0,0,70,0,236,0,188,0,194,0,222,0,133,0,28,0,0,0,58,0,48,0,0,0,0,0,168,0,91,0,184,0,82,0,108,0,11,0,3,0,182,0,0,0,147,0,208,0,191,0,0,0,177,0,0,0,110,0,169,0,0,0,40,0,73,0,1,0,60,0,0,0,153,0,120,0,214,0,0,0,176,0,45,0,234,0,194,0,0,0,0,0,3,0,51,0,213,0,102,0,252,0,136,0,4,0,165,0,220,0,243,0,250,0,0,0,0,0,115,0,213,0,203,0,175,0,30,0,0,0,13,0,242,0,13,0,26,0,142,0,115,0,33,0,201,0,172,0,123,0,100,0,86,0,103,0,0,0,205,0,16,0,161,0,24,0,104,0,8,0,38,0,110,0,0,0,45,0,0,0,151,0,45,0,20,0,0,0,195,0,250,0,109,0,129,0,160,0,0,0,0,0,8,0,0,0,188,0,114,0,163,0,34,0,214,0,0,0,115,0,108,0,99,0,0,0,150,0,29,0,160,0,194,0,20,0,55,0,253,0,117,0,60,0,0,0,0,0,14,0,152,0,151,0);
signal scenario_full  : scenario_type := (226,31,78,31,146,31,10,31,140,31,140,30,80,31,195,31,195,30,17,31,47,31,187,31,174,31,174,30,214,31,225,31,31,31,79,31,189,31,141,31,239,31,33,31,197,31,197,30,152,31,146,31,189,31,242,31,244,31,221,31,188,31,119,31,207,31,188,31,248,31,107,31,32,31,42,31,158,31,158,30,54,31,65,31,65,30,141,31,141,30,141,29,237,31,88,31,88,30,87,31,171,31,171,30,128,31,99,31,16,31,49,31,169,31,58,31,244,31,244,30,78,31,144,31,7,31,171,31,171,30,184,31,67,31,137,31,51,31,51,30,22,31,149,31,149,30,22,31,17,31,29,31,250,31,76,31,168,31,192,31,192,30,107,31,107,30,177,31,219,31,6,31,141,31,21,31,183,31,183,30,246,31,28,31,85,31,85,30,185,31,235,31,108,31,108,30,145,31,52,31,255,31,54,31,212,31,101,31,160,31,83,31,213,31,30,31,68,31,113,31,113,30,233,31,205,31,190,31,190,30,206,31,229,31,18,31,173,31,163,31,49,31,232,31,82,31,214,31,214,30,218,31,45,31,7,31,7,30,155,31,155,30,155,29,153,31,153,30,112,31,112,30,70,31,74,31,74,30,99,31,171,31,198,31,198,30,26,31,26,30,26,29,156,31,192,31,214,31,169,31,169,30,169,29,39,31,115,31,226,31,15,31,28,31,242,31,84,31,2,31,163,31,163,30,99,31,91,31,241,31,44,31,182,31,182,30,136,31,53,31,9,31,103,31,46,31,46,30,46,29,9,31,177,31,34,31,177,31,73,31,121,31,184,31,105,31,105,30,53,31,230,31,230,30,161,31,161,30,75,31,136,31,133,31,101,31,211,31,98,31,108,31,197,31,237,31,141,31,42,31,191,31,84,31,9,31,149,31,82,31,82,30,240,31,3,31,219,31,163,31,51,31,51,30,51,29,51,28,48,31,69,31,106,31,26,31,253,31,253,30,234,31,33,31,29,31,91,31,91,30,63,31,207,31,5,31,91,31,241,31,125,31,31,31,31,31,90,31,170,31,11,31,11,30,67,31,67,30,71,31,223,31,151,31,138,31,172,31,229,31,38,31,38,30,58,31,25,31,25,30,105,31,63,31,182,31,54,31,159,31,167,31,167,30,189,31,171,31,171,30,18,31,181,31,191,31,178,31,132,31,237,31,30,31,139,31,130,31,130,30,130,29,57,31,57,30,204,31,217,31,229,31,167,31,59,31,42,31,235,31,235,30,235,29,191,31,191,30,191,29,209,31,209,30,209,29,41,31,109,31,12,31,179,31,99,31,192,31,176,31,23,31,127,31,127,30,127,29,5,31,223,31,223,30,147,31,24,31,96,31,113,31,97,31,97,30,87,31,230,31,127,31,66,31,252,31,74,31,94,31,221,31,64,31,158,31,158,30,158,29,233,31,203,31,51,31,75,31,40,31,24,31,24,30,62,31,18,31,113,31,159,31,159,30,166,31,166,30,154,31,23,31,23,30,23,29,166,31,188,31,188,30,254,31,144,31,68,31,68,30,149,31,118,31,59,31,130,31,130,30,172,31,205,31,157,31,93,31,93,30,10,31,10,30,10,29,109,31,31,31,31,30,89,31,50,31,187,31,113,31,113,30,71,31,34,31,235,31,194,31,247,31,177,31,67,31,107,31,137,31,39,31,244,31,163,31,26,31,229,31,252,31,16,31,61,31,61,30,195,31,195,30,99,31,74,31,240,31,79,31,230,31,66,31,178,31,252,31,31,31,83,31,27,31,27,30,27,29,20,31,241,31,28,31,195,31,165,31,104,31,245,31,64,31,83,31,174,31,32,31,158,31,131,31,219,31,69,31,6,31,180,31,108,31,144,31,144,30,144,29,83,31,83,30,219,31,237,31,237,30,237,29,237,28,172,31,114,31,200,31,129,31,213,31,34,31,210,31,175,31,157,31,114,31,24,31,124,31,124,30,143,31,250,31,209,31,50,31,234,31,63,31,63,30,91,31,48,31,116,31,191,31,209,31,172,31,253,31,176,31,79,31,180,31,101,31,190,31,190,30,46,31,46,30,81,31,43,31,43,31,43,30,1,31,54,31,54,30,54,29,140,31,42,31,75,31,77,31,54,31,44,31,176,31,79,31,58,31,49,31,137,31,82,31,1,31,79,31,131,31,3,31,94,31,130,31,117,31,24,31,149,31,45,31,146,31,141,31,249,31,8,31,168,31,73,31,25,31,25,30,78,31,66,31,166,31,241,31,117,31,160,31,133,31,172,31,238,31,205,31,211,31,211,30,217,31,167,31,94,31,24,31,34,31,34,30,2,31,90,31,251,31,179,31,30,31,30,30,55,31,55,30,120,31,139,31,139,30,35,31,17,31,176,31,176,30,176,29,159,31,139,31,139,30,158,31,106,31,138,31,211,31,82,31,110,31,145,31,209,31,219,31,189,31,199,31,26,31,85,31,11,31,2,31,84,31,84,30,168,31,190,31,167,31,167,30,167,29,211,31,211,30,6,31,237,31,237,30,174,31,118,31,206,31,1,31,1,30,1,29,1,28,113,31,131,31,73,31,69,31,69,30,69,29,182,31,203,31,20,31,20,30,219,31,219,30,83,31,22,31,142,31,138,31,114,31,3,31,243,31,243,30,243,29,155,31,68,31,20,31,129,31,70,31,70,30,135,31,135,30,101,31,159,31,30,31,30,30,192,31,95,31,95,30,205,31,47,31,91,31,91,30,55,31,251,31,237,31,16,31,50,31,99,31,171,31,52,31,87,31,118,31,247,31,249,31,93,31,93,30,155,31,1,31,236,31,245,31,204,31,204,30,52,31,52,30,199,31,235,31,80,31,145,31,66,31,169,31,128,31,21,31,125,31,8,31,88,31,76,31,3,31,57,31,133,31,85,31,211,31,211,30,75,31,129,31,129,30,115,31,153,31,152,31,193,31,173,31,92,31,40,31,46,31,21,31,155,31,224,31,110,31,186,31,215,31,61,31,131,31,207,31,207,30,193,31,18,31,38,31,253,31,168,31,172,31,235,31,235,30,102,31,102,30,189,31,208,31,164,31,164,30,164,29,164,28,61,31,6,31,6,30,61,31,175,31,46,31,46,30,57,31,57,30,180,31,103,31,24,31,239,31,242,31,206,31,252,31,71,31,149,31,240,31,81,31,81,30,70,31,236,31,188,31,194,31,222,31,133,31,28,31,28,30,58,31,48,31,48,30,48,29,168,31,91,31,184,31,82,31,108,31,11,31,3,31,182,31,182,30,147,31,208,31,191,31,191,30,177,31,177,30,110,31,169,31,169,30,40,31,73,31,1,31,60,31,60,30,153,31,120,31,214,31,214,30,176,31,45,31,234,31,194,31,194,30,194,29,3,31,51,31,213,31,102,31,252,31,136,31,4,31,165,31,220,31,243,31,250,31,250,30,250,29,115,31,213,31,203,31,175,31,30,31,30,30,13,31,242,31,13,31,26,31,142,31,115,31,33,31,201,31,172,31,123,31,100,31,86,31,103,31,103,30,205,31,16,31,161,31,24,31,104,31,8,31,38,31,110,31,110,30,45,31,45,30,151,31,45,31,20,31,20,30,195,31,250,31,109,31,129,31,160,31,160,30,160,29,8,31,8,30,188,31,114,31,163,31,34,31,214,31,214,30,115,31,108,31,99,31,99,30,150,31,29,31,160,31,194,31,20,31,55,31,253,31,117,31,60,31,60,30,60,29,14,31,152,31,151,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
