-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 976;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (14,0,88,0,250,0,153,0,127,0,135,0,251,0,0,0,218,0,87,0,199,0,28,0,150,0,115,0,0,0,75,0,0,0,230,0,114,0,254,0,142,0,96,0,0,0,0,0,0,0,129,0,41,0,2,0,101,0,221,0,199,0,177,0,31,0,30,0,205,0,51,0,106,0,0,0,63,0,0,0,0,0,88,0,0,0,110,0,170,0,180,0,238,0,135,0,0,0,0,0,245,0,35,0,60,0,0,0,84,0,65,0,242,0,0,0,87,0,226,0,141,0,85,0,62,0,193,0,0,0,51,0,0,0,189,0,228,0,0,0,64,0,250,0,75,0,168,0,102,0,220,0,144,0,249,0,6,0,236,0,0,0,26,0,0,0,78,0,168,0,242,0,159,0,27,0,234,0,71,0,125,0,82,0,100,0,68,0,167,0,204,0,69,0,0,0,66,0,99,0,150,0,130,0,245,0,75,0,0,0,91,0,200,0,0,0,0,0,51,0,0,0,111,0,217,0,166,0,0,0,179,0,212,0,211,0,74,0,141,0,0,0,224,0,159,0,77,0,208,0,0,0,109,0,39,0,0,0,127,0,103,0,97,0,148,0,70,0,16,0,0,0,46,0,77,0,30,0,223,0,86,0,58,0,0,0,0,0,62,0,239,0,132,0,84,0,0,0,49,0,81,0,0,0,0,0,101,0,10,0,183,0,0,0,199,0,0,0,25,0,246,0,75,0,139,0,67,0,158,0,249,0,55,0,168,0,0,0,36,0,84,0,138,0,0,0,0,0,190,0,241,0,165,0,172,0,0,0,135,0,73,0,0,0,0,0,129,0,31,0,0,0,122,0,251,0,0,0,186,0,173,0,153,0,197,0,2,0,224,0,69,0,70,0,95,0,0,0,201,0,118,0,242,0,0,0,196,0,0,0,49,0,187,0,0,0,212,0,91,0,37,0,121,0,20,0,0,0,0,0,10,0,0,0,3,0,123,0,0,0,102,0,40,0,119,0,37,0,203,0,134,0,80,0,0,0,183,0,197,0,84,0,109,0,146,0,148,0,117,0,0,0,112,0,192,0,237,0,0,0,0,0,9,0,74,0,199,0,164,0,42,0,104,0,249,0,230,0,95,0,244,0,251,0,0,0,179,0,151,0,27,0,247,0,60,0,0,0,88,0,0,0,0,0,183,0,183,0,233,0,0,0,136,0,127,0,96,0,52,0,60,0,7,0,82,0,0,0,22,0,10,0,111,0,39,0,219,0,1,0,100,0,22,0,18,0,215,0,23,0,12,0,0,0,106,0,104,0,51,0,107,0,124,0,58,0,40,0,42,0,22,0,212,0,0,0,0,0,237,0,26,0,187,0,199,0,90,0,81,0,55,0,64,0,41,0,124,0,0,0,9,0,8,0,162,0,138,0,26,0,233,0,102,0,173,0,149,0,221,0,122,0,167,0,159,0,198,0,2,0,184,0,193,0,0,0,7,0,147,0,0,0,202,0,78,0,157,0,29,0,0,0,71,0,0,0,250,0,66,0,230,0,201,0,204,0,176,0,210,0,173,0,136,0,56,0,138,0,44,0,236,0,0,0,92,0,0,0,152,0,85,0,6,0,203,0,0,0,249,0,0,0,0,0,64,0,255,0,0,0,208,0,0,0,116,0,243,0,221,0,236,0,173,0,42,0,186,0,56,0,98,0,0,0,191,0,0,0,0,0,0,0,51,0,91,0,0,0,0,0,144,0,42,0,36,0,213,0,80,0,12,0,229,0,0,0,4,0,0,0,36,0,0,0,154,0,51,0,207,0,138,0,0,0,159,0,200,0,166,0,0,0,113,0,210,0,202,0,157,0,101,0,158,0,58,0,4,0,64,0,81,0,44,0,190,0,58,0,225,0,0,0,0,0,221,0,161,0,0,0,245,0,212,0,254,0,27,0,8,0,49,0,239,0,247,0,58,0,0,0,0,0,150,0,234,0,208,0,143,0,0,0,0,0,81,0,0,0,99,0,240,0,151,0,212,0,121,0,0,0,12,0,24,0,223,0,0,0,0,0,0,0,157,0,193,0,106,0,69,0,98,0,243,0,0,0,58,0,191,0,0,0,164,0,149,0,249,0,12,0,158,0,0,0,78,0,37,0,227,0,0,0,78,0,13,0,246,0,71,0,118,0,0,0,233,0,197,0,235,0,123,0,205,0,60,0,241,0,121,0,63,0,219,0,227,0,24,0,171,0,189,0,40,0,0,0,0,0,169,0,134,0,239,0,161,0,101,0,117,0,19,0,201,0,27,0,88,0,248,0,140,0,0,0,215,0,59,0,5,0,0,0,41,0,125,0,16,0,195,0,251,0,0,0,36,0,244,0,3,0,0,0,41,0,186,0,106,0,0,0,44,0,213,0,114,0,168,0,0,0,166,0,145,0,187,0,192,0,210,0,74,0,150,0,254,0,151,0,250,0,125,0,42,0,191,0,0,0,233,0,243,0,167,0,168,0,124,0,0,0,19,0,228,0,0,0,55,0,12,0,136,0,193,0,139,0,52,0,185,0,9,0,43,0,0,0,119,0,210,0,130,0,96,0,73,0,68,0,178,0,197,0,21,0,115,0,0,0,199,0,246,0,0,0,121,0,5,0,0,0,242,0,153,0,53,0,0,0,168,0,172,0,223,0,89,0,80,0,244,0,93,0,108,0,109,0,69,0,0,0,233,0,26,0,63,0,0,0,114,0,0,0,0,0,238,0,109,0,230,0,0,0,0,0,41,0,58,0,54,0,177,0,0,0,1,0,169,0,10,0,77,0,0,0,14,0,51,0,186,0,14,0,0,0,0,0,140,0,0,0,0,0,0,0,41,0,0,0,61,0,109,0,36,0,194,0,139,0,188,0,244,0,0,0,104,0,204,0,0,0,188,0,0,0,242,0,138,0,219,0,0,0,179,0,0,0,0,0,161,0,0,0,203,0,23,0,180,0,102,0,120,0,255,0,158,0,141,0,66,0,193,0,177,0,73,0,189,0,247,0,134,0,146,0,178,0,0,0,238,0,125,0,97,0,62,0,234,0,206,0,242,0,63,0,14,0,254,0,0,0,50,0,45,0,96,0,245,0,245,0,245,0,110,0,186,0,0,0,0,0,134,0,0,0,123,0,147,0,243,0,0,0,252,0,126,0,128,0,5,0,171,0,66,0,148,0,47,0,87,0,243,0,77,0,220,0,230,0,195,0,41,0,89,0,32,0,184,0,93,0,255,0,139,0,9,0,92,0,201,0,221,0,99,0,108,0,224,0,193,0,0,0,69,0,16,0,42,0,217,0,96,0,84,0,101,0,145,0,167,0,0,0,195,0,12,0,150,0,71,0,21,0,0,0,62,0,32,0,104,0,14,0,109,0,103,0,0,0,135,0,93,0,225,0,100,0,145,0,172,0,211,0,30,0,143,0,0,0,109,0,225,0,2,0,105,0,0,0,18,0,155,0,11,0,11,0,151,0,135,0,174,0,0,0,43,0,206,0,40,0,190,0,251,0,0,0,0,0,219,0,31,0,0,0,42,0,108,0,100,0,21,0,0,0,149,0,186,0,89,0,1,0,80,0,148,0,0,0,63,0,0,0,176,0,168,0,163,0,72,0,243,0,70,0,35,0,122,0,206,0,1,0,0,0,56,0,206,0,0,0,0,0,62,0,104,0,109,0,83,0,0,0,0,0,83,0,0,0,0,0,96,0,119,0,0,0,207,0,151,0,177,0,0,0,190,0,153,0,0,0,14,0,245,0,0,0,0,0,40,0,128,0,10,0,60,0,150,0,56,0,146,0,83,0,58,0,195,0,52,0,44,0,250,0,155,0,134,0,101,0,35,0,19,0,201,0,30,0,4,0,0,0,0,0,0,0,110,0,14,0,133,0,0,0,53,0,148,0,0,0,98,0,126,0,174,0,110,0,0,0,42,0,89,0,21,0,0,0,0,0,213,0,127,0,67,0,115,0,0,0,230,0,27,0,200,0,5,0,71,0,16,0,93,0,0,0,197,0,127,0,242,0,203,0,0,0,208,0,0,0,85,0,46,0,0,0,0,0,12,0,0,0,203,0,0,0,146,0,224,0,96,0,33,0,60,0,143,0,0,0,0,0,42,0,79,0,227,0,186,0,0,0,169,0,141,0,178,0,176,0,82,0,220,0,202,0,118,0,102,0,70,0,241,0,7,0,203,0,1,0,0,0,195,0,29,0,14,0,179,0,240,0,253,0,7,0,0,0,0,0,248,0,112,0,249,0,237,0,54,0,85,0,0,0,69,0,224,0,7,0,65,0,10,0,0,0,96,0,108,0,0,0,0,0,0,0,0,0,168,0,0,0,0,0,55,0,165,0,98,0,186,0,211,0,132,0,78,0,129,0,106,0);
signal scenario_full  : scenario_type := (14,31,88,31,250,31,153,31,127,31,135,31,251,31,251,30,218,31,87,31,199,31,28,31,150,31,115,31,115,30,75,31,75,30,230,31,114,31,254,31,142,31,96,31,96,30,96,29,96,28,129,31,41,31,2,31,101,31,221,31,199,31,177,31,31,31,30,31,205,31,51,31,106,31,106,30,63,31,63,30,63,29,88,31,88,30,110,31,170,31,180,31,238,31,135,31,135,30,135,29,245,31,35,31,60,31,60,30,84,31,65,31,242,31,242,30,87,31,226,31,141,31,85,31,62,31,193,31,193,30,51,31,51,30,189,31,228,31,228,30,64,31,250,31,75,31,168,31,102,31,220,31,144,31,249,31,6,31,236,31,236,30,26,31,26,30,78,31,168,31,242,31,159,31,27,31,234,31,71,31,125,31,82,31,100,31,68,31,167,31,204,31,69,31,69,30,66,31,99,31,150,31,130,31,245,31,75,31,75,30,91,31,200,31,200,30,200,29,51,31,51,30,111,31,217,31,166,31,166,30,179,31,212,31,211,31,74,31,141,31,141,30,224,31,159,31,77,31,208,31,208,30,109,31,39,31,39,30,127,31,103,31,97,31,148,31,70,31,16,31,16,30,46,31,77,31,30,31,223,31,86,31,58,31,58,30,58,29,62,31,239,31,132,31,84,31,84,30,49,31,81,31,81,30,81,29,101,31,10,31,183,31,183,30,199,31,199,30,25,31,246,31,75,31,139,31,67,31,158,31,249,31,55,31,168,31,168,30,36,31,84,31,138,31,138,30,138,29,190,31,241,31,165,31,172,31,172,30,135,31,73,31,73,30,73,29,129,31,31,31,31,30,122,31,251,31,251,30,186,31,173,31,153,31,197,31,2,31,224,31,69,31,70,31,95,31,95,30,201,31,118,31,242,31,242,30,196,31,196,30,49,31,187,31,187,30,212,31,91,31,37,31,121,31,20,31,20,30,20,29,10,31,10,30,3,31,123,31,123,30,102,31,40,31,119,31,37,31,203,31,134,31,80,31,80,30,183,31,197,31,84,31,109,31,146,31,148,31,117,31,117,30,112,31,192,31,237,31,237,30,237,29,9,31,74,31,199,31,164,31,42,31,104,31,249,31,230,31,95,31,244,31,251,31,251,30,179,31,151,31,27,31,247,31,60,31,60,30,88,31,88,30,88,29,183,31,183,31,233,31,233,30,136,31,127,31,96,31,52,31,60,31,7,31,82,31,82,30,22,31,10,31,111,31,39,31,219,31,1,31,100,31,22,31,18,31,215,31,23,31,12,31,12,30,106,31,104,31,51,31,107,31,124,31,58,31,40,31,42,31,22,31,212,31,212,30,212,29,237,31,26,31,187,31,199,31,90,31,81,31,55,31,64,31,41,31,124,31,124,30,9,31,8,31,162,31,138,31,26,31,233,31,102,31,173,31,149,31,221,31,122,31,167,31,159,31,198,31,2,31,184,31,193,31,193,30,7,31,147,31,147,30,202,31,78,31,157,31,29,31,29,30,71,31,71,30,250,31,66,31,230,31,201,31,204,31,176,31,210,31,173,31,136,31,56,31,138,31,44,31,236,31,236,30,92,31,92,30,152,31,85,31,6,31,203,31,203,30,249,31,249,30,249,29,64,31,255,31,255,30,208,31,208,30,116,31,243,31,221,31,236,31,173,31,42,31,186,31,56,31,98,31,98,30,191,31,191,30,191,29,191,28,51,31,91,31,91,30,91,29,144,31,42,31,36,31,213,31,80,31,12,31,229,31,229,30,4,31,4,30,36,31,36,30,154,31,51,31,207,31,138,31,138,30,159,31,200,31,166,31,166,30,113,31,210,31,202,31,157,31,101,31,158,31,58,31,4,31,64,31,81,31,44,31,190,31,58,31,225,31,225,30,225,29,221,31,161,31,161,30,245,31,212,31,254,31,27,31,8,31,49,31,239,31,247,31,58,31,58,30,58,29,150,31,234,31,208,31,143,31,143,30,143,29,81,31,81,30,99,31,240,31,151,31,212,31,121,31,121,30,12,31,24,31,223,31,223,30,223,29,223,28,157,31,193,31,106,31,69,31,98,31,243,31,243,30,58,31,191,31,191,30,164,31,149,31,249,31,12,31,158,31,158,30,78,31,37,31,227,31,227,30,78,31,13,31,246,31,71,31,118,31,118,30,233,31,197,31,235,31,123,31,205,31,60,31,241,31,121,31,63,31,219,31,227,31,24,31,171,31,189,31,40,31,40,30,40,29,169,31,134,31,239,31,161,31,101,31,117,31,19,31,201,31,27,31,88,31,248,31,140,31,140,30,215,31,59,31,5,31,5,30,41,31,125,31,16,31,195,31,251,31,251,30,36,31,244,31,3,31,3,30,41,31,186,31,106,31,106,30,44,31,213,31,114,31,168,31,168,30,166,31,145,31,187,31,192,31,210,31,74,31,150,31,254,31,151,31,250,31,125,31,42,31,191,31,191,30,233,31,243,31,167,31,168,31,124,31,124,30,19,31,228,31,228,30,55,31,12,31,136,31,193,31,139,31,52,31,185,31,9,31,43,31,43,30,119,31,210,31,130,31,96,31,73,31,68,31,178,31,197,31,21,31,115,31,115,30,199,31,246,31,246,30,121,31,5,31,5,30,242,31,153,31,53,31,53,30,168,31,172,31,223,31,89,31,80,31,244,31,93,31,108,31,109,31,69,31,69,30,233,31,26,31,63,31,63,30,114,31,114,30,114,29,238,31,109,31,230,31,230,30,230,29,41,31,58,31,54,31,177,31,177,30,1,31,169,31,10,31,77,31,77,30,14,31,51,31,186,31,14,31,14,30,14,29,140,31,140,30,140,29,140,28,41,31,41,30,61,31,109,31,36,31,194,31,139,31,188,31,244,31,244,30,104,31,204,31,204,30,188,31,188,30,242,31,138,31,219,31,219,30,179,31,179,30,179,29,161,31,161,30,203,31,23,31,180,31,102,31,120,31,255,31,158,31,141,31,66,31,193,31,177,31,73,31,189,31,247,31,134,31,146,31,178,31,178,30,238,31,125,31,97,31,62,31,234,31,206,31,242,31,63,31,14,31,254,31,254,30,50,31,45,31,96,31,245,31,245,31,245,31,110,31,186,31,186,30,186,29,134,31,134,30,123,31,147,31,243,31,243,30,252,31,126,31,128,31,5,31,171,31,66,31,148,31,47,31,87,31,243,31,77,31,220,31,230,31,195,31,41,31,89,31,32,31,184,31,93,31,255,31,139,31,9,31,92,31,201,31,221,31,99,31,108,31,224,31,193,31,193,30,69,31,16,31,42,31,217,31,96,31,84,31,101,31,145,31,167,31,167,30,195,31,12,31,150,31,71,31,21,31,21,30,62,31,32,31,104,31,14,31,109,31,103,31,103,30,135,31,93,31,225,31,100,31,145,31,172,31,211,31,30,31,143,31,143,30,109,31,225,31,2,31,105,31,105,30,18,31,155,31,11,31,11,31,151,31,135,31,174,31,174,30,43,31,206,31,40,31,190,31,251,31,251,30,251,29,219,31,31,31,31,30,42,31,108,31,100,31,21,31,21,30,149,31,186,31,89,31,1,31,80,31,148,31,148,30,63,31,63,30,176,31,168,31,163,31,72,31,243,31,70,31,35,31,122,31,206,31,1,31,1,30,56,31,206,31,206,30,206,29,62,31,104,31,109,31,83,31,83,30,83,29,83,31,83,30,83,29,96,31,119,31,119,30,207,31,151,31,177,31,177,30,190,31,153,31,153,30,14,31,245,31,245,30,245,29,40,31,128,31,10,31,60,31,150,31,56,31,146,31,83,31,58,31,195,31,52,31,44,31,250,31,155,31,134,31,101,31,35,31,19,31,201,31,30,31,4,31,4,30,4,29,4,28,110,31,14,31,133,31,133,30,53,31,148,31,148,30,98,31,126,31,174,31,110,31,110,30,42,31,89,31,21,31,21,30,21,29,213,31,127,31,67,31,115,31,115,30,230,31,27,31,200,31,5,31,71,31,16,31,93,31,93,30,197,31,127,31,242,31,203,31,203,30,208,31,208,30,85,31,46,31,46,30,46,29,12,31,12,30,203,31,203,30,146,31,224,31,96,31,33,31,60,31,143,31,143,30,143,29,42,31,79,31,227,31,186,31,186,30,169,31,141,31,178,31,176,31,82,31,220,31,202,31,118,31,102,31,70,31,241,31,7,31,203,31,1,31,1,30,195,31,29,31,14,31,179,31,240,31,253,31,7,31,7,30,7,29,248,31,112,31,249,31,237,31,54,31,85,31,85,30,69,31,224,31,7,31,65,31,10,31,10,30,96,31,108,31,108,30,108,29,108,28,108,27,168,31,168,30,168,29,55,31,165,31,98,31,186,31,211,31,132,31,78,31,129,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
