-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 797;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (80,0,117,0,96,0,17,0,214,0,251,0,148,0,150,0,123,0,0,0,40,0,93,0,65,0,253,0,217,0,22,0,210,0,166,0,0,0,72,0,0,0,53,0,178,0,20,0,243,0,112,0,15,0,194,0,69,0,217,0,0,0,216,0,0,0,0,0,219,0,196,0,155,0,195,0,90,0,0,0,94,0,38,0,120,0,37,0,66,0,230,0,156,0,0,0,104,0,0,0,139,0,190,0,0,0,205,0,14,0,238,0,0,0,147,0,9,0,0,0,11,0,192,0,0,0,194,0,170,0,0,0,0,0,60,0,68,0,227,0,0,0,61,0,133,0,0,0,0,0,0,0,254,0,148,0,55,0,97,0,33,0,17,0,110,0,250,0,216,0,117,0,143,0,0,0,147,0,42,0,202,0,0,0,146,0,102,0,162,0,19,0,0,0,74,0,48,0,43,0,81,0,107,0,0,0,0,0,150,0,0,0,0,0,29,0,211,0,209,0,70,0,37,0,60,0,243,0,0,0,66,0,74,0,30,0,80,0,247,0,251,0,178,0,96,0,210,0,106,0,181,0,200,0,191,0,93,0,18,0,191,0,0,0,41,0,73,0,0,0,255,0,59,0,175,0,235,0,98,0,0,0,230,0,251,0,0,0,197,0,51,0,0,0,95,0,0,0,229,0,254,0,0,0,196,0,0,0,255,0,48,0,58,0,201,0,69,0,49,0,151,0,118,0,0,0,149,0,206,0,0,0,0,0,23,0,0,0,0,0,69,0,0,0,114,0,118,0,0,0,0,0,105,0,0,0,183,0,77,0,13,0,53,0,198,0,148,0,0,0,25,0,13,0,220,0,115,0,19,0,61,0,0,0,0,0,229,0,118,0,21,0,219,0,161,0,37,0,38,0,109,0,58,0,0,0,30,0,215,0,192,0,0,0,183,0,187,0,0,0,159,0,204,0,220,0,0,0,48,0,242,0,18,0,234,0,107,0,184,0,232,0,101,0,0,0,27,0,75,0,154,0,77,0,34,0,0,0,77,0,141,0,250,0,239,0,124,0,0,0,0,0,115,0,70,0,81,0,139,0,130,0,34,0,129,0,213,0,46,0,200,0,110,0,32,0,84,0,0,0,206,0,163,0,27,0,149,0,0,0,223,0,28,0,165,0,171,0,0,0,83,0,182,0,143,0,196,0,31,0,226,0,146,0,0,0,0,0,0,0,160,0,208,0,174,0,121,0,155,0,0,0,93,0,140,0,74,0,73,0,175,0,21,0,0,0,0,0,185,0,148,0,151,0,180,0,35,0,0,0,109,0,41,0,16,0,136,0,117,0,210,0,132,0,0,0,9,0,27,0,245,0,155,0,194,0,0,0,48,0,180,0,126,0,13,0,221,0,0,0,34,0,167,0,0,0,77,0,138,0,0,0,211,0,117,0,156,0,58,0,83,0,183,0,198,0,63,0,0,0,98,0,89,0,0,0,0,0,254,0,85,0,224,0,68,0,209,0,45,0,69,0,238,0,102,0,124,0,7,0,7,0,0,0,113,0,0,0,31,0,214,0,5,0,32,0,162,0,196,0,65,0,28,0,209,0,189,0,0,0,0,0,71,0,99,0,97,0,123,0,246,0,72,0,0,0,244,0,164,0,0,0,122,0,48,0,118,0,211,0,238,0,40,0,175,0,8,0,0,0,0,0,89,0,75,0,0,0,114,0,237,0,0,0,132,0,123,0,30,0,195,0,178,0,0,0,213,0,0,0,165,0,0,0,173,0,235,0,169,0,205,0,127,0,76,0,24,0,52,0,220,0,112,0,0,0,48,0,31,0,242,0,224,0,0,0,226,0,22,0,232,0,142,0,128,0,117,0,196,0,0,0,0,0,142,0,142,0,111,0,0,0,231,0,158,0,253,0,77,0,154,0,243,0,0,0,0,0,53,0,126,0,101,0,97,0,121,0,127,0,60,0,243,0,23,0,14,0,0,0,141,0,0,0,80,0,160,0,165,0,204,0,0,0,188,0,198,0,228,0,161,0,62,0,111,0,139,0,0,0,0,0,175,0,0,0,145,0,62,0,6,0,153,0,42,0,65,0,159,0,0,0,0,0,8,0,128,0,85,0,156,0,209,0,236,0,122,0,249,0,158,0,99,0,172,0,0,0,57,0,0,0,95,0,0,0,0,0,0,0,102,0,225,0,115,0,234,0,133,0,49,0,86,0,134,0,152,0,170,0,149,0,249,0,23,0,47,0,0,0,17,0,194,0,238,0,0,0,197,0,124,0,239,0,23,0,95,0,0,0,162,0,170,0,163,0,35,0,0,0,174,0,0,0,32,0,97,0,160,0,0,0,127,0,251,0,190,0,55,0,83,0,100,0,36,0,160,0,135,0,0,0,0,0,63,0,106,0,117,0,6,0,216,0,45,0,35,0,33,0,146,0,137,0,92,0,0,0,56,0,10,0,166,0,74,0,178,0,0,0,185,0,0,0,38,0,0,0,203,0,2,0,187,0,0,0,0,0,117,0,213,0,19,0,21,0,175,0,51,0,128,0,167,0,0,0,93,0,22,0,0,0,152,0,0,0,12,0,154,0,95,0,96,0,157,0,57,0,243,0,223,0,12,0,0,0,143,0,99,0,0,0,0,0,150,0,235,0,139,0,56,0,170,0,108,0,185,0,0,0,248,0,0,0,151,0,45,0,26,0,238,0,142,0,159,0,185,0,233,0,0,0,169,0,0,0,193,0,186,0,0,0,148,0,112,0,165,0,112,0,67,0,38,0,99,0,94,0,0,0,0,0,55,0,68,0,184,0,136,0,157,0,0,0,152,0,178,0,7,0,240,0,0,0,83,0,122,0,99,0,156,0,164,0,59,0,108,0,151,0,7,0,141,0,4,0,248,0,56,0,93,0,0,0,189,0,13,0,0,0,216,0,98,0,81,0,0,0,0,0,149,0,231,0,170,0,240,0,44,0,226,0,11,0,133,0,151,0,91,0,9,0,75,0,251,0,75,0,235,0,0,0,0,0,0,0,162,0,0,0,195,0,0,0,0,0,0,0,0,0,62,0,202,0,0,0,252,0,172,0,196,0,223,0,0,0,220,0,1,0,147,0,137,0,145,0,0,0,0,0,0,0,51,0,85,0,21,0,196,0,236,0,0,0,0,0,102,0,0,0,0,0,12,0,141,0,135,0,207,0,204,0,104,0,8,0,6,0,62,0,142,0,67,0,0,0,70,0,0,0,84,0,4,0,0,0,2,0,117,0,0,0,0,0,137,0,51,0,17,0,56,0,214,0,0,0,140,0,136,0,209,0,227,0,0,0,203,0,250,0,241,0,209,0,152,0,11,0,98,0,0,0,0,0,221,0,35,0,42,0,0,0,42,0,199,0,196,0,24,0,57,0,0,0,181,0,191,0,129,0,237,0,22,0,238,0,217,0,180,0,38,0,63,0,193,0,0,0,165,0,241,0,225,0,163,0,75,0,190,0,34,0,209,0,24,0,44,0,188,0,0,0,52,0,29,0,198,0,0,0,144,0,73,0,249,0,0,0,0,0,73,0,225,0,145,0,0,0,195,0,0,0,119,0);
signal scenario_full  : scenario_type := (80,31,117,31,96,31,17,31,214,31,251,31,148,31,150,31,123,31,123,30,40,31,93,31,65,31,253,31,217,31,22,31,210,31,166,31,166,30,72,31,72,30,53,31,178,31,20,31,243,31,112,31,15,31,194,31,69,31,217,31,217,30,216,31,216,30,216,29,219,31,196,31,155,31,195,31,90,31,90,30,94,31,38,31,120,31,37,31,66,31,230,31,156,31,156,30,104,31,104,30,139,31,190,31,190,30,205,31,14,31,238,31,238,30,147,31,9,31,9,30,11,31,192,31,192,30,194,31,170,31,170,30,170,29,60,31,68,31,227,31,227,30,61,31,133,31,133,30,133,29,133,28,254,31,148,31,55,31,97,31,33,31,17,31,110,31,250,31,216,31,117,31,143,31,143,30,147,31,42,31,202,31,202,30,146,31,102,31,162,31,19,31,19,30,74,31,48,31,43,31,81,31,107,31,107,30,107,29,150,31,150,30,150,29,29,31,211,31,209,31,70,31,37,31,60,31,243,31,243,30,66,31,74,31,30,31,80,31,247,31,251,31,178,31,96,31,210,31,106,31,181,31,200,31,191,31,93,31,18,31,191,31,191,30,41,31,73,31,73,30,255,31,59,31,175,31,235,31,98,31,98,30,230,31,251,31,251,30,197,31,51,31,51,30,95,31,95,30,229,31,254,31,254,30,196,31,196,30,255,31,48,31,58,31,201,31,69,31,49,31,151,31,118,31,118,30,149,31,206,31,206,30,206,29,23,31,23,30,23,29,69,31,69,30,114,31,118,31,118,30,118,29,105,31,105,30,183,31,77,31,13,31,53,31,198,31,148,31,148,30,25,31,13,31,220,31,115,31,19,31,61,31,61,30,61,29,229,31,118,31,21,31,219,31,161,31,37,31,38,31,109,31,58,31,58,30,30,31,215,31,192,31,192,30,183,31,187,31,187,30,159,31,204,31,220,31,220,30,48,31,242,31,18,31,234,31,107,31,184,31,232,31,101,31,101,30,27,31,75,31,154,31,77,31,34,31,34,30,77,31,141,31,250,31,239,31,124,31,124,30,124,29,115,31,70,31,81,31,139,31,130,31,34,31,129,31,213,31,46,31,200,31,110,31,32,31,84,31,84,30,206,31,163,31,27,31,149,31,149,30,223,31,28,31,165,31,171,31,171,30,83,31,182,31,143,31,196,31,31,31,226,31,146,31,146,30,146,29,146,28,160,31,208,31,174,31,121,31,155,31,155,30,93,31,140,31,74,31,73,31,175,31,21,31,21,30,21,29,185,31,148,31,151,31,180,31,35,31,35,30,109,31,41,31,16,31,136,31,117,31,210,31,132,31,132,30,9,31,27,31,245,31,155,31,194,31,194,30,48,31,180,31,126,31,13,31,221,31,221,30,34,31,167,31,167,30,77,31,138,31,138,30,211,31,117,31,156,31,58,31,83,31,183,31,198,31,63,31,63,30,98,31,89,31,89,30,89,29,254,31,85,31,224,31,68,31,209,31,45,31,69,31,238,31,102,31,124,31,7,31,7,31,7,30,113,31,113,30,31,31,214,31,5,31,32,31,162,31,196,31,65,31,28,31,209,31,189,31,189,30,189,29,71,31,99,31,97,31,123,31,246,31,72,31,72,30,244,31,164,31,164,30,122,31,48,31,118,31,211,31,238,31,40,31,175,31,8,31,8,30,8,29,89,31,75,31,75,30,114,31,237,31,237,30,132,31,123,31,30,31,195,31,178,31,178,30,213,31,213,30,165,31,165,30,173,31,235,31,169,31,205,31,127,31,76,31,24,31,52,31,220,31,112,31,112,30,48,31,31,31,242,31,224,31,224,30,226,31,22,31,232,31,142,31,128,31,117,31,196,31,196,30,196,29,142,31,142,31,111,31,111,30,231,31,158,31,253,31,77,31,154,31,243,31,243,30,243,29,53,31,126,31,101,31,97,31,121,31,127,31,60,31,243,31,23,31,14,31,14,30,141,31,141,30,80,31,160,31,165,31,204,31,204,30,188,31,198,31,228,31,161,31,62,31,111,31,139,31,139,30,139,29,175,31,175,30,145,31,62,31,6,31,153,31,42,31,65,31,159,31,159,30,159,29,8,31,128,31,85,31,156,31,209,31,236,31,122,31,249,31,158,31,99,31,172,31,172,30,57,31,57,30,95,31,95,30,95,29,95,28,102,31,225,31,115,31,234,31,133,31,49,31,86,31,134,31,152,31,170,31,149,31,249,31,23,31,47,31,47,30,17,31,194,31,238,31,238,30,197,31,124,31,239,31,23,31,95,31,95,30,162,31,170,31,163,31,35,31,35,30,174,31,174,30,32,31,97,31,160,31,160,30,127,31,251,31,190,31,55,31,83,31,100,31,36,31,160,31,135,31,135,30,135,29,63,31,106,31,117,31,6,31,216,31,45,31,35,31,33,31,146,31,137,31,92,31,92,30,56,31,10,31,166,31,74,31,178,31,178,30,185,31,185,30,38,31,38,30,203,31,2,31,187,31,187,30,187,29,117,31,213,31,19,31,21,31,175,31,51,31,128,31,167,31,167,30,93,31,22,31,22,30,152,31,152,30,12,31,154,31,95,31,96,31,157,31,57,31,243,31,223,31,12,31,12,30,143,31,99,31,99,30,99,29,150,31,235,31,139,31,56,31,170,31,108,31,185,31,185,30,248,31,248,30,151,31,45,31,26,31,238,31,142,31,159,31,185,31,233,31,233,30,169,31,169,30,193,31,186,31,186,30,148,31,112,31,165,31,112,31,67,31,38,31,99,31,94,31,94,30,94,29,55,31,68,31,184,31,136,31,157,31,157,30,152,31,178,31,7,31,240,31,240,30,83,31,122,31,99,31,156,31,164,31,59,31,108,31,151,31,7,31,141,31,4,31,248,31,56,31,93,31,93,30,189,31,13,31,13,30,216,31,98,31,81,31,81,30,81,29,149,31,231,31,170,31,240,31,44,31,226,31,11,31,133,31,151,31,91,31,9,31,75,31,251,31,75,31,235,31,235,30,235,29,235,28,162,31,162,30,195,31,195,30,195,29,195,28,195,27,62,31,202,31,202,30,252,31,172,31,196,31,223,31,223,30,220,31,1,31,147,31,137,31,145,31,145,30,145,29,145,28,51,31,85,31,21,31,196,31,236,31,236,30,236,29,102,31,102,30,102,29,12,31,141,31,135,31,207,31,204,31,104,31,8,31,6,31,62,31,142,31,67,31,67,30,70,31,70,30,84,31,4,31,4,30,2,31,117,31,117,30,117,29,137,31,51,31,17,31,56,31,214,31,214,30,140,31,136,31,209,31,227,31,227,30,203,31,250,31,241,31,209,31,152,31,11,31,98,31,98,30,98,29,221,31,35,31,42,31,42,30,42,31,199,31,196,31,24,31,57,31,57,30,181,31,191,31,129,31,237,31,22,31,238,31,217,31,180,31,38,31,63,31,193,31,193,30,165,31,241,31,225,31,163,31,75,31,190,31,34,31,209,31,24,31,44,31,188,31,188,30,52,31,29,31,198,31,198,30,144,31,73,31,249,31,249,30,249,29,73,31,225,31,145,31,145,30,195,31,195,30,119,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
