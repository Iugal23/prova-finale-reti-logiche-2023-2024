-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_959 is
end project_tb_959;

architecture project_tb_arch_959 of project_tb_959 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 695;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,197,0,0,0,122,0,143,0,188,0,0,0,27,0,131,0,113,0,245,0,66,0,79,0,110,0,98,0,79,0,0,0,0,0,95,0,74,0,0,0,0,0,69,0,32,0,46,0,163,0,143,0,55,0,39,0,86,0,249,0,137,0,255,0,67,0,91,0,161,0,33,0,0,0,126,0,121,0,234,0,2,0,0,0,215,0,0,0,34,0,0,0,154,0,203,0,0,0,61,0,113,0,158,0,242,0,155,0,0,0,107,0,85,0,235,0,249,0,0,0,124,0,122,0,160,0,54,0,46,0,219,0,2,0,135,0,228,0,72,0,169,0,204,0,70,0,184,0,233,0,174,0,193,0,10,0,66,0,0,0,0,0,3,0,82,0,151,0,0,0,125,0,239,0,117,0,0,0,0,0,0,0,0,0,214,0,239,0,63,0,0,0,13,0,169,0,160,0,0,0,78,0,0,0,252,0,135,0,141,0,0,0,246,0,237,0,194,0,182,0,255,0,0,0,0,0,123,0,98,0,99,0,76,0,0,0,147,0,70,0,0,0,132,0,224,0,23,0,41,0,0,0,95,0,126,0,50,0,0,0,201,0,176,0,0,0,41,0,136,0,83,0,110,0,226,0,223,0,26,0,1,0,22,0,18,0,6,0,19,0,106,0,0,0,0,0,33,0,40,0,140,0,254,0,163,0,43,0,0,0,224,0,187,0,159,0,190,0,115,0,27,0,72,0,177,0,113,0,160,0,111,0,194,0,87,0,0,0,18,0,205,0,128,0,38,0,172,0,110,0,30,0,138,0,110,0,37,0,128,0,73,0,157,0,98,0,143,0,0,0,202,0,184,0,168,0,0,0,0,0,215,0,127,0,0,0,12,0,20,0,26,0,122,0,75,0,240,0,0,0,10,0,157,0,198,0,0,0,134,0,11,0,163,0,55,0,121,0,7,0,129,0,83,0,83,0,61,0,175,0,192,0,46,0,0,0,160,0,0,0,0,0,113,0,194,0,252,0,9,0,229,0,177,0,31,0,195,0,173,0,140,0,82,0,68,0,160,0,0,0,0,0,127,0,195,0,51,0,0,0,158,0,68,0,202,0,65,0,104,0,0,0,169,0,212,0,19,0,17,0,91,0,0,0,107,0,116,0,117,0,205,0,46,0,24,0,0,0,211,0,41,0,9,0,214,0,0,0,245,0,158,0,0,0,56,0,92,0,50,0,0,0,227,0,0,0,167,0,216,0,105,0,0,0,200,0,100,0,106,0,85,0,216,0,79,0,111,0,108,0,0,0,109,0,194,0,213,0,22,0,228,0,84,0,0,0,27,0,0,0,83,0,41,0,226,0,148,0,75,0,159,0,243,0,218,0,137,0,68,0,0,0,204,0,0,0,70,0,164,0,251,0,191,0,114,0,164,0,220,0,174,0,208,0,73,0,114,0,0,0,0,0,9,0,34,0,0,0,165,0,59,0,220,0,96,0,110,0,228,0,0,0,94,0,200,0,206,0,112,0,202,0,192,0,0,0,163,0,131,0,198,0,11,0,55,0,202,0,234,0,56,0,0,0,236,0,173,0,67,0,58,0,103,0,128,0,0,0,0,0,243,0,0,0,206,0,217,0,82,0,5,0,109,0,0,0,0,0,64,0,235,0,205,0,79,0,45,0,0,0,0,0,214,0,0,0,0,0,78,0,39,0,68,0,161,0,0,0,42,0,138,0,202,0,0,0,0,0,185,0,204,0,126,0,232,0,88,0,0,0,42,0,65,0,102,0,165,0,43,0,158,0,72,0,0,0,137,0,0,0,4,0,150,0,46,0,141,0,238,0,226,0,133,0,0,0,91,0,248,0,55,0,36,0,118,0,25,0,62,0,252,0,201,0,174,0,169,0,78,0,62,0,0,0,0,0,103,0,210,0,169,0,54,0,13,0,133,0,203,0,74,0,206,0,0,0,146,0,0,0,49,0,144,0,137,0,122,0,0,0,0,0,26,0,160,0,162,0,146,0,246,0,53,0,0,0,32,0,0,0,0,0,181,0,176,0,156,0,46,0,0,0,170,0,70,0,211,0,68,0,62,0,0,0,27,0,0,0,45,0,1,0,130,0,0,0,249,0,99,0,184,0,225,0,0,0,0,0,16,0,156,0,106,0,0,0,0,0,245,0,192,0,135,0,157,0,0,0,50,0,121,0,176,0,141,0,170,0,88,0,4,0,0,0,240,0,4,0,44,0,111,0,209,0,0,0,101,0,44,0,11,0,210,0,143,0,0,0,76,0,252,0,238,0,253,0,49,0,54,0,51,0,210,0,26,0,122,0,99,0,111,0,203,0,0,0,228,0,13,0,6,0,122,0,240,0,0,0,163,0,123,0,105,0,127,0,0,0,14,0,19,0,55,0,212,0,193,0,0,0,176,0,199,0,174,0,144,0,0,0,183,0,72,0,4,0,85,0,0,0,138,0,139,0,162,0,81,0,229,0,113,0,9,0,234,0,94,0,0,0,13,0,143,0,6,0,142,0,27,0,56,0,0,0,236,0,190,0,0,0,107,0,250,0,0,0,26,0,199,0,0,0,119,0,123,0,0,0,106,0,0,0,104,0,109,0,208,0,52,0,191,0,0,0,238,0,243,0,224,0,203,0,50,0,190,0,178,0,80,0,0,0,75,0,64,0,168,0,176,0,112,0,29,0,1,0,0,0,207,0,128,0,35,0,18,0,218,0,126,0,75,0,233,0,80,0,51,0,235,0,188,0,166,0,27,0,198,0,78,0,191,0,0,0,87,0,174,0,170,0,86,0,245,0,208,0,246,0,108,0,134,0,58,0,0,0,214,0,246,0,202,0,200,0,0,0,0,0,52,0,236,0,0,0,176,0,158,0,59,0,62,0,233,0,0,0,71,0,0,0,82,0,28,0,0,0,225,0,0,0,0,0,120,0,0,0,159,0,199,0,221,0,254,0,0,0,209,0,136,0,255,0,34,0,181,0,0,0,75,0,61,0,237,0,89,0,240,0,158,0,0,0,57,0,44,0,0,0,56,0,195,0,75,0,34,0,105,0,0,0,46,0,0,0,119,0,0,0,131,0,22,0,225,0,62,0,0,0,0,0,190,0,183,0,244,0,132,0);
signal scenario_full  : scenario_type := (0,0,197,31,197,30,122,31,143,31,188,31,188,30,27,31,131,31,113,31,245,31,66,31,79,31,110,31,98,31,79,31,79,30,79,29,95,31,74,31,74,30,74,29,69,31,32,31,46,31,163,31,143,31,55,31,39,31,86,31,249,31,137,31,255,31,67,31,91,31,161,31,33,31,33,30,126,31,121,31,234,31,2,31,2,30,215,31,215,30,34,31,34,30,154,31,203,31,203,30,61,31,113,31,158,31,242,31,155,31,155,30,107,31,85,31,235,31,249,31,249,30,124,31,122,31,160,31,54,31,46,31,219,31,2,31,135,31,228,31,72,31,169,31,204,31,70,31,184,31,233,31,174,31,193,31,10,31,66,31,66,30,66,29,3,31,82,31,151,31,151,30,125,31,239,31,117,31,117,30,117,29,117,28,117,27,214,31,239,31,63,31,63,30,13,31,169,31,160,31,160,30,78,31,78,30,252,31,135,31,141,31,141,30,246,31,237,31,194,31,182,31,255,31,255,30,255,29,123,31,98,31,99,31,76,31,76,30,147,31,70,31,70,30,132,31,224,31,23,31,41,31,41,30,95,31,126,31,50,31,50,30,201,31,176,31,176,30,41,31,136,31,83,31,110,31,226,31,223,31,26,31,1,31,22,31,18,31,6,31,19,31,106,31,106,30,106,29,33,31,40,31,140,31,254,31,163,31,43,31,43,30,224,31,187,31,159,31,190,31,115,31,27,31,72,31,177,31,113,31,160,31,111,31,194,31,87,31,87,30,18,31,205,31,128,31,38,31,172,31,110,31,30,31,138,31,110,31,37,31,128,31,73,31,157,31,98,31,143,31,143,30,202,31,184,31,168,31,168,30,168,29,215,31,127,31,127,30,12,31,20,31,26,31,122,31,75,31,240,31,240,30,10,31,157,31,198,31,198,30,134,31,11,31,163,31,55,31,121,31,7,31,129,31,83,31,83,31,61,31,175,31,192,31,46,31,46,30,160,31,160,30,160,29,113,31,194,31,252,31,9,31,229,31,177,31,31,31,195,31,173,31,140,31,82,31,68,31,160,31,160,30,160,29,127,31,195,31,51,31,51,30,158,31,68,31,202,31,65,31,104,31,104,30,169,31,212,31,19,31,17,31,91,31,91,30,107,31,116,31,117,31,205,31,46,31,24,31,24,30,211,31,41,31,9,31,214,31,214,30,245,31,158,31,158,30,56,31,92,31,50,31,50,30,227,31,227,30,167,31,216,31,105,31,105,30,200,31,100,31,106,31,85,31,216,31,79,31,111,31,108,31,108,30,109,31,194,31,213,31,22,31,228,31,84,31,84,30,27,31,27,30,83,31,41,31,226,31,148,31,75,31,159,31,243,31,218,31,137,31,68,31,68,30,204,31,204,30,70,31,164,31,251,31,191,31,114,31,164,31,220,31,174,31,208,31,73,31,114,31,114,30,114,29,9,31,34,31,34,30,165,31,59,31,220,31,96,31,110,31,228,31,228,30,94,31,200,31,206,31,112,31,202,31,192,31,192,30,163,31,131,31,198,31,11,31,55,31,202,31,234,31,56,31,56,30,236,31,173,31,67,31,58,31,103,31,128,31,128,30,128,29,243,31,243,30,206,31,217,31,82,31,5,31,109,31,109,30,109,29,64,31,235,31,205,31,79,31,45,31,45,30,45,29,214,31,214,30,214,29,78,31,39,31,68,31,161,31,161,30,42,31,138,31,202,31,202,30,202,29,185,31,204,31,126,31,232,31,88,31,88,30,42,31,65,31,102,31,165,31,43,31,158,31,72,31,72,30,137,31,137,30,4,31,150,31,46,31,141,31,238,31,226,31,133,31,133,30,91,31,248,31,55,31,36,31,118,31,25,31,62,31,252,31,201,31,174,31,169,31,78,31,62,31,62,30,62,29,103,31,210,31,169,31,54,31,13,31,133,31,203,31,74,31,206,31,206,30,146,31,146,30,49,31,144,31,137,31,122,31,122,30,122,29,26,31,160,31,162,31,146,31,246,31,53,31,53,30,32,31,32,30,32,29,181,31,176,31,156,31,46,31,46,30,170,31,70,31,211,31,68,31,62,31,62,30,27,31,27,30,45,31,1,31,130,31,130,30,249,31,99,31,184,31,225,31,225,30,225,29,16,31,156,31,106,31,106,30,106,29,245,31,192,31,135,31,157,31,157,30,50,31,121,31,176,31,141,31,170,31,88,31,4,31,4,30,240,31,4,31,44,31,111,31,209,31,209,30,101,31,44,31,11,31,210,31,143,31,143,30,76,31,252,31,238,31,253,31,49,31,54,31,51,31,210,31,26,31,122,31,99,31,111,31,203,31,203,30,228,31,13,31,6,31,122,31,240,31,240,30,163,31,123,31,105,31,127,31,127,30,14,31,19,31,55,31,212,31,193,31,193,30,176,31,199,31,174,31,144,31,144,30,183,31,72,31,4,31,85,31,85,30,138,31,139,31,162,31,81,31,229,31,113,31,9,31,234,31,94,31,94,30,13,31,143,31,6,31,142,31,27,31,56,31,56,30,236,31,190,31,190,30,107,31,250,31,250,30,26,31,199,31,199,30,119,31,123,31,123,30,106,31,106,30,104,31,109,31,208,31,52,31,191,31,191,30,238,31,243,31,224,31,203,31,50,31,190,31,178,31,80,31,80,30,75,31,64,31,168,31,176,31,112,31,29,31,1,31,1,30,207,31,128,31,35,31,18,31,218,31,126,31,75,31,233,31,80,31,51,31,235,31,188,31,166,31,27,31,198,31,78,31,191,31,191,30,87,31,174,31,170,31,86,31,245,31,208,31,246,31,108,31,134,31,58,31,58,30,214,31,246,31,202,31,200,31,200,30,200,29,52,31,236,31,236,30,176,31,158,31,59,31,62,31,233,31,233,30,71,31,71,30,82,31,28,31,28,30,225,31,225,30,225,29,120,31,120,30,159,31,199,31,221,31,254,31,254,30,209,31,136,31,255,31,34,31,181,31,181,30,75,31,61,31,237,31,89,31,240,31,158,31,158,30,57,31,44,31,44,30,56,31,195,31,75,31,34,31,105,31,105,30,46,31,46,30,119,31,119,30,131,31,22,31,225,31,62,31,62,30,62,29,190,31,183,31,244,31,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
