-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 837;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,0,0,37,0,232,0,144,0,73,0,0,0,0,0,199,0,101,0,161,0,243,0,0,0,167,0,20,0,184,0,0,0,221,0,96,0,74,0,154,0,86,0,0,0,0,0,79,0,91,0,237,0,200,0,0,0,30,0,0,0,163,0,80,0,149,0,255,0,3,0,11,0,105,0,148,0,3,0,52,0,146,0,67,0,0,0,220,0,149,0,13,0,175,0,194,0,108,0,106,0,98,0,7,0,28,0,159,0,125,0,230,0,200,0,74,0,204,0,110,0,60,0,165,0,193,0,72,0,199,0,175,0,123,0,0,0,236,0,248,0,58,0,123,0,0,0,38,0,192,0,217,0,0,0,156,0,133,0,239,0,227,0,153,0,75,0,0,0,0,0,0,0,183,0,0,0,201,0,0,0,28,0,0,0,41,0,70,0,70,0,192,0,47,0,108,0,132,0,119,0,92,0,0,0,75,0,97,0,16,0,108,0,0,0,60,0,95,0,42,0,215,0,188,0,79,0,0,0,216,0,239,0,0,0,0,0,107,0,159,0,219,0,0,0,172,0,16,0,219,0,206,0,29,0,125,0,157,0,0,0,116,0,0,0,112,0,47,0,228,0,170,0,0,0,0,0,105,0,0,0,0,0,28,0,54,0,174,0,177,0,0,0,221,0,0,0,168,0,248,0,0,0,35,0,216,0,142,0,125,0,144,0,0,0,131,0,0,0,194,0,96,0,50,0,0,0,193,0,0,0,68,0,0,0,13,0,0,0,142,0,255,0,36,0,190,0,248,0,2,0,38,0,0,0,216,0,98,0,229,0,0,0,60,0,90,0,225,0,31,0,163,0,247,0,140,0,241,0,0,0,0,0,215,0,168,0,205,0,0,0,0,0,134,0,109,0,0,0,0,0,0,0,228,0,0,0,107,0,152,0,23,0,92,0,145,0,168,0,88,0,57,0,79,0,114,0,16,0,0,0,0,0,160,0,221,0,150,0,119,0,0,0,159,0,67,0,205,0,255,0,0,0,80,0,188,0,52,0,174,0,187,0,95,0,200,0,102,0,145,0,71,0,56,0,45,0,209,0,133,0,81,0,242,0,0,0,152,0,247,0,116,0,56,0,82,0,27,0,0,0,51,0,66,0,14,0,55,0,215,0,128,0,175,0,197,0,6,0,5,0,176,0,41,0,36,0,250,0,43,0,46,0,249,0,80,0,88,0,0,0,92,0,120,0,0,0,173,0,0,0,56,0,246,0,251,0,6,0,82,0,113,0,150,0,94,0,193,0,62,0,0,0,141,0,183,0,27,0,162,0,22,0,0,0,150,0,192,0,159,0,36,0,235,0,0,0,13,0,26,0,57,0,1,0,65,0,0,0,213,0,192,0,74,0,214,0,0,0,236,0,52,0,226,0,71,0,145,0,0,0,164,0,221,0,236,0,74,0,143,0,0,0,216,0,245,0,53,0,182,0,0,0,78,0,11,0,0,0,107,0,75,0,41,0,0,0,67,0,58,0,234,0,66,0,0,0,0,0,193,0,0,0,238,0,163,0,196,0,166,0,206,0,102,0,130,0,190,0,202,0,0,0,0,0,0,0,149,0,83,0,3,0,0,0,65,0,178,0,82,0,214,0,148,0,0,0,0,0,0,0,0,0,46,0,216,0,0,0,13,0,247,0,0,0,135,0,155,0,66,0,192,0,234,0,63,0,1,0,122,0,195,0,2,0,7,0,197,0,0,0,115,0,23,0,36,0,0,0,26,0,106,0,53,0,111,0,21,0,96,0,18,0,55,0,103,0,222,0,61,0,0,0,206,0,7,0,191,0,51,0,191,0,0,0,136,0,158,0,173,0,32,0,0,0,174,0,0,0,26,0,54,0,7,0,232,0,116,0,141,0,229,0,1,0,0,0,63,0,19,0,0,0,148,0,0,0,173,0,236,0,104,0,0,0,51,0,139,0,0,0,119,0,0,0,0,0,240,0,73,0,67,0,0,0,133,0,132,0,143,0,151,0,209,0,186,0,118,0,0,0,182,0,23,0,50,0,236,0,45,0,164,0,237,0,37,0,149,0,13,0,0,0,46,0,139,0,34,0,201,0,46,0,0,0,67,0,170,0,42,0,89,0,113,0,0,0,74,0,0,0,0,0,106,0,247,0,0,0,18,0,227,0,200,0,241,0,119,0,139,0,0,0,0,0,92,0,0,0,223,0,56,0,0,0,0,0,195,0,0,0,28,0,169,0,153,0,143,0,0,0,190,0,32,0,115,0,78,0,121,0,0,0,192,0,0,0,0,0,144,0,79,0,102,0,113,0,0,0,100,0,56,0,113,0,101,0,52,0,252,0,201,0,205,0,208,0,52,0,20,0,233,0,109,0,0,0,41,0,237,0,83,0,90,0,129,0,53,0,247,0,6,0,199,0,103,0,111,0,18,0,83,0,87,0,217,0,21,0,102,0,0,0,125,0,135,0,242,0,136,0,105,0,84,0,168,0,242,0,237,0,1,0,0,0,128,0,105,0,0,0,169,0,0,0,51,0,98,0,0,0,0,0,208,0,8,0,131,0,136,0,217,0,106,0,213,0,242,0,94,0,114,0,85,0,79,0,0,0,0,0,208,0,26,0,102,0,0,0,224,0,71,0,206,0,0,0,0,0,179,0,186,0,173,0,20,0,0,0,232,0,0,0,231,0,47,0,125,0,54,0,119,0,255,0,0,0,241,0,139,0,123,0,99,0,73,0,120,0,0,0,246,0,115,0,18,0,120,0,208,0,212,0,92,0,233,0,89,0,107,0,183,0,0,0,16,0,218,0,56,0,62,0,78,0,45,0,135,0,110,0,245,0,226,0,0,0,222,0,179,0,171,0,221,0,163,0,0,0,54,0,97,0,84,0,0,0,0,0,213,0,0,0,0,0,238,0,53,0,146,0,0,0,117,0,167,0,8,0,0,0,4,0,160,0,77,0,45,0,141,0,73,0,0,0,164,0,0,0,143,0,0,0,118,0,132,0,179,0,42,0,89,0,0,0,225,0,67,0,181,0,0,0,249,0,81,0,57,0,180,0,215,0,0,0,207,0,132,0,202,0,239,0,170,0,123,0,124,0,29,0,3,0,191,0,243,0,85,0,171,0,12,0,159,0,0,0,3,0,0,0,103,0,0,0,220,0,236,0,247,0,191,0,0,0,184,0,174,0,234,0,135,0,0,0,192,0,243,0,0,0,122,0,95,0,123,0,127,0,217,0,39,0,120,0,111,0,120,0,8,0,0,0,167,0,33,0,166,0,75,0,26,0,0,0,0,0,206,0,218,0,24,0,111,0,240,0,102,0,0,0,10,0,122,0,4,0,75,0,164,0,49,0,19,0,0,0,69,0,218,0,61,0,0,0,80,0,23,0,0,0,230,0,73,0,121,0,39,0,0,0,83,0,0,0,1,0,156,0,101,0,66,0,151,0,113,0,0,0,4,0,0,0,66,0,238,0,33,0,204,0,247,0,232,0,77,0,69,0,95,0,46,0,103,0,200,0,64,0,216,0,15,0,162,0,0,0,253,0,0,0,58,0,153,0,176,0,5,0,0,0,5,0,118,0,88,0,9,0,5,0,148,0,184,0,189,0,101,0,216,0,20,0,45,0,179,0,0,0,16,0,226,0,44,0,0,0,151,0,48,0,240,0,0,0,5,0,0,0,4,0,232,0,162,0,159,0,0,0,7,0,222,0,71,0,0,0,43,0,32,0,72,0,112,0,98,0,255,0,159,0,58,0);
signal scenario_full  : scenario_type := (139,31,139,30,37,31,232,31,144,31,73,31,73,30,73,29,199,31,101,31,161,31,243,31,243,30,167,31,20,31,184,31,184,30,221,31,96,31,74,31,154,31,86,31,86,30,86,29,79,31,91,31,237,31,200,31,200,30,30,31,30,30,163,31,80,31,149,31,255,31,3,31,11,31,105,31,148,31,3,31,52,31,146,31,67,31,67,30,220,31,149,31,13,31,175,31,194,31,108,31,106,31,98,31,7,31,28,31,159,31,125,31,230,31,200,31,74,31,204,31,110,31,60,31,165,31,193,31,72,31,199,31,175,31,123,31,123,30,236,31,248,31,58,31,123,31,123,30,38,31,192,31,217,31,217,30,156,31,133,31,239,31,227,31,153,31,75,31,75,30,75,29,75,28,183,31,183,30,201,31,201,30,28,31,28,30,41,31,70,31,70,31,192,31,47,31,108,31,132,31,119,31,92,31,92,30,75,31,97,31,16,31,108,31,108,30,60,31,95,31,42,31,215,31,188,31,79,31,79,30,216,31,239,31,239,30,239,29,107,31,159,31,219,31,219,30,172,31,16,31,219,31,206,31,29,31,125,31,157,31,157,30,116,31,116,30,112,31,47,31,228,31,170,31,170,30,170,29,105,31,105,30,105,29,28,31,54,31,174,31,177,31,177,30,221,31,221,30,168,31,248,31,248,30,35,31,216,31,142,31,125,31,144,31,144,30,131,31,131,30,194,31,96,31,50,31,50,30,193,31,193,30,68,31,68,30,13,31,13,30,142,31,255,31,36,31,190,31,248,31,2,31,38,31,38,30,216,31,98,31,229,31,229,30,60,31,90,31,225,31,31,31,163,31,247,31,140,31,241,31,241,30,241,29,215,31,168,31,205,31,205,30,205,29,134,31,109,31,109,30,109,29,109,28,228,31,228,30,107,31,152,31,23,31,92,31,145,31,168,31,88,31,57,31,79,31,114,31,16,31,16,30,16,29,160,31,221,31,150,31,119,31,119,30,159,31,67,31,205,31,255,31,255,30,80,31,188,31,52,31,174,31,187,31,95,31,200,31,102,31,145,31,71,31,56,31,45,31,209,31,133,31,81,31,242,31,242,30,152,31,247,31,116,31,56,31,82,31,27,31,27,30,51,31,66,31,14,31,55,31,215,31,128,31,175,31,197,31,6,31,5,31,176,31,41,31,36,31,250,31,43,31,46,31,249,31,80,31,88,31,88,30,92,31,120,31,120,30,173,31,173,30,56,31,246,31,251,31,6,31,82,31,113,31,150,31,94,31,193,31,62,31,62,30,141,31,183,31,27,31,162,31,22,31,22,30,150,31,192,31,159,31,36,31,235,31,235,30,13,31,26,31,57,31,1,31,65,31,65,30,213,31,192,31,74,31,214,31,214,30,236,31,52,31,226,31,71,31,145,31,145,30,164,31,221,31,236,31,74,31,143,31,143,30,216,31,245,31,53,31,182,31,182,30,78,31,11,31,11,30,107,31,75,31,41,31,41,30,67,31,58,31,234,31,66,31,66,30,66,29,193,31,193,30,238,31,163,31,196,31,166,31,206,31,102,31,130,31,190,31,202,31,202,30,202,29,202,28,149,31,83,31,3,31,3,30,65,31,178,31,82,31,214,31,148,31,148,30,148,29,148,28,148,27,46,31,216,31,216,30,13,31,247,31,247,30,135,31,155,31,66,31,192,31,234,31,63,31,1,31,122,31,195,31,2,31,7,31,197,31,197,30,115,31,23,31,36,31,36,30,26,31,106,31,53,31,111,31,21,31,96,31,18,31,55,31,103,31,222,31,61,31,61,30,206,31,7,31,191,31,51,31,191,31,191,30,136,31,158,31,173,31,32,31,32,30,174,31,174,30,26,31,54,31,7,31,232,31,116,31,141,31,229,31,1,31,1,30,63,31,19,31,19,30,148,31,148,30,173,31,236,31,104,31,104,30,51,31,139,31,139,30,119,31,119,30,119,29,240,31,73,31,67,31,67,30,133,31,132,31,143,31,151,31,209,31,186,31,118,31,118,30,182,31,23,31,50,31,236,31,45,31,164,31,237,31,37,31,149,31,13,31,13,30,46,31,139,31,34,31,201,31,46,31,46,30,67,31,170,31,42,31,89,31,113,31,113,30,74,31,74,30,74,29,106,31,247,31,247,30,18,31,227,31,200,31,241,31,119,31,139,31,139,30,139,29,92,31,92,30,223,31,56,31,56,30,56,29,195,31,195,30,28,31,169,31,153,31,143,31,143,30,190,31,32,31,115,31,78,31,121,31,121,30,192,31,192,30,192,29,144,31,79,31,102,31,113,31,113,30,100,31,56,31,113,31,101,31,52,31,252,31,201,31,205,31,208,31,52,31,20,31,233,31,109,31,109,30,41,31,237,31,83,31,90,31,129,31,53,31,247,31,6,31,199,31,103,31,111,31,18,31,83,31,87,31,217,31,21,31,102,31,102,30,125,31,135,31,242,31,136,31,105,31,84,31,168,31,242,31,237,31,1,31,1,30,128,31,105,31,105,30,169,31,169,30,51,31,98,31,98,30,98,29,208,31,8,31,131,31,136,31,217,31,106,31,213,31,242,31,94,31,114,31,85,31,79,31,79,30,79,29,208,31,26,31,102,31,102,30,224,31,71,31,206,31,206,30,206,29,179,31,186,31,173,31,20,31,20,30,232,31,232,30,231,31,47,31,125,31,54,31,119,31,255,31,255,30,241,31,139,31,123,31,99,31,73,31,120,31,120,30,246,31,115,31,18,31,120,31,208,31,212,31,92,31,233,31,89,31,107,31,183,31,183,30,16,31,218,31,56,31,62,31,78,31,45,31,135,31,110,31,245,31,226,31,226,30,222,31,179,31,171,31,221,31,163,31,163,30,54,31,97,31,84,31,84,30,84,29,213,31,213,30,213,29,238,31,53,31,146,31,146,30,117,31,167,31,8,31,8,30,4,31,160,31,77,31,45,31,141,31,73,31,73,30,164,31,164,30,143,31,143,30,118,31,132,31,179,31,42,31,89,31,89,30,225,31,67,31,181,31,181,30,249,31,81,31,57,31,180,31,215,31,215,30,207,31,132,31,202,31,239,31,170,31,123,31,124,31,29,31,3,31,191,31,243,31,85,31,171,31,12,31,159,31,159,30,3,31,3,30,103,31,103,30,220,31,236,31,247,31,191,31,191,30,184,31,174,31,234,31,135,31,135,30,192,31,243,31,243,30,122,31,95,31,123,31,127,31,217,31,39,31,120,31,111,31,120,31,8,31,8,30,167,31,33,31,166,31,75,31,26,31,26,30,26,29,206,31,218,31,24,31,111,31,240,31,102,31,102,30,10,31,122,31,4,31,75,31,164,31,49,31,19,31,19,30,69,31,218,31,61,31,61,30,80,31,23,31,23,30,230,31,73,31,121,31,39,31,39,30,83,31,83,30,1,31,156,31,101,31,66,31,151,31,113,31,113,30,4,31,4,30,66,31,238,31,33,31,204,31,247,31,232,31,77,31,69,31,95,31,46,31,103,31,200,31,64,31,216,31,15,31,162,31,162,30,253,31,253,30,58,31,153,31,176,31,5,31,5,30,5,31,118,31,88,31,9,31,5,31,148,31,184,31,189,31,101,31,216,31,20,31,45,31,179,31,179,30,16,31,226,31,44,31,44,30,151,31,48,31,240,31,240,30,5,31,5,30,4,31,232,31,162,31,159,31,159,30,7,31,222,31,71,31,71,30,43,31,32,31,72,31,112,31,98,31,255,31,159,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
