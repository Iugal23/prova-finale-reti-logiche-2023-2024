-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_72 is
end project_tb_72;

architecture project_tb_arch_72 of project_tb_72 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 469;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,0,0,0,0,152,0,254,0,82,0,105,0,38,0,178,0,188,0,0,0,209,0,115,0,0,0,139,0,92,0,98,0,157,0,141,0,0,0,80,0,0,0,245,0,229,0,114,0,12,0,140,0,201,0,23,0,0,0,81,0,65,0,0,0,112,0,73,0,0,0,186,0,170,0,52,0,146,0,0,0,106,0,0,0,140,0,162,0,0,0,160,0,128,0,117,0,172,0,69,0,233,0,151,0,81,0,0,0,119,0,34,0,110,0,70,0,232,0,0,0,22,0,33,0,117,0,0,0,95,0,234,0,78,0,97,0,89,0,135,0,89,0,112,0,35,0,188,0,130,0,158,0,228,0,198,0,0,0,0,0,166,0,27,0,43,0,60,0,0,0,0,0,229,0,0,0,0,0,128,0,154,0,132,0,97,0,98,0,151,0,121,0,118,0,172,0,122,0,156,0,119,0,98,0,0,0,112,0,24,0,96,0,30,0,214,0,67,0,133,0,128,0,25,0,12,0,65,0,0,0,135,0,195,0,165,0,203,0,199,0,110,0,104,0,146,0,212,0,167,0,0,0,215,0,255,0,110,0,186,0,107,0,0,0,0,0,0,0,0,0,237,0,81,0,121,0,139,0,63,0,86,0,12,0,86,0,117,0,0,0,21,0,0,0,41,0,58,0,29,0,0,0,253,0,95,0,104,0,5,0,167,0,108,0,226,0,132,0,0,0,101,0,241,0,93,0,0,0,148,0,115,0,0,0,17,0,29,0,247,0,30,0,253,0,218,0,120,0,0,0,136,0,230,0,0,0,117,0,157,0,124,0,183,0,200,0,174,0,0,0,121,0,0,0,0,0,0,0,109,0,132,0,245,0,157,0,140,0,105,0,13,0,152,0,115,0,152,0,221,0,0,0,105,0,60,0,111,0,0,0,44,0,0,0,145,0,189,0,237,0,86,0,0,0,186,0,188,0,231,0,47,0,24,0,0,0,0,0,64,0,193,0,0,0,24,0,61,0,128,0,0,0,16,0,213,0,38,0,0,0,50,0,135,0,0,0,216,0,225,0,108,0,8,0,150,0,138,0,6,0,223,0,0,0,255,0,0,0,54,0,50,0,64,0,225,0,93,0,27,0,196,0,186,0,0,0,71,0,83,0,103,0,88,0,104,0,207,0,88,0,28,0,0,0,227,0,99,0,31,0,237,0,114,0,164,0,233,0,194,0,0,0,184,0,24,0,113,0,208,0,197,0,69,0,230,0,154,0,247,0,190,0,138,0,73,0,7,0,96,0,44,0,0,0,40,0,0,0,98,0,25,0,115,0,21,0,216,0,11,0,133,0,41,0,110,0,121,0,0,0,0,0,80,0,204,0,166,0,50,0,0,0,152,0,88,0,250,0,57,0,152,0,133,0,237,0,0,0,57,0,249,0,252,0,106,0,0,0,174,0,170,0,155,0,226,0,228,0,77,0,0,0,28,0,71,0,0,0,0,0,127,0,0,0,174,0,41,0,175,0,242,0,193,0,22,0,61,0,152,0,188,0,251,0,127,0,75,0,33,0,206,0,197,0,41,0,0,0,220,0,102,0,0,0,100,0,162,0,26,0,187,0,132,0,142,0,57,0,88,0,48,0,15,0,87,0,240,0,0,0,210,0,222,0,104,0,0,0,179,0,163,0,31,0,6,0,99,0,246,0,87,0,115,0,8,0,61,0,221,0,219,0,84,0,193,0,230,0,198,0,0,0,134,0,79,0,45,0,0,0,139,0,144,0,71,0,0,0,172,0,0,0,251,0,174,0,224,0,229,0,0,0,0,0,6,0,134,0,123,0,0,0,62,0,170,0,116,0,117,0,238,0,93,0,113,0,157,0,176,0,220,0,0,0,73,0,0,0,0,0,105,0,55,0,100,0,0,0,49,0,184,0,21,0,234,0,0,0,115,0,0,0,107,0,108,0,241,0,119,0,19,0,61,0,116,0,0,0,143,0,237,0,240,0,80,0,0,0,241,0,144,0,66,0,0,0,210,0,91,0,0,0,0,0,28,0,193,0,58,0,195,0,4,0,0,0,160,0,152,0,0,0,103,0,36,0,249,0,42,0,44,0,97,0,52,0);
signal scenario_full  : scenario_type := (169,31,169,30,169,29,152,31,254,31,82,31,105,31,38,31,178,31,188,31,188,30,209,31,115,31,115,30,139,31,92,31,98,31,157,31,141,31,141,30,80,31,80,30,245,31,229,31,114,31,12,31,140,31,201,31,23,31,23,30,81,31,65,31,65,30,112,31,73,31,73,30,186,31,170,31,52,31,146,31,146,30,106,31,106,30,140,31,162,31,162,30,160,31,128,31,117,31,172,31,69,31,233,31,151,31,81,31,81,30,119,31,34,31,110,31,70,31,232,31,232,30,22,31,33,31,117,31,117,30,95,31,234,31,78,31,97,31,89,31,135,31,89,31,112,31,35,31,188,31,130,31,158,31,228,31,198,31,198,30,198,29,166,31,27,31,43,31,60,31,60,30,60,29,229,31,229,30,229,29,128,31,154,31,132,31,97,31,98,31,151,31,121,31,118,31,172,31,122,31,156,31,119,31,98,31,98,30,112,31,24,31,96,31,30,31,214,31,67,31,133,31,128,31,25,31,12,31,65,31,65,30,135,31,195,31,165,31,203,31,199,31,110,31,104,31,146,31,212,31,167,31,167,30,215,31,255,31,110,31,186,31,107,31,107,30,107,29,107,28,107,27,237,31,81,31,121,31,139,31,63,31,86,31,12,31,86,31,117,31,117,30,21,31,21,30,41,31,58,31,29,31,29,30,253,31,95,31,104,31,5,31,167,31,108,31,226,31,132,31,132,30,101,31,241,31,93,31,93,30,148,31,115,31,115,30,17,31,29,31,247,31,30,31,253,31,218,31,120,31,120,30,136,31,230,31,230,30,117,31,157,31,124,31,183,31,200,31,174,31,174,30,121,31,121,30,121,29,121,28,109,31,132,31,245,31,157,31,140,31,105,31,13,31,152,31,115,31,152,31,221,31,221,30,105,31,60,31,111,31,111,30,44,31,44,30,145,31,189,31,237,31,86,31,86,30,186,31,188,31,231,31,47,31,24,31,24,30,24,29,64,31,193,31,193,30,24,31,61,31,128,31,128,30,16,31,213,31,38,31,38,30,50,31,135,31,135,30,216,31,225,31,108,31,8,31,150,31,138,31,6,31,223,31,223,30,255,31,255,30,54,31,50,31,64,31,225,31,93,31,27,31,196,31,186,31,186,30,71,31,83,31,103,31,88,31,104,31,207,31,88,31,28,31,28,30,227,31,99,31,31,31,237,31,114,31,164,31,233,31,194,31,194,30,184,31,24,31,113,31,208,31,197,31,69,31,230,31,154,31,247,31,190,31,138,31,73,31,7,31,96,31,44,31,44,30,40,31,40,30,98,31,25,31,115,31,21,31,216,31,11,31,133,31,41,31,110,31,121,31,121,30,121,29,80,31,204,31,166,31,50,31,50,30,152,31,88,31,250,31,57,31,152,31,133,31,237,31,237,30,57,31,249,31,252,31,106,31,106,30,174,31,170,31,155,31,226,31,228,31,77,31,77,30,28,31,71,31,71,30,71,29,127,31,127,30,174,31,41,31,175,31,242,31,193,31,22,31,61,31,152,31,188,31,251,31,127,31,75,31,33,31,206,31,197,31,41,31,41,30,220,31,102,31,102,30,100,31,162,31,26,31,187,31,132,31,142,31,57,31,88,31,48,31,15,31,87,31,240,31,240,30,210,31,222,31,104,31,104,30,179,31,163,31,31,31,6,31,99,31,246,31,87,31,115,31,8,31,61,31,221,31,219,31,84,31,193,31,230,31,198,31,198,30,134,31,79,31,45,31,45,30,139,31,144,31,71,31,71,30,172,31,172,30,251,31,174,31,224,31,229,31,229,30,229,29,6,31,134,31,123,31,123,30,62,31,170,31,116,31,117,31,238,31,93,31,113,31,157,31,176,31,220,31,220,30,73,31,73,30,73,29,105,31,55,31,100,31,100,30,49,31,184,31,21,31,234,31,234,30,115,31,115,30,107,31,108,31,241,31,119,31,19,31,61,31,116,31,116,30,143,31,237,31,240,31,80,31,80,30,241,31,144,31,66,31,66,30,210,31,91,31,91,30,91,29,28,31,193,31,58,31,195,31,4,31,4,30,160,31,152,31,152,30,103,31,36,31,249,31,42,31,44,31,97,31,52,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
