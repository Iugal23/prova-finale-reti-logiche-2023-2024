-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 722;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,88,0,0,0,172,0,13,0,119,0,32,0,164,0,112,0,65,0,194,0,0,0,116,0,170,0,99,0,173,0,0,0,253,0,74,0,226,0,126,0,233,0,122,0,202,0,198,0,0,0,22,0,95,0,47,0,117,0,0,0,83,0,249,0,177,0,212,0,119,0,240,0,141,0,0,0,225,0,161,0,100,0,254,0,253,0,0,0,97,0,254,0,233,0,246,0,142,0,0,0,194,0,191,0,156,0,39,0,73,0,0,0,0,0,0,0,204,0,86,0,0,0,33,0,57,0,162,0,136,0,99,0,33,0,142,0,89,0,123,0,0,0,152,0,95,0,76,0,151,0,0,0,99,0,212,0,119,0,113,0,185,0,169,0,200,0,0,0,240,0,183,0,46,0,153,0,174,0,160,0,0,0,4,0,124,0,154,0,75,0,148,0,242,0,29,0,240,0,121,0,12,0,166,0,247,0,168,0,16,0,81,0,172,0,103,0,164,0,138,0,217,0,175,0,122,0,219,0,0,0,1,0,116,0,104,0,1,0,152,0,215,0,202,0,34,0,0,0,0,0,211,0,0,0,33,0,118,0,221,0,135,0,16,0,234,0,56,0,197,0,189,0,18,0,143,0,188,0,189,0,0,0,213,0,17,0,0,0,196,0,206,0,147,0,0,0,210,0,182,0,192,0,0,0,209,0,41,0,170,0,21,0,53,0,48,0,101,0,170,0,99,0,194,0,0,0,0,0,12,0,0,0,44,0,0,0,239,0,138,0,0,0,182,0,0,0,14,0,0,0,89,0,129,0,37,0,101,0,0,0,111,0,58,0,0,0,227,0,32,0,95,0,186,0,15,0,15,0,192,0,96,0,33,0,50,0,188,0,92,0,127,0,204,0,15,0,16,0,168,0,171,0,146,0,46,0,0,0,39,0,80,0,134,0,0,0,27,0,0,0,0,0,90,0,23,0,0,0,2,0,79,0,0,0,94,0,0,0,0,0,165,0,0,0,8,0,0,0,105,0,39,0,94,0,238,0,34,0,0,0,112,0,0,0,17,0,221,0,14,0,0,0,247,0,37,0,101,0,0,0,221,0,194,0,221,0,0,0,60,0,239,0,131,0,47,0,22,0,0,0,16,0,109,0,239,0,180,0,252,0,24,0,220,0,30,0,252,0,16,0,202,0,162,0,59,0,228,0,0,0,172,0,155,0,50,0,249,0,11,0,0,0,0,0,111,0,223,0,182,0,51,0,253,0,166,0,137,0,34,0,42,0,239,0,25,0,233,0,43,0,0,0,17,0,0,0,77,0,231,0,0,0,121,0,70,0,0,0,0,0,225,0,118,0,98,0,0,0,0,0,85,0,36,0,0,0,200,0,115,0,144,0,217,0,246,0,0,0,131,0,241,0,69,0,76,0,0,0,199,0,119,0,141,0,0,0,97,0,239,0,211,0,50,0,228,0,93,0,121,0,69,0,189,0,126,0,34,0,144,0,228,0,0,0,163,0,145,0,16,0,228,0,51,0,191,0,181,0,231,0,21,0,11,0,213,0,0,0,0,0,24,0,141,0,41,0,0,0,50,0,0,0,175,0,199,0,0,0,255,0,56,0,0,0,200,0,101,0,73,0,25,0,90,0,53,0,80,0,129,0,111,0,199,0,149,0,84,0,0,0,0,0,227,0,144,0,220,0,152,0,1,0,206,0,0,0,0,0,146,0,0,0,88,0,56,0,85,0,15,0,62,0,107,0,0,0,231,0,0,0,19,0,162,0,0,0,0,0,53,0,224,0,38,0,114,0,21,0,0,0,156,0,14,0,0,0,62,0,235,0,0,0,62,0,110,0,202,0,191,0,16,0,225,0,202,0,0,0,0,0,122,0,108,0,0,0,0,0,29,0,0,0,55,0,173,0,242,0,127,0,18,0,41,0,52,0,164,0,75,0,22,0,36,0,53,0,0,0,169,0,0,0,0,0,126,0,226,0,0,0,0,0,117,0,100,0,199,0,81,0,0,0,18,0,41,0,164,0,97,0,0,0,94,0,0,0,21,0,136,0,0,0,255,0,142,0,12,0,0,0,15,0,164,0,154,0,70,0,0,0,144,0,254,0,0,0,74,0,34,0,169,0,225,0,0,0,241,0,3,0,3,0,79,0,248,0,162,0,120,0,0,0,242,0,103,0,0,0,0,0,101,0,217,0,87,0,0,0,234,0,253,0,139,0,160,0,167,0,237,0,186,0,49,0,55,0,33,0,30,0,120,0,196,0,231,0,171,0,134,0,111,0,187,0,66,0,47,0,0,0,101,0,237,0,89,0,91,0,95,0,0,0,180,0,200,0,3,0,0,0,0,0,59,0,36,0,136,0,169,0,103,0,160,0,29,0,0,0,0,0,0,0,82,0,0,0,0,0,13,0,114,0,255,0,0,0,30,0,153,0,64,0,162,0,0,0,180,0,0,0,254,0,12,0,42,0,54,0,0,0,145,0,179,0,119,0,116,0,237,0,145,0,0,0,38,0,203,0,89,0,33,0,187,0,149,0,107,0,0,0,0,0,199,0,0,0,243,0,0,0,18,0,233,0,125,0,194,0,0,0,88,0,179,0,154,0,48,0,190,0,203,0,229,0,117,0,227,0,0,0,199,0,184,0,0,0,133,0,112,0,101,0,49,0,45,0,21,0,78,0,234,0,32,0,0,0,229,0,126,0,178,0,209,0,0,0,60,0,38,0,191,0,65,0,0,0,243,0,155,0,69,0,110,0,133,0,241,0,15,0,64,0,95,0,227,0,75,0,42,0,182,0,146,0,209,0,95,0,116,0,119,0,0,0,2,0,253,0,0,0,69,0,90,0,216,0,127,0,250,0,192,0,209,0,250,0,190,0,0,0,34,0,175,0,0,0,0,0,34,0,68,0,0,0,48,0,72,0,40,0,4,0,44,0,0,0,182,0,128,0,196,0,38,0,192,0,237,0,245,0,84,0,156,0,139,0,105,0,0,0,252,0,174,0,139,0,0,0,134,0,155,0,0,0,39,0,206,0,197,0,84,0,221,0,0,0,91,0,49,0,23,0,228,0,247,0,153,0,235,0,12,0,98,0,41,0,0,0,176,0,151,0,104,0,124,0,0,0,165,0,76,0,129,0,42,0,57,0,188,0,227,0,0,0,56,0,0,0,128,0,244,0,238,0,180,0,130,0,127,0,0,0,0,0,249,0,0,0,129,0,67,0,205,0,162,0,0,0,111,0,0,0);
signal scenario_full  : scenario_type := (197,31,88,31,88,30,172,31,13,31,119,31,32,31,164,31,112,31,65,31,194,31,194,30,116,31,170,31,99,31,173,31,173,30,253,31,74,31,226,31,126,31,233,31,122,31,202,31,198,31,198,30,22,31,95,31,47,31,117,31,117,30,83,31,249,31,177,31,212,31,119,31,240,31,141,31,141,30,225,31,161,31,100,31,254,31,253,31,253,30,97,31,254,31,233,31,246,31,142,31,142,30,194,31,191,31,156,31,39,31,73,31,73,30,73,29,73,28,204,31,86,31,86,30,33,31,57,31,162,31,136,31,99,31,33,31,142,31,89,31,123,31,123,30,152,31,95,31,76,31,151,31,151,30,99,31,212,31,119,31,113,31,185,31,169,31,200,31,200,30,240,31,183,31,46,31,153,31,174,31,160,31,160,30,4,31,124,31,154,31,75,31,148,31,242,31,29,31,240,31,121,31,12,31,166,31,247,31,168,31,16,31,81,31,172,31,103,31,164,31,138,31,217,31,175,31,122,31,219,31,219,30,1,31,116,31,104,31,1,31,152,31,215,31,202,31,34,31,34,30,34,29,211,31,211,30,33,31,118,31,221,31,135,31,16,31,234,31,56,31,197,31,189,31,18,31,143,31,188,31,189,31,189,30,213,31,17,31,17,30,196,31,206,31,147,31,147,30,210,31,182,31,192,31,192,30,209,31,41,31,170,31,21,31,53,31,48,31,101,31,170,31,99,31,194,31,194,30,194,29,12,31,12,30,44,31,44,30,239,31,138,31,138,30,182,31,182,30,14,31,14,30,89,31,129,31,37,31,101,31,101,30,111,31,58,31,58,30,227,31,32,31,95,31,186,31,15,31,15,31,192,31,96,31,33,31,50,31,188,31,92,31,127,31,204,31,15,31,16,31,168,31,171,31,146,31,46,31,46,30,39,31,80,31,134,31,134,30,27,31,27,30,27,29,90,31,23,31,23,30,2,31,79,31,79,30,94,31,94,30,94,29,165,31,165,30,8,31,8,30,105,31,39,31,94,31,238,31,34,31,34,30,112,31,112,30,17,31,221,31,14,31,14,30,247,31,37,31,101,31,101,30,221,31,194,31,221,31,221,30,60,31,239,31,131,31,47,31,22,31,22,30,16,31,109,31,239,31,180,31,252,31,24,31,220,31,30,31,252,31,16,31,202,31,162,31,59,31,228,31,228,30,172,31,155,31,50,31,249,31,11,31,11,30,11,29,111,31,223,31,182,31,51,31,253,31,166,31,137,31,34,31,42,31,239,31,25,31,233,31,43,31,43,30,17,31,17,30,77,31,231,31,231,30,121,31,70,31,70,30,70,29,225,31,118,31,98,31,98,30,98,29,85,31,36,31,36,30,200,31,115,31,144,31,217,31,246,31,246,30,131,31,241,31,69,31,76,31,76,30,199,31,119,31,141,31,141,30,97,31,239,31,211,31,50,31,228,31,93,31,121,31,69,31,189,31,126,31,34,31,144,31,228,31,228,30,163,31,145,31,16,31,228,31,51,31,191,31,181,31,231,31,21,31,11,31,213,31,213,30,213,29,24,31,141,31,41,31,41,30,50,31,50,30,175,31,199,31,199,30,255,31,56,31,56,30,200,31,101,31,73,31,25,31,90,31,53,31,80,31,129,31,111,31,199,31,149,31,84,31,84,30,84,29,227,31,144,31,220,31,152,31,1,31,206,31,206,30,206,29,146,31,146,30,88,31,56,31,85,31,15,31,62,31,107,31,107,30,231,31,231,30,19,31,162,31,162,30,162,29,53,31,224,31,38,31,114,31,21,31,21,30,156,31,14,31,14,30,62,31,235,31,235,30,62,31,110,31,202,31,191,31,16,31,225,31,202,31,202,30,202,29,122,31,108,31,108,30,108,29,29,31,29,30,55,31,173,31,242,31,127,31,18,31,41,31,52,31,164,31,75,31,22,31,36,31,53,31,53,30,169,31,169,30,169,29,126,31,226,31,226,30,226,29,117,31,100,31,199,31,81,31,81,30,18,31,41,31,164,31,97,31,97,30,94,31,94,30,21,31,136,31,136,30,255,31,142,31,12,31,12,30,15,31,164,31,154,31,70,31,70,30,144,31,254,31,254,30,74,31,34,31,169,31,225,31,225,30,241,31,3,31,3,31,79,31,248,31,162,31,120,31,120,30,242,31,103,31,103,30,103,29,101,31,217,31,87,31,87,30,234,31,253,31,139,31,160,31,167,31,237,31,186,31,49,31,55,31,33,31,30,31,120,31,196,31,231,31,171,31,134,31,111,31,187,31,66,31,47,31,47,30,101,31,237,31,89,31,91,31,95,31,95,30,180,31,200,31,3,31,3,30,3,29,59,31,36,31,136,31,169,31,103,31,160,31,29,31,29,30,29,29,29,28,82,31,82,30,82,29,13,31,114,31,255,31,255,30,30,31,153,31,64,31,162,31,162,30,180,31,180,30,254,31,12,31,42,31,54,31,54,30,145,31,179,31,119,31,116,31,237,31,145,31,145,30,38,31,203,31,89,31,33,31,187,31,149,31,107,31,107,30,107,29,199,31,199,30,243,31,243,30,18,31,233,31,125,31,194,31,194,30,88,31,179,31,154,31,48,31,190,31,203,31,229,31,117,31,227,31,227,30,199,31,184,31,184,30,133,31,112,31,101,31,49,31,45,31,21,31,78,31,234,31,32,31,32,30,229,31,126,31,178,31,209,31,209,30,60,31,38,31,191,31,65,31,65,30,243,31,155,31,69,31,110,31,133,31,241,31,15,31,64,31,95,31,227,31,75,31,42,31,182,31,146,31,209,31,95,31,116,31,119,31,119,30,2,31,253,31,253,30,69,31,90,31,216,31,127,31,250,31,192,31,209,31,250,31,190,31,190,30,34,31,175,31,175,30,175,29,34,31,68,31,68,30,48,31,72,31,40,31,4,31,44,31,44,30,182,31,128,31,196,31,38,31,192,31,237,31,245,31,84,31,156,31,139,31,105,31,105,30,252,31,174,31,139,31,139,30,134,31,155,31,155,30,39,31,206,31,197,31,84,31,221,31,221,30,91,31,49,31,23,31,228,31,247,31,153,31,235,31,12,31,98,31,41,31,41,30,176,31,151,31,104,31,124,31,124,30,165,31,76,31,129,31,42,31,57,31,188,31,227,31,227,30,56,31,56,30,128,31,244,31,238,31,180,31,130,31,127,31,127,30,127,29,249,31,249,30,129,31,67,31,205,31,162,31,162,30,111,31,111,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
