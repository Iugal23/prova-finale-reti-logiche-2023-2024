-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 171;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (190,0,40,0,67,0,52,0,213,0,135,0,110,0,214,0,249,0,0,0,96,0,0,0,234,0,139,0,59,0,244,0,178,0,146,0,149,0,204,0,0,0,209,0,185,0,153,0,226,0,66,0,242,0,58,0,3,0,0,0,120,0,217,0,47,0,206,0,111,0,0,0,157,0,238,0,123,0,161,0,46,0,187,0,61,0,186,0,235,0,130,0,187,0,168,0,41,0,0,0,39,0,139,0,0,0,220,0,0,0,0,0,35,0,187,0,34,0,0,0,43,0,188,0,144,0,241,0,72,0,76,0,213,0,0,0,0,0,0,0,21,0,228,0,0,0,237,0,86,0,0,0,67,0,119,0,59,0,0,0,240,0,107,0,48,0,18,0,251,0,0,0,4,0,138,0,206,0,28,0,95,0,140,0,200,0,186,0,160,0,255,0,46,0,45,0,70,0,229,0,0,0,8,0,145,0,236,0,54,0,198,0,134,0,0,0,6,0,175,0,54,0,91,0,0,0,183,0,106,0,89,0,0,0,174,0,132,0,0,0,230,0,119,0,103,0,80,0,105,0,0,0,246,0,175,0,1,0,91,0,78,0,229,0,19,0,0,0,174,0,226,0,142,0,0,0,0,0,229,0,168,0,35,0,75,0,164,0,65,0,0,0,28,0,171,0,240,0,0,0,254,0,141,0,0,0,42,0,249,0,31,0,74,0,87,0,0,0,221,0,203,0,149,0,134,0,0,0,149,0,228,0,112,0,48,0,26,0,47,0,40,0);
signal scenario_full  : scenario_type := (190,31,40,31,67,31,52,31,213,31,135,31,110,31,214,31,249,31,249,30,96,31,96,30,234,31,139,31,59,31,244,31,178,31,146,31,149,31,204,31,204,30,209,31,185,31,153,31,226,31,66,31,242,31,58,31,3,31,3,30,120,31,217,31,47,31,206,31,111,31,111,30,157,31,238,31,123,31,161,31,46,31,187,31,61,31,186,31,235,31,130,31,187,31,168,31,41,31,41,30,39,31,139,31,139,30,220,31,220,30,220,29,35,31,187,31,34,31,34,30,43,31,188,31,144,31,241,31,72,31,76,31,213,31,213,30,213,29,213,28,21,31,228,31,228,30,237,31,86,31,86,30,67,31,119,31,59,31,59,30,240,31,107,31,48,31,18,31,251,31,251,30,4,31,138,31,206,31,28,31,95,31,140,31,200,31,186,31,160,31,255,31,46,31,45,31,70,31,229,31,229,30,8,31,145,31,236,31,54,31,198,31,134,31,134,30,6,31,175,31,54,31,91,31,91,30,183,31,106,31,89,31,89,30,174,31,132,31,132,30,230,31,119,31,103,31,80,31,105,31,105,30,246,31,175,31,1,31,91,31,78,31,229,31,19,31,19,30,174,31,226,31,142,31,142,30,142,29,229,31,168,31,35,31,75,31,164,31,65,31,65,30,28,31,171,31,240,31,240,30,254,31,141,31,141,30,42,31,249,31,31,31,74,31,87,31,87,30,221,31,203,31,149,31,134,31,134,30,149,31,228,31,112,31,48,31,26,31,47,31,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
