-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_780 is
end project_tb_780;

architecture project_tb_arch_780 of project_tb_780 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 587;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (3,0,233,0,59,0,246,0,40,0,198,0,240,0,212,0,194,0,0,0,0,0,197,0,0,0,0,0,1,0,0,0,89,0,59,0,143,0,36,0,223,0,140,0,105,0,55,0,254,0,88,0,230,0,0,0,245,0,0,0,3,0,0,0,48,0,0,0,68,0,104,0,238,0,0,0,224,0,165,0,7,0,0,0,39,0,244,0,225,0,92,0,202,0,231,0,114,0,22,0,164,0,103,0,80,0,209,0,185,0,48,0,0,0,157,0,39,0,4,0,59,0,30,0,133,0,144,0,214,0,0,0,209,0,106,0,121,0,174,0,95,0,26,0,242,0,249,0,102,0,0,0,149,0,74,0,106,0,0,0,17,0,220,0,187,0,178,0,49,0,172,0,127,0,65,0,45,0,100,0,0,0,44,0,44,0,67,0,236,0,0,0,171,0,23,0,220,0,70,0,223,0,95,0,59,0,238,0,124,0,0,0,0,0,55,0,20,0,130,0,215,0,86,0,0,0,132,0,201,0,39,0,143,0,172,0,4,0,94,0,228,0,81,0,0,0,125,0,0,0,204,0,179,0,212,0,117,0,110,0,117,0,74,0,81,0,212,0,62,0,201,0,118,0,139,0,0,0,0,0,179,0,30,0,0,0,23,0,248,0,180,0,187,0,0,0,54,0,0,0,116,0,209,0,0,0,128,0,126,0,0,0,0,0,233,0,46,0,114,0,0,0,58,0,0,0,0,0,0,0,40,0,0,0,115,0,252,0,0,0,98,0,223,0,0,0,87,0,215,0,37,0,152,0,207,0,201,0,0,0,210,0,0,0,122,0,0,0,198,0,208,0,152,0,203,0,0,0,109,0,203,0,250,0,25,0,0,0,53,0,232,0,120,0,108,0,235,0,0,0,0,0,222,0,0,0,108,0,0,0,113,0,65,0,95,0,143,0,196,0,176,0,0,0,209,0,199,0,83,0,82,0,74,0,0,0,181,0,179,0,229,0,0,0,0,0,76,0,132,0,0,0,85,0,0,0,161,0,132,0,3,0,118,0,213,0,96,0,70,0,6,0,248,0,0,0,240,0,0,0,117,0,65,0,147,0,0,0,22,0,134,0,61,0,112,0,0,0,170,0,0,0,233,0,240,0,0,0,87,0,78,0,0,0,177,0,16,0,16,0,115,0,199,0,23,0,17,0,189,0,32,0,15,0,0,0,227,0,128,0,0,0,29,0,230,0,106,0,13,0,205,0,234,0,81,0,95,0,254,0,150,0,201,0,0,0,133,0,203,0,162,0,69,0,36,0,76,0,141,0,0,0,14,0,21,0,57,0,12,0,0,0,115,0,217,0,212,0,0,0,0,0,151,0,190,0,27,0,180,0,190,0,166,0,250,0,19,0,188,0,162,0,85,0,234,0,14,0,78,0,95,0,113,0,0,0,0,0,0,0,162,0,192,0,0,0,0,0,251,0,119,0,10,0,191,0,131,0,228,0,205,0,92,0,0,0,0,0,0,0,224,0,169,0,134,0,117,0,125,0,127,0,0,0,238,0,234,0,148,0,34,0,186,0,135,0,96,0,249,0,44,0,106,0,171,0,92,0,113,0,0,0,0,0,0,0,1,0,160,0,224,0,237,0,0,0,0,0,5,0,137,0,43,0,207,0,237,0,0,0,102,0,0,0,139,0,0,0,11,0,0,0,245,0,129,0,200,0,156,0,52,0,212,0,0,0,152,0,60,0,32,0,85,0,208,0,55,0,195,0,123,0,46,0,0,0,161,0,0,0,217,0,168,0,23,0,219,0,147,0,203,0,19,0,127,0,212,0,0,0,128,0,173,0,109,0,84,0,86,0,63,0,76,0,29,0,154,0,37,0,0,0,237,0,164,0,167,0,167,0,219,0,95,0,0,0,142,0,0,0,9,0,99,0,67,0,0,0,147,0,0,0,236,0,64,0,6,0,149,0,28,0,61,0,166,0,134,0,42,0,64,0,56,0,254,0,35,0,26,0,177,0,58,0,156,0,0,0,0,0,222,0,151,0,0,0,211,0,178,0,69,0,75,0,199,0,101,0,0,0,0,0,162,0,0,0,0,0,144,0,18,0,149,0,148,0,224,0,0,0,0,0,121,0,147,0,0,0,87,0,0,0,50,0,150,0,54,0,231,0,245,0,231,0,23,0,179,0,2,0,125,0,125,0,176,0,0,0,114,0,59,0,0,0,91,0,43,0,144,0,238,0,230,0,9,0,229,0,122,0,207,0,175,0,208,0,0,0,143,0,0,0,128,0,69,0,205,0,0,0,149,0,0,0,127,0,157,0,69,0,109,0,0,0,116,0,251,0,125,0,136,0,0,0,208,0,99,0,212,0,197,0,120,0,116,0,26,0,223,0,174,0,222,0,113,0,0,0,97,0,169,0,0,0,0,0,131,0,0,0,98,0,175,0,0,0,94,0,222,0,226,0,0,0,147,0,173,0,164,0,0,0,0,0,189,0,0,0,130,0,101,0,0,0,152,0,173,0,167,0,0,0,0,0,38,0,0,0,171,0,171,0,0,0,213,0,67,0,238,0,157,0,22,0,190,0,84,0,91,0,0,0,151,0,185,0,190,0,0,0,144,0,197,0,73,0,136,0,92,0,209,0,132,0);
signal scenario_full  : scenario_type := (3,31,233,31,59,31,246,31,40,31,198,31,240,31,212,31,194,31,194,30,194,29,197,31,197,30,197,29,1,31,1,30,89,31,59,31,143,31,36,31,223,31,140,31,105,31,55,31,254,31,88,31,230,31,230,30,245,31,245,30,3,31,3,30,48,31,48,30,68,31,104,31,238,31,238,30,224,31,165,31,7,31,7,30,39,31,244,31,225,31,92,31,202,31,231,31,114,31,22,31,164,31,103,31,80,31,209,31,185,31,48,31,48,30,157,31,39,31,4,31,59,31,30,31,133,31,144,31,214,31,214,30,209,31,106,31,121,31,174,31,95,31,26,31,242,31,249,31,102,31,102,30,149,31,74,31,106,31,106,30,17,31,220,31,187,31,178,31,49,31,172,31,127,31,65,31,45,31,100,31,100,30,44,31,44,31,67,31,236,31,236,30,171,31,23,31,220,31,70,31,223,31,95,31,59,31,238,31,124,31,124,30,124,29,55,31,20,31,130,31,215,31,86,31,86,30,132,31,201,31,39,31,143,31,172,31,4,31,94,31,228,31,81,31,81,30,125,31,125,30,204,31,179,31,212,31,117,31,110,31,117,31,74,31,81,31,212,31,62,31,201,31,118,31,139,31,139,30,139,29,179,31,30,31,30,30,23,31,248,31,180,31,187,31,187,30,54,31,54,30,116,31,209,31,209,30,128,31,126,31,126,30,126,29,233,31,46,31,114,31,114,30,58,31,58,30,58,29,58,28,40,31,40,30,115,31,252,31,252,30,98,31,223,31,223,30,87,31,215,31,37,31,152,31,207,31,201,31,201,30,210,31,210,30,122,31,122,30,198,31,208,31,152,31,203,31,203,30,109,31,203,31,250,31,25,31,25,30,53,31,232,31,120,31,108,31,235,31,235,30,235,29,222,31,222,30,108,31,108,30,113,31,65,31,95,31,143,31,196,31,176,31,176,30,209,31,199,31,83,31,82,31,74,31,74,30,181,31,179,31,229,31,229,30,229,29,76,31,132,31,132,30,85,31,85,30,161,31,132,31,3,31,118,31,213,31,96,31,70,31,6,31,248,31,248,30,240,31,240,30,117,31,65,31,147,31,147,30,22,31,134,31,61,31,112,31,112,30,170,31,170,30,233,31,240,31,240,30,87,31,78,31,78,30,177,31,16,31,16,31,115,31,199,31,23,31,17,31,189,31,32,31,15,31,15,30,227,31,128,31,128,30,29,31,230,31,106,31,13,31,205,31,234,31,81,31,95,31,254,31,150,31,201,31,201,30,133,31,203,31,162,31,69,31,36,31,76,31,141,31,141,30,14,31,21,31,57,31,12,31,12,30,115,31,217,31,212,31,212,30,212,29,151,31,190,31,27,31,180,31,190,31,166,31,250,31,19,31,188,31,162,31,85,31,234,31,14,31,78,31,95,31,113,31,113,30,113,29,113,28,162,31,192,31,192,30,192,29,251,31,119,31,10,31,191,31,131,31,228,31,205,31,92,31,92,30,92,29,92,28,224,31,169,31,134,31,117,31,125,31,127,31,127,30,238,31,234,31,148,31,34,31,186,31,135,31,96,31,249,31,44,31,106,31,171,31,92,31,113,31,113,30,113,29,113,28,1,31,160,31,224,31,237,31,237,30,237,29,5,31,137,31,43,31,207,31,237,31,237,30,102,31,102,30,139,31,139,30,11,31,11,30,245,31,129,31,200,31,156,31,52,31,212,31,212,30,152,31,60,31,32,31,85,31,208,31,55,31,195,31,123,31,46,31,46,30,161,31,161,30,217,31,168,31,23,31,219,31,147,31,203,31,19,31,127,31,212,31,212,30,128,31,173,31,109,31,84,31,86,31,63,31,76,31,29,31,154,31,37,31,37,30,237,31,164,31,167,31,167,31,219,31,95,31,95,30,142,31,142,30,9,31,99,31,67,31,67,30,147,31,147,30,236,31,64,31,6,31,149,31,28,31,61,31,166,31,134,31,42,31,64,31,56,31,254,31,35,31,26,31,177,31,58,31,156,31,156,30,156,29,222,31,151,31,151,30,211,31,178,31,69,31,75,31,199,31,101,31,101,30,101,29,162,31,162,30,162,29,144,31,18,31,149,31,148,31,224,31,224,30,224,29,121,31,147,31,147,30,87,31,87,30,50,31,150,31,54,31,231,31,245,31,231,31,23,31,179,31,2,31,125,31,125,31,176,31,176,30,114,31,59,31,59,30,91,31,43,31,144,31,238,31,230,31,9,31,229,31,122,31,207,31,175,31,208,31,208,30,143,31,143,30,128,31,69,31,205,31,205,30,149,31,149,30,127,31,157,31,69,31,109,31,109,30,116,31,251,31,125,31,136,31,136,30,208,31,99,31,212,31,197,31,120,31,116,31,26,31,223,31,174,31,222,31,113,31,113,30,97,31,169,31,169,30,169,29,131,31,131,30,98,31,175,31,175,30,94,31,222,31,226,31,226,30,147,31,173,31,164,31,164,30,164,29,189,31,189,30,130,31,101,31,101,30,152,31,173,31,167,31,167,30,167,29,38,31,38,30,171,31,171,31,171,30,213,31,67,31,238,31,157,31,22,31,190,31,84,31,91,31,91,30,151,31,185,31,190,31,190,30,144,31,197,31,73,31,136,31,92,31,209,31,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
