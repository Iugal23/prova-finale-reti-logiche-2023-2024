-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 206;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,16,0,217,0,59,0,169,0,165,0,93,0,53,0,0,0,108,0,0,0,12,0,57,0,141,0,105,0,0,0,0,0,176,0,0,0,82,0,41,0,225,0,0,0,181,0,61,0,50,0,141,0,226,0,66,0,203,0,149,0,225,0,182,0,231,0,0,0,66,0,0,0,191,0,164,0,197,0,180,0,174,0,231,0,130,0,12,0,157,0,29,0,0,0,106,0,168,0,0,0,175,0,14,0,145,0,190,0,199,0,181,0,13,0,0,0,0,0,230,0,0,0,99,0,0,0,175,0,201,0,0,0,36,0,159,0,173,0,0,0,0,0,127,0,229,0,249,0,138,0,172,0,188,0,165,0,183,0,71,0,0,0,118,0,50,0,226,0,165,0,179,0,0,0,0,0,191,0,44,0,0,0,35,0,0,0,160,0,92,0,33,0,238,0,114,0,155,0,0,0,57,0,222,0,108,0,240,0,178,0,6,0,179,0,0,0,38,0,1,0,56,0,131,0,32,0,116,0,0,0,26,0,208,0,214,0,8,0,0,0,56,0,0,0,245,0,162,0,83,0,0,0,22,0,239,0,230,0,140,0,10,0,0,0,246,0,142,0,229,0,59,0,161,0,0,0,156,0,61,0,168,0,207,0,189,0,108,0,248,0,91,0,245,0,52,0,93,0,186,0,233,0,117,0,67,0,238,0,131,0,21,0,0,0,228,0,248,0,185,0,234,0,124,0,9,0,117,0,0,0,125,0,0,0,0,0,125,0,117,0,224,0,45,0,167,0,250,0,47,0,174,0,187,0,6,0,250,0,62,0,56,0,168,0,0,0,37,0,20,0,27,0,71,0,0,0,60,0,154,0,15,0,229,0,88,0,11,0,0,0,234,0,145,0,161,0,232,0,158,0,0,0,172,0,0,0,15,0,204,0);
signal scenario_full  : scenario_type := (0,0,16,31,217,31,59,31,169,31,165,31,93,31,53,31,53,30,108,31,108,30,12,31,57,31,141,31,105,31,105,30,105,29,176,31,176,30,82,31,41,31,225,31,225,30,181,31,61,31,50,31,141,31,226,31,66,31,203,31,149,31,225,31,182,31,231,31,231,30,66,31,66,30,191,31,164,31,197,31,180,31,174,31,231,31,130,31,12,31,157,31,29,31,29,30,106,31,168,31,168,30,175,31,14,31,145,31,190,31,199,31,181,31,13,31,13,30,13,29,230,31,230,30,99,31,99,30,175,31,201,31,201,30,36,31,159,31,173,31,173,30,173,29,127,31,229,31,249,31,138,31,172,31,188,31,165,31,183,31,71,31,71,30,118,31,50,31,226,31,165,31,179,31,179,30,179,29,191,31,44,31,44,30,35,31,35,30,160,31,92,31,33,31,238,31,114,31,155,31,155,30,57,31,222,31,108,31,240,31,178,31,6,31,179,31,179,30,38,31,1,31,56,31,131,31,32,31,116,31,116,30,26,31,208,31,214,31,8,31,8,30,56,31,56,30,245,31,162,31,83,31,83,30,22,31,239,31,230,31,140,31,10,31,10,30,246,31,142,31,229,31,59,31,161,31,161,30,156,31,61,31,168,31,207,31,189,31,108,31,248,31,91,31,245,31,52,31,93,31,186,31,233,31,117,31,67,31,238,31,131,31,21,31,21,30,228,31,248,31,185,31,234,31,124,31,9,31,117,31,117,30,125,31,125,30,125,29,125,31,117,31,224,31,45,31,167,31,250,31,47,31,174,31,187,31,6,31,250,31,62,31,56,31,168,31,168,30,37,31,20,31,27,31,71,31,71,30,60,31,154,31,15,31,229,31,88,31,11,31,11,30,234,31,145,31,161,31,232,31,158,31,158,30,172,31,172,30,15,31,204,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
