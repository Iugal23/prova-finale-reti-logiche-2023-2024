-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 744;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (77,0,202,0,70,0,0,0,0,0,228,0,243,0,33,0,252,0,130,0,0,0,19,0,207,0,147,0,47,0,244,0,25,0,39,0,168,0,224,0,0,0,82,0,27,0,78,0,172,0,52,0,4,0,89,0,243,0,95,0,0,0,146,0,236,0,229,0,56,0,171,0,198,0,0,0,117,0,0,0,27,0,90,0,0,0,0,0,103,0,115,0,0,0,81,0,202,0,1,0,211,0,0,0,3,0,0,0,93,0,6,0,196,0,0,0,116,0,0,0,63,0,6,0,0,0,131,0,172,0,197,0,219,0,0,0,191,0,43,0,0,0,0,0,58,0,178,0,227,0,0,0,31,0,167,0,215,0,186,0,74,0,68,0,0,0,233,0,203,0,44,0,129,0,223,0,69,0,0,0,35,0,164,0,94,0,197,0,115,0,170,0,40,0,0,0,94,0,113,0,0,0,242,0,214,0,200,0,15,0,210,0,90,0,40,0,0,0,30,0,84,0,0,0,0,0,168,0,8,0,136,0,225,0,229,0,0,0,0,0,41,0,22,0,0,0,28,0,237,0,84,0,61,0,37,0,235,0,0,0,228,0,125,0,33,0,9,0,209,0,165,0,0,0,186,0,0,0,204,0,255,0,19,0,140,0,238,0,0,0,100,0,68,0,0,0,193,0,0,0,195,0,153,0,175,0,102,0,28,0,0,0,218,0,61,0,0,0,12,0,120,0,195,0,0,0,0,0,67,0,78,0,187,0,191,0,0,0,133,0,0,0,94,0,62,0,24,0,35,0,0,0,0,0,93,0,52,0,0,0,0,0,176,0,246,0,0,0,76,0,198,0,76,0,111,0,3,0,0,0,145,0,0,0,97,0,229,0,56,0,123,0,0,0,179,0,163,0,0,0,174,0,232,0,0,0,38,0,83,0,0,0,148,0,145,0,90,0,105,0,140,0,26,0,138,0,26,0,0,0,0,0,0,0,17,0,58,0,26,0,14,0,0,0,91,0,46,0,0,0,190,0,165,0,0,0,203,0,40,0,176,0,131,0,196,0,242,0,102,0,202,0,146,0,28,0,0,0,248,0,245,0,40,0,160,0,0,0,140,0,32,0,141,0,210,0,0,0,98,0,56,0,125,0,0,0,65,0,126,0,0,0,200,0,0,0,159,0,251,0,184,0,88,0,82,0,81,0,38,0,0,0,239,0,144,0,192,0,167,0,235,0,132,0,0,0,149,0,92,0,173,0,0,0,188,0,116,0,43,0,18,0,116,0,0,0,0,0,37,0,159,0,86,0,0,0,96,0,158,0,209,0,229,0,67,0,245,0,161,0,121,0,148,0,118,0,243,0,0,0,167,0,231,0,163,0,91,0,255,0,175,0,206,0,129,0,156,0,0,0,186,0,239,0,230,0,103,0,3,0,199,0,184,0,76,0,9,0,65,0,94,0,10,0,0,0,110,0,133,0,218,0,182,0,169,0,40,0,180,0,0,0,16,0,185,0,153,0,222,0,202,0,103,0,46,0,118,0,234,0,121,0,225,0,72,0,173,0,239,0,174,0,181,0,64,0,193,0,0,0,5,0,29,0,0,0,205,0,217,0,83,0,202,0,141,0,0,0,13,0,100,0,37,0,156,0,0,0,21,0,238,0,107,0,189,0,0,0,111,0,35,0,177,0,90,0,235,0,70,0,42,0,37,0,49,0,0,0,200,0,148,0,111,0,199,0,125,0,39,0,0,0,32,0,242,0,75,0,0,0,163,0,190,0,138,0,111,0,155,0,115,0,0,0,170,0,213,0,0,0,3,0,229,0,1,0,150,0,50,0,157,0,136,0,0,0,234,0,0,0,102,0,255,0,191,0,65,0,146,0,20,0,0,0,158,0,46,0,0,0,114,0,0,0,208,0,131,0,94,0,0,0,0,0,0,0,60,0,58,0,0,0,0,0,201,0,218,0,53,0,0,0,14,0,195,0,23,0,9,0,0,0,2,0,96,0,33,0,203,0,86,0,160,0,126,0,239,0,0,0,189,0,202,0,0,0,60,0,247,0,192,0,139,0,0,0,106,0,209,0,241,0,156,0,0,0,36,0,42,0,38,0,0,0,0,0,88,0,38,0,11,0,115,0,36,0,145,0,211,0,120,0,0,0,5,0,11,0,77,0,66,0,241,0,126,0,112,0,45,0,109,0,10,0,132,0,129,0,214,0,167,0,0,0,0,0,202,0,114,0,76,0,0,0,141,0,139,0,0,0,35,0,22,0,0,0,29,0,20,0,33,0,0,0,0,0,125,0,96,0,0,0,153,0,50,0,0,0,192,0,96,0,199,0,144,0,91,0,0,0,102,0,207,0,94,0,137,0,0,0,176,0,248,0,151,0,127,0,0,0,54,0,229,0,223,0,0,0,154,0,184,0,56,0,249,0,154,0,28,0,0,0,216,0,13,0,119,0,92,0,49,0,0,0,218,0,82,0,112,0,219,0,0,0,174,0,0,0,35,0,0,0,4,0,190,0,226,0,192,0,236,0,125,0,19,0,87,0,109,0,206,0,147,0,194,0,166,0,252,0,19,0,86,0,89,0,230,0,222,0,0,0,200,0,209,0,0,0,196,0,32,0,82,0,98,0,41,0,147,0,0,0,42,0,29,0,136,0,49,0,204,0,0,0,0,0,103,0,38,0,252,0,149,0,59,0,0,0,253,0,237,0,0,0,0,0,75,0,0,0,128,0,0,0,0,0,242,0,201,0,146,0,0,0,244,0,120,0,44,0,114,0,166,0,234,0,133,0,180,0,73,0,247,0,185,0,143,0,35,0,37,0,137,0,39,0,183,0,2,0,36,0,203,0,0,0,247,0,201,0,122,0,0,0,124,0,157,0,205,0,0,0,106,0,202,0,41,0,161,0,0,0,157,0,0,0,0,0,181,0,226,0,0,0,37,0,0,0,133,0,76,0,170,0,194,0,0,0,215,0,0,0,117,0,176,0,0,0,174,0,0,0,17,0,186,0,228,0,0,0,0,0,41,0,237,0,133,0,198,0,215,0,68,0,42,0,0,0,187,0,0,0,0,0,104,0,22,0,174,0,247,0,102,0,158,0,220,0,150,0,0,0,184,0,189,0,0,0,0,0,67,0,8,0,219,0,0,0,0,0,0,0,157,0,182,0,0,0,153,0,219,0,15,0,149,0,149,0,190,0,110,0,36,0,0,0,67,0,82,0,14,0,0,0,23,0,64,0,89,0,72,0,92,0,140,0,0,0,208,0,151,0,170,0,206,0,0,0,251,0,14,0,116,0,241,0,74,0,227,0,210,0,252,0,212,0,242,0,7,0,0,0,243,0,151,0,50,0);
signal scenario_full  : scenario_type := (77,31,202,31,70,31,70,30,70,29,228,31,243,31,33,31,252,31,130,31,130,30,19,31,207,31,147,31,47,31,244,31,25,31,39,31,168,31,224,31,224,30,82,31,27,31,78,31,172,31,52,31,4,31,89,31,243,31,95,31,95,30,146,31,236,31,229,31,56,31,171,31,198,31,198,30,117,31,117,30,27,31,90,31,90,30,90,29,103,31,115,31,115,30,81,31,202,31,1,31,211,31,211,30,3,31,3,30,93,31,6,31,196,31,196,30,116,31,116,30,63,31,6,31,6,30,131,31,172,31,197,31,219,31,219,30,191,31,43,31,43,30,43,29,58,31,178,31,227,31,227,30,31,31,167,31,215,31,186,31,74,31,68,31,68,30,233,31,203,31,44,31,129,31,223,31,69,31,69,30,35,31,164,31,94,31,197,31,115,31,170,31,40,31,40,30,94,31,113,31,113,30,242,31,214,31,200,31,15,31,210,31,90,31,40,31,40,30,30,31,84,31,84,30,84,29,168,31,8,31,136,31,225,31,229,31,229,30,229,29,41,31,22,31,22,30,28,31,237,31,84,31,61,31,37,31,235,31,235,30,228,31,125,31,33,31,9,31,209,31,165,31,165,30,186,31,186,30,204,31,255,31,19,31,140,31,238,31,238,30,100,31,68,31,68,30,193,31,193,30,195,31,153,31,175,31,102,31,28,31,28,30,218,31,61,31,61,30,12,31,120,31,195,31,195,30,195,29,67,31,78,31,187,31,191,31,191,30,133,31,133,30,94,31,62,31,24,31,35,31,35,30,35,29,93,31,52,31,52,30,52,29,176,31,246,31,246,30,76,31,198,31,76,31,111,31,3,31,3,30,145,31,145,30,97,31,229,31,56,31,123,31,123,30,179,31,163,31,163,30,174,31,232,31,232,30,38,31,83,31,83,30,148,31,145,31,90,31,105,31,140,31,26,31,138,31,26,31,26,30,26,29,26,28,17,31,58,31,26,31,14,31,14,30,91,31,46,31,46,30,190,31,165,31,165,30,203,31,40,31,176,31,131,31,196,31,242,31,102,31,202,31,146,31,28,31,28,30,248,31,245,31,40,31,160,31,160,30,140,31,32,31,141,31,210,31,210,30,98,31,56,31,125,31,125,30,65,31,126,31,126,30,200,31,200,30,159,31,251,31,184,31,88,31,82,31,81,31,38,31,38,30,239,31,144,31,192,31,167,31,235,31,132,31,132,30,149,31,92,31,173,31,173,30,188,31,116,31,43,31,18,31,116,31,116,30,116,29,37,31,159,31,86,31,86,30,96,31,158,31,209,31,229,31,67,31,245,31,161,31,121,31,148,31,118,31,243,31,243,30,167,31,231,31,163,31,91,31,255,31,175,31,206,31,129,31,156,31,156,30,186,31,239,31,230,31,103,31,3,31,199,31,184,31,76,31,9,31,65,31,94,31,10,31,10,30,110,31,133,31,218,31,182,31,169,31,40,31,180,31,180,30,16,31,185,31,153,31,222,31,202,31,103,31,46,31,118,31,234,31,121,31,225,31,72,31,173,31,239,31,174,31,181,31,64,31,193,31,193,30,5,31,29,31,29,30,205,31,217,31,83,31,202,31,141,31,141,30,13,31,100,31,37,31,156,31,156,30,21,31,238,31,107,31,189,31,189,30,111,31,35,31,177,31,90,31,235,31,70,31,42,31,37,31,49,31,49,30,200,31,148,31,111,31,199,31,125,31,39,31,39,30,32,31,242,31,75,31,75,30,163,31,190,31,138,31,111,31,155,31,115,31,115,30,170,31,213,31,213,30,3,31,229,31,1,31,150,31,50,31,157,31,136,31,136,30,234,31,234,30,102,31,255,31,191,31,65,31,146,31,20,31,20,30,158,31,46,31,46,30,114,31,114,30,208,31,131,31,94,31,94,30,94,29,94,28,60,31,58,31,58,30,58,29,201,31,218,31,53,31,53,30,14,31,195,31,23,31,9,31,9,30,2,31,96,31,33,31,203,31,86,31,160,31,126,31,239,31,239,30,189,31,202,31,202,30,60,31,247,31,192,31,139,31,139,30,106,31,209,31,241,31,156,31,156,30,36,31,42,31,38,31,38,30,38,29,88,31,38,31,11,31,115,31,36,31,145,31,211,31,120,31,120,30,5,31,11,31,77,31,66,31,241,31,126,31,112,31,45,31,109,31,10,31,132,31,129,31,214,31,167,31,167,30,167,29,202,31,114,31,76,31,76,30,141,31,139,31,139,30,35,31,22,31,22,30,29,31,20,31,33,31,33,30,33,29,125,31,96,31,96,30,153,31,50,31,50,30,192,31,96,31,199,31,144,31,91,31,91,30,102,31,207,31,94,31,137,31,137,30,176,31,248,31,151,31,127,31,127,30,54,31,229,31,223,31,223,30,154,31,184,31,56,31,249,31,154,31,28,31,28,30,216,31,13,31,119,31,92,31,49,31,49,30,218,31,82,31,112,31,219,31,219,30,174,31,174,30,35,31,35,30,4,31,190,31,226,31,192,31,236,31,125,31,19,31,87,31,109,31,206,31,147,31,194,31,166,31,252,31,19,31,86,31,89,31,230,31,222,31,222,30,200,31,209,31,209,30,196,31,32,31,82,31,98,31,41,31,147,31,147,30,42,31,29,31,136,31,49,31,204,31,204,30,204,29,103,31,38,31,252,31,149,31,59,31,59,30,253,31,237,31,237,30,237,29,75,31,75,30,128,31,128,30,128,29,242,31,201,31,146,31,146,30,244,31,120,31,44,31,114,31,166,31,234,31,133,31,180,31,73,31,247,31,185,31,143,31,35,31,37,31,137,31,39,31,183,31,2,31,36,31,203,31,203,30,247,31,201,31,122,31,122,30,124,31,157,31,205,31,205,30,106,31,202,31,41,31,161,31,161,30,157,31,157,30,157,29,181,31,226,31,226,30,37,31,37,30,133,31,76,31,170,31,194,31,194,30,215,31,215,30,117,31,176,31,176,30,174,31,174,30,17,31,186,31,228,31,228,30,228,29,41,31,237,31,133,31,198,31,215,31,68,31,42,31,42,30,187,31,187,30,187,29,104,31,22,31,174,31,247,31,102,31,158,31,220,31,150,31,150,30,184,31,189,31,189,30,189,29,67,31,8,31,219,31,219,30,219,29,219,28,157,31,182,31,182,30,153,31,219,31,15,31,149,31,149,31,190,31,110,31,36,31,36,30,67,31,82,31,14,31,14,30,23,31,64,31,89,31,72,31,92,31,140,31,140,30,208,31,151,31,170,31,206,31,206,30,251,31,14,31,116,31,241,31,74,31,227,31,210,31,252,31,212,31,242,31,7,31,7,30,243,31,151,31,50,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
