-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_340 is
end project_tb_340;

architecture project_tb_arch_340 of project_tb_340 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 911;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (53,0,0,0,179,0,156,0,0,0,246,0,36,0,149,0,113,0,0,0,209,0,70,0,186,0,7,0,5,0,55,0,0,0,0,0,0,0,119,0,110,0,248,0,105,0,195,0,114,0,21,0,179,0,0,0,187,0,0,0,120,0,159,0,0,0,66,0,210,0,215,0,229,0,102,0,94,0,185,0,138,0,85,0,187,0,45,0,225,0,184,0,149,0,93,0,156,0,99,0,0,0,62,0,0,0,44,0,241,0,127,0,0,0,132,0,112,0,56,0,0,0,144,0,37,0,25,0,106,0,22,0,148,0,191,0,188,0,194,0,170,0,252,0,95,0,0,0,166,0,18,0,136,0,201,0,143,0,179,0,183,0,228,0,10,0,242,0,0,0,138,0,152,0,200,0,15,0,0,0,0,0,220,0,55,0,123,0,96,0,90,0,0,0,0,0,154,0,20,0,174,0,232,0,178,0,49,0,222,0,25,0,0,0,38,0,5,0,234,0,0,0,234,0,236,0,0,0,72,0,83,0,230,0,37,0,188,0,93,0,0,0,240,0,0,0,239,0,161,0,0,0,75,0,189,0,166,0,16,0,59,0,113,0,207,0,192,0,144,0,0,0,53,0,0,0,189,0,129,0,238,0,0,0,0,0,198,0,142,0,0,0,44,0,25,0,232,0,65,0,27,0,26,0,0,0,0,0,192,0,0,0,129,0,100,0,25,0,62,0,107,0,67,0,15,0,87,0,112,0,100,0,115,0,0,0,121,0,179,0,233,0,112,0,0,0,118,0,0,0,75,0,0,0,85,0,36,0,145,0,249,0,0,0,250,0,21,0,0,0,40,0,165,0,45,0,47,0,0,0,0,0,0,0,51,0,188,0,78,0,0,0,0,0,13,0,18,0,63,0,0,0,17,0,0,0,13,0,69,0,21,0,192,0,244,0,208,0,198,0,0,0,68,0,228,0,223,0,0,0,100,0,74,0,0,0,127,0,113,0,86,0,22,0,13,0,138,0,27,0,166,0,34,0,111,0,247,0,130,0,108,0,41,0,0,0,0,0,164,0,10,0,117,0,131,0,160,0,56,0,91,0,0,0,0,0,83,0,94,0,106,0,164,0,249,0,104,0,246,0,127,0,178,0,99,0,68,0,10,0,5,0,200,0,0,0,76,0,128,0,50,0,138,0,180,0,25,0,0,0,0,0,125,0,87,0,198,0,205,0,0,0,105,0,0,0,54,0,166,0,9,0,59,0,163,0,53,0,9,0,16,0,0,0,233,0,13,0,117,0,112,0,48,0,60,0,0,0,44,0,72,0,55,0,51,0,5,0,164,0,37,0,228,0,68,0,57,0,52,0,226,0,0,0,0,0,244,0,33,0,188,0,251,0,231,0,0,0,194,0,10,0,0,0,234,0,81,0,54,0,23,0,165,0,72,0,74,0,173,0,218,0,70,0,0,0,207,0,45,0,0,0,142,0,86,0,90,0,66,0,0,0,0,0,152,0,0,0,220,0,62,0,65,0,0,0,0,0,144,0,49,0,185,0,201,0,35,0,199,0,135,0,145,0,193,0,136,0,58,0,173,0,129,0,0,0,74,0,0,0,105,0,211,0,0,0,3,0,231,0,18,0,7,0,187,0,194,0,0,0,138,0,125,0,101,0,110,0,186,0,178,0,0,0,0,0,0,0,121,0,97,0,213,0,199,0,36,0,93,0,140,0,216,0,144,0,149,0,191,0,119,0,228,0,0,0,166,0,0,0,180,0,101,0,60,0,147,0,33,0,108,0,97,0,150,0,21,0,248,0,57,0,17,0,137,0,37,0,73,0,0,0,251,0,0,0,181,0,68,0,67,0,212,0,150,0,25,0,205,0,55,0,133,0,191,0,44,0,0,0,141,0,224,0,83,0,21,0,71,0,46,0,61,0,148,0,112,0,125,0,144,0,147,0,110,0,223,0,89,0,212,0,50,0,26,0,243,0,140,0,0,0,133,0,6,0,112,0,47,0,75,0,0,0,38,0,76,0,60,0,128,0,124,0,164,0,0,0,0,0,153,0,214,0,235,0,138,0,0,0,34,0,0,0,37,0,17,0,65,0,0,0,242,0,228,0,3,0,218,0,0,0,0,0,81,0,197,0,171,0,0,0,122,0,248,0,0,0,115,0,215,0,168,0,250,0,101,0,27,0,160,0,6,0,249,0,0,0,221,0,69,0,237,0,197,0,57,0,193,0,61,0,73,0,205,0,16,0,0,0,140,0,0,0,0,0,2,0,177,0,194,0,207,0,23,0,91,0,0,0,9,0,32,0,99,0,92,0,89,0,152,0,18,0,126,0,255,0,0,0,121,0,87,0,0,0,165,0,0,0,79,0,191,0,118,0,50,0,216,0,44,0,78,0,181,0,138,0,0,0,1,0,111,0,1,0,42,0,0,0,19,0,0,0,0,0,118,0,49,0,65,0,227,0,132,0,145,0,9,0,241,0,79,0,91,0,37,0,215,0,134,0,0,0,209,0,0,0,83,0,174,0,52,0,38,0,26,0,253,0,0,0,238,0,0,0,60,0,167,0,79,0,0,0,161,0,0,0,155,0,0,0,37,0,19,0,33,0,95,0,0,0,0,0,243,0,0,0,144,0,116,0,227,0,2,0,27,0,16,0,184,0,74,0,6,0,111,0,162,0,86,0,198,0,36,0,92,0,53,0,168,0,2,0,63,0,199,0,43,0,66,0,0,0,78,0,40,0,30,0,177,0,9,0,231,0,0,0,229,0,41,0,121,0,47,0,0,0,0,0,249,0,137,0,147,0,115,0,188,0,80,0,225,0,254,0,68,0,132,0,156,0,177,0,88,0,172,0,148,0,240,0,61,0,172,0,165,0,102,0,119,0,73,0,106,0,103,0,0,0,0,0,0,0,52,0,173,0,0,0,0,0,0,0,73,0,0,0,71,0,0,0,30,0,0,0,245,0,0,0,15,0,128,0,254,0,0,0,0,0,11,0,92,0,73,0,76,0,0,0,74,0,33,0,57,0,159,0,0,0,37,0,0,0,179,0,237,0,203,0,18,0,81,0,120,0,20,0,163,0,165,0,162,0,170,0,72,0,228,0,0,0,8,0,2,0,142,0,0,0,139,0,21,0,23,0,18,0,44,0,156,0,125,0,135,0,0,0,251,0,0,0,0,0,9,0,171,0,0,0,84,0,184,0,122,0,0,0,0,0,129,0,193,0,37,0,128,0,0,0,72,0,54,0,113,0,127,0,83,0,232,0,25,0,58,0,55,0,60,0,13,0,0,0,31,0,153,0,224,0,0,0,82,0,176,0,247,0,184,0,21,0,0,0,97,0,123,0,75,0,0,0,203,0,43,0,198,0,33,0,0,0,176,0,196,0,218,0,185,0,0,0,187,0,184,0,142,0,0,0,167,0,0,0,155,0,16,0,255,0,89,0,0,0,23,0,0,0,90,0,228,0,0,0,144,0,0,0,229,0,32,0,248,0,36,0,77,0,249,0,251,0,116,0,48,0,85,0,57,0,139,0,34,0,49,0,232,0,184,0,252,0,0,0,238,0,229,0,226,0,175,0,50,0,167,0,246,0,19,0,69,0,0,0,0,0,86,0,44,0,10,0,14,0,250,0,0,0,90,0,12,0,63,0,21,0,228,0,254,0,150,0,0,0,173,0,52,0,215,0,101,0,5,0,59,0,73,0,0,0,188,0,114,0,172,0,140,0,0,0,136,0,4,0,185,0,24,0,123,0,118,0,119,0,56,0,0,0,157,0,239,0,197,0,74,0,0,0,23,0,0,0,191,0,32,0,192,0,19,0,9,0,170,0,9,0,108,0,36,0,15,0,190,0,130,0,164,0,20,0,95,0,61,0,106,0,159,0,63,0,158,0,0,0,84,0,0,0,8,0,0,0,15,0,167,0,41,0,82,0,141,0,73,0,14,0,163,0,90,0,139,0,0,0,0,0,0,0,59,0,38,0,90,0,169,0,190,0,179,0,22,0,247,0,29,0,84,0,65,0,0,0,0,0,0,0,0,0,12,0,178,0,162,0,188,0,173,0,107,0,217,0,232,0,172,0,84,0,131,0,165,0);
signal scenario_full  : scenario_type := (53,31,53,30,179,31,156,31,156,30,246,31,36,31,149,31,113,31,113,30,209,31,70,31,186,31,7,31,5,31,55,31,55,30,55,29,55,28,119,31,110,31,248,31,105,31,195,31,114,31,21,31,179,31,179,30,187,31,187,30,120,31,159,31,159,30,66,31,210,31,215,31,229,31,102,31,94,31,185,31,138,31,85,31,187,31,45,31,225,31,184,31,149,31,93,31,156,31,99,31,99,30,62,31,62,30,44,31,241,31,127,31,127,30,132,31,112,31,56,31,56,30,144,31,37,31,25,31,106,31,22,31,148,31,191,31,188,31,194,31,170,31,252,31,95,31,95,30,166,31,18,31,136,31,201,31,143,31,179,31,183,31,228,31,10,31,242,31,242,30,138,31,152,31,200,31,15,31,15,30,15,29,220,31,55,31,123,31,96,31,90,31,90,30,90,29,154,31,20,31,174,31,232,31,178,31,49,31,222,31,25,31,25,30,38,31,5,31,234,31,234,30,234,31,236,31,236,30,72,31,83,31,230,31,37,31,188,31,93,31,93,30,240,31,240,30,239,31,161,31,161,30,75,31,189,31,166,31,16,31,59,31,113,31,207,31,192,31,144,31,144,30,53,31,53,30,189,31,129,31,238,31,238,30,238,29,198,31,142,31,142,30,44,31,25,31,232,31,65,31,27,31,26,31,26,30,26,29,192,31,192,30,129,31,100,31,25,31,62,31,107,31,67,31,15,31,87,31,112,31,100,31,115,31,115,30,121,31,179,31,233,31,112,31,112,30,118,31,118,30,75,31,75,30,85,31,36,31,145,31,249,31,249,30,250,31,21,31,21,30,40,31,165,31,45,31,47,31,47,30,47,29,47,28,51,31,188,31,78,31,78,30,78,29,13,31,18,31,63,31,63,30,17,31,17,30,13,31,69,31,21,31,192,31,244,31,208,31,198,31,198,30,68,31,228,31,223,31,223,30,100,31,74,31,74,30,127,31,113,31,86,31,22,31,13,31,138,31,27,31,166,31,34,31,111,31,247,31,130,31,108,31,41,31,41,30,41,29,164,31,10,31,117,31,131,31,160,31,56,31,91,31,91,30,91,29,83,31,94,31,106,31,164,31,249,31,104,31,246,31,127,31,178,31,99,31,68,31,10,31,5,31,200,31,200,30,76,31,128,31,50,31,138,31,180,31,25,31,25,30,25,29,125,31,87,31,198,31,205,31,205,30,105,31,105,30,54,31,166,31,9,31,59,31,163,31,53,31,9,31,16,31,16,30,233,31,13,31,117,31,112,31,48,31,60,31,60,30,44,31,72,31,55,31,51,31,5,31,164,31,37,31,228,31,68,31,57,31,52,31,226,31,226,30,226,29,244,31,33,31,188,31,251,31,231,31,231,30,194,31,10,31,10,30,234,31,81,31,54,31,23,31,165,31,72,31,74,31,173,31,218,31,70,31,70,30,207,31,45,31,45,30,142,31,86,31,90,31,66,31,66,30,66,29,152,31,152,30,220,31,62,31,65,31,65,30,65,29,144,31,49,31,185,31,201,31,35,31,199,31,135,31,145,31,193,31,136,31,58,31,173,31,129,31,129,30,74,31,74,30,105,31,211,31,211,30,3,31,231,31,18,31,7,31,187,31,194,31,194,30,138,31,125,31,101,31,110,31,186,31,178,31,178,30,178,29,178,28,121,31,97,31,213,31,199,31,36,31,93,31,140,31,216,31,144,31,149,31,191,31,119,31,228,31,228,30,166,31,166,30,180,31,101,31,60,31,147,31,33,31,108,31,97,31,150,31,21,31,248,31,57,31,17,31,137,31,37,31,73,31,73,30,251,31,251,30,181,31,68,31,67,31,212,31,150,31,25,31,205,31,55,31,133,31,191,31,44,31,44,30,141,31,224,31,83,31,21,31,71,31,46,31,61,31,148,31,112,31,125,31,144,31,147,31,110,31,223,31,89,31,212,31,50,31,26,31,243,31,140,31,140,30,133,31,6,31,112,31,47,31,75,31,75,30,38,31,76,31,60,31,128,31,124,31,164,31,164,30,164,29,153,31,214,31,235,31,138,31,138,30,34,31,34,30,37,31,17,31,65,31,65,30,242,31,228,31,3,31,218,31,218,30,218,29,81,31,197,31,171,31,171,30,122,31,248,31,248,30,115,31,215,31,168,31,250,31,101,31,27,31,160,31,6,31,249,31,249,30,221,31,69,31,237,31,197,31,57,31,193,31,61,31,73,31,205,31,16,31,16,30,140,31,140,30,140,29,2,31,177,31,194,31,207,31,23,31,91,31,91,30,9,31,32,31,99,31,92,31,89,31,152,31,18,31,126,31,255,31,255,30,121,31,87,31,87,30,165,31,165,30,79,31,191,31,118,31,50,31,216,31,44,31,78,31,181,31,138,31,138,30,1,31,111,31,1,31,42,31,42,30,19,31,19,30,19,29,118,31,49,31,65,31,227,31,132,31,145,31,9,31,241,31,79,31,91,31,37,31,215,31,134,31,134,30,209,31,209,30,83,31,174,31,52,31,38,31,26,31,253,31,253,30,238,31,238,30,60,31,167,31,79,31,79,30,161,31,161,30,155,31,155,30,37,31,19,31,33,31,95,31,95,30,95,29,243,31,243,30,144,31,116,31,227,31,2,31,27,31,16,31,184,31,74,31,6,31,111,31,162,31,86,31,198,31,36,31,92,31,53,31,168,31,2,31,63,31,199,31,43,31,66,31,66,30,78,31,40,31,30,31,177,31,9,31,231,31,231,30,229,31,41,31,121,31,47,31,47,30,47,29,249,31,137,31,147,31,115,31,188,31,80,31,225,31,254,31,68,31,132,31,156,31,177,31,88,31,172,31,148,31,240,31,61,31,172,31,165,31,102,31,119,31,73,31,106,31,103,31,103,30,103,29,103,28,52,31,173,31,173,30,173,29,173,28,73,31,73,30,71,31,71,30,30,31,30,30,245,31,245,30,15,31,128,31,254,31,254,30,254,29,11,31,92,31,73,31,76,31,76,30,74,31,33,31,57,31,159,31,159,30,37,31,37,30,179,31,237,31,203,31,18,31,81,31,120,31,20,31,163,31,165,31,162,31,170,31,72,31,228,31,228,30,8,31,2,31,142,31,142,30,139,31,21,31,23,31,18,31,44,31,156,31,125,31,135,31,135,30,251,31,251,30,251,29,9,31,171,31,171,30,84,31,184,31,122,31,122,30,122,29,129,31,193,31,37,31,128,31,128,30,72,31,54,31,113,31,127,31,83,31,232,31,25,31,58,31,55,31,60,31,13,31,13,30,31,31,153,31,224,31,224,30,82,31,176,31,247,31,184,31,21,31,21,30,97,31,123,31,75,31,75,30,203,31,43,31,198,31,33,31,33,30,176,31,196,31,218,31,185,31,185,30,187,31,184,31,142,31,142,30,167,31,167,30,155,31,16,31,255,31,89,31,89,30,23,31,23,30,90,31,228,31,228,30,144,31,144,30,229,31,32,31,248,31,36,31,77,31,249,31,251,31,116,31,48,31,85,31,57,31,139,31,34,31,49,31,232,31,184,31,252,31,252,30,238,31,229,31,226,31,175,31,50,31,167,31,246,31,19,31,69,31,69,30,69,29,86,31,44,31,10,31,14,31,250,31,250,30,90,31,12,31,63,31,21,31,228,31,254,31,150,31,150,30,173,31,52,31,215,31,101,31,5,31,59,31,73,31,73,30,188,31,114,31,172,31,140,31,140,30,136,31,4,31,185,31,24,31,123,31,118,31,119,31,56,31,56,30,157,31,239,31,197,31,74,31,74,30,23,31,23,30,191,31,32,31,192,31,19,31,9,31,170,31,9,31,108,31,36,31,15,31,190,31,130,31,164,31,20,31,95,31,61,31,106,31,159,31,63,31,158,31,158,30,84,31,84,30,8,31,8,30,15,31,167,31,41,31,82,31,141,31,73,31,14,31,163,31,90,31,139,31,139,30,139,29,139,28,59,31,38,31,90,31,169,31,190,31,179,31,22,31,247,31,29,31,84,31,65,31,65,30,65,29,65,28,65,27,12,31,178,31,162,31,188,31,173,31,107,31,217,31,232,31,172,31,84,31,131,31,165,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
