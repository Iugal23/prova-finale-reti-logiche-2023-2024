-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_909 is
end project_tb_909;

architecture project_tb_arch_909 of project_tb_909 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 802;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,151,0,0,0,242,0,180,0,0,0,107,0,169,0,68,0,36,0,226,0,193,0,39,0,207,0,11,0,0,0,198,0,89,0,0,0,0,0,177,0,43,0,21,0,14,0,90,0,29,0,208,0,241,0,93,0,230,0,70,0,229,0,212,0,77,0,42,0,216,0,0,0,13,0,175,0,3,0,73,0,121,0,0,0,0,0,226,0,141,0,0,0,169,0,226,0,30,0,18,0,44,0,66,0,78,0,77,0,106,0,152,0,43,0,33,0,236,0,0,0,9,0,242,0,119,0,233,0,75,0,223,0,191,0,68,0,191,0,197,0,35,0,30,0,175,0,28,0,0,0,116,0,148,0,0,0,0,0,92,0,245,0,0,0,66,0,121,0,45,0,0,0,82,0,63,0,77,0,201,0,200,0,0,0,201,0,217,0,81,0,0,0,207,0,212,0,0,0,121,0,67,0,156,0,0,0,172,0,135,0,21,0,6,0,245,0,39,0,187,0,72,0,0,0,105,0,223,0,148,0,252,0,118,0,44,0,0,0,117,0,55,0,17,0,174,0,190,0,0,0,93,0,0,0,92,0,0,0,125,0,0,0,0,0,152,0,130,0,153,0,57,0,0,0,0,0,63,0,231,0,0,0,0,0,174,0,63,0,202,0,44,0,169,0,0,0,235,0,137,0,80,0,210,0,183,0,126,0,53,0,3,0,191,0,176,0,240,0,207,0,30,0,173,0,190,0,129,0,127,0,118,0,0,0,28,0,211,0,245,0,0,0,61,0,15,0,141,0,232,0,168,0,57,0,18,0,214,0,222,0,247,0,162,0,170,0,41,0,9,0,0,0,24,0,68,0,92,0,198,0,0,0,227,0,0,0,179,0,0,0,169,0,0,0,0,0,76,0,174,0,0,0,193,0,174,0,0,0,248,0,0,0,60,0,82,0,147,0,181,0,123,0,19,0,108,0,236,0,114,0,1,0,28,0,0,0,127,0,5,0,72,0,233,0,177,0,37,0,0,0,121,0,28,0,101,0,0,0,117,0,198,0,185,0,158,0,0,0,179,0,0,0,123,0,165,0,64,0,196,0,118,0,181,0,60,0,115,0,188,0,108,0,196,0,245,0,177,0,249,0,141,0,0,0,94,0,228,0,228,0,120,0,50,0,232,0,6,0,140,0,96,0,65,0,181,0,137,0,76,0,26,0,0,0,72,0,33,0,213,0,109,0,0,0,44,0,102,0,100,0,146,0,0,0,162,0,33,0,253,0,11,0,248,0,0,0,130,0,0,0,0,0,130,0,0,0,0,0,16,0,229,0,251,0,22,0,0,0,232,0,87,0,0,0,2,0,192,0,252,0,216,0,0,0,79,0,0,0,89,0,140,0,241,0,108,0,103,0,79,0,91,0,19,0,26,0,147,0,124,0,161,0,0,0,210,0,167,0,213,0,2,0,37,0,12,0,82,0,96,0,0,0,252,0,255,0,166,0,103,0,175,0,122,0,198,0,111,0,24,0,69,0,224,0,0,0,0,0,188,0,0,0,155,0,142,0,0,0,128,0,16,0,107,0,108,0,69,0,238,0,154,0,31,0,247,0,91,0,117,0,244,0,23,0,226,0,127,0,218,0,140,0,13,0,170,0,72,0,14,0,139,0,244,0,30,0,153,0,30,0,0,0,52,0,48,0,0,0,124,0,0,0,43,0,199,0,54,0,170,0,95,0,224,0,51,0,0,0,69,0,81,0,181,0,0,0,222,0,218,0,169,0,225,0,180,0,140,0,0,0,0,0,84,0,32,0,29,0,0,0,109,0,17,0,88,0,152,0,0,0,110,0,171,0,10,0,102,0,165,0,44,0,47,0,46,0,26,0,1,0,194,0,104,0,235,0,11,0,0,0,202,0,115,0,94,0,49,0,185,0,165,0,0,0,125,0,6,0,192,0,0,0,180,0,178,0,223,0,204,0,156,0,44,0,119,0,0,0,91,0,0,0,45,0,2,0,225,0,182,0,194,0,247,0,187,0,77,0,102,0,3,0,250,0,72,0,240,0,0,0,102,0,12,0,109,0,121,0,201,0,239,0,85,0,210,0,4,0,207,0,169,0,22,0,251,0,177,0,248,0,240,0,0,0,0,0,0,0,127,0,217,0,103,0,129,0,71,0,148,0,8,0,0,0,48,0,59,0,138,0,0,0,135,0,19,0,0,0,187,0,23,0,169,0,39,0,0,0,64,0,255,0,198,0,20,0,125,0,225,0,29,0,137,0,18,0,254,0,251,0,200,0,58,0,42,0,16,0,114,0,0,0,200,0,232,0,226,0,177,0,58,0,0,0,16,0,190,0,89,0,16,0,0,0,242,0,3,0,150,0,114,0,0,0,82,0,168,0,0,0,0,0,192,0,0,0,89,0,242,0,0,0,70,0,249,0,0,0,0,0,126,0,76,0,29,0,90,0,64,0,0,0,0,0,26,0,55,0,0,0,141,0,34,0,0,0,0,0,89,0,137,0,186,0,133,0,43,0,0,0,69,0,22,0,34,0,228,0,27,0,56,0,189,0,123,0,111,0,116,0,141,0,82,0,161,0,228,0,17,0,59,0,0,0,54,0,0,0,223,0,196,0,0,0,152,0,69,0,79,0,0,0,214,0,10,0,79,0,239,0,121,0,57,0,36,0,102,0,0,0,200,0,230,0,35,0,0,0,72,0,240,0,121,0,94,0,161,0,2,0,196,0,79,0,133,0,50,0,172,0,62,0,2,0,117,0,123,0,86,0,21,0,194,0,57,0,254,0,80,0,126,0,244,0,80,0,0,0,0,0,59,0,45,0,128,0,173,0,34,0,204,0,59,0,254,0,140,0,72,0,54,0,46,0,142,0,184,0,205,0,229,0,0,0,87,0,4,0,203,0,26,0,192,0,246,0,177,0,164,0,179,0,110,0,70,0,196,0,207,0,186,0,172,0,49,0,42,0,77,0,26,0,110,0,8,0,123,0,36,0,15,0,137,0,117,0,118,0,251,0,168,0,59,0,95,0,187,0,85,0,95,0,187,0,0,0,0,0,74,0,0,0,98,0,0,0,104,0,121,0,127,0,74,0,0,0,227,0,157,0,236,0,0,0,42,0,116,0,0,0,47,0,135,0,0,0,223,0,246,0,202,0,189,0,0,0,220,0,0,0,0,0,101,0,79,0,191,0,87,0,0,0,0,0,0,0,252,0,11,0,101,0,67,0,151,0,136,0,0,0,117,0,175,0,133,0,19,0,13,0,38,0,27,0,0,0,0,0,0,0,0,0,18,0,0,0,34,0,223,0,36,0,57,0,132,0,0,0,129,0,194,0,0,0,0,0,108,0,215,0,136,0,238,0,225,0,168,0,126,0,191,0,86,0,0,0,51,0,0,0,129,0,170,0,152,0,0,0,51,0,68,0,128,0,0,0,0,0,216,0,177,0,67,0,253,0,0,0,56,0,237,0,46,0,187,0,240,0,243,0,31,0,28,0,223,0,175,0,179,0,5,0,143,0,219,0,58,0,201,0,28,0,120,0,106,0,210,0,133,0,142,0,193,0,62,0,109,0,206,0,200,0,178,0,0,0,31,0,218,0,25,0);
signal scenario_full  : scenario_type := (214,31,151,31,151,30,242,31,180,31,180,30,107,31,169,31,68,31,36,31,226,31,193,31,39,31,207,31,11,31,11,30,198,31,89,31,89,30,89,29,177,31,43,31,21,31,14,31,90,31,29,31,208,31,241,31,93,31,230,31,70,31,229,31,212,31,77,31,42,31,216,31,216,30,13,31,175,31,3,31,73,31,121,31,121,30,121,29,226,31,141,31,141,30,169,31,226,31,30,31,18,31,44,31,66,31,78,31,77,31,106,31,152,31,43,31,33,31,236,31,236,30,9,31,242,31,119,31,233,31,75,31,223,31,191,31,68,31,191,31,197,31,35,31,30,31,175,31,28,31,28,30,116,31,148,31,148,30,148,29,92,31,245,31,245,30,66,31,121,31,45,31,45,30,82,31,63,31,77,31,201,31,200,31,200,30,201,31,217,31,81,31,81,30,207,31,212,31,212,30,121,31,67,31,156,31,156,30,172,31,135,31,21,31,6,31,245,31,39,31,187,31,72,31,72,30,105,31,223,31,148,31,252,31,118,31,44,31,44,30,117,31,55,31,17,31,174,31,190,31,190,30,93,31,93,30,92,31,92,30,125,31,125,30,125,29,152,31,130,31,153,31,57,31,57,30,57,29,63,31,231,31,231,30,231,29,174,31,63,31,202,31,44,31,169,31,169,30,235,31,137,31,80,31,210,31,183,31,126,31,53,31,3,31,191,31,176,31,240,31,207,31,30,31,173,31,190,31,129,31,127,31,118,31,118,30,28,31,211,31,245,31,245,30,61,31,15,31,141,31,232,31,168,31,57,31,18,31,214,31,222,31,247,31,162,31,170,31,41,31,9,31,9,30,24,31,68,31,92,31,198,31,198,30,227,31,227,30,179,31,179,30,169,31,169,30,169,29,76,31,174,31,174,30,193,31,174,31,174,30,248,31,248,30,60,31,82,31,147,31,181,31,123,31,19,31,108,31,236,31,114,31,1,31,28,31,28,30,127,31,5,31,72,31,233,31,177,31,37,31,37,30,121,31,28,31,101,31,101,30,117,31,198,31,185,31,158,31,158,30,179,31,179,30,123,31,165,31,64,31,196,31,118,31,181,31,60,31,115,31,188,31,108,31,196,31,245,31,177,31,249,31,141,31,141,30,94,31,228,31,228,31,120,31,50,31,232,31,6,31,140,31,96,31,65,31,181,31,137,31,76,31,26,31,26,30,72,31,33,31,213,31,109,31,109,30,44,31,102,31,100,31,146,31,146,30,162,31,33,31,253,31,11,31,248,31,248,30,130,31,130,30,130,29,130,31,130,30,130,29,16,31,229,31,251,31,22,31,22,30,232,31,87,31,87,30,2,31,192,31,252,31,216,31,216,30,79,31,79,30,89,31,140,31,241,31,108,31,103,31,79,31,91,31,19,31,26,31,147,31,124,31,161,31,161,30,210,31,167,31,213,31,2,31,37,31,12,31,82,31,96,31,96,30,252,31,255,31,166,31,103,31,175,31,122,31,198,31,111,31,24,31,69,31,224,31,224,30,224,29,188,31,188,30,155,31,142,31,142,30,128,31,16,31,107,31,108,31,69,31,238,31,154,31,31,31,247,31,91,31,117,31,244,31,23,31,226,31,127,31,218,31,140,31,13,31,170,31,72,31,14,31,139,31,244,31,30,31,153,31,30,31,30,30,52,31,48,31,48,30,124,31,124,30,43,31,199,31,54,31,170,31,95,31,224,31,51,31,51,30,69,31,81,31,181,31,181,30,222,31,218,31,169,31,225,31,180,31,140,31,140,30,140,29,84,31,32,31,29,31,29,30,109,31,17,31,88,31,152,31,152,30,110,31,171,31,10,31,102,31,165,31,44,31,47,31,46,31,26,31,1,31,194,31,104,31,235,31,11,31,11,30,202,31,115,31,94,31,49,31,185,31,165,31,165,30,125,31,6,31,192,31,192,30,180,31,178,31,223,31,204,31,156,31,44,31,119,31,119,30,91,31,91,30,45,31,2,31,225,31,182,31,194,31,247,31,187,31,77,31,102,31,3,31,250,31,72,31,240,31,240,30,102,31,12,31,109,31,121,31,201,31,239,31,85,31,210,31,4,31,207,31,169,31,22,31,251,31,177,31,248,31,240,31,240,30,240,29,240,28,127,31,217,31,103,31,129,31,71,31,148,31,8,31,8,30,48,31,59,31,138,31,138,30,135,31,19,31,19,30,187,31,23,31,169,31,39,31,39,30,64,31,255,31,198,31,20,31,125,31,225,31,29,31,137,31,18,31,254,31,251,31,200,31,58,31,42,31,16,31,114,31,114,30,200,31,232,31,226,31,177,31,58,31,58,30,16,31,190,31,89,31,16,31,16,30,242,31,3,31,150,31,114,31,114,30,82,31,168,31,168,30,168,29,192,31,192,30,89,31,242,31,242,30,70,31,249,31,249,30,249,29,126,31,76,31,29,31,90,31,64,31,64,30,64,29,26,31,55,31,55,30,141,31,34,31,34,30,34,29,89,31,137,31,186,31,133,31,43,31,43,30,69,31,22,31,34,31,228,31,27,31,56,31,189,31,123,31,111,31,116,31,141,31,82,31,161,31,228,31,17,31,59,31,59,30,54,31,54,30,223,31,196,31,196,30,152,31,69,31,79,31,79,30,214,31,10,31,79,31,239,31,121,31,57,31,36,31,102,31,102,30,200,31,230,31,35,31,35,30,72,31,240,31,121,31,94,31,161,31,2,31,196,31,79,31,133,31,50,31,172,31,62,31,2,31,117,31,123,31,86,31,21,31,194,31,57,31,254,31,80,31,126,31,244,31,80,31,80,30,80,29,59,31,45,31,128,31,173,31,34,31,204,31,59,31,254,31,140,31,72,31,54,31,46,31,142,31,184,31,205,31,229,31,229,30,87,31,4,31,203,31,26,31,192,31,246,31,177,31,164,31,179,31,110,31,70,31,196,31,207,31,186,31,172,31,49,31,42,31,77,31,26,31,110,31,8,31,123,31,36,31,15,31,137,31,117,31,118,31,251,31,168,31,59,31,95,31,187,31,85,31,95,31,187,31,187,30,187,29,74,31,74,30,98,31,98,30,104,31,121,31,127,31,74,31,74,30,227,31,157,31,236,31,236,30,42,31,116,31,116,30,47,31,135,31,135,30,223,31,246,31,202,31,189,31,189,30,220,31,220,30,220,29,101,31,79,31,191,31,87,31,87,30,87,29,87,28,252,31,11,31,101,31,67,31,151,31,136,31,136,30,117,31,175,31,133,31,19,31,13,31,38,31,27,31,27,30,27,29,27,28,27,27,18,31,18,30,34,31,223,31,36,31,57,31,132,31,132,30,129,31,194,31,194,30,194,29,108,31,215,31,136,31,238,31,225,31,168,31,126,31,191,31,86,31,86,30,51,31,51,30,129,31,170,31,152,31,152,30,51,31,68,31,128,31,128,30,128,29,216,31,177,31,67,31,253,31,253,30,56,31,237,31,46,31,187,31,240,31,243,31,31,31,28,31,223,31,175,31,179,31,5,31,143,31,219,31,58,31,201,31,28,31,120,31,106,31,210,31,133,31,142,31,193,31,62,31,109,31,206,31,200,31,178,31,178,30,31,31,218,31,25,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
