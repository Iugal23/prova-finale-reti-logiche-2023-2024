-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_660 is
end project_tb_660;

architecture project_tb_arch_660 of project_tb_660 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 568;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (150,0,48,0,202,0,168,0,117,0,0,0,119,0,0,0,84,0,177,0,79,0,255,0,0,0,131,0,117,0,88,0,91,0,122,0,118,0,44,0,103,0,33,0,176,0,170,0,157,0,163,0,116,0,105,0,162,0,110,0,29,0,139,0,175,0,84,0,59,0,4,0,161,0,183,0,205,0,251,0,55,0,201,0,166,0,148,0,0,0,5,0,113,0,67,0,130,0,142,0,235,0,99,0,235,0,194,0,199,0,125,0,230,0,226,0,0,0,119,0,136,0,173,0,191,0,32,0,0,0,0,0,0,0,0,0,67,0,0,0,33,0,0,0,50,0,81,0,158,0,25,0,52,0,28,0,130,0,99,0,103,0,226,0,119,0,0,0,216,0,10,0,0,0,62,0,64,0,0,0,158,0,0,0,161,0,61,0,246,0,15,0,148,0,0,0,99,0,4,0,54,0,154,0,0,0,0,0,252,0,0,0,78,0,0,0,116,0,65,0,135,0,199,0,252,0,0,0,225,0,0,0,136,0,234,0,85,0,165,0,181,0,72,0,69,0,118,0,132,0,0,0,96,0,0,0,201,0,0,0,34,0,27,0,83,0,203,0,0,0,235,0,71,0,228,0,37,0,0,0,38,0,241,0,38,0,19,0,246,0,32,0,5,0,0,0,128,0,0,0,36,0,0,0,97,0,1,0,210,0,0,0,0,0,137,0,14,0,35,0,129,0,152,0,125,0,0,0,239,0,0,0,104,0,133,0,0,0,1,0,185,0,50,0,55,0,44,0,61,0,0,0,220,0,30,0,0,0,50,0,82,0,0,0,164,0,117,0,152,0,212,0,203,0,0,0,0,0,249,0,78,0,11,0,17,0,139,0,107,0,128,0,0,0,248,0,134,0,111,0,0,0,120,0,226,0,0,0,206,0,95,0,176,0,0,0,202,0,0,0,0,0,243,0,141,0,185,0,0,0,216,0,195,0,159,0,187,0,106,0,146,0,13,0,49,0,128,0,251,0,0,0,153,0,60,0,108,0,62,0,252,0,11,0,159,0,81,0,0,0,252,0,82,0,182,0,130,0,112,0,214,0,45,0,55,0,239,0,197,0,239,0,1,0,109,0,233,0,141,0,100,0,194,0,99,0,11,0,0,0,248,0,0,0,173,0,28,0,214,0,0,0,100,0,33,0,255,0,171,0,184,0,203,0,229,0,177,0,156,0,211,0,190,0,88,0,60,0,139,0,19,0,249,0,169,0,0,0,84,0,232,0,54,0,177,0,4,0,0,0,44,0,61,0,0,0,47,0,0,0,38,0,18,0,0,0,123,0,0,0,109,0,34,0,163,0,50,0,0,0,0,0,159,0,108,0,140,0,37,0,123,0,42,0,245,0,209,0,162,0,219,0,70,0,216,0,0,0,35,0,0,0,249,0,0,0,142,0,11,0,236,0,9,0,175,0,51,0,228,0,223,0,72,0,71,0,0,0,0,0,51,0,0,0,247,0,155,0,0,0,172,0,90,0,124,0,242,0,0,0,226,0,0,0,0,0,53,0,106,0,144,0,0,0,118,0,186,0,0,0,195,0,87,0,139,0,136,0,0,0,41,0,110,0,0,0,219,0,188,0,160,0,239,0,102,0,66,0,0,0,14,0,237,0,163,0,6,0,170,0,25,0,162,0,0,0,5,0,200,0,154,0,0,0,102,0,212,0,121,0,0,0,0,0,0,0,77,0,168,0,113,0,8,0,188,0,128,0,115,0,12,0,174,0,94,0,184,0,48,0,63,0,0,0,109,0,8,0,10,0,210,0,0,0,219,0,65,0,0,0,7,0,204,0,0,0,36,0,205,0,228,0,163,0,117,0,138,0,0,0,0,0,16,0,18,0,85,0,218,0,47,0,0,0,139,0,230,0,246,0,208,0,95,0,157,0,242,0,229,0,28,0,0,0,137,0,17,0,226,0,0,0,153,0,74,0,0,0,198,0,0,0,122,0,237,0,208,0,41,0,148,0,176,0,0,0,2,0,176,0,171,0,239,0,112,0,107,0,45,0,212,0,249,0,223,0,41,0,172,0,0,0,49,0,124,0,63,0,18,0,113,0,0,0,0,0,58,0,30,0,245,0,237,0,228,0,0,0,6,0,155,0,190,0,68,0,91,0,173,0,133,0,0,0,94,0,135,0,0,0,0,0,0,0,178,0,27,0,37,0,20,0,128,0,200,0,230,0,0,0,231,0,25,0,0,0,79,0,206,0,38,0,197,0,41,0,140,0,127,0,207,0,32,0,75,0,9,0,70,0,0,0,219,0,0,0,8,0,201,0,207,0,90,0,72,0,207,0,33,0,12,0,22,0,169,0,71,0,0,0,0,0,11,0,0,0,136,0,240,0,52,0,48,0,225,0,27,0,186,0,213,0,134,0,0,0,0,0,44,0,0,0,180,0,58,0,0,0,187,0,243,0,186,0,217,0,16,0,0,0,0,0,192,0,114,0,99,0,75,0,0,0,88,0,53,0,170,0,86,0,0,0,0,0,157,0,229,0,0,0,159,0,0,0,0,0);
signal scenario_full  : scenario_type := (150,31,48,31,202,31,168,31,117,31,117,30,119,31,119,30,84,31,177,31,79,31,255,31,255,30,131,31,117,31,88,31,91,31,122,31,118,31,44,31,103,31,33,31,176,31,170,31,157,31,163,31,116,31,105,31,162,31,110,31,29,31,139,31,175,31,84,31,59,31,4,31,161,31,183,31,205,31,251,31,55,31,201,31,166,31,148,31,148,30,5,31,113,31,67,31,130,31,142,31,235,31,99,31,235,31,194,31,199,31,125,31,230,31,226,31,226,30,119,31,136,31,173,31,191,31,32,31,32,30,32,29,32,28,32,27,67,31,67,30,33,31,33,30,50,31,81,31,158,31,25,31,52,31,28,31,130,31,99,31,103,31,226,31,119,31,119,30,216,31,10,31,10,30,62,31,64,31,64,30,158,31,158,30,161,31,61,31,246,31,15,31,148,31,148,30,99,31,4,31,54,31,154,31,154,30,154,29,252,31,252,30,78,31,78,30,116,31,65,31,135,31,199,31,252,31,252,30,225,31,225,30,136,31,234,31,85,31,165,31,181,31,72,31,69,31,118,31,132,31,132,30,96,31,96,30,201,31,201,30,34,31,27,31,83,31,203,31,203,30,235,31,71,31,228,31,37,31,37,30,38,31,241,31,38,31,19,31,246,31,32,31,5,31,5,30,128,31,128,30,36,31,36,30,97,31,1,31,210,31,210,30,210,29,137,31,14,31,35,31,129,31,152,31,125,31,125,30,239,31,239,30,104,31,133,31,133,30,1,31,185,31,50,31,55,31,44,31,61,31,61,30,220,31,30,31,30,30,50,31,82,31,82,30,164,31,117,31,152,31,212,31,203,31,203,30,203,29,249,31,78,31,11,31,17,31,139,31,107,31,128,31,128,30,248,31,134,31,111,31,111,30,120,31,226,31,226,30,206,31,95,31,176,31,176,30,202,31,202,30,202,29,243,31,141,31,185,31,185,30,216,31,195,31,159,31,187,31,106,31,146,31,13,31,49,31,128,31,251,31,251,30,153,31,60,31,108,31,62,31,252,31,11,31,159,31,81,31,81,30,252,31,82,31,182,31,130,31,112,31,214,31,45,31,55,31,239,31,197,31,239,31,1,31,109,31,233,31,141,31,100,31,194,31,99,31,11,31,11,30,248,31,248,30,173,31,28,31,214,31,214,30,100,31,33,31,255,31,171,31,184,31,203,31,229,31,177,31,156,31,211,31,190,31,88,31,60,31,139,31,19,31,249,31,169,31,169,30,84,31,232,31,54,31,177,31,4,31,4,30,44,31,61,31,61,30,47,31,47,30,38,31,18,31,18,30,123,31,123,30,109,31,34,31,163,31,50,31,50,30,50,29,159,31,108,31,140,31,37,31,123,31,42,31,245,31,209,31,162,31,219,31,70,31,216,31,216,30,35,31,35,30,249,31,249,30,142,31,11,31,236,31,9,31,175,31,51,31,228,31,223,31,72,31,71,31,71,30,71,29,51,31,51,30,247,31,155,31,155,30,172,31,90,31,124,31,242,31,242,30,226,31,226,30,226,29,53,31,106,31,144,31,144,30,118,31,186,31,186,30,195,31,87,31,139,31,136,31,136,30,41,31,110,31,110,30,219,31,188,31,160,31,239,31,102,31,66,31,66,30,14,31,237,31,163,31,6,31,170,31,25,31,162,31,162,30,5,31,200,31,154,31,154,30,102,31,212,31,121,31,121,30,121,29,121,28,77,31,168,31,113,31,8,31,188,31,128,31,115,31,12,31,174,31,94,31,184,31,48,31,63,31,63,30,109,31,8,31,10,31,210,31,210,30,219,31,65,31,65,30,7,31,204,31,204,30,36,31,205,31,228,31,163,31,117,31,138,31,138,30,138,29,16,31,18,31,85,31,218,31,47,31,47,30,139,31,230,31,246,31,208,31,95,31,157,31,242,31,229,31,28,31,28,30,137,31,17,31,226,31,226,30,153,31,74,31,74,30,198,31,198,30,122,31,237,31,208,31,41,31,148,31,176,31,176,30,2,31,176,31,171,31,239,31,112,31,107,31,45,31,212,31,249,31,223,31,41,31,172,31,172,30,49,31,124,31,63,31,18,31,113,31,113,30,113,29,58,31,30,31,245,31,237,31,228,31,228,30,6,31,155,31,190,31,68,31,91,31,173,31,133,31,133,30,94,31,135,31,135,30,135,29,135,28,178,31,27,31,37,31,20,31,128,31,200,31,230,31,230,30,231,31,25,31,25,30,79,31,206,31,38,31,197,31,41,31,140,31,127,31,207,31,32,31,75,31,9,31,70,31,70,30,219,31,219,30,8,31,201,31,207,31,90,31,72,31,207,31,33,31,12,31,22,31,169,31,71,31,71,30,71,29,11,31,11,30,136,31,240,31,52,31,48,31,225,31,27,31,186,31,213,31,134,31,134,30,134,29,44,31,44,30,180,31,58,31,58,30,187,31,243,31,186,31,217,31,16,31,16,30,16,29,192,31,114,31,99,31,75,31,75,30,88,31,53,31,170,31,86,31,86,30,86,29,157,31,229,31,229,30,159,31,159,30,159,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
