-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_363 is
end project_tb_363;

architecture project_tb_arch_363 of project_tb_363 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 489;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,102,0,174,0,142,0,15,0,239,0,196,0,11,0,177,0,132,0,0,0,187,0,0,0,35,0,156,0,125,0,204,0,147,0,93,0,186,0,0,0,54,0,216,0,0,0,0,0,83,0,27,0,54,0,87,0,168,0,34,0,0,0,4,0,0,0,0,0,246,0,0,0,186,0,0,0,127,0,180,0,84,0,100,0,72,0,55,0,237,0,145,0,0,0,206,0,199,0,106,0,178,0,215,0,29,0,86,0,143,0,120,0,202,0,185,0,54,0,0,0,44,0,14,0,225,0,148,0,9,0,238,0,146,0,35,0,31,0,67,0,130,0,0,0,80,0,251,0,159,0,224,0,223,0,0,0,0,0,51,0,156,0,111,0,78,0,69,0,79,0,141,0,88,0,104,0,82,0,0,0,0,0,142,0,41,0,0,0,220,0,76,0,191,0,255,0,225,0,149,0,0,0,220,0,28,0,11,0,34,0,181,0,0,0,23,0,0,0,197,0,158,0,14,0,182,0,16,0,0,0,109,0,78,0,186,0,0,0,124,0,91,0,82,0,26,0,161,0,249,0,118,0,123,0,27,0,60,0,220,0,8,0,190,0,0,0,165,0,246,0,209,0,0,0,118,0,0,0,189,0,50,0,142,0,75,0,0,0,0,0,205,0,155,0,214,0,153,0,177,0,165,0,209,0,67,0,0,0,172,0,0,0,72,0,151,0,0,0,31,0,95,0,126,0,68,0,171,0,144,0,237,0,110,0,242,0,252,0,136,0,255,0,48,0,244,0,180,0,163,0,107,0,225,0,169,0,0,0,66,0,168,0,224,0,32,0,17,0,216,0,80,0,77,0,229,0,115,0,161,0,24,0,174,0,44,0,145,0,0,0,24,0,223,0,20,0,64,0,0,0,138,0,0,0,66,0,62,0,5,0,91,0,186,0,69,0,0,0,253,0,236,0,16,0,183,0,138,0,142,0,0,0,0,0,156,0,210,0,8,0,200,0,109,0,156,0,0,0,25,0,14,0,129,0,175,0,150,0,57,0,122,0,38,0,60,0,56,0,97,0,79,0,0,0,0,0,147,0,0,0,0,0,85,0,10,0,0,0,104,0,0,0,48,0,43,0,102,0,81,0,204,0,58,0,161,0,0,0,0,0,0,0,25,0,135,0,131,0,198,0,0,0,19,0,0,0,97,0,149,0,1,0,55,0,14,0,160,0,217,0,148,0,90,0,141,0,82,0,0,0,236,0,0,0,0,0,0,0,196,0,43,0,0,0,232,0,0,0,0,0,4,0,16,0,48,0,222,0,0,0,76,0,6,0,181,0,173,0,243,0,32,0,158,0,0,0,123,0,152,0,250,0,0,0,200,0,0,0,248,0,236,0,105,0,118,0,0,0,0,0,175,0,161,0,0,0,20,0,0,0,123,0,189,0,0,0,28,0,77,0,0,0,0,0,114,0,161,0,25,0,121,0,79,0,217,0,210,0,164,0,246,0,113,0,83,0,127,0,93,0,109,0,19,0,0,0,211,0,2,0,0,0,0,0,192,0,0,0,126,0,161,0,203,0,123,0,0,0,74,0,221,0,167,0,140,0,54,0,50,0,46,0,209,0,192,0,69,0,17,0,122,0,106,0,164,0,0,0,86,0,83,0,73,0,232,0,0,0,88,0,245,0,157,0,41,0,0,0,240,0,0,0,191,0,214,0,97,0,0,0,0,0,152,0,115,0,77,0,154,0,0,0,185,0,143,0,44,0,156,0,0,0,103,0,141,0,27,0,48,0,197,0,65,0,135,0,240,0,29,0,58,0,18,0,0,0,178,0,0,0,0,0,24,0,0,0,100,0,96,0,57,0,114,0,28,0,52,0,168,0,15,0,78,0,198,0,0,0,51,0,97,0,163,0,177,0,72,0,152,0,8,0,231,0,0,0,126,0,0,0,132,0,194,0,128,0,246,0,239,0,122,0,1,0,0,0,233,0,82,0,226,0,0,0,49,0,0,0,0,0,122,0,225,0,12,0,133,0,194,0,59,0,95,0,204,0,88,0,192,0,138,0,108,0,190,0,197,0,119,0,0,0,72,0,112,0,35,0,21,0,46,0,0,0,0,0,33,0,155,0,110,0,176,0,32,0,205,0,7,0,112,0,0,0,0,0,12,0,105,0,108,0,133,0,117,0,124,0,250,0,29,0,183,0,0,0);
signal scenario_full  : scenario_type := (16,31,102,31,174,31,142,31,15,31,239,31,196,31,11,31,177,31,132,31,132,30,187,31,187,30,35,31,156,31,125,31,204,31,147,31,93,31,186,31,186,30,54,31,216,31,216,30,216,29,83,31,27,31,54,31,87,31,168,31,34,31,34,30,4,31,4,30,4,29,246,31,246,30,186,31,186,30,127,31,180,31,84,31,100,31,72,31,55,31,237,31,145,31,145,30,206,31,199,31,106,31,178,31,215,31,29,31,86,31,143,31,120,31,202,31,185,31,54,31,54,30,44,31,14,31,225,31,148,31,9,31,238,31,146,31,35,31,31,31,67,31,130,31,130,30,80,31,251,31,159,31,224,31,223,31,223,30,223,29,51,31,156,31,111,31,78,31,69,31,79,31,141,31,88,31,104,31,82,31,82,30,82,29,142,31,41,31,41,30,220,31,76,31,191,31,255,31,225,31,149,31,149,30,220,31,28,31,11,31,34,31,181,31,181,30,23,31,23,30,197,31,158,31,14,31,182,31,16,31,16,30,109,31,78,31,186,31,186,30,124,31,91,31,82,31,26,31,161,31,249,31,118,31,123,31,27,31,60,31,220,31,8,31,190,31,190,30,165,31,246,31,209,31,209,30,118,31,118,30,189,31,50,31,142,31,75,31,75,30,75,29,205,31,155,31,214,31,153,31,177,31,165,31,209,31,67,31,67,30,172,31,172,30,72,31,151,31,151,30,31,31,95,31,126,31,68,31,171,31,144,31,237,31,110,31,242,31,252,31,136,31,255,31,48,31,244,31,180,31,163,31,107,31,225,31,169,31,169,30,66,31,168,31,224,31,32,31,17,31,216,31,80,31,77,31,229,31,115,31,161,31,24,31,174,31,44,31,145,31,145,30,24,31,223,31,20,31,64,31,64,30,138,31,138,30,66,31,62,31,5,31,91,31,186,31,69,31,69,30,253,31,236,31,16,31,183,31,138,31,142,31,142,30,142,29,156,31,210,31,8,31,200,31,109,31,156,31,156,30,25,31,14,31,129,31,175,31,150,31,57,31,122,31,38,31,60,31,56,31,97,31,79,31,79,30,79,29,147,31,147,30,147,29,85,31,10,31,10,30,104,31,104,30,48,31,43,31,102,31,81,31,204,31,58,31,161,31,161,30,161,29,161,28,25,31,135,31,131,31,198,31,198,30,19,31,19,30,97,31,149,31,1,31,55,31,14,31,160,31,217,31,148,31,90,31,141,31,82,31,82,30,236,31,236,30,236,29,236,28,196,31,43,31,43,30,232,31,232,30,232,29,4,31,16,31,48,31,222,31,222,30,76,31,6,31,181,31,173,31,243,31,32,31,158,31,158,30,123,31,152,31,250,31,250,30,200,31,200,30,248,31,236,31,105,31,118,31,118,30,118,29,175,31,161,31,161,30,20,31,20,30,123,31,189,31,189,30,28,31,77,31,77,30,77,29,114,31,161,31,25,31,121,31,79,31,217,31,210,31,164,31,246,31,113,31,83,31,127,31,93,31,109,31,19,31,19,30,211,31,2,31,2,30,2,29,192,31,192,30,126,31,161,31,203,31,123,31,123,30,74,31,221,31,167,31,140,31,54,31,50,31,46,31,209,31,192,31,69,31,17,31,122,31,106,31,164,31,164,30,86,31,83,31,73,31,232,31,232,30,88,31,245,31,157,31,41,31,41,30,240,31,240,30,191,31,214,31,97,31,97,30,97,29,152,31,115,31,77,31,154,31,154,30,185,31,143,31,44,31,156,31,156,30,103,31,141,31,27,31,48,31,197,31,65,31,135,31,240,31,29,31,58,31,18,31,18,30,178,31,178,30,178,29,24,31,24,30,100,31,96,31,57,31,114,31,28,31,52,31,168,31,15,31,78,31,198,31,198,30,51,31,97,31,163,31,177,31,72,31,152,31,8,31,231,31,231,30,126,31,126,30,132,31,194,31,128,31,246,31,239,31,122,31,1,31,1,30,233,31,82,31,226,31,226,30,49,31,49,30,49,29,122,31,225,31,12,31,133,31,194,31,59,31,95,31,204,31,88,31,192,31,138,31,108,31,190,31,197,31,119,31,119,30,72,31,112,31,35,31,21,31,46,31,46,30,46,29,33,31,155,31,110,31,176,31,32,31,205,31,7,31,112,31,112,30,112,29,12,31,105,31,108,31,133,31,117,31,124,31,250,31,29,31,183,31,183,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
