-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 212;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,109,0,131,0,0,0,147,0,125,0,43,0,0,0,231,0,130,0,72,0,120,0,0,0,179,0,75,0,118,0,119,0,96,0,23,0,0,0,227,0,37,0,177,0,181,0,251,0,118,0,81,0,53,0,86,0,0,0,147,0,0,0,0,0,0,0,151,0,62,0,194,0,39,0,50,0,132,0,124,0,167,0,50,0,148,0,185,0,121,0,0,0,252,0,0,0,101,0,146,0,73,0,115,0,89,0,81,0,146,0,193,0,179,0,218,0,216,0,112,0,174,0,243,0,0,0,32,0,141,0,179,0,107,0,245,0,0,0,0,0,0,0,149,0,206,0,205,0,75,0,225,0,133,0,30,0,67,0,35,0,0,0,29,0,228,0,143,0,18,0,119,0,130,0,137,0,170,0,140,0,162,0,161,0,86,0,210,0,235,0,0,0,180,0,0,0,170,0,223,0,68,0,44,0,162,0,162,0,106,0,0,0,0,0,5,0,195,0,114,0,0,0,125,0,43,0,214,0,112,0,51,0,24,0,241,0,222,0,79,0,0,0,126,0,200,0,0,0,0,0,25,0,186,0,229,0,82,0,0,0,101,0,56,0,101,0,175,0,0,0,28,0,106,0,0,0,151,0,130,0,0,0,236,0,194,0,28,0,183,0,145,0,51,0,191,0,15,0,98,0,0,0,0,0,0,0,79,0,61,0,164,0,90,0,93,0,0,0,80,0,250,0,139,0,0,0,0,0,111,0,8,0,244,0,60,0,90,0,0,0,169,0,0,0,181,0,206,0,96,0,172,0,0,0,201,0,18,0,238,0,153,0,0,0,2,0,149,0,0,0,13,0,41,0,137,0,49,0,0,0,88,0,0,0,0,0,135,0,0,0,98,0,109,0,45,0,131,0,119,0,102,0,180,0,0,0,232,0,0,0,0,0,121,0,0,0,94,0,106,0,69,0);
signal scenario_full  : scenario_type := (128,31,109,31,131,31,131,30,147,31,125,31,43,31,43,30,231,31,130,31,72,31,120,31,120,30,179,31,75,31,118,31,119,31,96,31,23,31,23,30,227,31,37,31,177,31,181,31,251,31,118,31,81,31,53,31,86,31,86,30,147,31,147,30,147,29,147,28,151,31,62,31,194,31,39,31,50,31,132,31,124,31,167,31,50,31,148,31,185,31,121,31,121,30,252,31,252,30,101,31,146,31,73,31,115,31,89,31,81,31,146,31,193,31,179,31,218,31,216,31,112,31,174,31,243,31,243,30,32,31,141,31,179,31,107,31,245,31,245,30,245,29,245,28,149,31,206,31,205,31,75,31,225,31,133,31,30,31,67,31,35,31,35,30,29,31,228,31,143,31,18,31,119,31,130,31,137,31,170,31,140,31,162,31,161,31,86,31,210,31,235,31,235,30,180,31,180,30,170,31,223,31,68,31,44,31,162,31,162,31,106,31,106,30,106,29,5,31,195,31,114,31,114,30,125,31,43,31,214,31,112,31,51,31,24,31,241,31,222,31,79,31,79,30,126,31,200,31,200,30,200,29,25,31,186,31,229,31,82,31,82,30,101,31,56,31,101,31,175,31,175,30,28,31,106,31,106,30,151,31,130,31,130,30,236,31,194,31,28,31,183,31,145,31,51,31,191,31,15,31,98,31,98,30,98,29,98,28,79,31,61,31,164,31,90,31,93,31,93,30,80,31,250,31,139,31,139,30,139,29,111,31,8,31,244,31,60,31,90,31,90,30,169,31,169,30,181,31,206,31,96,31,172,31,172,30,201,31,18,31,238,31,153,31,153,30,2,31,149,31,149,30,13,31,41,31,137,31,49,31,49,30,88,31,88,30,88,29,135,31,135,30,98,31,109,31,45,31,131,31,119,31,102,31,180,31,180,30,232,31,232,30,232,29,121,31,121,30,94,31,106,31,69,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
