-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 413;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (61,0,9,0,191,0,142,0,0,0,0,0,135,0,0,0,64,0,0,0,42,0,251,0,148,0,0,0,113,0,0,0,66,0,29,0,0,0,0,0,21,0,93,0,78,0,159,0,214,0,250,0,131,0,233,0,32,0,86,0,139,0,201,0,72,0,46,0,223,0,0,0,129,0,39,0,96,0,3,0,219,0,0,0,27,0,148,0,206,0,170,0,42,0,0,0,101,0,0,0,0,0,0,0,203,0,66,0,77,0,197,0,125,0,24,0,214,0,0,0,239,0,0,0,6,0,211,0,39,0,0,0,7,0,140,0,133,0,46,0,87,0,0,0,135,0,45,0,0,0,137,0,157,0,160,0,235,0,218,0,225,0,190,0,90,0,60,0,0,0,89,0,138,0,178,0,31,0,0,0,216,0,39,0,201,0,3,0,212,0,0,0,220,0,17,0,121,0,0,0,197,0,129,0,32,0,39,0,251,0,140,0,112,0,0,0,0,0,32,0,177,0,27,0,0,0,134,0,216,0,249,0,131,0,92,0,203,0,191,0,80,0,206,0,4,0,179,0,235,0,227,0,72,0,38,0,149,0,16,0,90,0,85,0,238,0,120,0,174,0,0,0,241,0,0,0,218,0,56,0,35,0,0,0,0,0,110,0,24,0,140,0,143,0,42,0,41,0,181,0,127,0,47,0,215,0,152,0,112,0,0,0,79,0,199,0,100,0,27,0,33,0,236,0,57,0,0,0,208,0,161,0,210,0,189,0,250,0,64,0,5,0,0,0,0,0,0,0,141,0,202,0,80,0,0,0,16,0,74,0,0,0,189,0,204,0,57,0,238,0,0,0,0,0,68,0,124,0,173,0,0,0,83,0,0,0,22,0,0,0,127,0,246,0,85,0,133,0,36,0,7,0,0,0,189,0,157,0,144,0,96,0,234,0,0,0,86,0,196,0,91,0,0,0,21,0,107,0,0,0,140,0,165,0,213,0,0,0,0,0,204,0,91,0,0,0,215,0,180,0,197,0,87,0,205,0,222,0,0,0,0,0,106,0,31,0,129,0,41,0,0,0,0,0,255,0,13,0,217,0,0,0,138,0,78,0,58,0,236,0,196,0,0,0,33,0,188,0,216,0,67,0,0,0,88,0,0,0,248,0,48,0,86,0,57,0,0,0,57,0,79,0,133,0,204,0,157,0,179,0,34,0,0,0,108,0,150,0,82,0,203,0,225,0,144,0,25,0,15,0,81,0,197,0,74,0,12,0,80,0,189,0,81,0,0,0,0,0,8,0,187,0,111,0,31,0,142,0,25,0,238,0,43,0,169,0,51,0,86,0,246,0,0,0,117,0,197,0,156,0,37,0,59,0,0,0,194,0,74,0,39,0,0,0,152,0,233,0,151,0,91,0,0,0,211,0,108,0,120,0,228,0,104,0,0,0,174,0,35,0,0,0,91,0,0,0,9,0,149,0,92,0,0,0,0,0,222,0,95,0,25,0,228,0,0,0,188,0,198,0,7,0,229,0,0,0,253,0,0,0,40,0,180,0,213,0,179,0,240,0,187,0,178,0,51,0,155,0,0,0,226,0,166,0,0,0,69,0,0,0,133,0,100,0,0,0,5,0,54,0,0,0,127,0,121,0,0,0,177,0,100,0,142,0,163,0,0,0,122,0,75,0,20,0,77,0,21,0,0,0,201,0,216,0,220,0,181,0,12,0,79,0,248,0,84,0,128,0,249,0,178,0,168,0,135,0,0,0,0,0,165,0,0,0,162,0,0,0,65,0,29,0,0,0,179,0,79,0,0,0,144,0,0,0,188,0,133,0,110,0,0,0,187,0,0,0,252,0,70,0,14,0,56,0,41,0);
signal scenario_full  : scenario_type := (61,31,9,31,191,31,142,31,142,30,142,29,135,31,135,30,64,31,64,30,42,31,251,31,148,31,148,30,113,31,113,30,66,31,29,31,29,30,29,29,21,31,93,31,78,31,159,31,214,31,250,31,131,31,233,31,32,31,86,31,139,31,201,31,72,31,46,31,223,31,223,30,129,31,39,31,96,31,3,31,219,31,219,30,27,31,148,31,206,31,170,31,42,31,42,30,101,31,101,30,101,29,101,28,203,31,66,31,77,31,197,31,125,31,24,31,214,31,214,30,239,31,239,30,6,31,211,31,39,31,39,30,7,31,140,31,133,31,46,31,87,31,87,30,135,31,45,31,45,30,137,31,157,31,160,31,235,31,218,31,225,31,190,31,90,31,60,31,60,30,89,31,138,31,178,31,31,31,31,30,216,31,39,31,201,31,3,31,212,31,212,30,220,31,17,31,121,31,121,30,197,31,129,31,32,31,39,31,251,31,140,31,112,31,112,30,112,29,32,31,177,31,27,31,27,30,134,31,216,31,249,31,131,31,92,31,203,31,191,31,80,31,206,31,4,31,179,31,235,31,227,31,72,31,38,31,149,31,16,31,90,31,85,31,238,31,120,31,174,31,174,30,241,31,241,30,218,31,56,31,35,31,35,30,35,29,110,31,24,31,140,31,143,31,42,31,41,31,181,31,127,31,47,31,215,31,152,31,112,31,112,30,79,31,199,31,100,31,27,31,33,31,236,31,57,31,57,30,208,31,161,31,210,31,189,31,250,31,64,31,5,31,5,30,5,29,5,28,141,31,202,31,80,31,80,30,16,31,74,31,74,30,189,31,204,31,57,31,238,31,238,30,238,29,68,31,124,31,173,31,173,30,83,31,83,30,22,31,22,30,127,31,246,31,85,31,133,31,36,31,7,31,7,30,189,31,157,31,144,31,96,31,234,31,234,30,86,31,196,31,91,31,91,30,21,31,107,31,107,30,140,31,165,31,213,31,213,30,213,29,204,31,91,31,91,30,215,31,180,31,197,31,87,31,205,31,222,31,222,30,222,29,106,31,31,31,129,31,41,31,41,30,41,29,255,31,13,31,217,31,217,30,138,31,78,31,58,31,236,31,196,31,196,30,33,31,188,31,216,31,67,31,67,30,88,31,88,30,248,31,48,31,86,31,57,31,57,30,57,31,79,31,133,31,204,31,157,31,179,31,34,31,34,30,108,31,150,31,82,31,203,31,225,31,144,31,25,31,15,31,81,31,197,31,74,31,12,31,80,31,189,31,81,31,81,30,81,29,8,31,187,31,111,31,31,31,142,31,25,31,238,31,43,31,169,31,51,31,86,31,246,31,246,30,117,31,197,31,156,31,37,31,59,31,59,30,194,31,74,31,39,31,39,30,152,31,233,31,151,31,91,31,91,30,211,31,108,31,120,31,228,31,104,31,104,30,174,31,35,31,35,30,91,31,91,30,9,31,149,31,92,31,92,30,92,29,222,31,95,31,25,31,228,31,228,30,188,31,198,31,7,31,229,31,229,30,253,31,253,30,40,31,180,31,213,31,179,31,240,31,187,31,178,31,51,31,155,31,155,30,226,31,166,31,166,30,69,31,69,30,133,31,100,31,100,30,5,31,54,31,54,30,127,31,121,31,121,30,177,31,100,31,142,31,163,31,163,30,122,31,75,31,20,31,77,31,21,31,21,30,201,31,216,31,220,31,181,31,12,31,79,31,248,31,84,31,128,31,249,31,178,31,168,31,135,31,135,30,135,29,165,31,165,30,162,31,162,30,65,31,29,31,29,30,179,31,79,31,79,30,144,31,144,30,188,31,133,31,110,31,110,30,187,31,187,30,252,31,70,31,14,31,56,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
