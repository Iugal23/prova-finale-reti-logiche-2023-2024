-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 694;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (55,0,63,0,146,0,10,0,238,0,113,0,43,0,154,0,241,0,0,0,0,0,49,0,246,0,0,0,184,0,69,0,0,0,101,0,30,0,67,0,0,0,0,0,14,0,0,0,70,0,244,0,0,0,181,0,50,0,0,0,77,0,70,0,95,0,72,0,90,0,144,0,233,0,0,0,255,0,119,0,10,0,213,0,155,0,0,0,176,0,0,0,35,0,96,0,0,0,178,0,243,0,0,0,0,0,147,0,169,0,0,0,31,0,0,0,106,0,101,0,167,0,26,0,169,0,249,0,147,0,24,0,112,0,11,0,192,0,149,0,77,0,153,0,219,0,15,0,250,0,0,0,211,0,52,0,0,0,0,0,29,0,207,0,101,0,109,0,180,0,0,0,229,0,0,0,227,0,252,0,102,0,48,0,0,0,249,0,174,0,0,0,55,0,224,0,99,0,158,0,203,0,109,0,25,0,46,0,206,0,100,0,214,0,22,0,203,0,136,0,70,0,205,0,0,0,158,0,139,0,0,0,245,0,46,0,41,0,0,0,199,0,59,0,0,0,68,0,19,0,202,0,129,0,249,0,54,0,0,0,251,0,155,0,0,0,0,0,9,0,15,0,0,0,3,0,0,0,0,0,240,0,90,0,0,0,23,0,133,0,158,0,185,0,221,0,124,0,127,0,252,0,0,0,0,0,0,0,172,0,31,0,14,0,111,0,249,0,19,0,8,0,244,0,107,0,176,0,225,0,81,0,45,0,212,0,0,0,122,0,119,0,194,0,226,0,255,0,0,0,134,0,0,0,233,0,164,0,0,0,2,0,113,0,247,0,0,0,0,0,174,0,148,0,59,0,228,0,156,0,215,0,180,0,221,0,75,0,205,0,0,0,0,0,8,0,189,0,0,0,215,0,243,0,31,0,151,0,191,0,0,0,234,0,213,0,0,0,15,0,215,0,0,0,149,0,186,0,192,0,0,0,0,0,252,0,0,0,0,0,0,0,0,0,86,0,211,0,209,0,70,0,96,0,233,0,95,0,253,0,53,0,0,0,124,0,122,0,128,0,0,0,4,0,0,0,19,0,183,0,229,0,35,0,177,0,122,0,0,0,132,0,0,0,191,0,148,0,64,0,104,0,156,0,0,0,127,0,28,0,184,0,160,0,144,0,218,0,0,0,187,0,0,0,168,0,202,0,0,0,179,0,51,0,51,0,223,0,101,0,68,0,50,0,237,0,37,0,85,0,0,0,0,0,120,0,14,0,120,0,214,0,41,0,248,0,0,0,176,0,214,0,254,0,213,0,23,0,222,0,0,0,8,0,2,0,1,0,0,0,0,0,189,0,21,0,103,0,198,0,0,0,85,0,0,0,153,0,57,0,0,0,17,0,58,0,45,0,168,0,201,0,119,0,112,0,251,0,171,0,180,0,216,0,250,0,17,0,210,0,235,0,97,0,210,0,25,0,85,0,198,0,124,0,136,0,153,0,0,0,0,0,118,0,90,0,205,0,27,0,122,0,241,0,0,0,181,0,251,0,144,0,241,0,76,0,24,0,56,0,0,0,0,0,220,0,234,0,54,0,39,0,16,0,215,0,89,0,73,0,154,0,131,0,91,0,0,0,25,0,34,0,1,0,152,0,245,0,226,0,84,0,0,0,142,0,166,0,211,0,191,0,104,0,211,0,243,0,5,0,0,0,0,0,0,0,57,0,0,0,0,0,56,0,205,0,5,0,152,0,0,0,78,0,225,0,142,0,236,0,100,0,250,0,0,0,36,0,0,0,160,0,171,0,21,0,39,0,0,0,214,0,0,0,125,0,72,0,26,0,210,0,56,0,0,0,0,0,0,0,109,0,111,0,158,0,165,0,150,0,0,0,0,0,241,0,126,0,218,0,141,0,200,0,108,0,158,0,230,0,5,0,185,0,141,0,249,0,101,0,119,0,78,0,0,0,66,0,28,0,9,0,158,0,0,0,0,0,69,0,10,0,97,0,231,0,97,0,157,0,221,0,123,0,100,0,0,0,0,0,173,0,170,0,0,0,83,0,96,0,0,0,254,0,0,0,101,0,245,0,25,0,181,0,52,0,220,0,59,0,204,0,88,0,207,0,0,0,61,0,0,0,4,0,95,0,57,0,104,0,100,0,0,0,173,0,58,0,0,0,21,0,115,0,194,0,8,0,0,0,53,0,0,0,106,0,44,0,0,0,92,0,0,0,0,0,48,0,178,0,189,0,234,0,163,0,195,0,124,0,132,0,235,0,0,0,0,0,70,0,42,0,253,0,130,0,0,0,223,0,39,0,0,0,73,0,0,0,183,0,60,0,218,0,0,0,89,0,140,0,222,0,159,0,151,0,134,0,108,0,223,0,217,0,0,0,0,0,105,0,154,0,17,0,23,0,13,0,108,0,221,0,36,0,220,0,90,0,35,0,41,0,0,0,20,0,108,0,200,0,149,0,0,0,129,0,236,0,97,0,45,0,0,0,124,0,94,0,181,0,210,0,215,0,180,0,0,0,0,0,9,0,67,0,0,0,236,0,175,0,75,0,35,0,132,0,78,0,195,0,0,0,185,0,31,0,246,0,246,0,1,0,16,0,72,0,0,0,6,0,42,0,17,0,145,0,0,0,0,0,200,0,195,0,0,0,90,0,158,0,0,0,175,0,143,0,124,0,117,0,147,0,126,0,0,0,221,0,140,0,184,0,107,0,0,0,4,0,161,0,65,0,217,0,224,0,65,0,0,0,146,0,88,0,219,0,57,0,0,0,246,0,0,0,0,0,198,0,5,0,1,0,86,0,19,0,81,0,92,0,239,0,160,0,45,0,23,0,123,0,0,0,0,0,0,0,1,0,245,0,225,0,11,0,36,0,229,0,234,0,0,0,103,0,124,0,45,0,49,0,86,0,27,0,142,0,0,0,153,0,30,0,242,0,170,0,0,0,125,0,199,0,32,0,227,0,142,0,14,0,55,0,89,0,196,0,255,0,190,0,247,0,73,0,0,0,84,0,152,0,157,0,71,0,115,0,178,0,79,0,0,0,151,0,101,0,0,0,141,0,88,0,0,0,0,0,203,0,188,0,0,0,229,0,0,0,0,0,78,0,155,0,122,0,192,0,193,0);
signal scenario_full  : scenario_type := (55,31,63,31,146,31,10,31,238,31,113,31,43,31,154,31,241,31,241,30,241,29,49,31,246,31,246,30,184,31,69,31,69,30,101,31,30,31,67,31,67,30,67,29,14,31,14,30,70,31,244,31,244,30,181,31,50,31,50,30,77,31,70,31,95,31,72,31,90,31,144,31,233,31,233,30,255,31,119,31,10,31,213,31,155,31,155,30,176,31,176,30,35,31,96,31,96,30,178,31,243,31,243,30,243,29,147,31,169,31,169,30,31,31,31,30,106,31,101,31,167,31,26,31,169,31,249,31,147,31,24,31,112,31,11,31,192,31,149,31,77,31,153,31,219,31,15,31,250,31,250,30,211,31,52,31,52,30,52,29,29,31,207,31,101,31,109,31,180,31,180,30,229,31,229,30,227,31,252,31,102,31,48,31,48,30,249,31,174,31,174,30,55,31,224,31,99,31,158,31,203,31,109,31,25,31,46,31,206,31,100,31,214,31,22,31,203,31,136,31,70,31,205,31,205,30,158,31,139,31,139,30,245,31,46,31,41,31,41,30,199,31,59,31,59,30,68,31,19,31,202,31,129,31,249,31,54,31,54,30,251,31,155,31,155,30,155,29,9,31,15,31,15,30,3,31,3,30,3,29,240,31,90,31,90,30,23,31,133,31,158,31,185,31,221,31,124,31,127,31,252,31,252,30,252,29,252,28,172,31,31,31,14,31,111,31,249,31,19,31,8,31,244,31,107,31,176,31,225,31,81,31,45,31,212,31,212,30,122,31,119,31,194,31,226,31,255,31,255,30,134,31,134,30,233,31,164,31,164,30,2,31,113,31,247,31,247,30,247,29,174,31,148,31,59,31,228,31,156,31,215,31,180,31,221,31,75,31,205,31,205,30,205,29,8,31,189,31,189,30,215,31,243,31,31,31,151,31,191,31,191,30,234,31,213,31,213,30,15,31,215,31,215,30,149,31,186,31,192,31,192,30,192,29,252,31,252,30,252,29,252,28,252,27,86,31,211,31,209,31,70,31,96,31,233,31,95,31,253,31,53,31,53,30,124,31,122,31,128,31,128,30,4,31,4,30,19,31,183,31,229,31,35,31,177,31,122,31,122,30,132,31,132,30,191,31,148,31,64,31,104,31,156,31,156,30,127,31,28,31,184,31,160,31,144,31,218,31,218,30,187,31,187,30,168,31,202,31,202,30,179,31,51,31,51,31,223,31,101,31,68,31,50,31,237,31,37,31,85,31,85,30,85,29,120,31,14,31,120,31,214,31,41,31,248,31,248,30,176,31,214,31,254,31,213,31,23,31,222,31,222,30,8,31,2,31,1,31,1,30,1,29,189,31,21,31,103,31,198,31,198,30,85,31,85,30,153,31,57,31,57,30,17,31,58,31,45,31,168,31,201,31,119,31,112,31,251,31,171,31,180,31,216,31,250,31,17,31,210,31,235,31,97,31,210,31,25,31,85,31,198,31,124,31,136,31,153,31,153,30,153,29,118,31,90,31,205,31,27,31,122,31,241,31,241,30,181,31,251,31,144,31,241,31,76,31,24,31,56,31,56,30,56,29,220,31,234,31,54,31,39,31,16,31,215,31,89,31,73,31,154,31,131,31,91,31,91,30,25,31,34,31,1,31,152,31,245,31,226,31,84,31,84,30,142,31,166,31,211,31,191,31,104,31,211,31,243,31,5,31,5,30,5,29,5,28,57,31,57,30,57,29,56,31,205,31,5,31,152,31,152,30,78,31,225,31,142,31,236,31,100,31,250,31,250,30,36,31,36,30,160,31,171,31,21,31,39,31,39,30,214,31,214,30,125,31,72,31,26,31,210,31,56,31,56,30,56,29,56,28,109,31,111,31,158,31,165,31,150,31,150,30,150,29,241,31,126,31,218,31,141,31,200,31,108,31,158,31,230,31,5,31,185,31,141,31,249,31,101,31,119,31,78,31,78,30,66,31,28,31,9,31,158,31,158,30,158,29,69,31,10,31,97,31,231,31,97,31,157,31,221,31,123,31,100,31,100,30,100,29,173,31,170,31,170,30,83,31,96,31,96,30,254,31,254,30,101,31,245,31,25,31,181,31,52,31,220,31,59,31,204,31,88,31,207,31,207,30,61,31,61,30,4,31,95,31,57,31,104,31,100,31,100,30,173,31,58,31,58,30,21,31,115,31,194,31,8,31,8,30,53,31,53,30,106,31,44,31,44,30,92,31,92,30,92,29,48,31,178,31,189,31,234,31,163,31,195,31,124,31,132,31,235,31,235,30,235,29,70,31,42,31,253,31,130,31,130,30,223,31,39,31,39,30,73,31,73,30,183,31,60,31,218,31,218,30,89,31,140,31,222,31,159,31,151,31,134,31,108,31,223,31,217,31,217,30,217,29,105,31,154,31,17,31,23,31,13,31,108,31,221,31,36,31,220,31,90,31,35,31,41,31,41,30,20,31,108,31,200,31,149,31,149,30,129,31,236,31,97,31,45,31,45,30,124,31,94,31,181,31,210,31,215,31,180,31,180,30,180,29,9,31,67,31,67,30,236,31,175,31,75,31,35,31,132,31,78,31,195,31,195,30,185,31,31,31,246,31,246,31,1,31,16,31,72,31,72,30,6,31,42,31,17,31,145,31,145,30,145,29,200,31,195,31,195,30,90,31,158,31,158,30,175,31,143,31,124,31,117,31,147,31,126,31,126,30,221,31,140,31,184,31,107,31,107,30,4,31,161,31,65,31,217,31,224,31,65,31,65,30,146,31,88,31,219,31,57,31,57,30,246,31,246,30,246,29,198,31,5,31,1,31,86,31,19,31,81,31,92,31,239,31,160,31,45,31,23,31,123,31,123,30,123,29,123,28,1,31,245,31,225,31,11,31,36,31,229,31,234,31,234,30,103,31,124,31,45,31,49,31,86,31,27,31,142,31,142,30,153,31,30,31,242,31,170,31,170,30,125,31,199,31,32,31,227,31,142,31,14,31,55,31,89,31,196,31,255,31,190,31,247,31,73,31,73,30,84,31,152,31,157,31,71,31,115,31,178,31,79,31,79,30,151,31,101,31,101,30,141,31,88,31,88,30,88,29,203,31,188,31,188,30,229,31,229,30,229,29,78,31,155,31,122,31,192,31,193,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
