-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 360;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (233,0,116,0,82,0,54,0,154,0,144,0,174,0,145,0,0,0,0,0,191,0,27,0,189,0,185,0,206,0,0,0,0,0,24,0,127,0,70,0,0,0,188,0,0,0,132,0,150,0,231,0,18,0,54,0,206,0,239,0,243,0,242,0,46,0,0,0,69,0,7,0,165,0,74,0,253,0,19,0,181,0,35,0,207,0,0,0,134,0,0,0,89,0,0,0,0,0,40,0,13,0,0,0,62,0,124,0,153,0,160,0,154,0,0,0,192,0,24,0,34,0,59,0,16,0,0,0,200,0,201,0,41,0,83,0,214,0,111,0,177,0,0,0,174,0,219,0,9,0,229,0,83,0,18,0,170,0,27,0,36,0,70,0,188,0,193,0,240,0,162,0,208,0,82,0,90,0,21,0,165,0,58,0,75,0,0,0,211,0,0,0,20,0,232,0,9,0,2,0,200,0,0,0,37,0,61,0,200,0,0,0,213,0,0,0,0,0,27,0,0,0,0,0,82,0,230,0,44,0,228,0,0,0,158,0,170,0,0,0,0,0,165,0,199,0,117,0,108,0,102,0,98,0,252,0,137,0,0,0,0,0,240,0,190,0,222,0,5,0,0,0,0,0,104,0,0,0,119,0,159,0,165,0,81,0,118,0,28,0,78,0,0,0,0,0,235,0,0,0,0,0,0,0,151,0,210,0,15,0,55,0,54,0,185,0,78,0,0,0,3,0,223,0,30,0,84,0,68,0,9,0,0,0,161,0,217,0,26,0,14,0,0,0,97,0,0,0,111,0,195,0,219,0,252,0,213,0,71,0,226,0,0,0,107,0,121,0,81,0,146,0,121,0,0,0,188,0,19,0,203,0,0,0,82,0,0,0,102,0,89,0,215,0,200,0,46,0,202,0,0,0,133,0,0,0,0,0,0,0,78,0,0,0,24,0,62,0,46,0,0,0,55,0,0,0,210,0,166,0,174,0,0,0,79,0,86,0,0,0,215,0,154,0,245,0,176,0,204,0,49,0,125,0,28,0,237,0,52,0,199,0,242,0,65,0,42,0,200,0,31,0,0,0,230,0,252,0,0,0,64,0,85,0,51,0,101,0,0,0,94,0,0,0,166,0,149,0,140,0,183,0,0,0,185,0,200,0,0,0,0,0,203,0,74,0,184,0,0,0,0,0,0,0,250,0,62,0,0,0,0,0,175,0,223,0,165,0,235,0,119,0,113,0,220,0,122,0,0,0,160,0,220,0,16,0,183,0,157,0,246,0,47,0,0,0,0,0,214,0,126,0,136,0,42,0,99,0,0,0,194,0,187,0,76,0,58,0,158,0,201,0,22,0,10,0,33,0,224,0,45,0,0,0,223,0,168,0,132,0,255,0,98,0,0,0,151,0,0,0,105,0,246,0,60,0,179,0,113,0,63,0,37,0,0,0,37,0,141,0,156,0,0,0,162,0,0,0,209,0,193,0,242,0,53,0,0,0,157,0,84,0,78,0,94,0,32,0,196,0,155,0,21,0,17,0,77,0,129,0,0,0,0,0,0,0,0,0,38,0,38,0,98,0,229,0,18,0,94,0,157,0,206,0,116,0,0,0,7,0,47,0,14,0,50,0,114,0,108,0);
signal scenario_full  : scenario_type := (233,31,116,31,82,31,54,31,154,31,144,31,174,31,145,31,145,30,145,29,191,31,27,31,189,31,185,31,206,31,206,30,206,29,24,31,127,31,70,31,70,30,188,31,188,30,132,31,150,31,231,31,18,31,54,31,206,31,239,31,243,31,242,31,46,31,46,30,69,31,7,31,165,31,74,31,253,31,19,31,181,31,35,31,207,31,207,30,134,31,134,30,89,31,89,30,89,29,40,31,13,31,13,30,62,31,124,31,153,31,160,31,154,31,154,30,192,31,24,31,34,31,59,31,16,31,16,30,200,31,201,31,41,31,83,31,214,31,111,31,177,31,177,30,174,31,219,31,9,31,229,31,83,31,18,31,170,31,27,31,36,31,70,31,188,31,193,31,240,31,162,31,208,31,82,31,90,31,21,31,165,31,58,31,75,31,75,30,211,31,211,30,20,31,232,31,9,31,2,31,200,31,200,30,37,31,61,31,200,31,200,30,213,31,213,30,213,29,27,31,27,30,27,29,82,31,230,31,44,31,228,31,228,30,158,31,170,31,170,30,170,29,165,31,199,31,117,31,108,31,102,31,98,31,252,31,137,31,137,30,137,29,240,31,190,31,222,31,5,31,5,30,5,29,104,31,104,30,119,31,159,31,165,31,81,31,118,31,28,31,78,31,78,30,78,29,235,31,235,30,235,29,235,28,151,31,210,31,15,31,55,31,54,31,185,31,78,31,78,30,3,31,223,31,30,31,84,31,68,31,9,31,9,30,161,31,217,31,26,31,14,31,14,30,97,31,97,30,111,31,195,31,219,31,252,31,213,31,71,31,226,31,226,30,107,31,121,31,81,31,146,31,121,31,121,30,188,31,19,31,203,31,203,30,82,31,82,30,102,31,89,31,215,31,200,31,46,31,202,31,202,30,133,31,133,30,133,29,133,28,78,31,78,30,24,31,62,31,46,31,46,30,55,31,55,30,210,31,166,31,174,31,174,30,79,31,86,31,86,30,215,31,154,31,245,31,176,31,204,31,49,31,125,31,28,31,237,31,52,31,199,31,242,31,65,31,42,31,200,31,31,31,31,30,230,31,252,31,252,30,64,31,85,31,51,31,101,31,101,30,94,31,94,30,166,31,149,31,140,31,183,31,183,30,185,31,200,31,200,30,200,29,203,31,74,31,184,31,184,30,184,29,184,28,250,31,62,31,62,30,62,29,175,31,223,31,165,31,235,31,119,31,113,31,220,31,122,31,122,30,160,31,220,31,16,31,183,31,157,31,246,31,47,31,47,30,47,29,214,31,126,31,136,31,42,31,99,31,99,30,194,31,187,31,76,31,58,31,158,31,201,31,22,31,10,31,33,31,224,31,45,31,45,30,223,31,168,31,132,31,255,31,98,31,98,30,151,31,151,30,105,31,246,31,60,31,179,31,113,31,63,31,37,31,37,30,37,31,141,31,156,31,156,30,162,31,162,30,209,31,193,31,242,31,53,31,53,30,157,31,84,31,78,31,94,31,32,31,196,31,155,31,21,31,17,31,77,31,129,31,129,30,129,29,129,28,129,27,38,31,38,31,98,31,229,31,18,31,94,31,157,31,206,31,116,31,116,30,7,31,47,31,14,31,50,31,114,31,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
