-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 767;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (229,0,0,0,16,0,221,0,41,0,234,0,0,0,93,0,142,0,105,0,0,0,55,0,0,0,129,0,0,0,77,0,28,0,246,0,42,0,105,0,0,0,31,0,40,0,202,0,0,0,0,0,29,0,165,0,103,0,16,0,184,0,83,0,159,0,202,0,39,0,131,0,234,0,0,0,70,0,102,0,211,0,92,0,194,0,0,0,55,0,181,0,0,0,250,0,41,0,0,0,253,0,177,0,186,0,25,0,13,0,69,0,0,0,0,0,217,0,0,0,17,0,94,0,72,0,173,0,207,0,0,0,160,0,112,0,68,0,28,0,0,0,212,0,107,0,156,0,96,0,251,0,77,0,181,0,238,0,40,0,42,0,160,0,0,0,27,0,51,0,123,0,174,0,82,0,0,0,79,0,172,0,71,0,201,0,71,0,255,0,23,0,103,0,82,0,233,0,55,0,48,0,0,0,88,0,161,0,72,0,0,0,121,0,1,0,90,0,128,0,173,0,38,0,160,0,37,0,51,0,248,0,0,0,0,0,181,0,71,0,104,0,0,0,19,0,189,0,187,0,112,0,227,0,42,0,240,0,249,0,168,0,239,0,234,0,48,0,239,0,116,0,229,0,18,0,0,0,0,0,38,0,90,0,169,0,157,0,0,0,0,0,68,0,88,0,41,0,114,0,0,0,31,0,60,0,167,0,247,0,153,0,0,0,88,0,0,0,206,0,207,0,96,0,37,0,0,0,0,0,253,0,153,0,96,0,39,0,0,0,229,0,244,0,179,0,0,0,21,0,5,0,225,0,164,0,0,0,115,0,0,0,226,0,104,0,110,0,11,0,15,0,0,0,0,0,13,0,203,0,122,0,197,0,236,0,237,0,0,0,164,0,58,0,160,0,248,0,64,0,63,0,63,0,6,0,213,0,0,0,202,0,60,0,218,0,176,0,250,0,0,0,57,0,148,0,14,0,9,0,29,0,235,0,192,0,129,0,153,0,80,0,58,0,160,0,0,0,214,0,95,0,234,0,0,0,191,0,35,0,200,0,0,0,131,0,0,0,121,0,0,0,44,0,230,0,68,0,224,0,22,0,77,0,229,0,6,0,173,0,166,0,177,0,125,0,34,0,0,0,155,0,127,0,140,0,109,0,178,0,33,0,1,0,131,0,20,0,247,0,0,0,0,0,209,0,0,0,246,0,207,0,181,0,0,0,255,0,191,0,221,0,53,0,99,0,0,0,221,0,114,0,0,0,83,0,0,0,125,0,194,0,241,0,157,0,177,0,0,0,118,0,90,0,104,0,250,0,4,0,188,0,129,0,178,0,11,0,221,0,116,0,0,0,212,0,15,0,241,0,252,0,138,0,47,0,46,0,0,0,252,0,0,0,145,0,168,0,10,0,134,0,244,0,169,0,4,0,13,0,196,0,53,0,200,0,107,0,10,0,99,0,68,0,121,0,131,0,36,0,95,0,131,0,3,0,27,0,178,0,4,0,134,0,215,0,196,0,245,0,138,0,0,0,0,0,81,0,152,0,109,0,242,0,44,0,37,0,192,0,7,0,0,0,178,0,78,0,1,0,98,0,103,0,0,0,136,0,235,0,197,0,0,0,233,0,227,0,155,0,67,0,0,0,93,0,71,0,225,0,150,0,120,0,244,0,0,0,158,0,79,0,5,0,0,0,48,0,22,0,87,0,136,0,46,0,0,0,243,0,0,0,0,0,37,0,80,0,190,0,27,0,211,0,226,0,206,0,26,0,133,0,1,0,71,0,124,0,20,0,163,0,21,0,85,0,144,0,24,0,30,0,195,0,146,0,87,0,0,0,59,0,55,0,207,0,153,0,29,0,114,0,0,0,183,0,169,0,133,0,215,0,57,0,9,0,116,0,103,0,21,0,235,0,103,0,0,0,111,0,123,0,0,0,102,0,204,0,235,0,176,0,122,0,0,0,242,0,172,0,235,0,33,0,157,0,0,0,113,0,156,0,88,0,21,0,6,0,53,0,187,0,0,0,92,0,0,0,37,0,0,0,241,0,223,0,233,0,0,0,31,0,77,0,186,0,0,0,0,0,253,0,187,0,0,0,168,0,0,0,227,0,245,0,0,0,139,0,156,0,0,0,0,0,229,0,0,0,178,0,244,0,180,0,109,0,176,0,143,0,0,0,239,0,0,0,239,0,0,0,198,0,126,0,112,0,120,0,217,0,0,0,101,0,0,0,92,0,95,0,203,0,0,0,176,0,107,0,30,0,158,0,3,0,0,0,168,0,0,0,150,0,222,0,0,0,247,0,157,0,50,0,0,0,146,0,14,0,149,0,160,0,9,0,138,0,0,0,2,0,16,0,149,0,113,0,167,0,16,0,160,0,0,0,218,0,0,0,77,0,0,0,0,0,88,0,173,0,102,0,0,0,0,0,162,0,110,0,0,0,148,0,248,0,117,0,42,0,0,0,134,0,238,0,11,0,208,0,215,0,89,0,0,0,55,0,233,0,165,0,244,0,9,0,114,0,131,0,0,0,6,0,231,0,117,0,235,0,0,0,44,0,88,0,242,0,80,0,160,0,0,0,0,0,0,0,178,0,249,0,174,0,0,0,0,0,0,0,50,0,117,0,0,0,9,0,198,0,158,0,90,0,0,0,0,0,0,0,143,0,45,0,61,0,17,0,32,0,252,0,115,0,229,0,0,0,36,0,224,0,193,0,29,0,208,0,252,0,0,0,61,0,0,0,183,0,86,0,131,0,181,0,0,0,157,0,0,0,17,0,150,0,127,0,50,0,249,0,156,0,225,0,238,0,202,0,127,0,0,0,68,0,69,0,225,0,102,0,233,0,104,0,0,0,81,0,248,0,161,0,183,0,117,0,156,0,155,0,11,0,0,0,88,0,0,0,243,0,183,0,14,0,142,0,210,0,0,0,70,0,19,0,20,0,147,0,72,0,169,0,0,0,39,0,86,0,38,0,164,0,165,0,43,0,0,0,95,0,216,0,195,0,0,0,17,0,252,0,48,0,69,0,35,0,156,0,163,0,12,0,242,0,252,0,90,0,68,0,232,0,32,0,0,0,144,0,3,0,0,0,52,0,59,0,0,0,252,0,153,0,0,0,46,0,197,0,199,0,91,0,112,0,0,0,68,0,95,0,30,0,57,0,193,0,148,0,0,0,189,0,0,0,206,0,204,0,0,0,0,0,230,0,88,0,100,0,138,0,239,0,123,0,0,0,54,0,75,0,109,0,237,0,143,0,0,0,236,0,0,0,250,0,225,0,45,0,3,0,18,0,122,0,121,0,180,0,20,0,201,0,193,0,172,0,97,0,120,0,67,0,214,0,164,0,154,0,108,0,175,0,11,0,143,0,10,0,50,0,201,0,144,0,186,0,154,0,0,0,55,0,13,0,53,0,0,0,191,0,145,0,161,0,182,0,0,0,0,0,0,0,181,0,131,0);
signal scenario_full  : scenario_type := (229,31,229,30,16,31,221,31,41,31,234,31,234,30,93,31,142,31,105,31,105,30,55,31,55,30,129,31,129,30,77,31,28,31,246,31,42,31,105,31,105,30,31,31,40,31,202,31,202,30,202,29,29,31,165,31,103,31,16,31,184,31,83,31,159,31,202,31,39,31,131,31,234,31,234,30,70,31,102,31,211,31,92,31,194,31,194,30,55,31,181,31,181,30,250,31,41,31,41,30,253,31,177,31,186,31,25,31,13,31,69,31,69,30,69,29,217,31,217,30,17,31,94,31,72,31,173,31,207,31,207,30,160,31,112,31,68,31,28,31,28,30,212,31,107,31,156,31,96,31,251,31,77,31,181,31,238,31,40,31,42,31,160,31,160,30,27,31,51,31,123,31,174,31,82,31,82,30,79,31,172,31,71,31,201,31,71,31,255,31,23,31,103,31,82,31,233,31,55,31,48,31,48,30,88,31,161,31,72,31,72,30,121,31,1,31,90,31,128,31,173,31,38,31,160,31,37,31,51,31,248,31,248,30,248,29,181,31,71,31,104,31,104,30,19,31,189,31,187,31,112,31,227,31,42,31,240,31,249,31,168,31,239,31,234,31,48,31,239,31,116,31,229,31,18,31,18,30,18,29,38,31,90,31,169,31,157,31,157,30,157,29,68,31,88,31,41,31,114,31,114,30,31,31,60,31,167,31,247,31,153,31,153,30,88,31,88,30,206,31,207,31,96,31,37,31,37,30,37,29,253,31,153,31,96,31,39,31,39,30,229,31,244,31,179,31,179,30,21,31,5,31,225,31,164,31,164,30,115,31,115,30,226,31,104,31,110,31,11,31,15,31,15,30,15,29,13,31,203,31,122,31,197,31,236,31,237,31,237,30,164,31,58,31,160,31,248,31,64,31,63,31,63,31,6,31,213,31,213,30,202,31,60,31,218,31,176,31,250,31,250,30,57,31,148,31,14,31,9,31,29,31,235,31,192,31,129,31,153,31,80,31,58,31,160,31,160,30,214,31,95,31,234,31,234,30,191,31,35,31,200,31,200,30,131,31,131,30,121,31,121,30,44,31,230,31,68,31,224,31,22,31,77,31,229,31,6,31,173,31,166,31,177,31,125,31,34,31,34,30,155,31,127,31,140,31,109,31,178,31,33,31,1,31,131,31,20,31,247,31,247,30,247,29,209,31,209,30,246,31,207,31,181,31,181,30,255,31,191,31,221,31,53,31,99,31,99,30,221,31,114,31,114,30,83,31,83,30,125,31,194,31,241,31,157,31,177,31,177,30,118,31,90,31,104,31,250,31,4,31,188,31,129,31,178,31,11,31,221,31,116,31,116,30,212,31,15,31,241,31,252,31,138,31,47,31,46,31,46,30,252,31,252,30,145,31,168,31,10,31,134,31,244,31,169,31,4,31,13,31,196,31,53,31,200,31,107,31,10,31,99,31,68,31,121,31,131,31,36,31,95,31,131,31,3,31,27,31,178,31,4,31,134,31,215,31,196,31,245,31,138,31,138,30,138,29,81,31,152,31,109,31,242,31,44,31,37,31,192,31,7,31,7,30,178,31,78,31,1,31,98,31,103,31,103,30,136,31,235,31,197,31,197,30,233,31,227,31,155,31,67,31,67,30,93,31,71,31,225,31,150,31,120,31,244,31,244,30,158,31,79,31,5,31,5,30,48,31,22,31,87,31,136,31,46,31,46,30,243,31,243,30,243,29,37,31,80,31,190,31,27,31,211,31,226,31,206,31,26,31,133,31,1,31,71,31,124,31,20,31,163,31,21,31,85,31,144,31,24,31,30,31,195,31,146,31,87,31,87,30,59,31,55,31,207,31,153,31,29,31,114,31,114,30,183,31,169,31,133,31,215,31,57,31,9,31,116,31,103,31,21,31,235,31,103,31,103,30,111,31,123,31,123,30,102,31,204,31,235,31,176,31,122,31,122,30,242,31,172,31,235,31,33,31,157,31,157,30,113,31,156,31,88,31,21,31,6,31,53,31,187,31,187,30,92,31,92,30,37,31,37,30,241,31,223,31,233,31,233,30,31,31,77,31,186,31,186,30,186,29,253,31,187,31,187,30,168,31,168,30,227,31,245,31,245,30,139,31,156,31,156,30,156,29,229,31,229,30,178,31,244,31,180,31,109,31,176,31,143,31,143,30,239,31,239,30,239,31,239,30,198,31,126,31,112,31,120,31,217,31,217,30,101,31,101,30,92,31,95,31,203,31,203,30,176,31,107,31,30,31,158,31,3,31,3,30,168,31,168,30,150,31,222,31,222,30,247,31,157,31,50,31,50,30,146,31,14,31,149,31,160,31,9,31,138,31,138,30,2,31,16,31,149,31,113,31,167,31,16,31,160,31,160,30,218,31,218,30,77,31,77,30,77,29,88,31,173,31,102,31,102,30,102,29,162,31,110,31,110,30,148,31,248,31,117,31,42,31,42,30,134,31,238,31,11,31,208,31,215,31,89,31,89,30,55,31,233,31,165,31,244,31,9,31,114,31,131,31,131,30,6,31,231,31,117,31,235,31,235,30,44,31,88,31,242,31,80,31,160,31,160,30,160,29,160,28,178,31,249,31,174,31,174,30,174,29,174,28,50,31,117,31,117,30,9,31,198,31,158,31,90,31,90,30,90,29,90,28,143,31,45,31,61,31,17,31,32,31,252,31,115,31,229,31,229,30,36,31,224,31,193,31,29,31,208,31,252,31,252,30,61,31,61,30,183,31,86,31,131,31,181,31,181,30,157,31,157,30,17,31,150,31,127,31,50,31,249,31,156,31,225,31,238,31,202,31,127,31,127,30,68,31,69,31,225,31,102,31,233,31,104,31,104,30,81,31,248,31,161,31,183,31,117,31,156,31,155,31,11,31,11,30,88,31,88,30,243,31,183,31,14,31,142,31,210,31,210,30,70,31,19,31,20,31,147,31,72,31,169,31,169,30,39,31,86,31,38,31,164,31,165,31,43,31,43,30,95,31,216,31,195,31,195,30,17,31,252,31,48,31,69,31,35,31,156,31,163,31,12,31,242,31,252,31,90,31,68,31,232,31,32,31,32,30,144,31,3,31,3,30,52,31,59,31,59,30,252,31,153,31,153,30,46,31,197,31,199,31,91,31,112,31,112,30,68,31,95,31,30,31,57,31,193,31,148,31,148,30,189,31,189,30,206,31,204,31,204,30,204,29,230,31,88,31,100,31,138,31,239,31,123,31,123,30,54,31,75,31,109,31,237,31,143,31,143,30,236,31,236,30,250,31,225,31,45,31,3,31,18,31,122,31,121,31,180,31,20,31,201,31,193,31,172,31,97,31,120,31,67,31,214,31,164,31,154,31,108,31,175,31,11,31,143,31,10,31,50,31,201,31,144,31,186,31,154,31,154,30,55,31,13,31,53,31,53,30,191,31,145,31,161,31,182,31,182,30,182,29,182,28,181,31,131,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
