-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 232;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,105,0,47,0,61,0,63,0,134,0,86,0,88,0,50,0,116,0,29,0,0,0,172,0,30,0,89,0,134,0,136,0,0,0,0,0,34,0,0,0,146,0,212,0,0,0,109,0,0,0,189,0,84,0,0,0,203,0,183,0,188,0,15,0,139,0,0,0,164,0,124,0,209,0,140,0,221,0,16,0,0,0,0,0,46,0,47,0,241,0,0,0,245,0,32,0,84,0,250,0,92,0,168,0,0,0,176,0,160,0,94,0,235,0,0,0,235,0,195,0,0,0,217,0,38,0,167,0,244,0,229,0,37,0,0,0,0,0,242,0,23,0,174,0,137,0,244,0,141,0,170,0,0,0,0,0,155,0,195,0,44,0,60,0,0,0,206,0,115,0,225,0,159,0,32,0,206,0,0,0,12,0,0,0,62,0,0,0,0,0,0,0,96,0,216,0,33,0,138,0,145,0,1,0,99,0,155,0,0,0,140,0,66,0,31,0,0,0,229,0,209,0,0,0,196,0,36,0,225,0,0,0,90,0,202,0,0,0,192,0,225,0,242,0,133,0,0,0,131,0,211,0,0,0,38,0,0,0,80,0,0,0,132,0,0,0,108,0,17,0,204,0,181,0,0,0,42,0,0,0,114,0,135,0,87,0,128,0,26,0,212,0,0,0,24,0,74,0,24,0,203,0,220,0,46,0,92,0,153,0,121,0,74,0,112,0,189,0,69,0,210,0,6,0,69,0,109,0,28,0,245,0,28,0,191,0,32,0,35,0,14,0,154,0,0,0,62,0,185,0,221,0,17,0,184,0,233,0,0,0,82,0,0,0,182,0,221,0,5,0,167,0,249,0,154,0,0,0,201,0,188,0,144,0,219,0,5,0,30,0,129,0,155,0,180,0,45,0,6,0,93,0,34,0,96,0,44,0,180,0,72,0,78,0,247,0,0,0,2,0,81,0,12,0,6,0,45,0,71,0,47,0,230,0,246,0,185,0,245,0,0,0,16,0,66,0,27,0,0,0,0,0,109,0,0,0,241,0,113,0,0,0);
signal scenario_full  : scenario_type := (0,0,105,31,47,31,61,31,63,31,134,31,86,31,88,31,50,31,116,31,29,31,29,30,172,31,30,31,89,31,134,31,136,31,136,30,136,29,34,31,34,30,146,31,212,31,212,30,109,31,109,30,189,31,84,31,84,30,203,31,183,31,188,31,15,31,139,31,139,30,164,31,124,31,209,31,140,31,221,31,16,31,16,30,16,29,46,31,47,31,241,31,241,30,245,31,32,31,84,31,250,31,92,31,168,31,168,30,176,31,160,31,94,31,235,31,235,30,235,31,195,31,195,30,217,31,38,31,167,31,244,31,229,31,37,31,37,30,37,29,242,31,23,31,174,31,137,31,244,31,141,31,170,31,170,30,170,29,155,31,195,31,44,31,60,31,60,30,206,31,115,31,225,31,159,31,32,31,206,31,206,30,12,31,12,30,62,31,62,30,62,29,62,28,96,31,216,31,33,31,138,31,145,31,1,31,99,31,155,31,155,30,140,31,66,31,31,31,31,30,229,31,209,31,209,30,196,31,36,31,225,31,225,30,90,31,202,31,202,30,192,31,225,31,242,31,133,31,133,30,131,31,211,31,211,30,38,31,38,30,80,31,80,30,132,31,132,30,108,31,17,31,204,31,181,31,181,30,42,31,42,30,114,31,135,31,87,31,128,31,26,31,212,31,212,30,24,31,74,31,24,31,203,31,220,31,46,31,92,31,153,31,121,31,74,31,112,31,189,31,69,31,210,31,6,31,69,31,109,31,28,31,245,31,28,31,191,31,32,31,35,31,14,31,154,31,154,30,62,31,185,31,221,31,17,31,184,31,233,31,233,30,82,31,82,30,182,31,221,31,5,31,167,31,249,31,154,31,154,30,201,31,188,31,144,31,219,31,5,31,30,31,129,31,155,31,180,31,45,31,6,31,93,31,34,31,96,31,44,31,180,31,72,31,78,31,247,31,247,30,2,31,81,31,12,31,6,31,45,31,71,31,47,31,230,31,246,31,185,31,245,31,245,30,16,31,66,31,27,31,27,30,27,29,109,31,109,30,241,31,113,31,113,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
