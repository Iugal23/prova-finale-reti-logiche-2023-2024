-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 236;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,64,0,137,0,166,0,0,0,202,0,22,0,228,0,0,0,0,0,63,0,96,0,167,0,0,0,196,0,119,0,14,0,49,0,1,0,109,0,0,0,78,0,138,0,94,0,245,0,164,0,0,0,85,0,0,0,35,0,246,0,107,0,0,0,6,0,8,0,0,0,147,0,83,0,231,0,97,0,150,0,11,0,27,0,83,0,203,0,246,0,65,0,176,0,222,0,167,0,60,0,156,0,82,0,186,0,18,0,188,0,163,0,245,0,161,0,158,0,0,0,0,0,0,0,184,0,147,0,159,0,189,0,205,0,154,0,46,0,238,0,247,0,235,0,51,0,140,0,140,0,83,0,0,0,20,0,81,0,128,0,219,0,18,0,102,0,44,0,222,0,0,0,118,0,164,0,121,0,101,0,66,0,107,0,182,0,153,0,245,0,135,0,81,0,53,0,51,0,43,0,9,0,82,0,236,0,134,0,0,0,239,0,0,0,0,0,147,0,130,0,192,0,0,0,188,0,11,0,228,0,54,0,42,0,164,0,69,0,17,0,204,0,78,0,47,0,231,0,0,0,3,0,84,0,0,0,143,0,37,0,0,0,186,0,51,0,249,0,179,0,55,0,251,0,162,0,67,0,140,0,204,0,255,0,242,0,243,0,239,0,175,0,202,0,246,0,207,0,0,0,111,0,153,0,245,0,221,0,223,0,56,0,0,0,190,0,108,0,2,0,212,0,91,0,0,0,116,0,0,0,155,0,170,0,0,0,188,0,0,0,102,0,110,0,56,0,224,0,210,0,235,0,146,0,43,0,166,0,0,0,66,0,103,0,0,0,0,0,226,0,90,0,160,0,0,0,0,0,222,0,9,0,253,0,170,0,169,0,32,0,0,0,0,0,156,0,243,0,144,0,0,0,241,0,27,0,115,0,192,0,229,0,0,0,135,0,231,0,59,0,0,0,26,0,68,0,215,0,73,0,124,0,165,0,235,0,240,0,44,0,120,0,203,0,0,0,15,0,101,0,107,0,144,0,218,0,108,0,17,0,155,0,196,0,17,0,85,0,0,0);
signal scenario_full  : scenario_type := (134,31,64,31,137,31,166,31,166,30,202,31,22,31,228,31,228,30,228,29,63,31,96,31,167,31,167,30,196,31,119,31,14,31,49,31,1,31,109,31,109,30,78,31,138,31,94,31,245,31,164,31,164,30,85,31,85,30,35,31,246,31,107,31,107,30,6,31,8,31,8,30,147,31,83,31,231,31,97,31,150,31,11,31,27,31,83,31,203,31,246,31,65,31,176,31,222,31,167,31,60,31,156,31,82,31,186,31,18,31,188,31,163,31,245,31,161,31,158,31,158,30,158,29,158,28,184,31,147,31,159,31,189,31,205,31,154,31,46,31,238,31,247,31,235,31,51,31,140,31,140,31,83,31,83,30,20,31,81,31,128,31,219,31,18,31,102,31,44,31,222,31,222,30,118,31,164,31,121,31,101,31,66,31,107,31,182,31,153,31,245,31,135,31,81,31,53,31,51,31,43,31,9,31,82,31,236,31,134,31,134,30,239,31,239,30,239,29,147,31,130,31,192,31,192,30,188,31,11,31,228,31,54,31,42,31,164,31,69,31,17,31,204,31,78,31,47,31,231,31,231,30,3,31,84,31,84,30,143,31,37,31,37,30,186,31,51,31,249,31,179,31,55,31,251,31,162,31,67,31,140,31,204,31,255,31,242,31,243,31,239,31,175,31,202,31,246,31,207,31,207,30,111,31,153,31,245,31,221,31,223,31,56,31,56,30,190,31,108,31,2,31,212,31,91,31,91,30,116,31,116,30,155,31,170,31,170,30,188,31,188,30,102,31,110,31,56,31,224,31,210,31,235,31,146,31,43,31,166,31,166,30,66,31,103,31,103,30,103,29,226,31,90,31,160,31,160,30,160,29,222,31,9,31,253,31,170,31,169,31,32,31,32,30,32,29,156,31,243,31,144,31,144,30,241,31,27,31,115,31,192,31,229,31,229,30,135,31,231,31,59,31,59,30,26,31,68,31,215,31,73,31,124,31,165,31,235,31,240,31,44,31,120,31,203,31,203,30,15,31,101,31,107,31,144,31,218,31,108,31,17,31,155,31,196,31,17,31,85,31,85,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
