-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_585 is
end project_tb_585;

architecture project_tb_arch_585 of project_tb_585 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 414;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (53,0,42,0,0,0,41,0,239,0,205,0,0,0,12,0,199,0,154,0,83,0,50,0,109,0,0,0,202,0,94,0,202,0,0,0,207,0,74,0,153,0,196,0,115,0,0,0,49,0,0,0,201,0,136,0,45,0,0,0,129,0,157,0,0,0,175,0,50,0,66,0,50,0,60,0,60,0,171,0,82,0,248,0,123,0,103,0,105,0,0,0,107,0,0,0,172,0,220,0,241,0,0,0,198,0,33,0,26,0,154,0,69,0,111,0,35,0,167,0,116,0,0,0,66,0,187,0,0,0,193,0,130,0,113,0,48,0,234,0,194,0,0,0,0,0,22,0,0,0,111,0,0,0,143,0,167,0,49,0,253,0,198,0,0,0,222,0,34,0,236,0,65,0,153,0,0,0,37,0,221,0,208,0,0,0,145,0,96,0,133,0,224,0,169,0,96,0,53,0,218,0,79,0,246,0,236,0,3,0,215,0,235,0,203,0,228,0,244,0,85,0,72,0,14,0,72,0,0,0,14,0,0,0,0,0,204,0,125,0,227,0,169,0,118,0,166,0,0,0,230,0,159,0,3,0,161,0,146,0,231,0,0,0,32,0,163,0,234,0,49,0,147,0,48,0,17,0,80,0,242,0,155,0,8,0,147,0,233,0,176,0,0,0,0,0,137,0,118,0,115,0,0,0,0,0,36,0,98,0,0,0,0,0,187,0,185,0,14,0,200,0,175,0,239,0,214,0,57,0,180,0,122,0,255,0,0,0,165,0,0,0,0,0,97,0,213,0,189,0,37,0,246,0,211,0,58,0,92,0,212,0,197,0,126,0,161,0,140,0,180,0,21,0,14,0,41,0,21,0,0,0,133,0,158,0,74,0,81,0,0,0,168,0,180,0,241,0,0,0,0,0,73,0,25,0,35,0,0,0,28,0,0,0,23,0,234,0,152,0,250,0,191,0,19,0,0,0,0,0,125,0,0,0,148,0,144,0,104,0,243,0,111,0,78,0,122,0,0,0,109,0,81,0,13,0,64,0,242,0,8,0,91,0,202,0,32,0,178,0,221,0,54,0,218,0,210,0,248,0,2,0,222,0,144,0,232,0,198,0,105,0,112,0,171,0,30,0,137,0,220,0,0,0,55,0,35,0,0,0,0,0,144,0,0,0,217,0,201,0,89,0,59,0,171,0,13,0,227,0,157,0,0,0,62,0,23,0,241,0,0,0,197,0,156,0,196,0,103,0,87,0,226,0,199,0,122,0,148,0,0,0,75,0,96,0,13,0,0,0,134,0,235,0,44,0,0,0,77,0,73,0,60,0,0,0,235,0,84,0,6,0,14,0,114,0,129,0,0,0,24,0,0,0,213,0,122,0,154,0,250,0,152,0,73,0,0,0,126,0,60,0,88,0,126,0,18,0,132,0,236,0,105,0,129,0,51,0,120,0,171,0,167,0,0,0,85,0,206,0,25,0,156,0,17,0,184,0,157,0,39,0,248,0,0,0,0,0,227,0,25,0,0,0,94,0,221,0,167,0,40,0,217,0,70,0,165,0,212,0,0,0,0,0,230,0,126,0,100,0,91,0,245,0,142,0,196,0,32,0,28,0,0,0,185,0,226,0,37,0,84,0,116,0,254,0,115,0,184,0,0,0,0,0,11,0,150,0,121,0,97,0,95,0,203,0,46,0,13,0,30,0,8,0,187,0,236,0,59,0,0,0,0,0,0,0,0,0,52,0,72,0,25,0,0,0,216,0,0,0,112,0,9,0,255,0,157,0,243,0,233,0,0,0,98,0,92,0,0,0,0,0,57,0,0,0,223,0,185,0,76,0,220,0,56,0,1,0,36,0,64,0,0,0,0,0,95,0);
signal scenario_full  : scenario_type := (53,31,42,31,42,30,41,31,239,31,205,31,205,30,12,31,199,31,154,31,83,31,50,31,109,31,109,30,202,31,94,31,202,31,202,30,207,31,74,31,153,31,196,31,115,31,115,30,49,31,49,30,201,31,136,31,45,31,45,30,129,31,157,31,157,30,175,31,50,31,66,31,50,31,60,31,60,31,171,31,82,31,248,31,123,31,103,31,105,31,105,30,107,31,107,30,172,31,220,31,241,31,241,30,198,31,33,31,26,31,154,31,69,31,111,31,35,31,167,31,116,31,116,30,66,31,187,31,187,30,193,31,130,31,113,31,48,31,234,31,194,31,194,30,194,29,22,31,22,30,111,31,111,30,143,31,167,31,49,31,253,31,198,31,198,30,222,31,34,31,236,31,65,31,153,31,153,30,37,31,221,31,208,31,208,30,145,31,96,31,133,31,224,31,169,31,96,31,53,31,218,31,79,31,246,31,236,31,3,31,215,31,235,31,203,31,228,31,244,31,85,31,72,31,14,31,72,31,72,30,14,31,14,30,14,29,204,31,125,31,227,31,169,31,118,31,166,31,166,30,230,31,159,31,3,31,161,31,146,31,231,31,231,30,32,31,163,31,234,31,49,31,147,31,48,31,17,31,80,31,242,31,155,31,8,31,147,31,233,31,176,31,176,30,176,29,137,31,118,31,115,31,115,30,115,29,36,31,98,31,98,30,98,29,187,31,185,31,14,31,200,31,175,31,239,31,214,31,57,31,180,31,122,31,255,31,255,30,165,31,165,30,165,29,97,31,213,31,189,31,37,31,246,31,211,31,58,31,92,31,212,31,197,31,126,31,161,31,140,31,180,31,21,31,14,31,41,31,21,31,21,30,133,31,158,31,74,31,81,31,81,30,168,31,180,31,241,31,241,30,241,29,73,31,25,31,35,31,35,30,28,31,28,30,23,31,234,31,152,31,250,31,191,31,19,31,19,30,19,29,125,31,125,30,148,31,144,31,104,31,243,31,111,31,78,31,122,31,122,30,109,31,81,31,13,31,64,31,242,31,8,31,91,31,202,31,32,31,178,31,221,31,54,31,218,31,210,31,248,31,2,31,222,31,144,31,232,31,198,31,105,31,112,31,171,31,30,31,137,31,220,31,220,30,55,31,35,31,35,30,35,29,144,31,144,30,217,31,201,31,89,31,59,31,171,31,13,31,227,31,157,31,157,30,62,31,23,31,241,31,241,30,197,31,156,31,196,31,103,31,87,31,226,31,199,31,122,31,148,31,148,30,75,31,96,31,13,31,13,30,134,31,235,31,44,31,44,30,77,31,73,31,60,31,60,30,235,31,84,31,6,31,14,31,114,31,129,31,129,30,24,31,24,30,213,31,122,31,154,31,250,31,152,31,73,31,73,30,126,31,60,31,88,31,126,31,18,31,132,31,236,31,105,31,129,31,51,31,120,31,171,31,167,31,167,30,85,31,206,31,25,31,156,31,17,31,184,31,157,31,39,31,248,31,248,30,248,29,227,31,25,31,25,30,94,31,221,31,167,31,40,31,217,31,70,31,165,31,212,31,212,30,212,29,230,31,126,31,100,31,91,31,245,31,142,31,196,31,32,31,28,31,28,30,185,31,226,31,37,31,84,31,116,31,254,31,115,31,184,31,184,30,184,29,11,31,150,31,121,31,97,31,95,31,203,31,46,31,13,31,30,31,8,31,187,31,236,31,59,31,59,30,59,29,59,28,59,27,52,31,72,31,25,31,25,30,216,31,216,30,112,31,9,31,255,31,157,31,243,31,233,31,233,30,98,31,92,31,92,30,92,29,57,31,57,30,223,31,185,31,76,31,220,31,56,31,1,31,36,31,64,31,64,30,64,29,95,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
