-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_33 is
end project_tb_33;

architecture project_tb_arch_33 of project_tb_33 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 266;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (98,0,139,0,67,0,107,0,252,0,213,0,0,0,1,0,181,0,41,0,224,0,32,0,210,0,27,0,135,0,102,0,98,0,218,0,190,0,58,0,0,0,165,0,0,0,114,0,121,0,95,0,155,0,253,0,253,0,0,0,0,0,232,0,0,0,63,0,0,0,69,0,0,0,117,0,217,0,189,0,170,0,131,0,0,0,43,0,128,0,58,0,106,0,199,0,244,0,0,0,0,0,116,0,0,0,115,0,42,0,12,0,16,0,6,0,120,0,0,0,1,0,0,0,59,0,34,0,0,0,212,0,0,0,0,0,28,0,0,0,103,0,127,0,0,0,54,0,242,0,108,0,125,0,0,0,0,0,0,0,228,0,168,0,0,0,0,0,213,0,128,0,66,0,198,0,135,0,36,0,185,0,0,0,0,0,125,0,2,0,2,0,58,0,243,0,104,0,92,0,176,0,79,0,156,0,0,0,0,0,110,0,65,0,188,0,226,0,0,0,87,0,179,0,220,0,187,0,153,0,192,0,199,0,0,0,0,0,36,0,202,0,78,0,143,0,0,0,124,0,28,0,121,0,29,0,235,0,118,0,75,0,0,0,113,0,230,0,169,0,98,0,107,0,220,0,36,0,0,0,117,0,118,0,196,0,96,0,203,0,112,0,89,0,20,0,0,0,54,0,22,0,105,0,140,0,0,0,0,0,168,0,152,0,0,0,47,0,93,0,0,0,113,0,208,0,5,0,220,0,36,0,205,0,224,0,212,0,187,0,124,0,239,0,79,0,170,0,52,0,108,0,0,0,190,0,242,0,65,0,22,0,109,0,228,0,252,0,184,0,187,0,49,0,75,0,149,0,152,0,156,0,3,0,0,0,129,0,99,0,82,0,33,0,109,0,172,0,0,0,33,0,101,0,0,0,226,0,75,0,141,0,77,0,208,0,0,0,120,0,236,0,231,0,181,0,184,0,172,0,242,0,43,0,58,0,128,0,26,0,196,0,244,0,134,0,175,0,214,0,0,0,0,0,131,0,73,0,194,0,98,0,29,0,215,0,0,0,145,0,0,0,164,0,94,0,0,0,0,0,0,0,156,0,0,0,172,0,96,0,61,0,60,0,199,0,121,0,50,0,137,0,6,0,23,0,5,0,116,0,48,0,9,0,46,0,0,0,164,0,211,0,0,0,0,0,0,0,131,0,153,0);
signal scenario_full  : scenario_type := (98,31,139,31,67,31,107,31,252,31,213,31,213,30,1,31,181,31,41,31,224,31,32,31,210,31,27,31,135,31,102,31,98,31,218,31,190,31,58,31,58,30,165,31,165,30,114,31,121,31,95,31,155,31,253,31,253,31,253,30,253,29,232,31,232,30,63,31,63,30,69,31,69,30,117,31,217,31,189,31,170,31,131,31,131,30,43,31,128,31,58,31,106,31,199,31,244,31,244,30,244,29,116,31,116,30,115,31,42,31,12,31,16,31,6,31,120,31,120,30,1,31,1,30,59,31,34,31,34,30,212,31,212,30,212,29,28,31,28,30,103,31,127,31,127,30,54,31,242,31,108,31,125,31,125,30,125,29,125,28,228,31,168,31,168,30,168,29,213,31,128,31,66,31,198,31,135,31,36,31,185,31,185,30,185,29,125,31,2,31,2,31,58,31,243,31,104,31,92,31,176,31,79,31,156,31,156,30,156,29,110,31,65,31,188,31,226,31,226,30,87,31,179,31,220,31,187,31,153,31,192,31,199,31,199,30,199,29,36,31,202,31,78,31,143,31,143,30,124,31,28,31,121,31,29,31,235,31,118,31,75,31,75,30,113,31,230,31,169,31,98,31,107,31,220,31,36,31,36,30,117,31,118,31,196,31,96,31,203,31,112,31,89,31,20,31,20,30,54,31,22,31,105,31,140,31,140,30,140,29,168,31,152,31,152,30,47,31,93,31,93,30,113,31,208,31,5,31,220,31,36,31,205,31,224,31,212,31,187,31,124,31,239,31,79,31,170,31,52,31,108,31,108,30,190,31,242,31,65,31,22,31,109,31,228,31,252,31,184,31,187,31,49,31,75,31,149,31,152,31,156,31,3,31,3,30,129,31,99,31,82,31,33,31,109,31,172,31,172,30,33,31,101,31,101,30,226,31,75,31,141,31,77,31,208,31,208,30,120,31,236,31,231,31,181,31,184,31,172,31,242,31,43,31,58,31,128,31,26,31,196,31,244,31,134,31,175,31,214,31,214,30,214,29,131,31,73,31,194,31,98,31,29,31,215,31,215,30,145,31,145,30,164,31,94,31,94,30,94,29,94,28,156,31,156,30,172,31,96,31,61,31,60,31,199,31,121,31,50,31,137,31,6,31,23,31,5,31,116,31,48,31,9,31,46,31,46,30,164,31,211,31,211,30,211,29,211,28,131,31,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
