-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_662 is
end project_tb_662;

architecture project_tb_arch_662 of project_tb_662 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 439;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,61,0,151,0,69,0,112,0,170,0,97,0,0,0,246,0,28,0,222,0,0,0,186,0,220,0,82,0,219,0,55,0,223,0,54,0,179,0,249,0,53,0,0,0,105,0,237,0,0,0,191,0,104,0,100,0,0,0,62,0,59,0,82,0,245,0,5,0,107,0,252,0,153,0,0,0,105,0,180,0,86,0,172,0,62,0,160,0,254,0,0,0,218,0,180,0,0,0,0,0,0,0,0,0,0,0,120,0,47,0,61,0,67,0,168,0,255,0,151,0,104,0,20,0,169,0,61,0,51,0,40,0,203,0,0,0,0,0,32,0,242,0,0,0,185,0,35,0,243,0,121,0,239,0,101,0,38,0,237,0,30,0,12,0,208,0,12,0,238,0,0,0,79,0,243,0,38,0,0,0,25,0,0,0,0,0,56,0,4,0,76,0,160,0,0,0,154,0,178,0,29,0,0,0,46,0,124,0,63,0,172,0,0,0,131,0,56,0,221,0,125,0,83,0,55,0,145,0,0,0,4,0,198,0,218,0,4,0,252,0,158,0,139,0,44,0,54,0,142,0,207,0,0,0,192,0,136,0,189,0,155,0,71,0,33,0,214,0,128,0,99,0,211,0,191,0,0,0,28,0,0,0,69,0,102,0,213,0,0,0,0,0,137,0,0,0,0,0,78,0,172,0,183,0,244,0,122,0,0,0,192,0,179,0,65,0,2,0,0,0,131,0,15,0,158,0,0,0,224,0,10,0,0,0,143,0,236,0,0,0,223,0,139,0,173,0,95,0,226,0,151,0,119,0,0,0,106,0,135,0,119,0,67,0,0,0,44,0,150,0,149,0,0,0,212,0,0,0,111,0,121,0,227,0,0,0,248,0,2,0,172,0,221,0,0,0,152,0,27,0,220,0,82,0,0,0,230,0,234,0,81,0,241,0,141,0,159,0,19,0,21,0,243,0,0,0,123,0,0,0,211,0,137,0,0,0,251,0,62,0,214,0,0,0,94,0,0,0,237,0,0,0,59,0,48,0,86,0,35,0,0,0,78,0,229,0,0,0,0,0,0,0,4,0,167,0,88,0,243,0,126,0,99,0,232,0,232,0,0,0,56,0,132,0,184,0,72,0,0,0,23,0,131,0,129,0,243,0,47,0,0,0,157,0,0,0,69,0,0,0,58,0,93,0,245,0,0,0,148,0,0,0,0,0,250,0,0,0,175,0,0,0,160,0,0,0,253,0,0,0,182,0,236,0,0,0,0,0,197,0,63,0,84,0,70,0,33,0,8,0,0,0,106,0,198,0,6,0,0,0,27,0,156,0,143,0,208,0,52,0,0,0,168,0,71,0,27,0,84,0,0,0,222,0,1,0,218,0,192,0,0,0,0,0,73,0,0,0,15,0,101,0,188,0,94,0,143,0,51,0,180,0,89,0,100,0,0,0,200,0,217,0,54,0,148,0,243,0,80,0,149,0,165,0,118,0,0,0,44,0,15,0,239,0,57,0,129,0,0,0,108,0,34,0,0,0,9,0,244,0,108,0,8,0,174,0,148,0,1,0,187,0,121,0,20,0,60,0,80,0,0,0,92,0,246,0,0,0,87,0,143,0,100,0,25,0,83,0,0,0,61,0,228,0,1,0,113,0,0,0,81,0,0,0,8,0,97,0,0,0,165,0,132,0,0,0,150,0,93,0,205,0,0,0,121,0,87,0,0,0,0,0,0,0,0,0,0,0,70,0,48,0,0,0,0,0,162,0,0,0,12,0,109,0,0,0,232,0,68,0,220,0,97,0,0,0,0,0,163,0,161,0,0,0,204,0,0,0,123,0,0,0,100,0,129,0,0,0,178,0,123,0,0,0,0,0,0,0,188,0,69,0,65,0,121,0,0,0,25,0,229,0,0,0,216,0,180,0,151,0,24,0,238,0,0,0,90,0,141,0,66,0,246,0,0,0,126,0,1,0,0,0,0,0,124,0);
signal scenario_full  : scenario_type := (0,0,61,31,151,31,69,31,112,31,170,31,97,31,97,30,246,31,28,31,222,31,222,30,186,31,220,31,82,31,219,31,55,31,223,31,54,31,179,31,249,31,53,31,53,30,105,31,237,31,237,30,191,31,104,31,100,31,100,30,62,31,59,31,82,31,245,31,5,31,107,31,252,31,153,31,153,30,105,31,180,31,86,31,172,31,62,31,160,31,254,31,254,30,218,31,180,31,180,30,180,29,180,28,180,27,180,26,120,31,47,31,61,31,67,31,168,31,255,31,151,31,104,31,20,31,169,31,61,31,51,31,40,31,203,31,203,30,203,29,32,31,242,31,242,30,185,31,35,31,243,31,121,31,239,31,101,31,38,31,237,31,30,31,12,31,208,31,12,31,238,31,238,30,79,31,243,31,38,31,38,30,25,31,25,30,25,29,56,31,4,31,76,31,160,31,160,30,154,31,178,31,29,31,29,30,46,31,124,31,63,31,172,31,172,30,131,31,56,31,221,31,125,31,83,31,55,31,145,31,145,30,4,31,198,31,218,31,4,31,252,31,158,31,139,31,44,31,54,31,142,31,207,31,207,30,192,31,136,31,189,31,155,31,71,31,33,31,214,31,128,31,99,31,211,31,191,31,191,30,28,31,28,30,69,31,102,31,213,31,213,30,213,29,137,31,137,30,137,29,78,31,172,31,183,31,244,31,122,31,122,30,192,31,179,31,65,31,2,31,2,30,131,31,15,31,158,31,158,30,224,31,10,31,10,30,143,31,236,31,236,30,223,31,139,31,173,31,95,31,226,31,151,31,119,31,119,30,106,31,135,31,119,31,67,31,67,30,44,31,150,31,149,31,149,30,212,31,212,30,111,31,121,31,227,31,227,30,248,31,2,31,172,31,221,31,221,30,152,31,27,31,220,31,82,31,82,30,230,31,234,31,81,31,241,31,141,31,159,31,19,31,21,31,243,31,243,30,123,31,123,30,211,31,137,31,137,30,251,31,62,31,214,31,214,30,94,31,94,30,237,31,237,30,59,31,48,31,86,31,35,31,35,30,78,31,229,31,229,30,229,29,229,28,4,31,167,31,88,31,243,31,126,31,99,31,232,31,232,31,232,30,56,31,132,31,184,31,72,31,72,30,23,31,131,31,129,31,243,31,47,31,47,30,157,31,157,30,69,31,69,30,58,31,93,31,245,31,245,30,148,31,148,30,148,29,250,31,250,30,175,31,175,30,160,31,160,30,253,31,253,30,182,31,236,31,236,30,236,29,197,31,63,31,84,31,70,31,33,31,8,31,8,30,106,31,198,31,6,31,6,30,27,31,156,31,143,31,208,31,52,31,52,30,168,31,71,31,27,31,84,31,84,30,222,31,1,31,218,31,192,31,192,30,192,29,73,31,73,30,15,31,101,31,188,31,94,31,143,31,51,31,180,31,89,31,100,31,100,30,200,31,217,31,54,31,148,31,243,31,80,31,149,31,165,31,118,31,118,30,44,31,15,31,239,31,57,31,129,31,129,30,108,31,34,31,34,30,9,31,244,31,108,31,8,31,174,31,148,31,1,31,187,31,121,31,20,31,60,31,80,31,80,30,92,31,246,31,246,30,87,31,143,31,100,31,25,31,83,31,83,30,61,31,228,31,1,31,113,31,113,30,81,31,81,30,8,31,97,31,97,30,165,31,132,31,132,30,150,31,93,31,205,31,205,30,121,31,87,31,87,30,87,29,87,28,87,27,87,26,70,31,48,31,48,30,48,29,162,31,162,30,12,31,109,31,109,30,232,31,68,31,220,31,97,31,97,30,97,29,163,31,161,31,161,30,204,31,204,30,123,31,123,30,100,31,129,31,129,30,178,31,123,31,123,30,123,29,123,28,188,31,69,31,65,31,121,31,121,30,25,31,229,31,229,30,216,31,180,31,151,31,24,31,238,31,238,30,90,31,141,31,66,31,246,31,246,30,126,31,1,31,1,30,1,29,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
