-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 519;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (192,0,0,0,207,0,0,0,8,0,0,0,245,0,30,0,101,0,94,0,236,0,4,0,227,0,216,0,38,0,85,0,227,0,188,0,92,0,88,0,0,0,169,0,37,0,59,0,0,0,221,0,114,0,214,0,34,0,34,0,150,0,182,0,0,0,219,0,172,0,204,0,220,0,127,0,79,0,197,0,0,0,12,0,56,0,20,0,87,0,83,0,0,0,6,0,224,0,171,0,64,0,157,0,188,0,238,0,111,0,204,0,14,0,0,0,132,0,186,0,55,0,27,0,84,0,116,0,162,0,166,0,0,0,239,0,137,0,158,0,131,0,90,0,158,0,0,0,224,0,0,0,0,0,0,0,226,0,172,0,67,0,72,0,117,0,0,0,114,0,74,0,87,0,30,0,134,0,204,0,176,0,0,0,219,0,141,0,236,0,169,0,81,0,28,0,61,0,14,0,0,0,0,0,158,0,77,0,231,0,105,0,234,0,0,0,85,0,0,0,0,0,0,0,0,0,70,0,238,0,0,0,3,0,184,0,0,0,238,0,253,0,167,0,219,0,0,0,0,0,235,0,0,0,56,0,30,0,0,0,63,0,63,0,186,0,14,0,239,0,234,0,0,0,0,0,0,0,26,0,230,0,22,0,0,0,249,0,95,0,217,0,2,0,0,0,202,0,183,0,75,0,168,0,232,0,215,0,80,0,0,0,12,0,190,0,0,0,0,0,237,0,89,0,179,0,213,0,205,0,244,0,107,0,228,0,150,0,217,0,127,0,66,0,0,0,0,0,225,0,22,0,236,0,69,0,188,0,26,0,62,0,49,0,0,0,50,0,217,0,88,0,233,0,82,0,160,0,36,0,248,0,0,0,70,0,20,0,239,0,0,0,0,0,24,0,224,0,0,0,0,0,0,0,198,0,196,0,250,0,231,0,134,0,89,0,220,0,227,0,54,0,197,0,193,0,204,0,0,0,241,0,23,0,195,0,0,0,33,0,2,0,73,0,66,0,41,0,0,0,171,0,72,0,72,0,0,0,1,0,123,0,75,0,0,0,13,0,140,0,0,0,0,0,73,0,72,0,84,0,0,0,212,0,83,0,232,0,67,0,51,0,120,0,39,0,1,0,4,0,0,0,164,0,58,0,0,0,162,0,3,0,0,0,48,0,143,0,0,0,229,0,125,0,101,0,115,0,0,0,35,0,0,0,0,0,89,0,46,0,32,0,92,0,130,0,50,0,80,0,51,0,182,0,0,0,0,0,163,0,171,0,0,0,28,0,101,0,173,0,185,0,0,0,245,0,151,0,0,0,86,0,1,0,165,0,0,0,180,0,192,0,0,0,18,0,53,0,41,0,203,0,214,0,187,0,111,0,127,0,124,0,47,0,91,0,198,0,168,0,79,0,78,0,0,0,26,0,102,0,137,0,42,0,91,0,0,0,159,0,144,0,247,0,5,0,184,0,163,0,232,0,22,0,0,0,27,0,0,0,251,0,11,0,0,0,246,0,12,0,63,0,240,0,222,0,45,0,16,0,0,0,0,0,0,0,133,0,0,0,250,0,233,0,0,0,122,0,0,0,0,0,254,0,196,0,220,0,106,0,0,0,83,0,175,0,172,0,227,0,0,0,237,0,84,0,24,0,183,0,2,0,173,0,0,0,116,0,168,0,181,0,140,0,23,0,0,0,0,0,163,0,50,0,121,0,0,0,0,0,170,0,133,0,255,0,214,0,141,0,244,0,129,0,174,0,195,0,0,0,0,0,7,0,0,0,26,0,0,0,56,0,237,0,0,0,246,0,88,0,169,0,112,0,240,0,0,0,235,0,254,0,202,0,0,0,0,0,42,0,0,0,142,0,135,0,73,0,188,0,0,0,0,0,188,0,248,0,135,0,75,0,192,0,65,0,0,0,21,0,197,0,0,0,0,0,163,0,46,0,75,0,29,0,61,0,190,0,189,0,63,0,60,0,84,0,121,0,0,0,61,0,238,0,120,0,58,0,32,0,114,0,8,0,148,0,205,0,162,0,112,0,0,0,251,0,0,0,204,0,63,0,214,0,60,0,229,0,0,0,131,0,104,0,145,0,0,0,153,0,27,0,0,0,0,0,39,0,195,0,170,0,0,0,0,0,182,0,128,0,120,0,13,0,109,0,116,0,0,0,163,0,0,0,62,0,255,0,0,0,0,0,107,0,190,0,0,0,0,0,53,0,0,0,20,0,0,0,38,0,219,0,216,0,144,0,61,0,93,0,77,0,87,0,75,0,200,0,145,0,9,0,144,0,154,0,170,0,212,0,78,0,100,0,213,0,94,0,83,0,6,0,0,0,65,0,129,0);
signal scenario_full  : scenario_type := (192,31,192,30,207,31,207,30,8,31,8,30,245,31,30,31,101,31,94,31,236,31,4,31,227,31,216,31,38,31,85,31,227,31,188,31,92,31,88,31,88,30,169,31,37,31,59,31,59,30,221,31,114,31,214,31,34,31,34,31,150,31,182,31,182,30,219,31,172,31,204,31,220,31,127,31,79,31,197,31,197,30,12,31,56,31,20,31,87,31,83,31,83,30,6,31,224,31,171,31,64,31,157,31,188,31,238,31,111,31,204,31,14,31,14,30,132,31,186,31,55,31,27,31,84,31,116,31,162,31,166,31,166,30,239,31,137,31,158,31,131,31,90,31,158,31,158,30,224,31,224,30,224,29,224,28,226,31,172,31,67,31,72,31,117,31,117,30,114,31,74,31,87,31,30,31,134,31,204,31,176,31,176,30,219,31,141,31,236,31,169,31,81,31,28,31,61,31,14,31,14,30,14,29,158,31,77,31,231,31,105,31,234,31,234,30,85,31,85,30,85,29,85,28,85,27,70,31,238,31,238,30,3,31,184,31,184,30,238,31,253,31,167,31,219,31,219,30,219,29,235,31,235,30,56,31,30,31,30,30,63,31,63,31,186,31,14,31,239,31,234,31,234,30,234,29,234,28,26,31,230,31,22,31,22,30,249,31,95,31,217,31,2,31,2,30,202,31,183,31,75,31,168,31,232,31,215,31,80,31,80,30,12,31,190,31,190,30,190,29,237,31,89,31,179,31,213,31,205,31,244,31,107,31,228,31,150,31,217,31,127,31,66,31,66,30,66,29,225,31,22,31,236,31,69,31,188,31,26,31,62,31,49,31,49,30,50,31,217,31,88,31,233,31,82,31,160,31,36,31,248,31,248,30,70,31,20,31,239,31,239,30,239,29,24,31,224,31,224,30,224,29,224,28,198,31,196,31,250,31,231,31,134,31,89,31,220,31,227,31,54,31,197,31,193,31,204,31,204,30,241,31,23,31,195,31,195,30,33,31,2,31,73,31,66,31,41,31,41,30,171,31,72,31,72,31,72,30,1,31,123,31,75,31,75,30,13,31,140,31,140,30,140,29,73,31,72,31,84,31,84,30,212,31,83,31,232,31,67,31,51,31,120,31,39,31,1,31,4,31,4,30,164,31,58,31,58,30,162,31,3,31,3,30,48,31,143,31,143,30,229,31,125,31,101,31,115,31,115,30,35,31,35,30,35,29,89,31,46,31,32,31,92,31,130,31,50,31,80,31,51,31,182,31,182,30,182,29,163,31,171,31,171,30,28,31,101,31,173,31,185,31,185,30,245,31,151,31,151,30,86,31,1,31,165,31,165,30,180,31,192,31,192,30,18,31,53,31,41,31,203,31,214,31,187,31,111,31,127,31,124,31,47,31,91,31,198,31,168,31,79,31,78,31,78,30,26,31,102,31,137,31,42,31,91,31,91,30,159,31,144,31,247,31,5,31,184,31,163,31,232,31,22,31,22,30,27,31,27,30,251,31,11,31,11,30,246,31,12,31,63,31,240,31,222,31,45,31,16,31,16,30,16,29,16,28,133,31,133,30,250,31,233,31,233,30,122,31,122,30,122,29,254,31,196,31,220,31,106,31,106,30,83,31,175,31,172,31,227,31,227,30,237,31,84,31,24,31,183,31,2,31,173,31,173,30,116,31,168,31,181,31,140,31,23,31,23,30,23,29,163,31,50,31,121,31,121,30,121,29,170,31,133,31,255,31,214,31,141,31,244,31,129,31,174,31,195,31,195,30,195,29,7,31,7,30,26,31,26,30,56,31,237,31,237,30,246,31,88,31,169,31,112,31,240,31,240,30,235,31,254,31,202,31,202,30,202,29,42,31,42,30,142,31,135,31,73,31,188,31,188,30,188,29,188,31,248,31,135,31,75,31,192,31,65,31,65,30,21,31,197,31,197,30,197,29,163,31,46,31,75,31,29,31,61,31,190,31,189,31,63,31,60,31,84,31,121,31,121,30,61,31,238,31,120,31,58,31,32,31,114,31,8,31,148,31,205,31,162,31,112,31,112,30,251,31,251,30,204,31,63,31,214,31,60,31,229,31,229,30,131,31,104,31,145,31,145,30,153,31,27,31,27,30,27,29,39,31,195,31,170,31,170,30,170,29,182,31,128,31,120,31,13,31,109,31,116,31,116,30,163,31,163,30,62,31,255,31,255,30,255,29,107,31,190,31,190,30,190,29,53,31,53,30,20,31,20,30,38,31,219,31,216,31,144,31,61,31,93,31,77,31,87,31,75,31,200,31,145,31,9,31,144,31,154,31,170,31,212,31,78,31,100,31,213,31,94,31,83,31,6,31,6,30,65,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
