-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 753;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,196,0,32,0,181,0,31,0,248,0,232,0,0,0,0,0,0,0,0,0,0,0,0,0,112,0,33,0,38,0,22,0,44,0,15,0,0,0,45,0,19,0,184,0,188,0,0,0,153,0,97,0,30,0,0,0,61,0,1,0,81,0,83,0,0,0,144,0,59,0,102,0,153,0,179,0,17,0,69,0,215,0,0,0,0,0,0,0,166,0,130,0,240,0,252,0,135,0,84,0,80,0,7,0,87,0,96,0,117,0,75,0,29,0,42,0,176,0,175,0,101,0,136,0,44,0,86,0,213,0,232,0,45,0,69,0,232,0,30,0,28,0,172,0,25,0,0,0,58,0,239,0,105,0,217,0,0,0,125,0,0,0,35,0,102,0,30,0,249,0,18,0,18,0,91,0,89,0,61,0,124,0,0,0,11,0,123,0,107,0,137,0,128,0,176,0,32,0,141,0,32,0,0,0,109,0,39,0,252,0,246,0,90,0,203,0,198,0,236,0,3,0,159,0,79,0,219,0,203,0,96,0,237,0,0,0,137,0,0,0,24,0,0,0,5,0,0,0,0,0,82,0,54,0,107,0,1,0,50,0,0,0,44,0,91,0,224,0,58,0,165,0,162,0,0,0,88,0,37,0,85,0,27,0,64,0,194,0,220,0,59,0,36,0,101,0,248,0,0,0,0,0,0,0,96,0,83,0,33,0,26,0,177,0,46,0,0,0,241,0,232,0,100,0,160,0,0,0,91,0,212,0,0,0,155,0,208,0,98,0,229,0,0,0,27,0,0,0,65,0,0,0,252,0,100,0,166,0,0,0,183,0,188,0,141,0,0,0,216,0,137,0,136,0,0,0,124,0,92,0,218,0,219,0,5,0,241,0,34,0,110,0,238,0,0,0,86,0,181,0,219,0,134,0,28,0,153,0,194,0,51,0,131,0,233,0,146,0,0,0,109,0,28,0,205,0,0,0,68,0,6,0,51,0,0,0,0,0,0,0,191,0,127,0,0,0,0,0,47,0,231,0,179,0,171,0,233,0,222,0,158,0,144,0,84,0,157,0,54,0,99,0,185,0,185,0,226,0,58,0,35,0,174,0,181,0,249,0,205,0,185,0,7,0,10,0,0,0,1,0,87,0,76,0,131,0,194,0,198,0,6,0,53,0,57,0,233,0,83,0,221,0,197,0,89,0,0,0,84,0,240,0,186,0,227,0,0,0,14,0,209,0,253,0,10,0,66,0,226,0,232,0,0,0,0,0,172,0,151,0,86,0,37,0,99,0,28,0,166,0,0,0,0,0,19,0,0,0,48,0,94,0,164,0,66,0,188,0,120,0,210,0,198,0,0,0,0,0,241,0,243,0,228,0,211,0,163,0,130,0,0,0,150,0,69,0,203,0,247,0,130,0,140,0,0,0,2,0,20,0,88,0,158,0,107,0,17,0,79,0,160,0,25,0,0,0,85,0,240,0,233,0,0,0,0,0,0,0,222,0,97,0,0,0,140,0,222,0,101,0,73,0,236,0,80,0,110,0,23,0,182,0,245,0,0,0,102,0,0,0,0,0,129,0,230,0,96,0,0,0,0,0,160,0,0,0,0,0,100,0,82,0,216,0,196,0,129,0,182,0,248,0,218,0,5,0,194,0,60,0,226,0,37,0,98,0,237,0,0,0,140,0,20,0,172,0,124,0,167,0,135,0,74,0,1,0,248,0,62,0,32,0,123,0,252,0,0,0,0,0,8,0,45,0,90,0,26,0,142,0,125,0,84,0,0,0,190,0,0,0,16,0,0,0,117,0,179,0,193,0,144,0,6,0,153,0,112,0,176,0,122,0,0,0,42,0,0,0,0,0,222,0,172,0,30,0,106,0,82,0,3,0,213,0,52,0,243,0,0,0,27,0,0,0,177,0,0,0,105,0,18,0,250,0,4,0,29,0,0,0,63,0,213,0,0,0,116,0,31,0,118,0,123,0,145,0,219,0,0,0,69,0,107,0,230,0,89,0,227,0,0,0,18,0,107,0,0,0,220,0,76,0,116,0,78,0,58,0,33,0,176,0,12,0,78,0,0,0,168,0,175,0,103,0,43,0,0,0,124,0,77,0,59,0,158,0,107,0,0,0,218,0,125,0,189,0,198,0,0,0,0,0,94,0,13,0,199,0,12,0,72,0,50,0,76,0,161,0,65,0,0,0,159,0,0,0,216,0,183,0,46,0,0,0,131,0,146,0,0,0,20,0,104,0,123,0,174,0,0,0,44,0,26,0,110,0,0,0,0,0,195,0,200,0,155,0,150,0,152,0,110,0,242,0,195,0,251,0,0,0,253,0,220,0,0,0,28,0,11,0,0,0,140,0,0,0,171,0,185,0,161,0,0,0,163,0,0,0,128,0,29,0,146,0,206,0,0,0,94,0,8,0,101,0,0,0,165,0,195,0,172,0,150,0,0,0,119,0,144,0,188,0,75,0,35,0,37,0,216,0,75,0,202,0,189,0,40,0,120,0,252,0,238,0,171,0,238,0,107,0,32,0,0,0,0,0,154,0,72,0,246,0,15,0,190,0,200,0,0,0,0,0,138,0,168,0,130,0,149,0,50,0,167,0,120,0,247,0,0,0,0,0,71,0,0,0,36,0,112,0,101,0,177,0,156,0,0,0,195,0,238,0,203,0,183,0,0,0,0,0,0,0,0,0,252,0,123,0,219,0,153,0,215,0,209,0,10,0,153,0,132,0,239,0,85,0,218,0,103,0,0,0,242,0,240,0,33,0,194,0,118,0,13,0,0,0,241,0,163,0,114,0,0,0,107,0,0,0,232,0,143,0,173,0,107,0,97,0,137,0,0,0,115,0,190,0,41,0,68,0,12,0,112,0,76,0,174,0,84,0,212,0,90,0,120,0,234,0,233,0,157,0,73,0,237,0,120,0,0,0,200,0,10,0,62,0,15,0,245,0,115,0,21,0,139,0,53,0,206,0,208,0,148,0,227,0,255,0,159,0,64,0,135,0,75,0,31,0,164,0,77,0,139,0,85,0,95,0,0,0,155,0,33,0,0,0,62,0,27,0,0,0,135,0,19,0,181,0,125,0,154,0,195,0,89,0,176,0,214,0,233,0,174,0,49,0,0,0,205,0,57,0,172,0,196,0,214,0,134,0,67,0,195,0,163,0,159,0,25,0,0,0,91,0,234,0,63,0,169,0,0,0,96,0,23,0,46,0,244,0,74,0,48,0,221,0,238,0,30,0,77,0,194,0,200,0,151,0,224,0,228,0,209,0,99,0,197,0,162,0,254,0,16,0,0,0,43,0,212,0,79,0,215,0,10,0,0,0,39,0,99,0,0,0,150,0,8,0,0,0,207,0,203,0,0,0,0,0,0,0,7,0,0,0);
signal scenario_full  : scenario_type := (0,0,196,31,32,31,181,31,31,31,248,31,232,31,232,30,232,29,232,28,232,27,232,26,232,25,112,31,33,31,38,31,22,31,44,31,15,31,15,30,45,31,19,31,184,31,188,31,188,30,153,31,97,31,30,31,30,30,61,31,1,31,81,31,83,31,83,30,144,31,59,31,102,31,153,31,179,31,17,31,69,31,215,31,215,30,215,29,215,28,166,31,130,31,240,31,252,31,135,31,84,31,80,31,7,31,87,31,96,31,117,31,75,31,29,31,42,31,176,31,175,31,101,31,136,31,44,31,86,31,213,31,232,31,45,31,69,31,232,31,30,31,28,31,172,31,25,31,25,30,58,31,239,31,105,31,217,31,217,30,125,31,125,30,35,31,102,31,30,31,249,31,18,31,18,31,91,31,89,31,61,31,124,31,124,30,11,31,123,31,107,31,137,31,128,31,176,31,32,31,141,31,32,31,32,30,109,31,39,31,252,31,246,31,90,31,203,31,198,31,236,31,3,31,159,31,79,31,219,31,203,31,96,31,237,31,237,30,137,31,137,30,24,31,24,30,5,31,5,30,5,29,82,31,54,31,107,31,1,31,50,31,50,30,44,31,91,31,224,31,58,31,165,31,162,31,162,30,88,31,37,31,85,31,27,31,64,31,194,31,220,31,59,31,36,31,101,31,248,31,248,30,248,29,248,28,96,31,83,31,33,31,26,31,177,31,46,31,46,30,241,31,232,31,100,31,160,31,160,30,91,31,212,31,212,30,155,31,208,31,98,31,229,31,229,30,27,31,27,30,65,31,65,30,252,31,100,31,166,31,166,30,183,31,188,31,141,31,141,30,216,31,137,31,136,31,136,30,124,31,92,31,218,31,219,31,5,31,241,31,34,31,110,31,238,31,238,30,86,31,181,31,219,31,134,31,28,31,153,31,194,31,51,31,131,31,233,31,146,31,146,30,109,31,28,31,205,31,205,30,68,31,6,31,51,31,51,30,51,29,51,28,191,31,127,31,127,30,127,29,47,31,231,31,179,31,171,31,233,31,222,31,158,31,144,31,84,31,157,31,54,31,99,31,185,31,185,31,226,31,58,31,35,31,174,31,181,31,249,31,205,31,185,31,7,31,10,31,10,30,1,31,87,31,76,31,131,31,194,31,198,31,6,31,53,31,57,31,233,31,83,31,221,31,197,31,89,31,89,30,84,31,240,31,186,31,227,31,227,30,14,31,209,31,253,31,10,31,66,31,226,31,232,31,232,30,232,29,172,31,151,31,86,31,37,31,99,31,28,31,166,31,166,30,166,29,19,31,19,30,48,31,94,31,164,31,66,31,188,31,120,31,210,31,198,31,198,30,198,29,241,31,243,31,228,31,211,31,163,31,130,31,130,30,150,31,69,31,203,31,247,31,130,31,140,31,140,30,2,31,20,31,88,31,158,31,107,31,17,31,79,31,160,31,25,31,25,30,85,31,240,31,233,31,233,30,233,29,233,28,222,31,97,31,97,30,140,31,222,31,101,31,73,31,236,31,80,31,110,31,23,31,182,31,245,31,245,30,102,31,102,30,102,29,129,31,230,31,96,31,96,30,96,29,160,31,160,30,160,29,100,31,82,31,216,31,196,31,129,31,182,31,248,31,218,31,5,31,194,31,60,31,226,31,37,31,98,31,237,31,237,30,140,31,20,31,172,31,124,31,167,31,135,31,74,31,1,31,248,31,62,31,32,31,123,31,252,31,252,30,252,29,8,31,45,31,90,31,26,31,142,31,125,31,84,31,84,30,190,31,190,30,16,31,16,30,117,31,179,31,193,31,144,31,6,31,153,31,112,31,176,31,122,31,122,30,42,31,42,30,42,29,222,31,172,31,30,31,106,31,82,31,3,31,213,31,52,31,243,31,243,30,27,31,27,30,177,31,177,30,105,31,18,31,250,31,4,31,29,31,29,30,63,31,213,31,213,30,116,31,31,31,118,31,123,31,145,31,219,31,219,30,69,31,107,31,230,31,89,31,227,31,227,30,18,31,107,31,107,30,220,31,76,31,116,31,78,31,58,31,33,31,176,31,12,31,78,31,78,30,168,31,175,31,103,31,43,31,43,30,124,31,77,31,59,31,158,31,107,31,107,30,218,31,125,31,189,31,198,31,198,30,198,29,94,31,13,31,199,31,12,31,72,31,50,31,76,31,161,31,65,31,65,30,159,31,159,30,216,31,183,31,46,31,46,30,131,31,146,31,146,30,20,31,104,31,123,31,174,31,174,30,44,31,26,31,110,31,110,30,110,29,195,31,200,31,155,31,150,31,152,31,110,31,242,31,195,31,251,31,251,30,253,31,220,31,220,30,28,31,11,31,11,30,140,31,140,30,171,31,185,31,161,31,161,30,163,31,163,30,128,31,29,31,146,31,206,31,206,30,94,31,8,31,101,31,101,30,165,31,195,31,172,31,150,31,150,30,119,31,144,31,188,31,75,31,35,31,37,31,216,31,75,31,202,31,189,31,40,31,120,31,252,31,238,31,171,31,238,31,107,31,32,31,32,30,32,29,154,31,72,31,246,31,15,31,190,31,200,31,200,30,200,29,138,31,168,31,130,31,149,31,50,31,167,31,120,31,247,31,247,30,247,29,71,31,71,30,36,31,112,31,101,31,177,31,156,31,156,30,195,31,238,31,203,31,183,31,183,30,183,29,183,28,183,27,252,31,123,31,219,31,153,31,215,31,209,31,10,31,153,31,132,31,239,31,85,31,218,31,103,31,103,30,242,31,240,31,33,31,194,31,118,31,13,31,13,30,241,31,163,31,114,31,114,30,107,31,107,30,232,31,143,31,173,31,107,31,97,31,137,31,137,30,115,31,190,31,41,31,68,31,12,31,112,31,76,31,174,31,84,31,212,31,90,31,120,31,234,31,233,31,157,31,73,31,237,31,120,31,120,30,200,31,10,31,62,31,15,31,245,31,115,31,21,31,139,31,53,31,206,31,208,31,148,31,227,31,255,31,159,31,64,31,135,31,75,31,31,31,164,31,77,31,139,31,85,31,95,31,95,30,155,31,33,31,33,30,62,31,27,31,27,30,135,31,19,31,181,31,125,31,154,31,195,31,89,31,176,31,214,31,233,31,174,31,49,31,49,30,205,31,57,31,172,31,196,31,214,31,134,31,67,31,195,31,163,31,159,31,25,31,25,30,91,31,234,31,63,31,169,31,169,30,96,31,23,31,46,31,244,31,74,31,48,31,221,31,238,31,30,31,77,31,194,31,200,31,151,31,224,31,228,31,209,31,99,31,197,31,162,31,254,31,16,31,16,30,43,31,212,31,79,31,215,31,10,31,10,30,39,31,99,31,99,30,150,31,8,31,8,30,207,31,203,31,203,30,203,29,203,28,7,31,7,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
