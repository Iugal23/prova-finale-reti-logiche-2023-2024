-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 197;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (54,0,173,0,0,0,60,0,0,0,0,0,30,0,229,0,142,0,229,0,54,0,0,0,0,0,36,0,185,0,153,0,191,0,216,0,13,0,0,0,53,0,0,0,140,0,0,0,93,0,152,0,149,0,113,0,207,0,30,0,159,0,22,0,0,0,158,0,234,0,127,0,113,0,0,0,7,0,140,0,0,0,178,0,0,0,74,0,225,0,236,0,0,0,0,0,17,0,0,0,94,0,166,0,0,0,28,0,0,0,219,0,167,0,0,0,39,0,151,0,95,0,162,0,28,0,228,0,253,0,0,0,43,0,0,0,114,0,182,0,155,0,0,0,127,0,202,0,61,0,218,0,66,0,121,0,82,0,23,0,174,0,12,0,142,0,0,0,169,0,200,0,81,0,0,0,230,0,5,0,0,0,245,0,150,0,9,0,55,0,0,0,86,0,0,0,10,0,209,0,0,0,0,0,251,0,202,0,206,0,114,0,199,0,206,0,0,0,69,0,208,0,38,0,153,0,0,0,122,0,73,0,42,0,87,0,0,0,0,0,245,0,0,0,21,0,135,0,92,0,0,0,0,0,23,0,160,0,0,0,72,0,0,0,127,0,102,0,211,0,192,0,38,0,205,0,166,0,0,0,89,0,0,0,220,0,0,0,152,0,28,0,78,0,0,0,183,0,11,0,182,0,0,0,246,0,162,0,70,0,96,0,69,0,228,0,28,0,118,0,80,0,189,0,242,0,198,0,123,0,178,0,64,0,15,0,0,0,162,0,223,0,200,0,158,0,0,0,209,0,180,0,50,0,208,0,43,0,11,0,41,0,216,0,191,0,30,0,124,0,149,0,0,0,53,0,219,0,200,0,69,0,202,0,169,0,249,0,203,0,0,0,174,0);
signal scenario_full  : scenario_type := (54,31,173,31,173,30,60,31,60,30,60,29,30,31,229,31,142,31,229,31,54,31,54,30,54,29,36,31,185,31,153,31,191,31,216,31,13,31,13,30,53,31,53,30,140,31,140,30,93,31,152,31,149,31,113,31,207,31,30,31,159,31,22,31,22,30,158,31,234,31,127,31,113,31,113,30,7,31,140,31,140,30,178,31,178,30,74,31,225,31,236,31,236,30,236,29,17,31,17,30,94,31,166,31,166,30,28,31,28,30,219,31,167,31,167,30,39,31,151,31,95,31,162,31,28,31,228,31,253,31,253,30,43,31,43,30,114,31,182,31,155,31,155,30,127,31,202,31,61,31,218,31,66,31,121,31,82,31,23,31,174,31,12,31,142,31,142,30,169,31,200,31,81,31,81,30,230,31,5,31,5,30,245,31,150,31,9,31,55,31,55,30,86,31,86,30,10,31,209,31,209,30,209,29,251,31,202,31,206,31,114,31,199,31,206,31,206,30,69,31,208,31,38,31,153,31,153,30,122,31,73,31,42,31,87,31,87,30,87,29,245,31,245,30,21,31,135,31,92,31,92,30,92,29,23,31,160,31,160,30,72,31,72,30,127,31,102,31,211,31,192,31,38,31,205,31,166,31,166,30,89,31,89,30,220,31,220,30,152,31,28,31,78,31,78,30,183,31,11,31,182,31,182,30,246,31,162,31,70,31,96,31,69,31,228,31,28,31,118,31,80,31,189,31,242,31,198,31,123,31,178,31,64,31,15,31,15,30,162,31,223,31,200,31,158,31,158,30,209,31,180,31,50,31,208,31,43,31,11,31,41,31,216,31,191,31,30,31,124,31,149,31,149,30,53,31,219,31,200,31,69,31,202,31,169,31,249,31,203,31,203,30,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
