-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 166;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,230,0,182,0,14,0,179,0,220,0,229,0,131,0,138,0,210,0,0,0,160,0,90,0,252,0,0,0,81,0,204,0,41,0,84,0,235,0,252,0,84,0,236,0,244,0,219,0,71,0,104,0,14,0,47,0,217,0,143,0,242,0,131,0,170,0,0,0,203,0,254,0,13,0,46,0,15,0,51,0,3,0,20,0,82,0,46,0,94,0,188,0,37,0,121,0,137,0,181,0,0,0,195,0,0,0,107,0,99,0,58,0,44,0,201,0,195,0,243,0,0,0,23,0,45,0,139,0,87,0,44,0,254,0,0,0,74,0,0,0,231,0,214,0,0,0,152,0,75,0,249,0,45,0,252,0,90,0,195,0,43,0,86,0,221,0,150,0,0,0,0,0,0,0,186,0,164,0,5,0,152,0,236,0,43,0,35,0,10,0,32,0,225,0,162,0,0,0,183,0,188,0,153,0,247,0,0,0,17,0,170,0,0,0,0,0,220,0,112,0,43,0,108,0,86,0,134,0,0,0,38,0,139,0,50,0,0,0,0,0,241,0,117,0,0,0,242,0,27,0,0,0,180,0,0,0,0,0,96,0,0,0,142,0,178,0,0,0,3,0,0,0,145,0,164,0,28,0,233,0,236,0,205,0,193,0,3,0,0,0,115,0,212,0,202,0,94,0,64,0,197,0,156,0,32,0,38,0,41,0,181,0,117,0,87,0,206,0,253,0,23,0,129,0,40,0,232,0,208,0);
signal scenario_full  : scenario_type := (34,31,230,31,182,31,14,31,179,31,220,31,229,31,131,31,138,31,210,31,210,30,160,31,90,31,252,31,252,30,81,31,204,31,41,31,84,31,235,31,252,31,84,31,236,31,244,31,219,31,71,31,104,31,14,31,47,31,217,31,143,31,242,31,131,31,170,31,170,30,203,31,254,31,13,31,46,31,15,31,51,31,3,31,20,31,82,31,46,31,94,31,188,31,37,31,121,31,137,31,181,31,181,30,195,31,195,30,107,31,99,31,58,31,44,31,201,31,195,31,243,31,243,30,23,31,45,31,139,31,87,31,44,31,254,31,254,30,74,31,74,30,231,31,214,31,214,30,152,31,75,31,249,31,45,31,252,31,90,31,195,31,43,31,86,31,221,31,150,31,150,30,150,29,150,28,186,31,164,31,5,31,152,31,236,31,43,31,35,31,10,31,32,31,225,31,162,31,162,30,183,31,188,31,153,31,247,31,247,30,17,31,170,31,170,30,170,29,220,31,112,31,43,31,108,31,86,31,134,31,134,30,38,31,139,31,50,31,50,30,50,29,241,31,117,31,117,30,242,31,27,31,27,30,180,31,180,30,180,29,96,31,96,30,142,31,178,31,178,30,3,31,3,30,145,31,164,31,28,31,233,31,236,31,205,31,193,31,3,31,3,30,115,31,212,31,202,31,94,31,64,31,197,31,156,31,32,31,38,31,41,31,181,31,117,31,87,31,206,31,253,31,23,31,129,31,40,31,232,31,208,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
