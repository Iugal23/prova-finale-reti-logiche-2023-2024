-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 321;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,188,0,86,0,43,0,53,0,146,0,237,0,134,0,91,0,206,0,47,0,38,0,7,0,240,0,186,0,228,0,53,0,126,0,245,0,0,0,67,0,123,0,0,0,213,0,131,0,148,0,13,0,176,0,0,0,88,0,61,0,0,0,197,0,109,0,195,0,146,0,44,0,0,0,0,0,250,0,39,0,149,0,0,0,116,0,0,0,198,0,56,0,186,0,56,0,182,0,77,0,143,0,67,0,0,0,177,0,92,0,0,0,159,0,105,0,233,0,102,0,167,0,38,0,167,0,0,0,188,0,12,0,0,0,0,0,0,0,190,0,70,0,96,0,0,0,181,0,93,0,67,0,104,0,9,0,246,0,0,0,119,0,196,0,17,0,125,0,7,0,0,0,44,0,240,0,79,0,158,0,104,0,0,0,228,0,4,0,47,0,100,0,85,0,207,0,231,0,42,0,31,0,67,0,167,0,235,0,203,0,81,0,204,0,157,0,48,0,115,0,14,0,34,0,222,0,28,0,109,0,73,0,0,0,199,0,72,0,0,0,94,0,66,0,88,0,153,0,0,0,188,0,134,0,227,0,0,0,173,0,147,0,0,0,92,0,239,0,5,0,254,0,209,0,247,0,50,0,11,0,193,0,94,0,230,0,134,0,84,0,139,0,153,0,0,0,243,0,242,0,0,0,0,0,205,0,229,0,173,0,104,0,34,0,245,0,6,0,45,0,0,0,158,0,164,0,46,0,0,0,129,0,49,0,129,0,224,0,0,0,68,0,234,0,118,0,224,0,118,0,241,0,195,0,83,0,107,0,228,0,55,0,185,0,115,0,201,0,8,0,231,0,136,0,13,0,127,0,119,0,105,0,229,0,101,0,160,0,4,0,219,0,0,0,89,0,238,0,211,0,93,0,0,0,42,0,0,0,0,0,0,0,0,0,156,0,0,0,206,0,0,0,0,0,180,0,0,0,27,0,133,0,167,0,157,0,9,0,0,0,0,0,0,0,148,0,94,0,220,0,235,0,0,0,98,0,91,0,230,0,188,0,8,0,216,0,251,0,106,0,101,0,56,0,212,0,0,0,0,0,38,0,106,0,162,0,86,0,198,0,182,0,0,0,74,0,14,0,0,0,0,0,0,0,188,0,250,0,205,0,82,0,200,0,121,0,56,0,217,0,101,0,131,0,0,0,0,0,231,0,249,0,198,0,103,0,98,0,0,0,157,0,149,0,188,0,134,0,50,0,201,0,166,0,0,0,235,0,183,0,233,0,252,0,21,0,11,0,0,0,202,0,116,0,181,0,132,0,190,0,144,0,0,0,84,0,167,0,0,0,13,0,2,0,0,0,0,0,0,0,27,0,81,0,0,0,0,0,0,0,141,0,0,0,0,0,0,0,120,0,245,0,253,0,194,0,199,0,0,0,225,0,0,0,151,0,0,0,0,0);
signal scenario_full  : scenario_type := (232,31,188,31,86,31,43,31,53,31,146,31,237,31,134,31,91,31,206,31,47,31,38,31,7,31,240,31,186,31,228,31,53,31,126,31,245,31,245,30,67,31,123,31,123,30,213,31,131,31,148,31,13,31,176,31,176,30,88,31,61,31,61,30,197,31,109,31,195,31,146,31,44,31,44,30,44,29,250,31,39,31,149,31,149,30,116,31,116,30,198,31,56,31,186,31,56,31,182,31,77,31,143,31,67,31,67,30,177,31,92,31,92,30,159,31,105,31,233,31,102,31,167,31,38,31,167,31,167,30,188,31,12,31,12,30,12,29,12,28,190,31,70,31,96,31,96,30,181,31,93,31,67,31,104,31,9,31,246,31,246,30,119,31,196,31,17,31,125,31,7,31,7,30,44,31,240,31,79,31,158,31,104,31,104,30,228,31,4,31,47,31,100,31,85,31,207,31,231,31,42,31,31,31,67,31,167,31,235,31,203,31,81,31,204,31,157,31,48,31,115,31,14,31,34,31,222,31,28,31,109,31,73,31,73,30,199,31,72,31,72,30,94,31,66,31,88,31,153,31,153,30,188,31,134,31,227,31,227,30,173,31,147,31,147,30,92,31,239,31,5,31,254,31,209,31,247,31,50,31,11,31,193,31,94,31,230,31,134,31,84,31,139,31,153,31,153,30,243,31,242,31,242,30,242,29,205,31,229,31,173,31,104,31,34,31,245,31,6,31,45,31,45,30,158,31,164,31,46,31,46,30,129,31,49,31,129,31,224,31,224,30,68,31,234,31,118,31,224,31,118,31,241,31,195,31,83,31,107,31,228,31,55,31,185,31,115,31,201,31,8,31,231,31,136,31,13,31,127,31,119,31,105,31,229,31,101,31,160,31,4,31,219,31,219,30,89,31,238,31,211,31,93,31,93,30,42,31,42,30,42,29,42,28,42,27,156,31,156,30,206,31,206,30,206,29,180,31,180,30,27,31,133,31,167,31,157,31,9,31,9,30,9,29,9,28,148,31,94,31,220,31,235,31,235,30,98,31,91,31,230,31,188,31,8,31,216,31,251,31,106,31,101,31,56,31,212,31,212,30,212,29,38,31,106,31,162,31,86,31,198,31,182,31,182,30,74,31,14,31,14,30,14,29,14,28,188,31,250,31,205,31,82,31,200,31,121,31,56,31,217,31,101,31,131,31,131,30,131,29,231,31,249,31,198,31,103,31,98,31,98,30,157,31,149,31,188,31,134,31,50,31,201,31,166,31,166,30,235,31,183,31,233,31,252,31,21,31,11,31,11,30,202,31,116,31,181,31,132,31,190,31,144,31,144,30,84,31,167,31,167,30,13,31,2,31,2,30,2,29,2,28,27,31,81,31,81,30,81,29,81,28,141,31,141,30,141,29,141,28,120,31,245,31,253,31,194,31,199,31,199,30,225,31,225,30,151,31,151,30,151,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
