-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_411 is
end project_tb_411;

architecture project_tb_arch_411 of project_tb_411 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 271;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,176,0,242,0,0,0,63,0,210,0,3,0,66,0,176,0,54,0,127,0,204,0,0,0,204,0,0,0,1,0,144,0,13,0,0,0,54,0,61,0,178,0,0,0,108,0,8,0,87,0,165,0,190,0,0,0,183,0,58,0,0,0,112,0,208,0,0,0,0,0,137,0,17,0,207,0,189,0,236,0,43,0,254,0,32,0,0,0,0,0,48,0,244,0,4,0,202,0,24,0,215,0,255,0,0,0,44,0,123,0,0,0,237,0,24,0,57,0,142,0,19,0,172,0,8,0,62,0,47,0,0,0,16,0,211,0,0,0,0,0,213,0,203,0,0,0,236,0,0,0,249,0,222,0,166,0,0,0,52,0,199,0,0,0,0,0,135,0,22,0,236,0,126,0,0,0,45,0,247,0,1,0,12,0,41,0,1,0,103,0,22,0,0,0,0,0,228,0,187,0,166,0,145,0,126,0,21,0,250,0,0,0,120,0,0,0,20,0,40,0,160,0,199,0,192,0,36,0,151,0,87,0,55,0,194,0,0,0,4,0,217,0,27,0,122,0,157,0,85,0,243,0,0,0,72,0,193,0,151,0,81,0,226,0,0,0,0,0,240,0,129,0,229,0,76,0,11,0,226,0,191,0,118,0,44,0,237,0,105,0,79,0,0,0,19,0,41,0,74,0,0,0,90,0,170,0,207,0,13,0,146,0,142,0,0,0,0,0,51,0,198,0,8,0,0,0,194,0,87,0,125,0,0,0,0,0,70,0,36,0,148,0,242,0,204,0,0,0,74,0,68,0,51,0,192,0,107,0,0,0,148,0,190,0,199,0,15,0,119,0,25,0,61,0,59,0,44,0,205,0,181,0,0,0,120,0,0,0,95,0,18,0,0,0,87,0,241,0,53,0,88,0,188,0,53,0,47,0,0,0,159,0,92,0,218,0,13,0,46,0,39,0,79,0,44,0,0,0,44,0,182,0,113,0,86,0,218,0,83,0,44,0,216,0,53,0,0,0,253,0,50,0,53,0,160,0,67,0,181,0,175,0,151,0,93,0,63,0,230,0,97,0,53,0,254,0,211,0,197,0,0,0,0,0,252,0,39,0,11,0,0,0,243,0,254,0,0,0,8,0,142,0,185,0,11,0,106,0,249,0,231,0,205,0,251,0,242,0,107,0,252,0,44,0,188,0,4,0,0,0,0,0,0,0,0,0,0,0,60,0);
signal scenario_full  : scenario_type := (0,0,176,31,242,31,242,30,63,31,210,31,3,31,66,31,176,31,54,31,127,31,204,31,204,30,204,31,204,30,1,31,144,31,13,31,13,30,54,31,61,31,178,31,178,30,108,31,8,31,87,31,165,31,190,31,190,30,183,31,58,31,58,30,112,31,208,31,208,30,208,29,137,31,17,31,207,31,189,31,236,31,43,31,254,31,32,31,32,30,32,29,48,31,244,31,4,31,202,31,24,31,215,31,255,31,255,30,44,31,123,31,123,30,237,31,24,31,57,31,142,31,19,31,172,31,8,31,62,31,47,31,47,30,16,31,211,31,211,30,211,29,213,31,203,31,203,30,236,31,236,30,249,31,222,31,166,31,166,30,52,31,199,31,199,30,199,29,135,31,22,31,236,31,126,31,126,30,45,31,247,31,1,31,12,31,41,31,1,31,103,31,22,31,22,30,22,29,228,31,187,31,166,31,145,31,126,31,21,31,250,31,250,30,120,31,120,30,20,31,40,31,160,31,199,31,192,31,36,31,151,31,87,31,55,31,194,31,194,30,4,31,217,31,27,31,122,31,157,31,85,31,243,31,243,30,72,31,193,31,151,31,81,31,226,31,226,30,226,29,240,31,129,31,229,31,76,31,11,31,226,31,191,31,118,31,44,31,237,31,105,31,79,31,79,30,19,31,41,31,74,31,74,30,90,31,170,31,207,31,13,31,146,31,142,31,142,30,142,29,51,31,198,31,8,31,8,30,194,31,87,31,125,31,125,30,125,29,70,31,36,31,148,31,242,31,204,31,204,30,74,31,68,31,51,31,192,31,107,31,107,30,148,31,190,31,199,31,15,31,119,31,25,31,61,31,59,31,44,31,205,31,181,31,181,30,120,31,120,30,95,31,18,31,18,30,87,31,241,31,53,31,88,31,188,31,53,31,47,31,47,30,159,31,92,31,218,31,13,31,46,31,39,31,79,31,44,31,44,30,44,31,182,31,113,31,86,31,218,31,83,31,44,31,216,31,53,31,53,30,253,31,50,31,53,31,160,31,67,31,181,31,175,31,151,31,93,31,63,31,230,31,97,31,53,31,254,31,211,31,197,31,197,30,197,29,252,31,39,31,11,31,11,30,243,31,254,31,254,30,8,31,142,31,185,31,11,31,106,31,249,31,231,31,205,31,251,31,242,31,107,31,252,31,44,31,188,31,4,31,4,30,4,29,4,28,4,27,4,26,60,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
