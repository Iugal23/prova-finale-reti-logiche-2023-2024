-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 637;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,51,0,129,0,52,0,218,0,83,0,122,0,255,0,0,0,239,0,76,0,124,0,0,0,46,0,81,0,204,0,222,0,0,0,22,0,189,0,166,0,65,0,62,0,199,0,0,0,41,0,41,0,23,0,244,0,196,0,134,0,0,0,17,0,0,0,0,0,0,0,0,0,214,0,192,0,108,0,29,0,148,0,170,0,205,0,114,0,104,0,224,0,145,0,100,0,220,0,193,0,132,0,62,0,4,0,70,0,55,0,0,0,50,0,20,0,0,0,178,0,153,0,0,0,146,0,170,0,6,0,0,0,30,0,28,0,16,0,0,0,134,0,0,0,16,0,188,0,138,0,120,0,55,0,251,0,84,0,0,0,245,0,55,0,98,0,61,0,88,0,179,0,145,0,241,0,0,0,0,0,237,0,180,0,56,0,0,0,5,0,139,0,0,0,0,0,197,0,158,0,206,0,136,0,167,0,161,0,51,0,114,0,0,0,69,0,47,0,83,0,30,0,129,0,0,0,46,0,0,0,87,0,249,0,161,0,36,0,53,0,51,0,121,0,0,0,158,0,83,0,194,0,81,0,197,0,106,0,170,0,2,0,206,0,241,0,7,0,169,0,191,0,165,0,95,0,141,0,240,0,38,0,110,0,129,0,0,0,109,0,0,0,128,0,0,0,55,0,196,0,189,0,30,0,250,0,0,0,55,0,0,0,0,0,42,0,240,0,201,0,42,0,104,0,100,0,120,0,230,0,197,0,0,0,41,0,162,0,133,0,29,0,167,0,86,0,48,0,175,0,0,0,115,0,134,0,85,0,251,0,12,0,91,0,191,0,236,0,0,0,212,0,141,0,99,0,164,0,72,0,177,0,203,0,165,0,45,0,183,0,0,0,0,0,195,0,17,0,5,0,10,0,0,0,0,0,120,0,0,0,0,0,84,0,0,0,73,0,58,0,74,0,0,0,157,0,0,0,171,0,0,0,135,0,39,0,212,0,0,0,88,0,10,0,0,0,64,0,74,0,79,0,27,0,0,0,11,0,0,0,0,0,55,0,255,0,86,0,0,0,106,0,45,0,136,0,182,0,17,0,255,0,36,0,248,0,216,0,0,0,0,0,0,0,125,0,211,0,0,0,246,0,182,0,20,0,186,0,0,0,70,0,0,0,252,0,135,0,0,0,144,0,0,0,0,0,80,0,0,0,109,0,9,0,25,0,0,0,19,0,51,0,134,0,103,0,0,0,70,0,132,0,0,0,183,0,173,0,130,0,50,0,0,0,0,0,183,0,83,0,230,0,134,0,240,0,228,0,29,0,205,0,107,0,101,0,0,0,173,0,0,0,26,0,55,0,19,0,108,0,222,0,52,0,235,0,234,0,60,0,155,0,167,0,78,0,78,0,241,0,152,0,230,0,55,0,180,0,9,0,63,0,67,0,105,0,56,0,0,0,198,0,8,0,0,0,184,0,0,0,0,0,127,0,10,0,186,0,92,0,142,0,133,0,79,0,160,0,84,0,46,0,28,0,173,0,0,0,134,0,147,0,95,0,94,0,179,0,109,0,71,0,0,0,58,0,0,0,82,0,0,0,5,0,69,0,201,0,25,0,0,0,105,0,110,0,53,0,149,0,159,0,0,0,2,0,171,0,195,0,177,0,166,0,40,0,28,0,80,0,21,0,179,0,30,0,150,0,138,0,44,0,0,0,8,0,229,0,0,0,220,0,132,0,0,0,0,0,26,0,0,0,4,0,239,0,116,0,170,0,0,0,90,0,105,0,84,0,70,0,110,0,118,0,151,0,0,0,27,0,41,0,251,0,0,0,169,0,50,0,141,0,203,0,222,0,117,0,97,0,146,0,0,0,209,0,22,0,170,0,0,0,154,0,204,0,252,0,206,0,0,0,139,0,0,0,231,0,171,0,128,0,249,0,118,0,30,0,70,0,0,0,0,0,238,0,194,0,12,0,136,0,138,0,0,0,26,0,157,0,49,0,0,0,232,0,41,0,0,0,243,0,106,0,116,0,82,0,62,0,46,0,104,0,228,0,149,0,27,0,62,0,213,0,11,0,168,0,108,0,149,0,223,0,98,0,166,0,98,0,57,0,123,0,168,0,89,0,150,0,56,0,183,0,32,0,246,0,69,0,205,0,18,0,189,0,0,0,204,0,0,0,0,0,252,0,72,0,165,0,235,0,0,0,161,0,18,0,0,0,183,0,94,0,176,0,0,0,183,0,28,0,249,0,141,0,18,0,0,0,207,0,221,0,235,0,128,0,66,0,59,0,38,0,0,0,0,0,111,0,0,0,151,0,0,0,221,0,58,0,0,0,198,0,22,0,223,0,149,0,57,0,142,0,0,0,232,0,0,0,119,0,253,0,213,0,201,0,64,0,241,0,96,0,177,0,188,0,243,0,9,0,85,0,230,0,187,0,124,0,0,0,174,0,0,0,178,0,177,0,1,0,0,0,90,0,42,0,64,0,159,0,0,0,0,0,245,0,108,0,102,0,0,0,104,0,84,0,113,0,69,0,181,0,0,0,32,0,179,0,207,0,194,0,245,0,101,0,0,0,59,0,0,0,158,0,108,0,0,0,209,0,209,0,204,0,0,0,0,0,0,0,239,0,16,0,224,0,81,0,9,0,0,0,16,0,205,0,243,0,30,0,46,0,0,0,20,0,88,0,42,0,0,0,0,0,97,0,148,0,36,0,0,0,173,0,234,0,64,0,237,0,99,0,81,0,226,0,183,0,188,0,93,0,0,0,13,0,38,0,51,0,86,0,252,0,114,0,0,0,8,0,241,0,139,0,123,0,103,0,91,0,165,0,28,0,88,0,67,0,158,0,9,0,98,0,0,0,167,0,0,0);
signal scenario_full  : scenario_type := (181,31,51,31,129,31,52,31,218,31,83,31,122,31,255,31,255,30,239,31,76,31,124,31,124,30,46,31,81,31,204,31,222,31,222,30,22,31,189,31,166,31,65,31,62,31,199,31,199,30,41,31,41,31,23,31,244,31,196,31,134,31,134,30,17,31,17,30,17,29,17,28,17,27,214,31,192,31,108,31,29,31,148,31,170,31,205,31,114,31,104,31,224,31,145,31,100,31,220,31,193,31,132,31,62,31,4,31,70,31,55,31,55,30,50,31,20,31,20,30,178,31,153,31,153,30,146,31,170,31,6,31,6,30,30,31,28,31,16,31,16,30,134,31,134,30,16,31,188,31,138,31,120,31,55,31,251,31,84,31,84,30,245,31,55,31,98,31,61,31,88,31,179,31,145,31,241,31,241,30,241,29,237,31,180,31,56,31,56,30,5,31,139,31,139,30,139,29,197,31,158,31,206,31,136,31,167,31,161,31,51,31,114,31,114,30,69,31,47,31,83,31,30,31,129,31,129,30,46,31,46,30,87,31,249,31,161,31,36,31,53,31,51,31,121,31,121,30,158,31,83,31,194,31,81,31,197,31,106,31,170,31,2,31,206,31,241,31,7,31,169,31,191,31,165,31,95,31,141,31,240,31,38,31,110,31,129,31,129,30,109,31,109,30,128,31,128,30,55,31,196,31,189,31,30,31,250,31,250,30,55,31,55,30,55,29,42,31,240,31,201,31,42,31,104,31,100,31,120,31,230,31,197,31,197,30,41,31,162,31,133,31,29,31,167,31,86,31,48,31,175,31,175,30,115,31,134,31,85,31,251,31,12,31,91,31,191,31,236,31,236,30,212,31,141,31,99,31,164,31,72,31,177,31,203,31,165,31,45,31,183,31,183,30,183,29,195,31,17,31,5,31,10,31,10,30,10,29,120,31,120,30,120,29,84,31,84,30,73,31,58,31,74,31,74,30,157,31,157,30,171,31,171,30,135,31,39,31,212,31,212,30,88,31,10,31,10,30,64,31,74,31,79,31,27,31,27,30,11,31,11,30,11,29,55,31,255,31,86,31,86,30,106,31,45,31,136,31,182,31,17,31,255,31,36,31,248,31,216,31,216,30,216,29,216,28,125,31,211,31,211,30,246,31,182,31,20,31,186,31,186,30,70,31,70,30,252,31,135,31,135,30,144,31,144,30,144,29,80,31,80,30,109,31,9,31,25,31,25,30,19,31,51,31,134,31,103,31,103,30,70,31,132,31,132,30,183,31,173,31,130,31,50,31,50,30,50,29,183,31,83,31,230,31,134,31,240,31,228,31,29,31,205,31,107,31,101,31,101,30,173,31,173,30,26,31,55,31,19,31,108,31,222,31,52,31,235,31,234,31,60,31,155,31,167,31,78,31,78,31,241,31,152,31,230,31,55,31,180,31,9,31,63,31,67,31,105,31,56,31,56,30,198,31,8,31,8,30,184,31,184,30,184,29,127,31,10,31,186,31,92,31,142,31,133,31,79,31,160,31,84,31,46,31,28,31,173,31,173,30,134,31,147,31,95,31,94,31,179,31,109,31,71,31,71,30,58,31,58,30,82,31,82,30,5,31,69,31,201,31,25,31,25,30,105,31,110,31,53,31,149,31,159,31,159,30,2,31,171,31,195,31,177,31,166,31,40,31,28,31,80,31,21,31,179,31,30,31,150,31,138,31,44,31,44,30,8,31,229,31,229,30,220,31,132,31,132,30,132,29,26,31,26,30,4,31,239,31,116,31,170,31,170,30,90,31,105,31,84,31,70,31,110,31,118,31,151,31,151,30,27,31,41,31,251,31,251,30,169,31,50,31,141,31,203,31,222,31,117,31,97,31,146,31,146,30,209,31,22,31,170,31,170,30,154,31,204,31,252,31,206,31,206,30,139,31,139,30,231,31,171,31,128,31,249,31,118,31,30,31,70,31,70,30,70,29,238,31,194,31,12,31,136,31,138,31,138,30,26,31,157,31,49,31,49,30,232,31,41,31,41,30,243,31,106,31,116,31,82,31,62,31,46,31,104,31,228,31,149,31,27,31,62,31,213,31,11,31,168,31,108,31,149,31,223,31,98,31,166,31,98,31,57,31,123,31,168,31,89,31,150,31,56,31,183,31,32,31,246,31,69,31,205,31,18,31,189,31,189,30,204,31,204,30,204,29,252,31,72,31,165,31,235,31,235,30,161,31,18,31,18,30,183,31,94,31,176,31,176,30,183,31,28,31,249,31,141,31,18,31,18,30,207,31,221,31,235,31,128,31,66,31,59,31,38,31,38,30,38,29,111,31,111,30,151,31,151,30,221,31,58,31,58,30,198,31,22,31,223,31,149,31,57,31,142,31,142,30,232,31,232,30,119,31,253,31,213,31,201,31,64,31,241,31,96,31,177,31,188,31,243,31,9,31,85,31,230,31,187,31,124,31,124,30,174,31,174,30,178,31,177,31,1,31,1,30,90,31,42,31,64,31,159,31,159,30,159,29,245,31,108,31,102,31,102,30,104,31,84,31,113,31,69,31,181,31,181,30,32,31,179,31,207,31,194,31,245,31,101,31,101,30,59,31,59,30,158,31,108,31,108,30,209,31,209,31,204,31,204,30,204,29,204,28,239,31,16,31,224,31,81,31,9,31,9,30,16,31,205,31,243,31,30,31,46,31,46,30,20,31,88,31,42,31,42,30,42,29,97,31,148,31,36,31,36,30,173,31,234,31,64,31,237,31,99,31,81,31,226,31,183,31,188,31,93,31,93,30,13,31,38,31,51,31,86,31,252,31,114,31,114,30,8,31,241,31,139,31,123,31,103,31,91,31,165,31,28,31,88,31,67,31,158,31,9,31,98,31,98,30,167,31,167,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
