-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_764 is
end project_tb_764;

architecture project_tb_arch_764 of project_tb_764 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 433;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (163,0,11,0,51,0,0,0,128,0,98,0,241,0,15,0,148,0,145,0,0,0,254,0,143,0,184,0,101,0,19,0,0,0,19,0,0,0,45,0,147,0,0,0,0,0,105,0,231,0,0,0,225,0,158,0,0,0,209,0,0,0,149,0,126,0,59,0,0,0,224,0,222,0,37,0,117,0,0,0,187,0,213,0,0,0,170,0,253,0,0,0,2,0,57,0,0,0,109,0,0,0,0,0,12,0,0,0,53,0,11,0,199,0,91,0,227,0,0,0,58,0,89,0,132,0,217,0,134,0,0,0,138,0,67,0,0,0,0,0,13,0,0,0,0,0,209,0,154,0,176,0,169,0,13,0,163,0,122,0,2,0,178,0,210,0,73,0,75,0,0,0,28,0,243,0,135,0,212,0,226,0,102,0,69,0,151,0,62,0,32,0,90,0,160,0,0,0,245,0,0,0,7,0,0,0,148,0,29,0,21,0,0,0,184,0,209,0,153,0,0,0,35,0,172,0,235,0,0,0,56,0,0,0,129,0,59,0,233,0,0,0,155,0,149,0,94,0,0,0,165,0,137,0,246,0,199,0,140,0,49,0,0,0,52,0,149,0,74,0,198,0,131,0,102,0,22,0,199,0,190,0,0,0,29,0,62,0,41,0,59,0,0,0,3,0,130,0,196,0,0,0,0,0,187,0,157,0,68,0,83,0,112,0,116,0,193,0,2,0,227,0,113,0,173,0,85,0,228,0,191,0,88,0,0,0,172,0,255,0,181,0,225,0,123,0,27,0,137,0,15,0,31,0,107,0,190,0,120,0,162,0,222,0,77,0,35,0,121,0,78,0,162,0,66,0,28,0,27,0,0,0,126,0,25,0,138,0,60,0,0,0,174,0,204,0,0,0,0,0,111,0,40,0,192,0,165,0,0,0,0,0,10,0,0,0,128,0,172,0,241,0,0,0,247,0,0,0,38,0,58,0,64,0,246,0,229,0,30,0,7,0,239,0,115,0,0,0,216,0,0,0,245,0,18,0,0,0,145,0,197,0,34,0,225,0,255,0,198,0,0,0,60,0,9,0,63,0,93,0,74,0,170,0,125,0,202,0,138,0,0,0,19,0,236,0,95,0,64,0,178,0,0,0,211,0,149,0,109,0,255,0,0,0,84,0,170,0,142,0,142,0,219,0,0,0,0,0,168,0,23,0,189,0,0,0,0,0,200,0,191,0,0,0,0,0,0,0,115,0,5,0,16,0,219,0,115,0,150,0,140,0,0,0,252,0,0,0,95,0,47,0,0,0,0,0,0,0,184,0,146,0,118,0,65,0,231,0,0,0,227,0,58,0,247,0,166,0,99,0,0,0,0,0,225,0,190,0,0,0,165,0,252,0,21,0,149,0,35,0,252,0,0,0,171,0,218,0,0,0,142,0,31,0,0,0,18,0,0,0,0,0,0,0,187,0,70,0,7,0,0,0,148,0,40,0,0,0,172,0,105,0,200,0,89,0,140,0,240,0,221,0,29,0,189,0,106,0,64,0,0,0,118,0,36,0,107,0,135,0,91,0,155,0,0,0,0,0,218,0,65,0,0,0,239,0,99,0,200,0,0,0,0,0,200,0,143,0,124,0,105,0,237,0,223,0,0,0,0,0,224,0,163,0,70,0,200,0,189,0,0,0,47,0,73,0,87,0,34,0,52,0,210,0,0,0,3,0,0,0,128,0,0,0,161,0,0,0,0,0,0,0,142,0,0,0,250,0,249,0,60,0,227,0,209,0,131,0,120,0,1,0,0,0,155,0,241,0,7,0,184,0,0,0,190,0,69,0,0,0,29,0,243,0,0,0,0,0,96,0,134,0,68,0,222,0,0,0,0,0,168,0,64,0,254,0,192,0,4,0,93,0,0,0,0,0,219,0,241,0,0,0,153,0,0,0,196,0,0,0,42,0,0,0,115,0);
signal scenario_full  : scenario_type := (163,31,11,31,51,31,51,30,128,31,98,31,241,31,15,31,148,31,145,31,145,30,254,31,143,31,184,31,101,31,19,31,19,30,19,31,19,30,45,31,147,31,147,30,147,29,105,31,231,31,231,30,225,31,158,31,158,30,209,31,209,30,149,31,126,31,59,31,59,30,224,31,222,31,37,31,117,31,117,30,187,31,213,31,213,30,170,31,253,31,253,30,2,31,57,31,57,30,109,31,109,30,109,29,12,31,12,30,53,31,11,31,199,31,91,31,227,31,227,30,58,31,89,31,132,31,217,31,134,31,134,30,138,31,67,31,67,30,67,29,13,31,13,30,13,29,209,31,154,31,176,31,169,31,13,31,163,31,122,31,2,31,178,31,210,31,73,31,75,31,75,30,28,31,243,31,135,31,212,31,226,31,102,31,69,31,151,31,62,31,32,31,90,31,160,31,160,30,245,31,245,30,7,31,7,30,148,31,29,31,21,31,21,30,184,31,209,31,153,31,153,30,35,31,172,31,235,31,235,30,56,31,56,30,129,31,59,31,233,31,233,30,155,31,149,31,94,31,94,30,165,31,137,31,246,31,199,31,140,31,49,31,49,30,52,31,149,31,74,31,198,31,131,31,102,31,22,31,199,31,190,31,190,30,29,31,62,31,41,31,59,31,59,30,3,31,130,31,196,31,196,30,196,29,187,31,157,31,68,31,83,31,112,31,116,31,193,31,2,31,227,31,113,31,173,31,85,31,228,31,191,31,88,31,88,30,172,31,255,31,181,31,225,31,123,31,27,31,137,31,15,31,31,31,107,31,190,31,120,31,162,31,222,31,77,31,35,31,121,31,78,31,162,31,66,31,28,31,27,31,27,30,126,31,25,31,138,31,60,31,60,30,174,31,204,31,204,30,204,29,111,31,40,31,192,31,165,31,165,30,165,29,10,31,10,30,128,31,172,31,241,31,241,30,247,31,247,30,38,31,58,31,64,31,246,31,229,31,30,31,7,31,239,31,115,31,115,30,216,31,216,30,245,31,18,31,18,30,145,31,197,31,34,31,225,31,255,31,198,31,198,30,60,31,9,31,63,31,93,31,74,31,170,31,125,31,202,31,138,31,138,30,19,31,236,31,95,31,64,31,178,31,178,30,211,31,149,31,109,31,255,31,255,30,84,31,170,31,142,31,142,31,219,31,219,30,219,29,168,31,23,31,189,31,189,30,189,29,200,31,191,31,191,30,191,29,191,28,115,31,5,31,16,31,219,31,115,31,150,31,140,31,140,30,252,31,252,30,95,31,47,31,47,30,47,29,47,28,184,31,146,31,118,31,65,31,231,31,231,30,227,31,58,31,247,31,166,31,99,31,99,30,99,29,225,31,190,31,190,30,165,31,252,31,21,31,149,31,35,31,252,31,252,30,171,31,218,31,218,30,142,31,31,31,31,30,18,31,18,30,18,29,18,28,187,31,70,31,7,31,7,30,148,31,40,31,40,30,172,31,105,31,200,31,89,31,140,31,240,31,221,31,29,31,189,31,106,31,64,31,64,30,118,31,36,31,107,31,135,31,91,31,155,31,155,30,155,29,218,31,65,31,65,30,239,31,99,31,200,31,200,30,200,29,200,31,143,31,124,31,105,31,237,31,223,31,223,30,223,29,224,31,163,31,70,31,200,31,189,31,189,30,47,31,73,31,87,31,34,31,52,31,210,31,210,30,3,31,3,30,128,31,128,30,161,31,161,30,161,29,161,28,142,31,142,30,250,31,249,31,60,31,227,31,209,31,131,31,120,31,1,31,1,30,155,31,241,31,7,31,184,31,184,30,190,31,69,31,69,30,29,31,243,31,243,30,243,29,96,31,134,31,68,31,222,31,222,30,222,29,168,31,64,31,254,31,192,31,4,31,93,31,93,30,93,29,219,31,241,31,241,30,153,31,153,30,196,31,196,30,42,31,42,30,115,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
