-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_571 is
end project_tb_571;

architecture project_tb_arch_571 of project_tb_571 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 874;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,38,0,198,0,234,0,164,0,0,0,142,0,169,0,183,0,232,0,200,0,44,0,8,0,74,0,101,0,98,0,12,0,225,0,65,0,119,0,77,0,254,0,69,0,196,0,125,0,105,0,232,0,159,0,28,0,0,0,21,0,120,0,159,0,118,0,90,0,0,0,254,0,0,0,230,0,189,0,15,0,76,0,237,0,137,0,0,0,227,0,148,0,21,0,187,0,230,0,136,0,33,0,82,0,0,0,216,0,59,0,0,0,161,0,27,0,0,0,225,0,150,0,147,0,179,0,0,0,34,0,15,0,31,0,0,0,85,0,0,0,116,0,187,0,0,0,238,0,233,0,101,0,239,0,154,0,234,0,178,0,218,0,209,0,0,0,199,0,245,0,34,0,0,0,140,0,113,0,45,0,108,0,0,0,3,0,0,0,55,0,218,0,0,0,0,0,134,0,132,0,10,0,193,0,146,0,178,0,236,0,146,0,0,0,66,0,184,0,5,0,19,0,0,0,180,0,233,0,59,0,234,0,22,0,209,0,224,0,162,0,0,0,75,0,177,0,225,0,206,0,178,0,11,0,49,0,0,0,0,0,5,0,200,0,131,0,118,0,159,0,0,0,13,0,0,0,26,0,181,0,165,0,75,0,208,0,156,0,0,0,149,0,212,0,25,0,244,0,0,0,240,0,214,0,0,0,0,0,0,0,0,0,7,0,0,0,201,0,117,0,184,0,47,0,132,0,85,0,194,0,225,0,112,0,32,0,48,0,229,0,0,0,20,0,84,0,214,0,98,0,165,0,102,0,20,0,85,0,104,0,140,0,0,0,125,0,75,0,0,0,232,0,16,0,244,0,171,0,137,0,0,0,242,0,8,0,0,0,76,0,0,0,131,0,170,0,224,0,94,0,0,0,103,0,127,0,183,0,125,0,83,0,161,0,148,0,217,0,184,0,185,0,21,0,0,0,0,0,0,0,197,0,71,0,153,0,196,0,228,0,33,0,213,0,52,0,247,0,196,0,0,0,245,0,0,0,210,0,0,0,244,0,163,0,164,0,16,0,207,0,36,0,0,0,0,0,177,0,64,0,151,0,13,0,22,0,0,0,0,0,0,0,248,0,88,0,103,0,59,0,83,0,47,0,156,0,131,0,43,0,120,0,0,0,192,0,0,0,73,0,221,0,0,0,233,0,204,0,20,0,76,0,219,0,167,0,31,0,121,0,192,0,0,0,226,0,0,0,97,0,146,0,231,0,62,0,0,0,47,0,0,0,237,0,111,0,60,0,2,0,157,0,160,0,0,0,0,0,173,0,145,0,95,0,0,0,0,0,253,0,183,0,226,0,115,0,204,0,141,0,140,0,80,0,0,0,120,0,177,0,0,0,0,0,242,0,25,0,83,0,212,0,29,0,0,0,29,0,108,0,198,0,217,0,129,0,0,0,0,0,0,0,221,0,120,0,114,0,18,0,0,0,231,0,97,0,0,0,220,0,170,0,206,0,14,0,211,0,0,0,76,0,0,0,238,0,216,0,19,0,169,0,241,0,150,0,110,0,3,0,188,0,38,0,126,0,108,0,250,0,125,0,102,0,0,0,182,0,55,0,0,0,187,0,8,0,117,0,231,0,85,0,0,0,70,0,141,0,20,0,130,0,193,0,109,0,46,0,69,0,165,0,74,0,207,0,0,0,6,0,130,0,104,0,184,0,69,0,18,0,181,0,123,0,250,0,0,0,253,0,68,0,153,0,35,0,56,0,214,0,231,0,90,0,143,0,240,0,98,0,51,0,0,0,70,0,0,0,0,0,0,0,138,0,154,0,207,0,0,0,84,0,0,0,0,0,140,0,0,0,86,0,170,0,41,0,201,0,104,0,17,0,14,0,0,0,149,0,213,0,29,0,33,0,82,0,0,0,17,0,91,0,0,0,8,0,112,0,0,0,57,0,38,0,110,0,0,0,214,0,80,0,125,0,250,0,0,0,28,0,194,0,0,0,81,0,100,0,216,0,82,0,59,0,0,0,157,0,71,0,0,0,0,0,68,0,1,0,184,0,120,0,214,0,0,0,112,0,223,0,37,0,198,0,114,0,222,0,114,0,0,0,20,0,0,0,48,0,0,0,236,0,102,0,246,0,74,0,62,0,194,0,92,0,0,0,32,0,237,0,0,0,0,0,163,0,121,0,0,0,152,0,69,0,143,0,189,0,0,0,18,0,176,0,150,0,41,0,217,0,175,0,234,0,35,0,124,0,137,0,0,0,249,0,200,0,95,0,0,0,199,0,41,0,0,0,0,0,131,0,0,0,223,0,28,0,134,0,98,0,214,0,0,0,178,0,172,0,242,0,186,0,57,0,169,0,150,0,0,0,166,0,218,0,0,0,0,0,140,0,134,0,4,0,69,0,205,0,228,0,180,0,126,0,61,0,156,0,18,0,127,0,0,0,28,0,145,0,173,0,85,0,126,0,249,0,115,0,253,0,211,0,71,0,93,0,217,0,197,0,11,0,38,0,0,0,0,0,0,0,111,0,0,0,0,0,241,0,195,0,224,0,0,0,5,0,84,0,154,0,0,0,94,0,157,0,97,0,201,0,80,0,186,0,0,0,158,0,54,0,197,0,71,0,76,0,0,0,139,0,50,0,162,0,111,0,90,0,179,0,2,0,0,0,0,0,118,0,117,0,0,0,72,0,133,0,16,0,0,0,54,0,135,0,225,0,142,0,86,0,191,0,142,0,227,0,51,0,54,0,0,0,127,0,0,0,129,0,166,0,0,0,120,0,24,0,110,0,138,0,99,0,64,0,26,0,33,0,70,0,0,0,91,0,2,0,183,0,199,0,249,0,253,0,47,0,57,0,0,0,67,0,236,0,116,0,53,0,134,0,193,0,0,0,127,0,202,0,160,0,0,0,0,0,144,0,0,0,0,0,135,0,72,0,113,0,212,0,51,0,121,0,0,0,130,0,151,0,60,0,0,0,0,0,42,0,219,0,0,0,182,0,125,0,115,0,184,0,43,0,238,0,146,0,149,0,0,0,214,0,0,0,78,0,252,0,218,0,171,0,87,0,22,0,220,0,229,0,126,0,73,0,169,0,0,0,174,0,45,0,131,0,0,0,47,0,96,0,54,0,17,0,111,0,70,0,66,0,90,0,31,0,0,0,117,0,51,0,96,0,117,0,0,0,0,0,93,0,43,0,0,0,46,0,124,0,152,0,234,0,73,0,185,0,0,0,63,0,148,0,223,0,16,0,73,0,206,0,203,0,77,0,74,0,55,0,208,0,78,0,84,0,169,0,22,0,87,0,77,0,240,0,0,0,0,0,249,0,160,0,0,0,0,0,133,0,162,0,137,0,42,0,0,0,158,0,221,0,233,0,241,0,218,0,0,0,193,0,229,0,13,0,39,0,0,0,152,0,47,0,82,0,0,0,75,0,0,0,157,0,70,0,39,0,124,0,0,0,254,0,177,0,148,0,59,0,0,0,233,0,0,0,0,0,0,0,255,0,0,0,0,0,0,0,6,0,30,0,18,0,5,0,26,0,0,0,205,0,118,0,103,0,117,0,130,0,102,0,16,0,233,0,145,0,217,0,152,0,16,0,230,0,203,0,164,0,141,0,161,0,0,0,0,0,0,0,171,0,162,0,68,0,0,0,114,0,11,0,205,0,97,0,0,0,73,0,140,0,89,0,70,0,166,0,74,0,0,0,64,0,211,0,10,0,157,0,174,0,168,0,15,0,202,0,0,0,100,0,64,0,137,0,102,0,233,0,46,0,108,0,0,0,12,0,53,0,249,0,52,0,112,0,0,0,253,0,93,0,54,0,142,0,243,0,0,0,143,0,208,0,128,0,223,0,57,0,0,0,50,0,232,0,144,0,192,0,0,0,131,0,0,0,110,0,234,0,37,0,11,0,201,0,154,0,0,0);
signal scenario_full  : scenario_type := (0,0,38,31,198,31,234,31,164,31,164,30,142,31,169,31,183,31,232,31,200,31,44,31,8,31,74,31,101,31,98,31,12,31,225,31,65,31,119,31,77,31,254,31,69,31,196,31,125,31,105,31,232,31,159,31,28,31,28,30,21,31,120,31,159,31,118,31,90,31,90,30,254,31,254,30,230,31,189,31,15,31,76,31,237,31,137,31,137,30,227,31,148,31,21,31,187,31,230,31,136,31,33,31,82,31,82,30,216,31,59,31,59,30,161,31,27,31,27,30,225,31,150,31,147,31,179,31,179,30,34,31,15,31,31,31,31,30,85,31,85,30,116,31,187,31,187,30,238,31,233,31,101,31,239,31,154,31,234,31,178,31,218,31,209,31,209,30,199,31,245,31,34,31,34,30,140,31,113,31,45,31,108,31,108,30,3,31,3,30,55,31,218,31,218,30,218,29,134,31,132,31,10,31,193,31,146,31,178,31,236,31,146,31,146,30,66,31,184,31,5,31,19,31,19,30,180,31,233,31,59,31,234,31,22,31,209,31,224,31,162,31,162,30,75,31,177,31,225,31,206,31,178,31,11,31,49,31,49,30,49,29,5,31,200,31,131,31,118,31,159,31,159,30,13,31,13,30,26,31,181,31,165,31,75,31,208,31,156,31,156,30,149,31,212,31,25,31,244,31,244,30,240,31,214,31,214,30,214,29,214,28,214,27,7,31,7,30,201,31,117,31,184,31,47,31,132,31,85,31,194,31,225,31,112,31,32,31,48,31,229,31,229,30,20,31,84,31,214,31,98,31,165,31,102,31,20,31,85,31,104,31,140,31,140,30,125,31,75,31,75,30,232,31,16,31,244,31,171,31,137,31,137,30,242,31,8,31,8,30,76,31,76,30,131,31,170,31,224,31,94,31,94,30,103,31,127,31,183,31,125,31,83,31,161,31,148,31,217,31,184,31,185,31,21,31,21,30,21,29,21,28,197,31,71,31,153,31,196,31,228,31,33,31,213,31,52,31,247,31,196,31,196,30,245,31,245,30,210,31,210,30,244,31,163,31,164,31,16,31,207,31,36,31,36,30,36,29,177,31,64,31,151,31,13,31,22,31,22,30,22,29,22,28,248,31,88,31,103,31,59,31,83,31,47,31,156,31,131,31,43,31,120,31,120,30,192,31,192,30,73,31,221,31,221,30,233,31,204,31,20,31,76,31,219,31,167,31,31,31,121,31,192,31,192,30,226,31,226,30,97,31,146,31,231,31,62,31,62,30,47,31,47,30,237,31,111,31,60,31,2,31,157,31,160,31,160,30,160,29,173,31,145,31,95,31,95,30,95,29,253,31,183,31,226,31,115,31,204,31,141,31,140,31,80,31,80,30,120,31,177,31,177,30,177,29,242,31,25,31,83,31,212,31,29,31,29,30,29,31,108,31,198,31,217,31,129,31,129,30,129,29,129,28,221,31,120,31,114,31,18,31,18,30,231,31,97,31,97,30,220,31,170,31,206,31,14,31,211,31,211,30,76,31,76,30,238,31,216,31,19,31,169,31,241,31,150,31,110,31,3,31,188,31,38,31,126,31,108,31,250,31,125,31,102,31,102,30,182,31,55,31,55,30,187,31,8,31,117,31,231,31,85,31,85,30,70,31,141,31,20,31,130,31,193,31,109,31,46,31,69,31,165,31,74,31,207,31,207,30,6,31,130,31,104,31,184,31,69,31,18,31,181,31,123,31,250,31,250,30,253,31,68,31,153,31,35,31,56,31,214,31,231,31,90,31,143,31,240,31,98,31,51,31,51,30,70,31,70,30,70,29,70,28,138,31,154,31,207,31,207,30,84,31,84,30,84,29,140,31,140,30,86,31,170,31,41,31,201,31,104,31,17,31,14,31,14,30,149,31,213,31,29,31,33,31,82,31,82,30,17,31,91,31,91,30,8,31,112,31,112,30,57,31,38,31,110,31,110,30,214,31,80,31,125,31,250,31,250,30,28,31,194,31,194,30,81,31,100,31,216,31,82,31,59,31,59,30,157,31,71,31,71,30,71,29,68,31,1,31,184,31,120,31,214,31,214,30,112,31,223,31,37,31,198,31,114,31,222,31,114,31,114,30,20,31,20,30,48,31,48,30,236,31,102,31,246,31,74,31,62,31,194,31,92,31,92,30,32,31,237,31,237,30,237,29,163,31,121,31,121,30,152,31,69,31,143,31,189,31,189,30,18,31,176,31,150,31,41,31,217,31,175,31,234,31,35,31,124,31,137,31,137,30,249,31,200,31,95,31,95,30,199,31,41,31,41,30,41,29,131,31,131,30,223,31,28,31,134,31,98,31,214,31,214,30,178,31,172,31,242,31,186,31,57,31,169,31,150,31,150,30,166,31,218,31,218,30,218,29,140,31,134,31,4,31,69,31,205,31,228,31,180,31,126,31,61,31,156,31,18,31,127,31,127,30,28,31,145,31,173,31,85,31,126,31,249,31,115,31,253,31,211,31,71,31,93,31,217,31,197,31,11,31,38,31,38,30,38,29,38,28,111,31,111,30,111,29,241,31,195,31,224,31,224,30,5,31,84,31,154,31,154,30,94,31,157,31,97,31,201,31,80,31,186,31,186,30,158,31,54,31,197,31,71,31,76,31,76,30,139,31,50,31,162,31,111,31,90,31,179,31,2,31,2,30,2,29,118,31,117,31,117,30,72,31,133,31,16,31,16,30,54,31,135,31,225,31,142,31,86,31,191,31,142,31,227,31,51,31,54,31,54,30,127,31,127,30,129,31,166,31,166,30,120,31,24,31,110,31,138,31,99,31,64,31,26,31,33,31,70,31,70,30,91,31,2,31,183,31,199,31,249,31,253,31,47,31,57,31,57,30,67,31,236,31,116,31,53,31,134,31,193,31,193,30,127,31,202,31,160,31,160,30,160,29,144,31,144,30,144,29,135,31,72,31,113,31,212,31,51,31,121,31,121,30,130,31,151,31,60,31,60,30,60,29,42,31,219,31,219,30,182,31,125,31,115,31,184,31,43,31,238,31,146,31,149,31,149,30,214,31,214,30,78,31,252,31,218,31,171,31,87,31,22,31,220,31,229,31,126,31,73,31,169,31,169,30,174,31,45,31,131,31,131,30,47,31,96,31,54,31,17,31,111,31,70,31,66,31,90,31,31,31,31,30,117,31,51,31,96,31,117,31,117,30,117,29,93,31,43,31,43,30,46,31,124,31,152,31,234,31,73,31,185,31,185,30,63,31,148,31,223,31,16,31,73,31,206,31,203,31,77,31,74,31,55,31,208,31,78,31,84,31,169,31,22,31,87,31,77,31,240,31,240,30,240,29,249,31,160,31,160,30,160,29,133,31,162,31,137,31,42,31,42,30,158,31,221,31,233,31,241,31,218,31,218,30,193,31,229,31,13,31,39,31,39,30,152,31,47,31,82,31,82,30,75,31,75,30,157,31,70,31,39,31,124,31,124,30,254,31,177,31,148,31,59,31,59,30,233,31,233,30,233,29,233,28,255,31,255,30,255,29,255,28,6,31,30,31,18,31,5,31,26,31,26,30,205,31,118,31,103,31,117,31,130,31,102,31,16,31,233,31,145,31,217,31,152,31,16,31,230,31,203,31,164,31,141,31,161,31,161,30,161,29,161,28,171,31,162,31,68,31,68,30,114,31,11,31,205,31,97,31,97,30,73,31,140,31,89,31,70,31,166,31,74,31,74,30,64,31,211,31,10,31,157,31,174,31,168,31,15,31,202,31,202,30,100,31,64,31,137,31,102,31,233,31,46,31,108,31,108,30,12,31,53,31,249,31,52,31,112,31,112,30,253,31,93,31,54,31,142,31,243,31,243,30,143,31,208,31,128,31,223,31,57,31,57,30,50,31,232,31,144,31,192,31,192,30,131,31,131,30,110,31,234,31,37,31,11,31,201,31,154,31,154,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
