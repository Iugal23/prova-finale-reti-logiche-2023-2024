-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 774;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,216,0,181,0,206,0,135,0,44,0,245,0,54,0,112,0,0,0,245,0,232,0,193,0,109,0,147,0,181,0,227,0,0,0,213,0,0,0,119,0,170,0,12,0,2,0,4,0,0,0,214,0,64,0,191,0,42,0,0,0,196,0,158,0,0,0,63,0,38,0,115,0,239,0,74,0,0,0,147,0,46,0,0,0,0,0,218,0,187,0,44,0,32,0,29,0,0,0,223,0,61,0,57,0,0,0,0,0,92,0,29,0,0,0,0,0,0,0,54,0,164,0,157,0,227,0,129,0,67,0,244,0,123,0,155,0,249,0,9,0,71,0,70,0,98,0,136,0,17,0,0,0,28,0,43,0,23,0,250,0,178,0,132,0,193,0,184,0,242,0,65,0,138,0,250,0,106,0,0,0,124,0,59,0,111,0,28,0,43,0,0,0,0,0,190,0,182,0,48,0,183,0,102,0,129,0,143,0,186,0,0,0,99,0,115,0,140,0,117,0,94,0,9,0,50,0,0,0,238,0,115,0,183,0,0,0,117,0,183,0,60,0,184,0,0,0,240,0,129,0,254,0,0,0,248,0,194,0,251,0,17,0,131,0,104,0,0,0,94,0,201,0,0,0,250,0,154,0,155,0,79,0,46,0,203,0,0,0,143,0,224,0,0,0,252,0,0,0,254,0,2,0,131,0,104,0,165,0,166,0,0,0,211,0,0,0,106,0,250,0,90,0,83,0,243,0,0,0,173,0,107,0,222,0,114,0,216,0,0,0,0,0,34,0,75,0,0,0,42,0,35,0,0,0,0,0,109,0,182,0,94,0,196,0,196,0,171,0,10,0,182,0,0,0,185,0,61,0,82,0,252,0,189,0,0,0,31,0,1,0,132,0,0,0,172,0,4,0,156,0,229,0,133,0,146,0,43,0,21,0,153,0,159,0,0,0,68,0,209,0,71,0,71,0,103,0,70,0,182,0,0,0,147,0,240,0,23,0,0,0,95,0,187,0,135,0,82,0,117,0,0,0,0,0,17,0,232,0,192,0,0,0,103,0,0,0,255,0,81,0,243,0,123,0,166,0,173,0,0,0,12,0,1,0,212,0,0,0,76,0,175,0,84,0,100,0,29,0,29,0,37,0,0,0,78,0,139,0,0,0,211,0,0,0,109,0,196,0,139,0,62,0,103,0,200,0,239,0,231,0,242,0,222,0,233,0,227,0,205,0,72,0,0,0,0,0,229,0,122,0,72,0,91,0,155,0,168,0,161,0,0,0,227,0,63,0,0,0,74,0,110,0,191,0,172,0,53,0,229,0,0,0,49,0,196,0,173,0,0,0,0,0,93,0,46,0,215,0,211,0,91,0,232,0,71,0,72,0,143,0,166,0,0,0,0,0,183,0,62,0,20,0,145,0,79,0,223,0,241,0,0,0,183,0,234,0,190,0,32,0,71,0,0,0,42,0,115,0,50,0,0,0,149,0,151,0,109,0,113,0,1,0,165,0,0,0,48,0,56,0,243,0,76,0,0,0,149,0,214,0,137,0,4,0,18,0,221,0,69,0,109,0,15,0,170,0,45,0,234,0,185,0,236,0,191,0,13,0,96,0,0,0,140,0,55,0,70,0,216,0,134,0,106,0,119,0,22,0,34,0,0,0,0,0,209,0,76,0,72,0,73,0,39,0,0,0,0,0,215,0,113,0,128,0,167,0,28,0,151,0,52,0,9,0,67,0,124,0,117,0,111,0,227,0,100,0,91,0,4,0,14,0,0,0,66,0,184,0,0,0,0,0,0,0,13,0,123,0,247,0,0,0,0,0,98,0,217,0,239,0,0,0,223,0,197,0,243,0,251,0,251,0,4,0,171,0,161,0,180,0,0,0,116,0,207,0,59,0,211,0,0,0,114,0,0,0,239,0,222,0,21,0,109,0,208,0,199,0,0,0,66,0,0,0,199,0,40,0,0,0,107,0,132,0,236,0,105,0,0,0,163,0,161,0,179,0,156,0,5,0,0,0,91,0,31,0,129,0,116,0,128,0,202,0,131,0,31,0,206,0,54,0,122,0,236,0,0,0,71,0,147,0,101,0,118,0,131,0,214,0,177,0,84,0,167,0,191,0,239,0,0,0,0,0,0,0,0,0,139,0,220,0,223,0,93,0,0,0,212,0,23,0,115,0,142,0,0,0,163,0,131,0,56,0,0,0,16,0,247,0,232,0,89,0,217,0,10,0,19,0,105,0,237,0,0,0,0,0,218,0,101,0,229,0,161,0,246,0,0,0,77,0,205,0,93,0,26,0,0,0,0,0,18,0,35,0,60,0,86,0,0,0,41,0,60,0,104,0,160,0,0,0,186,0,199,0,101,0,19,0,18,0,106,0,178,0,0,0,0,0,49,0,0,0,178,0,170,0,225,0,222,0,154,0,189,0,181,0,249,0,128,0,81,0,120,0,228,0,75,0,27,0,0,0,139,0,0,0,0,0,0,0,1,0,108,0,241,0,177,0,143,0,0,0,55,0,195,0,246,0,193,0,62,0,225,0,12,0,0,0,238,0,0,0,79,0,96,0,115,0,209,0,153,0,50,0,194,0,164,0,103,0,60,0,252,0,5,0,130,0,148,0,82,0,234,0,230,0,224,0,240,0,13,0,8,0,219,0,7,0,0,0,0,0,21,0,75,0,222,0,0,0,155,0,222,0,189,0,55,0,204,0,25,0,140,0,56,0,0,0,201,0,223,0,0,0,76,0,159,0,72,0,71,0,104,0,50,0,0,0,0,0,0,0,0,0,75,0,15,0,36,0,106,0,34,0,126,0,129,0,17,0,187,0,182,0,248,0,0,0,112,0,39,0,195,0,129,0,248,0,71,0,85,0,53,0,204,0,239,0,43,0,23,0,0,0,0,0,148,0,0,0,217,0,127,0,157,0,0,0,163,0,89,0,0,0,191,0,87,0,50,0,0,0,181,0,211,0,205,0,186,0,127,0,45,0,0,0,225,0,208,0,47,0,120,0,223,0,155,0,0,0,84,0,162,0,104,0,234,0,146,0,161,0,66,0,0,0,56,0,175,0,235,0,63,0,50,0,117,0,232,0,76,0,0,0,28,0,69,0,228,0,97,0,237,0,0,0,125,0,213,0,0,0,165,0,0,0,143,0,132,0,0,0,249,0,205,0,0,0,132,0,110,0,118,0,0,0,56,0,182,0,153,0,0,0,174,0,249,0,239,0,71,0,0,0,202,0,168,0,197,0,109,0,116,0,139,0,24,0,38,0,252,0,244,0,219,0,172,0,248,0,0,0,226,0,45,0,92,0,67,0,0,0,21,0,0,0,104,0,0,0,61,0,148,0,154,0,173,0,166,0,90,0,74,0,53,0,11,0,227,0,47,0,32,0,97,0,73,0,243,0,93,0,246,0,187,0,135,0,129,0,184,0,0,0,0,0,0,0,0,0,103,0,77,0,174,0,0,0,255,0,15,0,143,0);
signal scenario_full  : scenario_type := (0,0,216,31,181,31,206,31,135,31,44,31,245,31,54,31,112,31,112,30,245,31,232,31,193,31,109,31,147,31,181,31,227,31,227,30,213,31,213,30,119,31,170,31,12,31,2,31,4,31,4,30,214,31,64,31,191,31,42,31,42,30,196,31,158,31,158,30,63,31,38,31,115,31,239,31,74,31,74,30,147,31,46,31,46,30,46,29,218,31,187,31,44,31,32,31,29,31,29,30,223,31,61,31,57,31,57,30,57,29,92,31,29,31,29,30,29,29,29,28,54,31,164,31,157,31,227,31,129,31,67,31,244,31,123,31,155,31,249,31,9,31,71,31,70,31,98,31,136,31,17,31,17,30,28,31,43,31,23,31,250,31,178,31,132,31,193,31,184,31,242,31,65,31,138,31,250,31,106,31,106,30,124,31,59,31,111,31,28,31,43,31,43,30,43,29,190,31,182,31,48,31,183,31,102,31,129,31,143,31,186,31,186,30,99,31,115,31,140,31,117,31,94,31,9,31,50,31,50,30,238,31,115,31,183,31,183,30,117,31,183,31,60,31,184,31,184,30,240,31,129,31,254,31,254,30,248,31,194,31,251,31,17,31,131,31,104,31,104,30,94,31,201,31,201,30,250,31,154,31,155,31,79,31,46,31,203,31,203,30,143,31,224,31,224,30,252,31,252,30,254,31,2,31,131,31,104,31,165,31,166,31,166,30,211,31,211,30,106,31,250,31,90,31,83,31,243,31,243,30,173,31,107,31,222,31,114,31,216,31,216,30,216,29,34,31,75,31,75,30,42,31,35,31,35,30,35,29,109,31,182,31,94,31,196,31,196,31,171,31,10,31,182,31,182,30,185,31,61,31,82,31,252,31,189,31,189,30,31,31,1,31,132,31,132,30,172,31,4,31,156,31,229,31,133,31,146,31,43,31,21,31,153,31,159,31,159,30,68,31,209,31,71,31,71,31,103,31,70,31,182,31,182,30,147,31,240,31,23,31,23,30,95,31,187,31,135,31,82,31,117,31,117,30,117,29,17,31,232,31,192,31,192,30,103,31,103,30,255,31,81,31,243,31,123,31,166,31,173,31,173,30,12,31,1,31,212,31,212,30,76,31,175,31,84,31,100,31,29,31,29,31,37,31,37,30,78,31,139,31,139,30,211,31,211,30,109,31,196,31,139,31,62,31,103,31,200,31,239,31,231,31,242,31,222,31,233,31,227,31,205,31,72,31,72,30,72,29,229,31,122,31,72,31,91,31,155,31,168,31,161,31,161,30,227,31,63,31,63,30,74,31,110,31,191,31,172,31,53,31,229,31,229,30,49,31,196,31,173,31,173,30,173,29,93,31,46,31,215,31,211,31,91,31,232,31,71,31,72,31,143,31,166,31,166,30,166,29,183,31,62,31,20,31,145,31,79,31,223,31,241,31,241,30,183,31,234,31,190,31,32,31,71,31,71,30,42,31,115,31,50,31,50,30,149,31,151,31,109,31,113,31,1,31,165,31,165,30,48,31,56,31,243,31,76,31,76,30,149,31,214,31,137,31,4,31,18,31,221,31,69,31,109,31,15,31,170,31,45,31,234,31,185,31,236,31,191,31,13,31,96,31,96,30,140,31,55,31,70,31,216,31,134,31,106,31,119,31,22,31,34,31,34,30,34,29,209,31,76,31,72,31,73,31,39,31,39,30,39,29,215,31,113,31,128,31,167,31,28,31,151,31,52,31,9,31,67,31,124,31,117,31,111,31,227,31,100,31,91,31,4,31,14,31,14,30,66,31,184,31,184,30,184,29,184,28,13,31,123,31,247,31,247,30,247,29,98,31,217,31,239,31,239,30,223,31,197,31,243,31,251,31,251,31,4,31,171,31,161,31,180,31,180,30,116,31,207,31,59,31,211,31,211,30,114,31,114,30,239,31,222,31,21,31,109,31,208,31,199,31,199,30,66,31,66,30,199,31,40,31,40,30,107,31,132,31,236,31,105,31,105,30,163,31,161,31,179,31,156,31,5,31,5,30,91,31,31,31,129,31,116,31,128,31,202,31,131,31,31,31,206,31,54,31,122,31,236,31,236,30,71,31,147,31,101,31,118,31,131,31,214,31,177,31,84,31,167,31,191,31,239,31,239,30,239,29,239,28,239,27,139,31,220,31,223,31,93,31,93,30,212,31,23,31,115,31,142,31,142,30,163,31,131,31,56,31,56,30,16,31,247,31,232,31,89,31,217,31,10,31,19,31,105,31,237,31,237,30,237,29,218,31,101,31,229,31,161,31,246,31,246,30,77,31,205,31,93,31,26,31,26,30,26,29,18,31,35,31,60,31,86,31,86,30,41,31,60,31,104,31,160,31,160,30,186,31,199,31,101,31,19,31,18,31,106,31,178,31,178,30,178,29,49,31,49,30,178,31,170,31,225,31,222,31,154,31,189,31,181,31,249,31,128,31,81,31,120,31,228,31,75,31,27,31,27,30,139,31,139,30,139,29,139,28,1,31,108,31,241,31,177,31,143,31,143,30,55,31,195,31,246,31,193,31,62,31,225,31,12,31,12,30,238,31,238,30,79,31,96,31,115,31,209,31,153,31,50,31,194,31,164,31,103,31,60,31,252,31,5,31,130,31,148,31,82,31,234,31,230,31,224,31,240,31,13,31,8,31,219,31,7,31,7,30,7,29,21,31,75,31,222,31,222,30,155,31,222,31,189,31,55,31,204,31,25,31,140,31,56,31,56,30,201,31,223,31,223,30,76,31,159,31,72,31,71,31,104,31,50,31,50,30,50,29,50,28,50,27,75,31,15,31,36,31,106,31,34,31,126,31,129,31,17,31,187,31,182,31,248,31,248,30,112,31,39,31,195,31,129,31,248,31,71,31,85,31,53,31,204,31,239,31,43,31,23,31,23,30,23,29,148,31,148,30,217,31,127,31,157,31,157,30,163,31,89,31,89,30,191,31,87,31,50,31,50,30,181,31,211,31,205,31,186,31,127,31,45,31,45,30,225,31,208,31,47,31,120,31,223,31,155,31,155,30,84,31,162,31,104,31,234,31,146,31,161,31,66,31,66,30,56,31,175,31,235,31,63,31,50,31,117,31,232,31,76,31,76,30,28,31,69,31,228,31,97,31,237,31,237,30,125,31,213,31,213,30,165,31,165,30,143,31,132,31,132,30,249,31,205,31,205,30,132,31,110,31,118,31,118,30,56,31,182,31,153,31,153,30,174,31,249,31,239,31,71,31,71,30,202,31,168,31,197,31,109,31,116,31,139,31,24,31,38,31,252,31,244,31,219,31,172,31,248,31,248,30,226,31,45,31,92,31,67,31,67,30,21,31,21,30,104,31,104,30,61,31,148,31,154,31,173,31,166,31,90,31,74,31,53,31,11,31,227,31,47,31,32,31,97,31,73,31,243,31,93,31,246,31,187,31,135,31,129,31,184,31,184,30,184,29,184,28,184,27,103,31,77,31,174,31,174,30,255,31,15,31,143,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
