-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_6 is
end project_tb_6;

architecture project_tb_arch_6 of project_tb_6 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 761;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (143,0,108,0,174,0,0,0,147,0,23,0,142,0,115,0,0,0,138,0,0,0,86,0,166,0,7,0,165,0,123,0,115,0,207,0,226,0,209,0,71,0,183,0,0,0,0,0,193,0,0,0,238,0,192,0,235,0,0,0,0,0,15,0,0,0,45,0,153,0,0,0,0,0,0,0,138,0,244,0,198,0,134,0,62,0,103,0,0,0,46,0,4,0,83,0,183,0,184,0,0,0,0,0,99,0,72,0,61,0,204,0,196,0,145,0,117,0,42,0,226,0,118,0,198,0,181,0,111,0,206,0,5,0,36,0,133,0,234,0,145,0,179,0,89,0,2,0,38,0,164,0,7,0,122,0,0,0,102,0,89,0,48,0,165,0,63,0,144,0,211,0,0,0,241,0,230,0,165,0,52,0,197,0,237,0,51,0,77,0,82,0,180,0,147,0,0,0,5,0,250,0,84,0,13,0,235,0,0,0,185,0,88,0,112,0,162,0,33,0,161,0,234,0,0,0,7,0,103,0,125,0,169,0,188,0,188,0,83,0,19,0,136,0,4,0,224,0,63,0,40,0,133,0,21,0,94,0,203,0,246,0,127,0,52,0,179,0,73,0,0,0,31,0,121,0,47,0,0,0,127,0,42,0,236,0,97,0,0,0,113,0,9,0,195,0,251,0,0,0,245,0,40,0,47,0,0,0,149,0,249,0,41,0,27,0,77,0,112,0,242,0,19,0,224,0,244,0,0,0,251,0,32,0,100,0,125,0,0,0,35,0,126,0,66,0,211,0,235,0,26,0,0,0,244,0,252,0,117,0,0,0,175,0,20,0,182,0,50,0,170,0,241,0,163,0,0,0,30,0,156,0,241,0,3,0,92,0,0,0,46,0,76,0,2,0,131,0,0,0,7,0,29,0,210,0,133,0,88,0,221,0,180,0,29,0,50,0,112,0,49,0,79,0,51,0,0,0,0,0,28,0,187,0,110,0,155,0,102,0,56,0,249,0,139,0,0,0,16,0,175,0,60,0,0,0,49,0,58,0,183,0,87,0,2,0,0,0,45,0,0,0,213,0,65,0,0,0,143,0,201,0,0,0,101,0,83,0,0,0,108,0,217,0,61,0,24,0,44,0,202,0,0,0,152,0,101,0,167,0,204,0,182,0,170,0,36,0,178,0,0,0,141,0,243,0,0,0,0,0,204,0,0,0,100,0,177,0,248,0,192,0,0,0,143,0,0,0,179,0,27,0,140,0,79,0,23,0,210,0,8,0,186,0,107,0,133,0,224,0,19,0,0,0,74,0,122,0,144,0,242,0,234,0,0,0,0,0,61,0,0,0,121,0,210,0,115,0,234,0,229,0,44,0,162,0,145,0,51,0,187,0,207,0,52,0,47,0,186,0,153,0,194,0,154,0,177,0,206,0,165,0,0,0,248,0,233,0,236,0,0,0,62,0,43,0,21,0,0,0,55,0,79,0,17,0,0,0,165,0,14,0,24,0,242,0,227,0,91,0,0,0,146,0,147,0,0,0,230,0,198,0,218,0,91,0,168,0,189,0,59,0,82,0,99,0,137,0,228,0,73,0,112,0,91,0,25,0,0,0,207,0,248,0,112,0,242,0,190,0,225,0,172,0,181,0,52,0,213,0,20,0,20,0,38,0,131,0,16,0,172,0,0,0,0,0,112,0,138,0,21,0,135,0,192,0,0,0,33,0,235,0,129,0,103,0,218,0,134,0,17,0,241,0,168,0,204,0,246,0,37,0,128,0,144,0,0,0,0,0,64,0,0,0,118,0,0,0,179,0,97,0,229,0,119,0,0,0,143,0,27,0,218,0,28,0,8,0,77,0,46,0,190,0,108,0,57,0,191,0,174,0,254,0,119,0,97,0,154,0,203,0,222,0,0,0,28,0,97,0,125,0,93,0,32,0,30,0,126,0,40,0,0,0,169,0,105,0,83,0,0,0,132,0,0,0,0,0,154,0,50,0,0,0,221,0,0,0,160,0,92,0,111,0,4,0,228,0,39,0,101,0,161,0,111,0,107,0,118,0,0,0,102,0,75,0,197,0,0,0,44,0,199,0,67,0,31,0,207,0,0,0,0,0,236,0,205,0,175,0,233,0,0,0,42,0,101,0,106,0,186,0,112,0,49,0,0,0,50,0,206,0,252,0,201,0,204,0,128,0,88,0,53,0,0,0,189,0,211,0,14,0,184,0,0,0,102,0,57,0,239,0,111,0,0,0,98,0,170,0,159,0,173,0,125,0,249,0,79,0,229,0,97,0,0,0,63,0,0,0,0,0,23,0,182,0,200,0,196,0,0,0,190,0,103,0,139,0,214,0,30,0,192,0,45,0,75,0,0,0,49,0,44,0,0,0,147,0,152,0,94,0,0,0,97,0,0,0,165,0,0,0,253,0,162,0,161,0,94,0,0,0,0,0,172,0,189,0,14,0,0,0,51,0,97,0,118,0,54,0,0,0,104,0,26,0,38,0,0,0,149,0,102,0,0,0,161,0,0,0,206,0,220,0,0,0,18,0,43,0,133,0,100,0,0,0,81,0,0,0,222,0,27,0,0,0,54,0,180,0,0,0,0,0,117,0,177,0,151,0,0,0,41,0,21,0,0,0,55,0,76,0,224,0,107,0,23,0,126,0,133,0,34,0,180,0,176,0,0,0,0,0,0,0,150,0,0,0,123,0,0,0,23,0,0,0,79,0,18,0,195,0,0,0,93,0,50,0,0,0,173,0,121,0,108,0,229,0,193,0,0,0,58,0,118,0,154,0,47,0,16,0,195,0,143,0,167,0,31,0,109,0,45,0,71,0,76,0,217,0,0,0,102,0,54,0,0,0,0,0,74,0,0,0,0,0,84,0,225,0,242,0,99,0,108,0,171,0,149,0,0,0,155,0,90,0,0,0,123,0,49,0,253,0,0,0,88,0,0,0,133,0,203,0,0,0,9,0,63,0,0,0,0,0,23,0,188,0,66,0,138,0,105,0,121,0,99,0,237,0,0,0,56,0,242,0,0,0,77,0,247,0,47,0,238,0,254,0,196,0,247,0,243,0,198,0,95,0,215,0,0,0,0,0,202,0,49,0,171,0,234,0,16,0,103,0,59,0,66,0,122,0,133,0,0,0,206,0,0,0,45,0,197,0,0,0,73,0,116,0,75,0,0,0,176,0,0,0,254,0,0,0,116,0,137,0,173,0,255,0,0,0,9,0,0,0,141,0,0,0,133,0,78,0,79,0,45,0,0,0,183,0,146,0,220,0,0,0,58,0,152,0,251,0,222,0,201,0,222,0,0,0,176,0,60,0,0,0,225,0,125,0,237,0,78,0,74,0,0,0,60,0,164,0,0,0,208,0,109,0,113,0,201,0,99,0,182,0,197,0,205,0,0,0,146,0,0,0,143,0,107,0);
signal scenario_full  : scenario_type := (143,31,108,31,174,31,174,30,147,31,23,31,142,31,115,31,115,30,138,31,138,30,86,31,166,31,7,31,165,31,123,31,115,31,207,31,226,31,209,31,71,31,183,31,183,30,183,29,193,31,193,30,238,31,192,31,235,31,235,30,235,29,15,31,15,30,45,31,153,31,153,30,153,29,153,28,138,31,244,31,198,31,134,31,62,31,103,31,103,30,46,31,4,31,83,31,183,31,184,31,184,30,184,29,99,31,72,31,61,31,204,31,196,31,145,31,117,31,42,31,226,31,118,31,198,31,181,31,111,31,206,31,5,31,36,31,133,31,234,31,145,31,179,31,89,31,2,31,38,31,164,31,7,31,122,31,122,30,102,31,89,31,48,31,165,31,63,31,144,31,211,31,211,30,241,31,230,31,165,31,52,31,197,31,237,31,51,31,77,31,82,31,180,31,147,31,147,30,5,31,250,31,84,31,13,31,235,31,235,30,185,31,88,31,112,31,162,31,33,31,161,31,234,31,234,30,7,31,103,31,125,31,169,31,188,31,188,31,83,31,19,31,136,31,4,31,224,31,63,31,40,31,133,31,21,31,94,31,203,31,246,31,127,31,52,31,179,31,73,31,73,30,31,31,121,31,47,31,47,30,127,31,42,31,236,31,97,31,97,30,113,31,9,31,195,31,251,31,251,30,245,31,40,31,47,31,47,30,149,31,249,31,41,31,27,31,77,31,112,31,242,31,19,31,224,31,244,31,244,30,251,31,32,31,100,31,125,31,125,30,35,31,126,31,66,31,211,31,235,31,26,31,26,30,244,31,252,31,117,31,117,30,175,31,20,31,182,31,50,31,170,31,241,31,163,31,163,30,30,31,156,31,241,31,3,31,92,31,92,30,46,31,76,31,2,31,131,31,131,30,7,31,29,31,210,31,133,31,88,31,221,31,180,31,29,31,50,31,112,31,49,31,79,31,51,31,51,30,51,29,28,31,187,31,110,31,155,31,102,31,56,31,249,31,139,31,139,30,16,31,175,31,60,31,60,30,49,31,58,31,183,31,87,31,2,31,2,30,45,31,45,30,213,31,65,31,65,30,143,31,201,31,201,30,101,31,83,31,83,30,108,31,217,31,61,31,24,31,44,31,202,31,202,30,152,31,101,31,167,31,204,31,182,31,170,31,36,31,178,31,178,30,141,31,243,31,243,30,243,29,204,31,204,30,100,31,177,31,248,31,192,31,192,30,143,31,143,30,179,31,27,31,140,31,79,31,23,31,210,31,8,31,186,31,107,31,133,31,224,31,19,31,19,30,74,31,122,31,144,31,242,31,234,31,234,30,234,29,61,31,61,30,121,31,210,31,115,31,234,31,229,31,44,31,162,31,145,31,51,31,187,31,207,31,52,31,47,31,186,31,153,31,194,31,154,31,177,31,206,31,165,31,165,30,248,31,233,31,236,31,236,30,62,31,43,31,21,31,21,30,55,31,79,31,17,31,17,30,165,31,14,31,24,31,242,31,227,31,91,31,91,30,146,31,147,31,147,30,230,31,198,31,218,31,91,31,168,31,189,31,59,31,82,31,99,31,137,31,228,31,73,31,112,31,91,31,25,31,25,30,207,31,248,31,112,31,242,31,190,31,225,31,172,31,181,31,52,31,213,31,20,31,20,31,38,31,131,31,16,31,172,31,172,30,172,29,112,31,138,31,21,31,135,31,192,31,192,30,33,31,235,31,129,31,103,31,218,31,134,31,17,31,241,31,168,31,204,31,246,31,37,31,128,31,144,31,144,30,144,29,64,31,64,30,118,31,118,30,179,31,97,31,229,31,119,31,119,30,143,31,27,31,218,31,28,31,8,31,77,31,46,31,190,31,108,31,57,31,191,31,174,31,254,31,119,31,97,31,154,31,203,31,222,31,222,30,28,31,97,31,125,31,93,31,32,31,30,31,126,31,40,31,40,30,169,31,105,31,83,31,83,30,132,31,132,30,132,29,154,31,50,31,50,30,221,31,221,30,160,31,92,31,111,31,4,31,228,31,39,31,101,31,161,31,111,31,107,31,118,31,118,30,102,31,75,31,197,31,197,30,44,31,199,31,67,31,31,31,207,31,207,30,207,29,236,31,205,31,175,31,233,31,233,30,42,31,101,31,106,31,186,31,112,31,49,31,49,30,50,31,206,31,252,31,201,31,204,31,128,31,88,31,53,31,53,30,189,31,211,31,14,31,184,31,184,30,102,31,57,31,239,31,111,31,111,30,98,31,170,31,159,31,173,31,125,31,249,31,79,31,229,31,97,31,97,30,63,31,63,30,63,29,23,31,182,31,200,31,196,31,196,30,190,31,103,31,139,31,214,31,30,31,192,31,45,31,75,31,75,30,49,31,44,31,44,30,147,31,152,31,94,31,94,30,97,31,97,30,165,31,165,30,253,31,162,31,161,31,94,31,94,30,94,29,172,31,189,31,14,31,14,30,51,31,97,31,118,31,54,31,54,30,104,31,26,31,38,31,38,30,149,31,102,31,102,30,161,31,161,30,206,31,220,31,220,30,18,31,43,31,133,31,100,31,100,30,81,31,81,30,222,31,27,31,27,30,54,31,180,31,180,30,180,29,117,31,177,31,151,31,151,30,41,31,21,31,21,30,55,31,76,31,224,31,107,31,23,31,126,31,133,31,34,31,180,31,176,31,176,30,176,29,176,28,150,31,150,30,123,31,123,30,23,31,23,30,79,31,18,31,195,31,195,30,93,31,50,31,50,30,173,31,121,31,108,31,229,31,193,31,193,30,58,31,118,31,154,31,47,31,16,31,195,31,143,31,167,31,31,31,109,31,45,31,71,31,76,31,217,31,217,30,102,31,54,31,54,30,54,29,74,31,74,30,74,29,84,31,225,31,242,31,99,31,108,31,171,31,149,31,149,30,155,31,90,31,90,30,123,31,49,31,253,31,253,30,88,31,88,30,133,31,203,31,203,30,9,31,63,31,63,30,63,29,23,31,188,31,66,31,138,31,105,31,121,31,99,31,237,31,237,30,56,31,242,31,242,30,77,31,247,31,47,31,238,31,254,31,196,31,247,31,243,31,198,31,95,31,215,31,215,30,215,29,202,31,49,31,171,31,234,31,16,31,103,31,59,31,66,31,122,31,133,31,133,30,206,31,206,30,45,31,197,31,197,30,73,31,116,31,75,31,75,30,176,31,176,30,254,31,254,30,116,31,137,31,173,31,255,31,255,30,9,31,9,30,141,31,141,30,133,31,78,31,79,31,45,31,45,30,183,31,146,31,220,31,220,30,58,31,152,31,251,31,222,31,201,31,222,31,222,30,176,31,60,31,60,30,225,31,125,31,237,31,78,31,74,31,74,30,60,31,164,31,164,30,208,31,109,31,113,31,201,31,99,31,182,31,197,31,205,31,205,30,146,31,146,30,143,31,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
