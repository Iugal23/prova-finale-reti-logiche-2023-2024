-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_282 is
end project_tb_282;

architecture project_tb_arch_282 of project_tb_282 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 296;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,253,0,193,0,185,0,226,0,0,0,0,0,89,0,9,0,0,0,152,0,28,0,0,0,245,0,171,0,0,0,209,0,86,0,5,0,155,0,0,0,147,0,240,0,0,0,35,0,48,0,166,0,80,0,169,0,127,0,3,0,0,0,205,0,17,0,31,0,57,0,70,0,3,0,32,0,224,0,5,0,168,0,228,0,89,0,125,0,134,0,105,0,0,0,0,0,132,0,190,0,52,0,253,0,210,0,80,0,255,0,35,0,201,0,198,0,236,0,82,0,177,0,33,0,132,0,60,0,202,0,68,0,196,0,128,0,151,0,69,0,0,0,0,0,94,0,102,0,0,0,210,0,142,0,0,0,142,0,171,0,0,0,144,0,0,0,246,0,109,0,116,0,245,0,51,0,70,0,217,0,160,0,252,0,17,0,174,0,0,0,236,0,241,0,53,0,81,0,176,0,0,0,174,0,51,0,160,0,0,0,62,0,0,0,117,0,0,0,7,0,250,0,129,0,0,0,212,0,54,0,45,0,151,0,175,0,0,0,175,0,0,0,122,0,52,0,212,0,0,0,154,0,41,0,181,0,207,0,66,0,32,0,250,0,170,0,83,0,189,0,122,0,90,0,73,0,248,0,191,0,87,0,166,0,0,0,154,0,132,0,242,0,51,0,97,0,12,0,134,0,0,0,161,0,194,0,172,0,107,0,226,0,69,0,1,0,213,0,179,0,250,0,0,0,189,0,158,0,5,0,60,0,71,0,48,0,46,0,0,0,72,0,133,0,191,0,21,0,137,0,104,0,20,0,222,0,0,0,15,0,40,0,0,0,204,0,107,0,125,0,0,0,0,0,255,0,0,0,33,0,44,0,113,0,144,0,238,0,0,0,0,0,24,0,209,0,0,0,94,0,39,0,0,0,32,0,113,0,0,0,37,0,64,0,0,0,93,0,0,0,180,0,0,0,0,0,79,0,0,0,62,0,119,0,0,0,82,0,202,0,198,0,172,0,54,0,84,0,222,0,49,0,228,0,57,0,0,0,58,0,1,0,241,0,200,0,100,0,123,0,223,0,205,0,231,0,243,0,128,0,0,0,43,0,244,0,132,0,79,0,0,0,46,0,219,0,212,0,188,0,181,0,3,0,50,0,143,0,20,0,22,0,0,0,97,0,8,0,86,0,248,0,178,0,112,0,0,0,161,0,221,0,145,0,56,0,187,0,80,0,112,0,118,0,198,0,100,0,0,0,90,0,62,0,112,0,119,0,0,0,34,0,5,0,0,0,194,0,0,0,49,0,60,0,249,0,35,0,97,0,42,0,180,0,3,0,218,0,0,0);
signal scenario_full  : scenario_type := (0,0,253,31,193,31,185,31,226,31,226,30,226,29,89,31,9,31,9,30,152,31,28,31,28,30,245,31,171,31,171,30,209,31,86,31,5,31,155,31,155,30,147,31,240,31,240,30,35,31,48,31,166,31,80,31,169,31,127,31,3,31,3,30,205,31,17,31,31,31,57,31,70,31,3,31,32,31,224,31,5,31,168,31,228,31,89,31,125,31,134,31,105,31,105,30,105,29,132,31,190,31,52,31,253,31,210,31,80,31,255,31,35,31,201,31,198,31,236,31,82,31,177,31,33,31,132,31,60,31,202,31,68,31,196,31,128,31,151,31,69,31,69,30,69,29,94,31,102,31,102,30,210,31,142,31,142,30,142,31,171,31,171,30,144,31,144,30,246,31,109,31,116,31,245,31,51,31,70,31,217,31,160,31,252,31,17,31,174,31,174,30,236,31,241,31,53,31,81,31,176,31,176,30,174,31,51,31,160,31,160,30,62,31,62,30,117,31,117,30,7,31,250,31,129,31,129,30,212,31,54,31,45,31,151,31,175,31,175,30,175,31,175,30,122,31,52,31,212,31,212,30,154,31,41,31,181,31,207,31,66,31,32,31,250,31,170,31,83,31,189,31,122,31,90,31,73,31,248,31,191,31,87,31,166,31,166,30,154,31,132,31,242,31,51,31,97,31,12,31,134,31,134,30,161,31,194,31,172,31,107,31,226,31,69,31,1,31,213,31,179,31,250,31,250,30,189,31,158,31,5,31,60,31,71,31,48,31,46,31,46,30,72,31,133,31,191,31,21,31,137,31,104,31,20,31,222,31,222,30,15,31,40,31,40,30,204,31,107,31,125,31,125,30,125,29,255,31,255,30,33,31,44,31,113,31,144,31,238,31,238,30,238,29,24,31,209,31,209,30,94,31,39,31,39,30,32,31,113,31,113,30,37,31,64,31,64,30,93,31,93,30,180,31,180,30,180,29,79,31,79,30,62,31,119,31,119,30,82,31,202,31,198,31,172,31,54,31,84,31,222,31,49,31,228,31,57,31,57,30,58,31,1,31,241,31,200,31,100,31,123,31,223,31,205,31,231,31,243,31,128,31,128,30,43,31,244,31,132,31,79,31,79,30,46,31,219,31,212,31,188,31,181,31,3,31,50,31,143,31,20,31,22,31,22,30,97,31,8,31,86,31,248,31,178,31,112,31,112,30,161,31,221,31,145,31,56,31,187,31,80,31,112,31,118,31,198,31,100,31,100,30,90,31,62,31,112,31,119,31,119,30,34,31,5,31,5,30,194,31,194,30,49,31,60,31,249,31,35,31,97,31,42,31,180,31,3,31,218,31,218,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
