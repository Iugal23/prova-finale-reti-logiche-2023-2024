-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 896;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (85,0,25,0,225,0,158,0,0,0,160,0,246,0,20,0,126,0,67,0,160,0,128,0,158,0,0,0,1,0,45,0,38,0,199,0,173,0,65,0,249,0,210,0,0,0,0,0,0,0,169,0,87,0,228,0,255,0,139,0,194,0,18,0,18,0,240,0,123,0,0,0,243,0,29,0,170,0,0,0,188,0,0,0,203,0,160,0,62,0,32,0,90,0,0,0,92,0,249,0,66,0,62,0,73,0,149,0,57,0,230,0,82,0,15,0,158,0,0,0,0,0,50,0,0,0,48,0,27,0,157,0,0,0,241,0,1,0,117,0,0,0,12,0,52,0,170,0,191,0,159,0,82,0,140,0,74,0,3,0,4,0,190,0,253,0,137,0,174,0,101,0,136,0,68,0,84,0,159,0,127,0,39,0,172,0,76,0,0,0,214,0,19,0,73,0,0,0,207,0,88,0,41,0,226,0,0,0,186,0,242,0,13,0,81,0,203,0,241,0,109,0,158,0,108,0,0,0,173,0,18,0,0,0,0,0,183,0,205,0,174,0,166,0,216,0,115,0,248,0,147,0,184,0,109,0,96,0,25,0,74,0,27,0,0,0,0,0,0,0,0,0,183,0,0,0,192,0,63,0,82,0,191,0,78,0,33,0,0,0,0,0,23,0,0,0,141,0,83,0,0,0,0,0,222,0,36,0,0,0,173,0,75,0,212,0,36,0,249,0,163,0,21,0,76,0,0,0,46,0,184,0,147,0,252,0,0,0,0,0,0,0,0,0,0,0,208,0,196,0,15,0,0,0,219,0,146,0,85,0,32,0,178,0,0,0,15,0,33,0,103,0,211,0,17,0,0,0,133,0,0,0,206,0,64,0,218,0,170,0,4,0,165,0,84,0,0,0,72,0,14,0,59,0,0,0,79,0,8,0,227,0,0,0,209,0,9,0,121,0,84,0,116,0,0,0,0,0,212,0,152,0,56,0,0,0,60,0,70,0,109,0,0,0,60,0,122,0,188,0,107,0,223,0,170,0,69,0,0,0,11,0,130,0,158,0,136,0,106,0,113,0,210,0,0,0,55,0,183,0,157,0,179,0,0,0,77,0,200,0,0,0,11,0,0,0,89,0,246,0,225,0,203,0,203,0,0,0,144,0,221,0,183,0,216,0,160,0,83,0,0,0,85,0,0,0,58,0,0,0,37,0,5,0,148,0,0,0,22,0,33,0,92,0,0,0,0,0,46,0,131,0,169,0,30,0,170,0,0,0,10,0,114,0,234,0,172,0,0,0,232,0,0,0,10,0,160,0,89,0,198,0,23,0,222,0,128,0,67,0,205,0,77,0,206,0,205,0,221,0,44,0,4,0,217,0,188,0,113,0,37,0,0,0,200,0,144,0,0,0,70,0,193,0,7,0,162,0,36,0,155,0,51,0,211,0,97,0,196,0,246,0,20,0,246,0,0,0,180,0,48,0,222,0,34,0,0,0,179,0,87,0,7,0,233,0,225,0,226,0,174,0,99,0,175,0,94,0,22,0,110,0,27,0,163,0,156,0,78,0,51,0,55,0,144,0,200,0,18,0,3,0,0,0,22,0,0,0,0,0,247,0,0,0,89,0,0,0,139,0,94,0,87,0,0,0,0,0,106,0,67,0,19,0,208,0,0,0,209,0,212,0,58,0,246,0,144,0,31,0,153,0,0,0,157,0,205,0,0,0,9,0,195,0,126,0,198,0,0,0,50,0,77,0,0,0,139,0,18,0,125,0,0,0,102,0,254,0,134,0,129,0,172,0,0,0,205,0,0,0,94,0,1,0,162,0,18,0,0,0,193,0,27,0,63,0,197,0,153,0,39,0,95,0,161,0,207,0,142,0,96,0,137,0,74,0,100,0,204,0,0,0,251,0,231,0,0,0,146,0,44,0,200,0,42,0,170,0,177,0,183,0,189,0,245,0,0,0,227,0,65,0,125,0,70,0,246,0,224,0,0,0,40,0,0,0,147,0,254,0,208,0,129,0,7,0,251,0,121,0,57,0,35,0,78,0,14,0,0,0,198,0,151,0,0,0,120,0,2,0,34,0,85,0,99,0,4,0,164,0,8,0,240,0,0,0,0,0,248,0,54,0,178,0,188,0,225,0,149,0,212,0,204,0,85,0,96,0,37,0,208,0,27,0,10,0,206,0,219,0,76,0,0,0,0,0,235,0,146,0,80,0,0,0,0,0,38,0,0,0,0,0,118,0,0,0,0,0,181,0,152,0,91,0,96,0,62,0,0,0,0,0,126,0,0,0,155,0,73,0,141,0,44,0,134,0,227,0,107,0,147,0,174,0,104,0,175,0,29,0,91,0,130,0,182,0,0,0,45,0,55,0,42,0,67,0,135,0,10,0,81,0,150,0,174,0,228,0,22,0,237,0,203,0,160,0,209,0,0,0,0,0,207,0,83,0,25,0,97,0,147,0,13,0,3,0,142,0,0,0,145,0,220,0,109,0,56,0,82,0,41,0,119,0,0,0,0,0,231,0,29,0,0,0,160,0,158,0,48,0,55,0,0,0,92,0,0,0,0,0,134,0,255,0,68,0,34,0,129,0,216,0,12,0,248,0,144,0,0,0,101,0,163,0,0,0,29,0,230,0,0,0,0,0,227,0,156,0,192,0,0,0,189,0,27,0,0,0,92,0,221,0,147,0,36,0,81,0,2,0,0,0,34,0,124,0,36,0,0,0,179,0,234,0,8,0,245,0,0,0,13,0,0,0,171,0,115,0,0,0,0,0,89,0,91,0,61,0,29,0,83,0,178,0,164,0,91,0,25,0,36,0,180,0,2,0,76,0,238,0,0,0,222,0,193,0,72,0,38,0,91,0,140,0,133,0,208,0,148,0,144,0,78,0,237,0,23,0,139,0,172,0,245,0,38,0,168,0,18,0,185,0,188,0,0,0,113,0,202,0,50,0,116,0,195,0,60,0,153,0,45,0,158,0,0,0,0,0,230,0,162,0,142,0,194,0,32,0,169,0,0,0,220,0,146,0,3,0,113,0,167,0,46,0,0,0,44,0,0,0,213,0,108,0,88,0,87,0,209,0,233,0,219,0,87,0,7,0,59,0,0,0,126,0,60,0,226,0,0,0,82,0,187,0,10,0,0,0,136,0,161,0,85,0,0,0,40,0,0,0,165,0,0,0,46,0,0,0,13,0,0,0,114,0,213,0,4,0,59,0,195,0,170,0,0,0,10,0,26,0,153,0,142,0,0,0,0,0,0,0,167,0,238,0,254,0,67,0,156,0,203,0,0,0,57,0,61,0,0,0,181,0,133,0,0,0,68,0,0,0,152,0,44,0,97,0,81,0,82,0,93,0,56,0,232,0,76,0,88,0,0,0,0,0,216,0,92,0,0,0,95,0,26,0,0,0,0,0,247,0,79,0,89,0,180,0,17,0,0,0,159,0,168,0,93,0,56,0,72,0,68,0,59,0,171,0,0,0,197,0,108,0,0,0,253,0,169,0,184,0,23,0,66,0,183,0,52,0,55,0,127,0,225,0,186,0,39,0,44,0,0,0,174,0,235,0,95,0,0,0,65,0,89,0,102,0,0,0,112,0,251,0,47,0,62,0,250,0,190,0,106,0,208,0,0,0,0,0,197,0,219,0,3,0,11,0,39,0,95,0,0,0,121,0,225,0,80,0,52,0,188,0,1,0,116,0,103,0,28,0,0,0,169,0,77,0,0,0,4,0,29,0,171,0,0,0,69,0,238,0,208,0,12,0,79,0,248,0,0,0,150,0,0,0,0,0,211,0,43,0,0,0,189,0,95,0,67,0,89,0,0,0,227,0,7,0,0,0,0,0,0,0,149,0,0,0,0,0,92,0,205,0,0,0,0,0,119,0,219,0,111,0,0,0,248,0,46,0,186,0,138,0,66,0,198,0,242,0,42,0,0,0,0,0,237,0,169,0,229,0,225,0,183,0,29,0,47,0,6,0,253,0,61,0,0,0,249,0,5,0,69,0,101,0,0,0,0,0,184,0,44,0);
signal scenario_full  : scenario_type := (85,31,25,31,225,31,158,31,158,30,160,31,246,31,20,31,126,31,67,31,160,31,128,31,158,31,158,30,1,31,45,31,38,31,199,31,173,31,65,31,249,31,210,31,210,30,210,29,210,28,169,31,87,31,228,31,255,31,139,31,194,31,18,31,18,31,240,31,123,31,123,30,243,31,29,31,170,31,170,30,188,31,188,30,203,31,160,31,62,31,32,31,90,31,90,30,92,31,249,31,66,31,62,31,73,31,149,31,57,31,230,31,82,31,15,31,158,31,158,30,158,29,50,31,50,30,48,31,27,31,157,31,157,30,241,31,1,31,117,31,117,30,12,31,52,31,170,31,191,31,159,31,82,31,140,31,74,31,3,31,4,31,190,31,253,31,137,31,174,31,101,31,136,31,68,31,84,31,159,31,127,31,39,31,172,31,76,31,76,30,214,31,19,31,73,31,73,30,207,31,88,31,41,31,226,31,226,30,186,31,242,31,13,31,81,31,203,31,241,31,109,31,158,31,108,31,108,30,173,31,18,31,18,30,18,29,183,31,205,31,174,31,166,31,216,31,115,31,248,31,147,31,184,31,109,31,96,31,25,31,74,31,27,31,27,30,27,29,27,28,27,27,183,31,183,30,192,31,63,31,82,31,191,31,78,31,33,31,33,30,33,29,23,31,23,30,141,31,83,31,83,30,83,29,222,31,36,31,36,30,173,31,75,31,212,31,36,31,249,31,163,31,21,31,76,31,76,30,46,31,184,31,147,31,252,31,252,30,252,29,252,28,252,27,252,26,208,31,196,31,15,31,15,30,219,31,146,31,85,31,32,31,178,31,178,30,15,31,33,31,103,31,211,31,17,31,17,30,133,31,133,30,206,31,64,31,218,31,170,31,4,31,165,31,84,31,84,30,72,31,14,31,59,31,59,30,79,31,8,31,227,31,227,30,209,31,9,31,121,31,84,31,116,31,116,30,116,29,212,31,152,31,56,31,56,30,60,31,70,31,109,31,109,30,60,31,122,31,188,31,107,31,223,31,170,31,69,31,69,30,11,31,130,31,158,31,136,31,106,31,113,31,210,31,210,30,55,31,183,31,157,31,179,31,179,30,77,31,200,31,200,30,11,31,11,30,89,31,246,31,225,31,203,31,203,31,203,30,144,31,221,31,183,31,216,31,160,31,83,31,83,30,85,31,85,30,58,31,58,30,37,31,5,31,148,31,148,30,22,31,33,31,92,31,92,30,92,29,46,31,131,31,169,31,30,31,170,31,170,30,10,31,114,31,234,31,172,31,172,30,232,31,232,30,10,31,160,31,89,31,198,31,23,31,222,31,128,31,67,31,205,31,77,31,206,31,205,31,221,31,44,31,4,31,217,31,188,31,113,31,37,31,37,30,200,31,144,31,144,30,70,31,193,31,7,31,162,31,36,31,155,31,51,31,211,31,97,31,196,31,246,31,20,31,246,31,246,30,180,31,48,31,222,31,34,31,34,30,179,31,87,31,7,31,233,31,225,31,226,31,174,31,99,31,175,31,94,31,22,31,110,31,27,31,163,31,156,31,78,31,51,31,55,31,144,31,200,31,18,31,3,31,3,30,22,31,22,30,22,29,247,31,247,30,89,31,89,30,139,31,94,31,87,31,87,30,87,29,106,31,67,31,19,31,208,31,208,30,209,31,212,31,58,31,246,31,144,31,31,31,153,31,153,30,157,31,205,31,205,30,9,31,195,31,126,31,198,31,198,30,50,31,77,31,77,30,139,31,18,31,125,31,125,30,102,31,254,31,134,31,129,31,172,31,172,30,205,31,205,30,94,31,1,31,162,31,18,31,18,30,193,31,27,31,63,31,197,31,153,31,39,31,95,31,161,31,207,31,142,31,96,31,137,31,74,31,100,31,204,31,204,30,251,31,231,31,231,30,146,31,44,31,200,31,42,31,170,31,177,31,183,31,189,31,245,31,245,30,227,31,65,31,125,31,70,31,246,31,224,31,224,30,40,31,40,30,147,31,254,31,208,31,129,31,7,31,251,31,121,31,57,31,35,31,78,31,14,31,14,30,198,31,151,31,151,30,120,31,2,31,34,31,85,31,99,31,4,31,164,31,8,31,240,31,240,30,240,29,248,31,54,31,178,31,188,31,225,31,149,31,212,31,204,31,85,31,96,31,37,31,208,31,27,31,10,31,206,31,219,31,76,31,76,30,76,29,235,31,146,31,80,31,80,30,80,29,38,31,38,30,38,29,118,31,118,30,118,29,181,31,152,31,91,31,96,31,62,31,62,30,62,29,126,31,126,30,155,31,73,31,141,31,44,31,134,31,227,31,107,31,147,31,174,31,104,31,175,31,29,31,91,31,130,31,182,31,182,30,45,31,55,31,42,31,67,31,135,31,10,31,81,31,150,31,174,31,228,31,22,31,237,31,203,31,160,31,209,31,209,30,209,29,207,31,83,31,25,31,97,31,147,31,13,31,3,31,142,31,142,30,145,31,220,31,109,31,56,31,82,31,41,31,119,31,119,30,119,29,231,31,29,31,29,30,160,31,158,31,48,31,55,31,55,30,92,31,92,30,92,29,134,31,255,31,68,31,34,31,129,31,216,31,12,31,248,31,144,31,144,30,101,31,163,31,163,30,29,31,230,31,230,30,230,29,227,31,156,31,192,31,192,30,189,31,27,31,27,30,92,31,221,31,147,31,36,31,81,31,2,31,2,30,34,31,124,31,36,31,36,30,179,31,234,31,8,31,245,31,245,30,13,31,13,30,171,31,115,31,115,30,115,29,89,31,91,31,61,31,29,31,83,31,178,31,164,31,91,31,25,31,36,31,180,31,2,31,76,31,238,31,238,30,222,31,193,31,72,31,38,31,91,31,140,31,133,31,208,31,148,31,144,31,78,31,237,31,23,31,139,31,172,31,245,31,38,31,168,31,18,31,185,31,188,31,188,30,113,31,202,31,50,31,116,31,195,31,60,31,153,31,45,31,158,31,158,30,158,29,230,31,162,31,142,31,194,31,32,31,169,31,169,30,220,31,146,31,3,31,113,31,167,31,46,31,46,30,44,31,44,30,213,31,108,31,88,31,87,31,209,31,233,31,219,31,87,31,7,31,59,31,59,30,126,31,60,31,226,31,226,30,82,31,187,31,10,31,10,30,136,31,161,31,85,31,85,30,40,31,40,30,165,31,165,30,46,31,46,30,13,31,13,30,114,31,213,31,4,31,59,31,195,31,170,31,170,30,10,31,26,31,153,31,142,31,142,30,142,29,142,28,167,31,238,31,254,31,67,31,156,31,203,31,203,30,57,31,61,31,61,30,181,31,133,31,133,30,68,31,68,30,152,31,44,31,97,31,81,31,82,31,93,31,56,31,232,31,76,31,88,31,88,30,88,29,216,31,92,31,92,30,95,31,26,31,26,30,26,29,247,31,79,31,89,31,180,31,17,31,17,30,159,31,168,31,93,31,56,31,72,31,68,31,59,31,171,31,171,30,197,31,108,31,108,30,253,31,169,31,184,31,23,31,66,31,183,31,52,31,55,31,127,31,225,31,186,31,39,31,44,31,44,30,174,31,235,31,95,31,95,30,65,31,89,31,102,31,102,30,112,31,251,31,47,31,62,31,250,31,190,31,106,31,208,31,208,30,208,29,197,31,219,31,3,31,11,31,39,31,95,31,95,30,121,31,225,31,80,31,52,31,188,31,1,31,116,31,103,31,28,31,28,30,169,31,77,31,77,30,4,31,29,31,171,31,171,30,69,31,238,31,208,31,12,31,79,31,248,31,248,30,150,31,150,30,150,29,211,31,43,31,43,30,189,31,95,31,67,31,89,31,89,30,227,31,7,31,7,30,7,29,7,28,149,31,149,30,149,29,92,31,205,31,205,30,205,29,119,31,219,31,111,31,111,30,248,31,46,31,186,31,138,31,66,31,198,31,242,31,42,31,42,30,42,29,237,31,169,31,229,31,225,31,183,31,29,31,47,31,6,31,253,31,61,31,61,30,249,31,5,31,69,31,101,31,101,30,101,29,184,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
