-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_493 is
end project_tb_493;

architecture project_tb_arch_493 of project_tb_493 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 157;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (21,0,57,0,164,0,35,0,231,0,183,0,107,0,1,0,113,0,161,0,212,0,147,0,0,0,232,0,155,0,34,0,210,0,253,0,0,0,172,0,84,0,73,0,74,0,231,0,119,0,74,0,191,0,0,0,0,0,139,0,0,0,248,0,70,0,242,0,228,0,191,0,110,0,21,0,108,0,95,0,0,0,247,0,134,0,220,0,6,0,0,0,41,0,58,0,66,0,77,0,61,0,228,0,0,0,254,0,78,0,241,0,0,0,191,0,0,0,106,0,209,0,23,0,247,0,145,0,150,0,59,0,170,0,75,0,0,0,183,0,155,0,171,0,0,0,200,0,44,0,251,0,192,0,183,0,174,0,152,0,45,0,227,0,79,0,2,0,162,0,250,0,0,0,150,0,66,0,121,0,91,0,50,0,199,0,144,0,34,0,104,0,129,0,32,0,187,0,0,0,157,0,0,0,51,0,0,0,0,0,133,0,252,0,0,0,116,0,52,0,72,0,172,0,0,0,206,0,130,0,241,0,21,0,248,0,0,0,135,0,56,0,137,0,0,0,64,0,49,0,0,0,20,0,185,0,212,0,19,0,96,0,0,0,226,0,244,0,202,0,28,0,18,0,216,0,86,0,228,0,105,0,24,0,220,0,113,0,40,0,0,0,175,0,0,0,236,0,111,0,114,0,0,0,0,0,118,0,202,0,0,0,45,0);
signal scenario_full  : scenario_type := (21,31,57,31,164,31,35,31,231,31,183,31,107,31,1,31,113,31,161,31,212,31,147,31,147,30,232,31,155,31,34,31,210,31,253,31,253,30,172,31,84,31,73,31,74,31,231,31,119,31,74,31,191,31,191,30,191,29,139,31,139,30,248,31,70,31,242,31,228,31,191,31,110,31,21,31,108,31,95,31,95,30,247,31,134,31,220,31,6,31,6,30,41,31,58,31,66,31,77,31,61,31,228,31,228,30,254,31,78,31,241,31,241,30,191,31,191,30,106,31,209,31,23,31,247,31,145,31,150,31,59,31,170,31,75,31,75,30,183,31,155,31,171,31,171,30,200,31,44,31,251,31,192,31,183,31,174,31,152,31,45,31,227,31,79,31,2,31,162,31,250,31,250,30,150,31,66,31,121,31,91,31,50,31,199,31,144,31,34,31,104,31,129,31,32,31,187,31,187,30,157,31,157,30,51,31,51,30,51,29,133,31,252,31,252,30,116,31,52,31,72,31,172,31,172,30,206,31,130,31,241,31,21,31,248,31,248,30,135,31,56,31,137,31,137,30,64,31,49,31,49,30,20,31,185,31,212,31,19,31,96,31,96,30,226,31,244,31,202,31,28,31,18,31,216,31,86,31,228,31,105,31,24,31,220,31,113,31,40,31,40,30,175,31,175,30,236,31,111,31,114,31,114,30,114,29,118,31,202,31,202,30,45,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
