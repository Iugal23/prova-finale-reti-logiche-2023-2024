-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_922 is
end project_tb_922;

architecture project_tb_arch_922 of project_tb_922 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (46,0,0,0,0,0,245,0,48,0,45,0,141,0,39,0,0,0,20,0,14,0,50,0,43,0,0,0,135,0,0,0,85,0,141,0,131,0,151,0,73,0,145,0,137,0,88,0,0,0,9,0,186,0,145,0,0,0,21,0,0,0,229,0,0,0,0,0,99,0,243,0,60,0,233,0,188,0,153,0,29,0,0,0,0,0,157,0,48,0,0,0,83,0,104,0,195,0,164,0,151,0,0,0,218,0,68,0,85,0,202,0,77,0,116,0,156,0,82,0,10,0,169,0,142,0,0,0,73,0,27,0,0,0,7,0,32,0,89,0,230,0,191,0,85,0,225,0,0,0,0,0,41,0,205,0,107,0,167,0,0,0,0,0,241,0,122,0,187,0,159,0,69,0,0,0,110,0,0,0,109,0,140,0,0,0,0,0,137,0,88,0,0,0,130,0,56,0,123,0,10,0,194,0,236,0,102,0,200,0,0,0,152,0,162,0,30,0,144,0,186,0,160,0,252,0,251,0,242,0,0,0,56,0,218,0,97,0,171,0,0,0,142,0,208,0,221,0,0,0,0,0,158,0,125,0,0,0,252,0,97,0,0,0,170,0,7,0,105,0,199,0,190,0,0,0,0,0,138,0,135,0,72,0,69,0,218,0,18,0,9,0,128,0,96,0,0,0,19,0,0,0,248,0,13,0,149,0,0,0,91,0,0,0,129,0,179,0,162,0,114,0,177,0,157,0,0,0,74,0,240,0,178,0,0,0,86,0,210,0,192,0,209,0,0,0,62,0,240,0,31,0,0,0,0,0,112,0,55,0,0,0,143,0,77,0,67,0,46,0,0,0,239,0,119,0,82,0,253,0,100,0,208,0,85,0,33,0,182,0,46,0,184,0,0,0,197,0,53,0,0,0,0,0,218,0,105,0,202,0,22,0,193,0,40,0,177,0,241,0,0,0,202,0,208,0,24,0,235,0,76,0,107,0,130,0,184,0,249,0,52,0,58,0,139,0,58,0,205,0,0,0,114,0,47,0,241,0,147,0,96,0,230,0,246,0,218,0,0,0,151,0,205,0,0,0,189,0,0,0,165,0,70,0,162,0,135,0,246,0,165,0,102,0,133,0,132,0,104,0,0,0,53,0,180,0,159,0,225,0,69,0,0,0,0,0,210,0,13,0,69,0,58,0,209,0,87,0,0,0,0,0,0,0,105,0,17,0,163,0,0,0,0,0,3,0,90,0,220,0,225,0,75,0,238,0,160,0,107,0,45,0,0,0,0,0,235,0,168,0,241,0,69,0,97,0,182,0,6,0,54,0,0,0,0,0,236,0,35,0,51,0,0,0,4,0,0,0,188,0,46,0,24,0,48,0,232,0,211,0,45,0,122,0,222,0,216,0,0,0,196,0,0,0,121,0,0,0,27,0,243,0,77,0,48,0,242,0,164,0,0,0,207,0,0,0,0,0,167,0,28,0,239,0,223,0,62,0,223,0,221,0,180,0,158,0,20,0,0,0,52,0,113,0,125,0,126,0,7,0,245,0,138,0,14,0,152,0,149,0,40,0,159,0,14,0,44,0,199,0,248,0,180,0,15,0,0,0,116,0,0,0,171,0,209,0,76,0,48,0,222,0,188,0,120,0,0,0,107,0,145,0,0,0,36,0,30,0,0,0,175,0,0,0,204,0,109,0,106,0,31,0,103,0,0,0,77,0,0,0,0,0,8,0,245,0,0,0,0,0,0,0,143,0,95,0,111,0,132,0,210,0,0,0,234,0,0,0,182,0,65,0,0,0,118,0,52,0,209,0,240,0,198,0,180,0,230,0,114,0,181,0,246,0,239,0,122,0,226,0,229,0,113,0,135,0,223,0,26,0,0,0,221,0,81,0,41,0,28,0,235,0,122,0,186,0,203,0,239,0,43,0,28,0,126,0,0,0,24,0,248,0,251,0,68,0,127,0,50,0,48,0,0,0,21,0,0,0,0,0,62,0,43,0,0,0,102,0,35,0,131,0,149,0,85,0,0,0,241,0,76,0,109,0,71,0,244,0,0,0,116,0,97,0,15,0,130,0,89,0,27,0,15,0,128,0,253,0,56,0,239,0,185,0,255,0,221,0,0,0,238,0,244,0,40,0,90,0,144,0,89,0,112,0,151,0,192,0,169,0,93,0,186,0,124,0,21,0,239,0,195,0,0,0,0,0,151,0,193,0,178,0,221,0,225,0,0,0,7,0,200,0,0,0,60,0,168,0,203,0,0,0,112,0,225,0,236,0,231,0,113,0,147,0,241,0,134,0,0,0,120,0,0,0,128,0,56,0,30,0,197,0,222,0,37,0,199,0,71,0,203,0,0,0,229,0,195,0,188,0,13,0,236,0,194,0,123,0,129,0,205,0,86,0,210,0,218,0,105,0,0,0,0,0,214,0,0,0,86,0,125,0,207,0,18,0,215,0,49,0,22,0,237,0,245,0,0,0,0,0,61,0,0,0,37,0,105,0,64,0,100,0,14,0,36,0,60,0,43,0,0,0,1,0,234,0,111,0,0,0,98,0,228,0,78,0,0,0,118,0,23,0,0,0,0,0,104,0,0,0,0,0,168,0,35,0,137,0,8,0,181,0,0,0,91,0,68,0,0,0,103,0,0,0,183,0,179,0,104,0,0,0,0,0,113,0,219,0,68,0,155,0,194,0,153,0,175,0,198,0,4,0,0,0,85,0,148,0,246,0,81,0,235,0,200,0,67,0,172,0,191,0,178,0,199,0,236,0,15,0,255,0,23,0,164,0,0,0,13,0,45,0,0,0,0,0,193,0,35,0,229,0,8,0,247,0,0,0,154,0,81,0,236,0,38,0,0,0,119,0,0,0,5,0,131,0,0,0,201,0,95,0,232,0,251,0,34,0,215,0,29,0,0,0,37,0,117,0,229,0,195,0,194,0,146,0,0,0,251,0,47,0,108,0,101,0,0,0,176,0,232,0,0,0,216,0,202,0,0,0,98,0,0,0,171,0,95,0,179,0,166,0,0,0,0,0,207,0,187,0,121,0,212,0,100,0,0,0,0,0,158,0,86,0,66,0,0,0,184,0,253,0,178,0,0,0,252,0,247,0,87,0,149,0,111,0,167,0,236,0,107,0,235,0,164,0,120,0,72,0,12,0,121,0,235,0,2,0,0,0,217,0,88,0,193,0,249,0,75,0,0,0,100,0,178,0,0,0,96,0,219,0,119,0,58,0,98,0,174,0,248,0,21,0,0,0,0,0,99,0,93,0,181,0,0,0,0,0,0,0,218,0,168,0,159,0,243,0,223,0,98,0,50,0,150,0,82,0,167,0,0,0,152,0,194,0,17,0,243,0,236,0,124,0,0,0,131,0,52,0,0,0,11,0,243,0,124,0,128,0,250,0,88,0,248,0,28,0,147,0,223,0,12,0,126,0,98,0,134,0,0,0,0,0,102,0,203,0,34,0,160,0,196,0,22,0,5,0,175,0,0,0,0,0,222,0,233,0,163,0,100,0,238,0,199,0,74,0,0,0,32,0,229,0,196,0,198,0,115,0,171,0,83,0,23,0,54,0,27,0,161,0,238,0,254,0,187,0,0,0,174,0,144,0,233,0,25,0,246,0,55,0,8,0,185,0,24,0,85,0,0,0,0,0,0,0,0,0,88,0,0,0,160,0,19,0,100,0,215,0,28,0,165,0,0,0,192,0,244,0,231,0,20,0,0,0,210,0,0,0,94,0,34,0,0,0,135,0,11,0,100,0,42,0,191,0,156,0,0,0,105,0,108,0,99,0,48,0,178,0,0,0,121,0,0,0,0,0,20,0,0,0,101,0,37,0,0,0,81,0,0,0,0,0,178,0,153,0,132,0,180,0,156,0,46,0,0,0,190,0,6,0,126,0,186,0,116,0,52,0,149,0,0,0,70,0,0,0,29,0,0,0,103,0,0,0,186,0,194,0,240,0,95,0,180,0,96,0,140,0,93,0,0,0,253,0,184,0,23,0,46,0,168,0,204,0,180,0,20,0,196,0,194,0,158,0,210,0,0,0,0,0,48,0,0,0,253,0,78,0,0,0,183,0,147,0,122,0,0,0,65,0,99,0,0,0,0,0,0,0,38,0,241,0,0,0,189,0,0,0,184,0,163,0,107,0,215,0,6,0,239,0,16,0,9,0,61,0,102,0,218,0,60,0,213,0,42,0,231,0,150,0,0,0,0,0,153,0,250,0,233,0,0,0,90,0,202,0,140,0,85,0,156,0,162,0,0,0,127,0,191,0,0,0,0,0,0,0,0,0,34,0,25,0,142,0,34,0,0,0,49,0,254,0,67,0,0,0,0,0,0,0,52,0,231,0,114,0,232,0,0,0,0,0,250,0,0,0,7,0);
signal scenario_full  : scenario_type := (46,31,46,30,46,29,245,31,48,31,45,31,141,31,39,31,39,30,20,31,14,31,50,31,43,31,43,30,135,31,135,30,85,31,141,31,131,31,151,31,73,31,145,31,137,31,88,31,88,30,9,31,186,31,145,31,145,30,21,31,21,30,229,31,229,30,229,29,99,31,243,31,60,31,233,31,188,31,153,31,29,31,29,30,29,29,157,31,48,31,48,30,83,31,104,31,195,31,164,31,151,31,151,30,218,31,68,31,85,31,202,31,77,31,116,31,156,31,82,31,10,31,169,31,142,31,142,30,73,31,27,31,27,30,7,31,32,31,89,31,230,31,191,31,85,31,225,31,225,30,225,29,41,31,205,31,107,31,167,31,167,30,167,29,241,31,122,31,187,31,159,31,69,31,69,30,110,31,110,30,109,31,140,31,140,30,140,29,137,31,88,31,88,30,130,31,56,31,123,31,10,31,194,31,236,31,102,31,200,31,200,30,152,31,162,31,30,31,144,31,186,31,160,31,252,31,251,31,242,31,242,30,56,31,218,31,97,31,171,31,171,30,142,31,208,31,221,31,221,30,221,29,158,31,125,31,125,30,252,31,97,31,97,30,170,31,7,31,105,31,199,31,190,31,190,30,190,29,138,31,135,31,72,31,69,31,218,31,18,31,9,31,128,31,96,31,96,30,19,31,19,30,248,31,13,31,149,31,149,30,91,31,91,30,129,31,179,31,162,31,114,31,177,31,157,31,157,30,74,31,240,31,178,31,178,30,86,31,210,31,192,31,209,31,209,30,62,31,240,31,31,31,31,30,31,29,112,31,55,31,55,30,143,31,77,31,67,31,46,31,46,30,239,31,119,31,82,31,253,31,100,31,208,31,85,31,33,31,182,31,46,31,184,31,184,30,197,31,53,31,53,30,53,29,218,31,105,31,202,31,22,31,193,31,40,31,177,31,241,31,241,30,202,31,208,31,24,31,235,31,76,31,107,31,130,31,184,31,249,31,52,31,58,31,139,31,58,31,205,31,205,30,114,31,47,31,241,31,147,31,96,31,230,31,246,31,218,31,218,30,151,31,205,31,205,30,189,31,189,30,165,31,70,31,162,31,135,31,246,31,165,31,102,31,133,31,132,31,104,31,104,30,53,31,180,31,159,31,225,31,69,31,69,30,69,29,210,31,13,31,69,31,58,31,209,31,87,31,87,30,87,29,87,28,105,31,17,31,163,31,163,30,163,29,3,31,90,31,220,31,225,31,75,31,238,31,160,31,107,31,45,31,45,30,45,29,235,31,168,31,241,31,69,31,97,31,182,31,6,31,54,31,54,30,54,29,236,31,35,31,51,31,51,30,4,31,4,30,188,31,46,31,24,31,48,31,232,31,211,31,45,31,122,31,222,31,216,31,216,30,196,31,196,30,121,31,121,30,27,31,243,31,77,31,48,31,242,31,164,31,164,30,207,31,207,30,207,29,167,31,28,31,239,31,223,31,62,31,223,31,221,31,180,31,158,31,20,31,20,30,52,31,113,31,125,31,126,31,7,31,245,31,138,31,14,31,152,31,149,31,40,31,159,31,14,31,44,31,199,31,248,31,180,31,15,31,15,30,116,31,116,30,171,31,209,31,76,31,48,31,222,31,188,31,120,31,120,30,107,31,145,31,145,30,36,31,30,31,30,30,175,31,175,30,204,31,109,31,106,31,31,31,103,31,103,30,77,31,77,30,77,29,8,31,245,31,245,30,245,29,245,28,143,31,95,31,111,31,132,31,210,31,210,30,234,31,234,30,182,31,65,31,65,30,118,31,52,31,209,31,240,31,198,31,180,31,230,31,114,31,181,31,246,31,239,31,122,31,226,31,229,31,113,31,135,31,223,31,26,31,26,30,221,31,81,31,41,31,28,31,235,31,122,31,186,31,203,31,239,31,43,31,28,31,126,31,126,30,24,31,248,31,251,31,68,31,127,31,50,31,48,31,48,30,21,31,21,30,21,29,62,31,43,31,43,30,102,31,35,31,131,31,149,31,85,31,85,30,241,31,76,31,109,31,71,31,244,31,244,30,116,31,97,31,15,31,130,31,89,31,27,31,15,31,128,31,253,31,56,31,239,31,185,31,255,31,221,31,221,30,238,31,244,31,40,31,90,31,144,31,89,31,112,31,151,31,192,31,169,31,93,31,186,31,124,31,21,31,239,31,195,31,195,30,195,29,151,31,193,31,178,31,221,31,225,31,225,30,7,31,200,31,200,30,60,31,168,31,203,31,203,30,112,31,225,31,236,31,231,31,113,31,147,31,241,31,134,31,134,30,120,31,120,30,128,31,56,31,30,31,197,31,222,31,37,31,199,31,71,31,203,31,203,30,229,31,195,31,188,31,13,31,236,31,194,31,123,31,129,31,205,31,86,31,210,31,218,31,105,31,105,30,105,29,214,31,214,30,86,31,125,31,207,31,18,31,215,31,49,31,22,31,237,31,245,31,245,30,245,29,61,31,61,30,37,31,105,31,64,31,100,31,14,31,36,31,60,31,43,31,43,30,1,31,234,31,111,31,111,30,98,31,228,31,78,31,78,30,118,31,23,31,23,30,23,29,104,31,104,30,104,29,168,31,35,31,137,31,8,31,181,31,181,30,91,31,68,31,68,30,103,31,103,30,183,31,179,31,104,31,104,30,104,29,113,31,219,31,68,31,155,31,194,31,153,31,175,31,198,31,4,31,4,30,85,31,148,31,246,31,81,31,235,31,200,31,67,31,172,31,191,31,178,31,199,31,236,31,15,31,255,31,23,31,164,31,164,30,13,31,45,31,45,30,45,29,193,31,35,31,229,31,8,31,247,31,247,30,154,31,81,31,236,31,38,31,38,30,119,31,119,30,5,31,131,31,131,30,201,31,95,31,232,31,251,31,34,31,215,31,29,31,29,30,37,31,117,31,229,31,195,31,194,31,146,31,146,30,251,31,47,31,108,31,101,31,101,30,176,31,232,31,232,30,216,31,202,31,202,30,98,31,98,30,171,31,95,31,179,31,166,31,166,30,166,29,207,31,187,31,121,31,212,31,100,31,100,30,100,29,158,31,86,31,66,31,66,30,184,31,253,31,178,31,178,30,252,31,247,31,87,31,149,31,111,31,167,31,236,31,107,31,235,31,164,31,120,31,72,31,12,31,121,31,235,31,2,31,2,30,217,31,88,31,193,31,249,31,75,31,75,30,100,31,178,31,178,30,96,31,219,31,119,31,58,31,98,31,174,31,248,31,21,31,21,30,21,29,99,31,93,31,181,31,181,30,181,29,181,28,218,31,168,31,159,31,243,31,223,31,98,31,50,31,150,31,82,31,167,31,167,30,152,31,194,31,17,31,243,31,236,31,124,31,124,30,131,31,52,31,52,30,11,31,243,31,124,31,128,31,250,31,88,31,248,31,28,31,147,31,223,31,12,31,126,31,98,31,134,31,134,30,134,29,102,31,203,31,34,31,160,31,196,31,22,31,5,31,175,31,175,30,175,29,222,31,233,31,163,31,100,31,238,31,199,31,74,31,74,30,32,31,229,31,196,31,198,31,115,31,171,31,83,31,23,31,54,31,27,31,161,31,238,31,254,31,187,31,187,30,174,31,144,31,233,31,25,31,246,31,55,31,8,31,185,31,24,31,85,31,85,30,85,29,85,28,85,27,88,31,88,30,160,31,19,31,100,31,215,31,28,31,165,31,165,30,192,31,244,31,231,31,20,31,20,30,210,31,210,30,94,31,34,31,34,30,135,31,11,31,100,31,42,31,191,31,156,31,156,30,105,31,108,31,99,31,48,31,178,31,178,30,121,31,121,30,121,29,20,31,20,30,101,31,37,31,37,30,81,31,81,30,81,29,178,31,153,31,132,31,180,31,156,31,46,31,46,30,190,31,6,31,126,31,186,31,116,31,52,31,149,31,149,30,70,31,70,30,29,31,29,30,103,31,103,30,186,31,194,31,240,31,95,31,180,31,96,31,140,31,93,31,93,30,253,31,184,31,23,31,46,31,168,31,204,31,180,31,20,31,196,31,194,31,158,31,210,31,210,30,210,29,48,31,48,30,253,31,78,31,78,30,183,31,147,31,122,31,122,30,65,31,99,31,99,30,99,29,99,28,38,31,241,31,241,30,189,31,189,30,184,31,163,31,107,31,215,31,6,31,239,31,16,31,9,31,61,31,102,31,218,31,60,31,213,31,42,31,231,31,150,31,150,30,150,29,153,31,250,31,233,31,233,30,90,31,202,31,140,31,85,31,156,31,162,31,162,30,127,31,191,31,191,30,191,29,191,28,191,27,34,31,25,31,142,31,34,31,34,30,49,31,254,31,67,31,67,30,67,29,67,28,52,31,231,31,114,31,232,31,232,30,232,29,250,31,250,30,7,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
