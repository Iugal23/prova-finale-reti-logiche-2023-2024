-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 898;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,223,0,25,0,125,0,25,0,138,0,4,0,0,0,195,0,141,0,230,0,132,0,0,0,161,0,153,0,248,0,107,0,204,0,225,0,0,0,217,0,160,0,120,0,0,0,16,0,241,0,172,0,242,0,0,0,0,0,105,0,202,0,249,0,163,0,116,0,164,0,120,0,37,0,0,0,133,0,89,0,19,0,55,0,155,0,113,0,0,0,86,0,190,0,123,0,237,0,82,0,0,0,173,0,139,0,126,0,0,0,121,0,17,0,174,0,132,0,194,0,0,0,193,0,87,0,214,0,36,0,67,0,208,0,1,0,0,0,60,0,238,0,154,0,68,0,20,0,125,0,173,0,160,0,177,0,0,0,17,0,0,0,230,0,94,0,43,0,223,0,0,0,222,0,0,0,201,0,38,0,0,0,87,0,31,0,12,0,34,0,198,0,164,0,41,0,55,0,233,0,53,0,0,0,0,0,15,0,191,0,0,0,204,0,59,0,183,0,200,0,232,0,113,0,66,0,5,0,195,0,0,0,229,0,0,0,102,0,0,0,192,0,225,0,115,0,182,0,241,0,61,0,0,0,193,0,0,0,130,0,0,0,21,0,248,0,254,0,40,0,123,0,221,0,22,0,191,0,0,0,141,0,0,0,18,0,0,0,162,0,45,0,0,0,171,0,0,0,73,0,91,0,48,0,181,0,0,0,0,0,14,0,0,0,85,0,197,0,0,0,45,0,248,0,0,0,0,0,0,0,0,0,63,0,0,0,53,0,0,0,188,0,252,0,58,0,166,0,0,0,60,0,13,0,0,0,0,0,116,0,89,0,0,0,0,0,36,0,229,0,15,0,40,0,59,0,208,0,20,0,0,0,253,0,0,0,44,0,62,0,243,0,167,0,0,0,0,0,160,0,54,0,147,0,128,0,116,0,108,0,0,0,114,0,235,0,104,0,15,0,103,0,13,0,246,0,124,0,0,0,18,0,0,0,203,0,75,0,54,0,251,0,0,0,0,0,151,0,30,0,18,0,0,0,192,0,223,0,124,0,86,0,245,0,149,0,109,0,0,0,106,0,0,0,110,0,102,0,17,0,35,0,177,0,17,0,117,0,135,0,95,0,189,0,181,0,221,0,28,0,159,0,228,0,104,0,253,0,0,0,127,0,95,0,0,0,73,0,152,0,244,0,145,0,0,0,0,0,145,0,0,0,161,0,0,0,0,0,50,0,0,0,0,0,0,0,72,0,74,0,209,0,99,0,165,0,0,0,0,0,97,0,101,0,55,0,192,0,196,0,48,0,0,0,0,0,71,0,200,0,0,0,161,0,47,0,199,0,210,0,190,0,0,0,96,0,86,0,30,0,75,0,77,0,127,0,149,0,0,0,0,0,37,0,15,0,144,0,226,0,18,0,120,0,0,0,180,0,75,0,104,0,142,0,163,0,0,0,0,0,234,0,0,0,116,0,163,0,0,0,58,0,126,0,8,0,0,0,0,0,67,0,0,0,89,0,52,0,60,0,112,0,135,0,163,0,108,0,73,0,253,0,0,0,214,0,179,0,197,0,37,0,0,0,0,0,244,0,110,0,95,0,53,0,212,0,213,0,26,0,172,0,32,0,0,0,172,0,157,0,55,0,73,0,163,0,138,0,106,0,139,0,113,0,142,0,145,0,109,0,81,0,168,0,118,0,69,0,152,0,192,0,52,0,0,0,164,0,225,0,46,0,0,0,8,0,169,0,171,0,122,0,189,0,234,0,210,0,214,0,99,0,0,0,80,0,247,0,190,0,240,0,237,0,33,0,249,0,152,0,91,0,162,0,85,0,0,0,44,0,78,0,113,0,238,0,255,0,183,0,0,0,50,0,0,0,192,0,131,0,95,0,154,0,0,0,18,0,187,0,152,0,109,0,101,0,33,0,120,0,137,0,0,0,69,0,57,0,198,0,0,0,211,0,11,0,37,0,247,0,0,0,100,0,173,0,62,0,208,0,5,0,15,0,19,0,0,0,0,0,120,0,219,0,185,0,45,0,209,0,113,0,66,0,238,0,24,0,0,0,218,0,75,0,59,0,84,0,164,0,1,0,0,0,175,0,166,0,165,0,0,0,71,0,154,0,128,0,37,0,0,0,81,0,133,0,0,0,182,0,100,0,136,0,40,0,222,0,0,0,189,0,36,0,0,0,108,0,141,0,25,0,100,0,86,0,0,0,99,0,130,0,109,0,26,0,0,0,14,0,69,0,135,0,125,0,55,0,134,0,92,0,0,0,159,0,216,0,165,0,0,0,105,0,166,0,0,0,224,0,6,0,153,0,0,0,253,0,81,0,143,0,68,0,194,0,71,0,0,0,178,0,0,0,219,0,0,0,54,0,85,0,46,0,0,0,60,0,0,0,150,0,70,0,146,0,244,0,173,0,115,0,204,0,85,0,70,0,11,0,137,0,24,0,172,0,126,0,55,0,156,0,49,0,105,0,99,0,212,0,71,0,0,0,170,0,45,0,100,0,246,0,51,0,210,0,142,0,188,0,154,0,79,0,180,0,39,0,64,0,21,0,251,0,0,0,156,0,122,0,66,0,75,0,135,0,41,0,27,0,117,0,125,0,110,0,245,0,0,0,37,0,34,0,161,0,134,0,55,0,208,0,85,0,200,0,134,0,0,0,88,0,181,0,61,0,232,0,134,0,168,0,217,0,68,0,60,0,153,0,54,0,0,0,121,0,17,0,0,0,56,0,75,0,42,0,76,0,98,0,190,0,167,0,0,0,218,0,0,0,113,0,152,0,13,0,227,0,0,0,231,0,0,0,94,0,69,0,0,0,240,0,7,0,197,0,112,0,0,0,52,0,18,0,0,0,0,0,225,0,162,0,206,0,108,0,221,0,58,0,228,0,224,0,48,0,114,0,111,0,31,0,153,0,0,0,0,0,14,0,111,0,200,0,34,0,87,0,236,0,82,0,6,0,249,0,27,0,9,0,0,0,0,0,80,0,49,0,94,0,78,0,0,0,13,0,175,0,139,0,193,0,130,0,0,0,5,0,213,0,0,0,86,0,0,0,28,0,0,0,249,0,0,0,122,0,107,0,38,0,222,0,246,0,57,0,124,0,119,0,99,0,202,0,101,0,124,0,55,0,170,0,0,0,226,0,0,0,92,0,27,0,87,0,166,0,0,0,13,0,202,0,114,0,8,0,4,0,169,0,218,0,40,0,172,0,98,0,79,0,145,0,0,0,0,0,249,0,0,0,12,0,248,0,0,0,250,0,140,0,0,0,140,0,96,0,200,0,14,0,86,0,0,0,227,0,255,0,152,0,29,0,251,0,42,0,161,0,203,0,10,0,0,0,39,0,0,0,168,0,34,0,45,0,35,0,254,0,244,0,251,0,48,0,154,0,100,0,0,0,174,0,142,0,119,0,232,0,44,0,24,0,231,0,49,0,0,0,71,0,149,0,111,0,190,0,42,0,79,0,210,0,236,0,67,0,0,0,165,0,111,0,147,0,141,0,253,0,130,0,168,0,23,0,193,0,0,0,199,0,0,0,91,0,185,0,23,0,167,0,52,0,0,0,0,0,109,0,68,0,216,0,146,0,33,0,122,0,0,0,70,0,188,0,127,0,0,0,0,0,120,0,153,0,108,0,57,0,227,0,170,0,172,0,196,0,0,0,0,0,249,0,0,0,17,0,126,0,204,0,0,0,28,0,174,0,162,0,0,0,221,0,246,0,0,0,127,0,242,0,215,0,0,0,61,0,180,0,0,0,79,0,115,0,137,0,5,0,122,0,0,0,52,0,64,0,0,0,85,0,249,0,12,0,100,0,0,0,170,0,117,0,24,0,181,0,209,0,131,0,83,0,179,0,4,0,134,0,21,0,163,0,154,0,0,0,1,0,0,0,214,0,19,0,95,0,226,0,4,0,249,0,87,0,238,0,197,0,154,0,244,0,184,0,0,0,0,0,0,0,0,0,232,0,166,0,62,0,123,0,109,0,0,0,84,0,0,0,0,0,0,0,0,0,0,0,112,0,158,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,223,31,25,31,125,31,25,31,138,31,4,31,4,30,195,31,141,31,230,31,132,31,132,30,161,31,153,31,248,31,107,31,204,31,225,31,225,30,217,31,160,31,120,31,120,30,16,31,241,31,172,31,242,31,242,30,242,29,105,31,202,31,249,31,163,31,116,31,164,31,120,31,37,31,37,30,133,31,89,31,19,31,55,31,155,31,113,31,113,30,86,31,190,31,123,31,237,31,82,31,82,30,173,31,139,31,126,31,126,30,121,31,17,31,174,31,132,31,194,31,194,30,193,31,87,31,214,31,36,31,67,31,208,31,1,31,1,30,60,31,238,31,154,31,68,31,20,31,125,31,173,31,160,31,177,31,177,30,17,31,17,30,230,31,94,31,43,31,223,31,223,30,222,31,222,30,201,31,38,31,38,30,87,31,31,31,12,31,34,31,198,31,164,31,41,31,55,31,233,31,53,31,53,30,53,29,15,31,191,31,191,30,204,31,59,31,183,31,200,31,232,31,113,31,66,31,5,31,195,31,195,30,229,31,229,30,102,31,102,30,192,31,225,31,115,31,182,31,241,31,61,31,61,30,193,31,193,30,130,31,130,30,21,31,248,31,254,31,40,31,123,31,221,31,22,31,191,31,191,30,141,31,141,30,18,31,18,30,162,31,45,31,45,30,171,31,171,30,73,31,91,31,48,31,181,31,181,30,181,29,14,31,14,30,85,31,197,31,197,30,45,31,248,31,248,30,248,29,248,28,248,27,63,31,63,30,53,31,53,30,188,31,252,31,58,31,166,31,166,30,60,31,13,31,13,30,13,29,116,31,89,31,89,30,89,29,36,31,229,31,15,31,40,31,59,31,208,31,20,31,20,30,253,31,253,30,44,31,62,31,243,31,167,31,167,30,167,29,160,31,54,31,147,31,128,31,116,31,108,31,108,30,114,31,235,31,104,31,15,31,103,31,13,31,246,31,124,31,124,30,18,31,18,30,203,31,75,31,54,31,251,31,251,30,251,29,151,31,30,31,18,31,18,30,192,31,223,31,124,31,86,31,245,31,149,31,109,31,109,30,106,31,106,30,110,31,102,31,17,31,35,31,177,31,17,31,117,31,135,31,95,31,189,31,181,31,221,31,28,31,159,31,228,31,104,31,253,31,253,30,127,31,95,31,95,30,73,31,152,31,244,31,145,31,145,30,145,29,145,31,145,30,161,31,161,30,161,29,50,31,50,30,50,29,50,28,72,31,74,31,209,31,99,31,165,31,165,30,165,29,97,31,101,31,55,31,192,31,196,31,48,31,48,30,48,29,71,31,200,31,200,30,161,31,47,31,199,31,210,31,190,31,190,30,96,31,86,31,30,31,75,31,77,31,127,31,149,31,149,30,149,29,37,31,15,31,144,31,226,31,18,31,120,31,120,30,180,31,75,31,104,31,142,31,163,31,163,30,163,29,234,31,234,30,116,31,163,31,163,30,58,31,126,31,8,31,8,30,8,29,67,31,67,30,89,31,52,31,60,31,112,31,135,31,163,31,108,31,73,31,253,31,253,30,214,31,179,31,197,31,37,31,37,30,37,29,244,31,110,31,95,31,53,31,212,31,213,31,26,31,172,31,32,31,32,30,172,31,157,31,55,31,73,31,163,31,138,31,106,31,139,31,113,31,142,31,145,31,109,31,81,31,168,31,118,31,69,31,152,31,192,31,52,31,52,30,164,31,225,31,46,31,46,30,8,31,169,31,171,31,122,31,189,31,234,31,210,31,214,31,99,31,99,30,80,31,247,31,190,31,240,31,237,31,33,31,249,31,152,31,91,31,162,31,85,31,85,30,44,31,78,31,113,31,238,31,255,31,183,31,183,30,50,31,50,30,192,31,131,31,95,31,154,31,154,30,18,31,187,31,152,31,109,31,101,31,33,31,120,31,137,31,137,30,69,31,57,31,198,31,198,30,211,31,11,31,37,31,247,31,247,30,100,31,173,31,62,31,208,31,5,31,15,31,19,31,19,30,19,29,120,31,219,31,185,31,45,31,209,31,113,31,66,31,238,31,24,31,24,30,218,31,75,31,59,31,84,31,164,31,1,31,1,30,175,31,166,31,165,31,165,30,71,31,154,31,128,31,37,31,37,30,81,31,133,31,133,30,182,31,100,31,136,31,40,31,222,31,222,30,189,31,36,31,36,30,108,31,141,31,25,31,100,31,86,31,86,30,99,31,130,31,109,31,26,31,26,30,14,31,69,31,135,31,125,31,55,31,134,31,92,31,92,30,159,31,216,31,165,31,165,30,105,31,166,31,166,30,224,31,6,31,153,31,153,30,253,31,81,31,143,31,68,31,194,31,71,31,71,30,178,31,178,30,219,31,219,30,54,31,85,31,46,31,46,30,60,31,60,30,150,31,70,31,146,31,244,31,173,31,115,31,204,31,85,31,70,31,11,31,137,31,24,31,172,31,126,31,55,31,156,31,49,31,105,31,99,31,212,31,71,31,71,30,170,31,45,31,100,31,246,31,51,31,210,31,142,31,188,31,154,31,79,31,180,31,39,31,64,31,21,31,251,31,251,30,156,31,122,31,66,31,75,31,135,31,41,31,27,31,117,31,125,31,110,31,245,31,245,30,37,31,34,31,161,31,134,31,55,31,208,31,85,31,200,31,134,31,134,30,88,31,181,31,61,31,232,31,134,31,168,31,217,31,68,31,60,31,153,31,54,31,54,30,121,31,17,31,17,30,56,31,75,31,42,31,76,31,98,31,190,31,167,31,167,30,218,31,218,30,113,31,152,31,13,31,227,31,227,30,231,31,231,30,94,31,69,31,69,30,240,31,7,31,197,31,112,31,112,30,52,31,18,31,18,30,18,29,225,31,162,31,206,31,108,31,221,31,58,31,228,31,224,31,48,31,114,31,111,31,31,31,153,31,153,30,153,29,14,31,111,31,200,31,34,31,87,31,236,31,82,31,6,31,249,31,27,31,9,31,9,30,9,29,80,31,49,31,94,31,78,31,78,30,13,31,175,31,139,31,193,31,130,31,130,30,5,31,213,31,213,30,86,31,86,30,28,31,28,30,249,31,249,30,122,31,107,31,38,31,222,31,246,31,57,31,124,31,119,31,99,31,202,31,101,31,124,31,55,31,170,31,170,30,226,31,226,30,92,31,27,31,87,31,166,31,166,30,13,31,202,31,114,31,8,31,4,31,169,31,218,31,40,31,172,31,98,31,79,31,145,31,145,30,145,29,249,31,249,30,12,31,248,31,248,30,250,31,140,31,140,30,140,31,96,31,200,31,14,31,86,31,86,30,227,31,255,31,152,31,29,31,251,31,42,31,161,31,203,31,10,31,10,30,39,31,39,30,168,31,34,31,45,31,35,31,254,31,244,31,251,31,48,31,154,31,100,31,100,30,174,31,142,31,119,31,232,31,44,31,24,31,231,31,49,31,49,30,71,31,149,31,111,31,190,31,42,31,79,31,210,31,236,31,67,31,67,30,165,31,111,31,147,31,141,31,253,31,130,31,168,31,23,31,193,31,193,30,199,31,199,30,91,31,185,31,23,31,167,31,52,31,52,30,52,29,109,31,68,31,216,31,146,31,33,31,122,31,122,30,70,31,188,31,127,31,127,30,127,29,120,31,153,31,108,31,57,31,227,31,170,31,172,31,196,31,196,30,196,29,249,31,249,30,17,31,126,31,204,31,204,30,28,31,174,31,162,31,162,30,221,31,246,31,246,30,127,31,242,31,215,31,215,30,61,31,180,31,180,30,79,31,115,31,137,31,5,31,122,31,122,30,52,31,64,31,64,30,85,31,249,31,12,31,100,31,100,30,170,31,117,31,24,31,181,31,209,31,131,31,83,31,179,31,4,31,134,31,21,31,163,31,154,31,154,30,1,31,1,30,214,31,19,31,95,31,226,31,4,31,249,31,87,31,238,31,197,31,154,31,244,31,184,31,184,30,184,29,184,28,184,27,232,31,166,31,62,31,123,31,109,31,109,30,84,31,84,30,84,29,84,28,84,27,84,26,112,31,158,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
