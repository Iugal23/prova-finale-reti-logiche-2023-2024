-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_620 is
end project_tb_620;

architecture project_tb_arch_620 of project_tb_620 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1001;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,192,0,0,0,0,0,23,0,139,0,46,0,42,0,103,0,220,0,221,0,44,0,0,0,91,0,0,0,31,0,0,0,168,0,220,0,251,0,126,0,103,0,74,0,0,0,63,0,0,0,246,0,61,0,0,0,162,0,0,0,0,0,101,0,97,0,195,0,121,0,80,0,154,0,0,0,0,0,0,0,191,0,41,0,27,0,0,0,25,0,171,0,237,0,84,0,214,0,252,0,110,0,240,0,195,0,20,0,251,0,189,0,0,0,64,0,129,0,0,0,60,0,57,0,78,0,0,0,255,0,0,0,118,0,210,0,113,0,0,0,6,0,30,0,172,0,208,0,211,0,15,0,76,0,0,0,0,0,58,0,86,0,22,0,0,0,122,0,223,0,45,0,238,0,134,0,114,0,9,0,225,0,5,0,110,0,151,0,11,0,0,0,0,0,86,0,165,0,217,0,96,0,41,0,0,0,204,0,97,0,145,0,81,0,242,0,196,0,152,0,89,0,103,0,136,0,221,0,251,0,76,0,136,0,163,0,154,0,234,0,85,0,196,0,0,0,3,0,182,0,156,0,146,0,222,0,16,0,193,0,215,0,134,0,191,0,235,0,0,0,222,0,80,0,44,0,145,0,94,0,226,0,178,0,229,0,28,0,79,0,240,0,149,0,181,0,0,0,173,0,0,0,14,0,64,0,184,0,241,0,156,0,0,0,252,0,114,0,175,0,144,0,141,0,0,0,48,0,93,0,75,0,3,0,179,0,6,0,253,0,34,0,136,0,148,0,0,0,121,0,1,0,90,0,20,0,235,0,134,0,16,0,0,0,181,0,0,0,120,0,0,0,0,0,0,0,94,0,108,0,0,0,144,0,183,0,243,0,202,0,163,0,37,0,82,0,120,0,155,0,126,0,207,0,0,0,65,0,53,0,243,0,0,0,123,0,241,0,95,0,86,0,51,0,154,0,154,0,59,0,93,0,47,0,234,0,0,0,149,0,162,0,0,0,0,0,117,0,130,0,170,0,159,0,63,0,46,0,54,0,2,0,0,0,205,0,83,0,61,0,209,0,52,0,23,0,241,0,58,0,125,0,0,0,0,0,43,0,107,0,252,0,94,0,137,0,137,0,134,0,164,0,161,0,199,0,0,0,0,0,242,0,27,0,206,0,0,0,27,0,54,0,57,0,220,0,44,0,0,0,130,0,239,0,176,0,139,0,0,0,111,0,78,0,203,0,0,0,171,0,148,0,11,0,161,0,119,0,0,0,85,0,95,0,218,0,0,0,151,0,133,0,182,0,116,0,38,0,0,0,165,0,73,0,8,0,146,0,3,0,0,0,251,0,104,0,0,0,107,0,66,0,216,0,40,0,107,0,217,0,184,0,189,0,234,0,0,0,204,0,106,0,179,0,13,0,0,0,253,0,12,0,36,0,52,0,226,0,82,0,247,0,44,0,0,0,161,0,248,0,76,0,176,0,12,0,0,0,0,0,128,0,162,0,131,0,2,0,97,0,0,0,0,0,23,0,138,0,131,0,0,0,0,0,27,0,51,0,134,0,122,0,207,0,34,0,0,0,252,0,169,0,0,0,221,0,208,0,95,0,64,0,139,0,218,0,127,0,51,0,0,0,241,0,0,0,156,0,84,0,0,0,21,0,0,0,51,0,128,0,112,0,65,0,75,0,96,0,0,0,0,0,241,0,71,0,136,0,75,0,0,0,26,0,51,0,105,0,0,0,75,0,19,0,17,0,229,0,100,0,151,0,88,0,99,0,190,0,0,0,0,0,75,0,15,0,215,0,167,0,72,0,130,0,0,0,171,0,52,0,158,0,0,0,179,0,252,0,37,0,128,0,204,0,230,0,0,0,0,0,0,0,225,0,70,0,64,0,79,0,165,0,0,0,0,0,0,0,229,0,187,0,155,0,246,0,68,0,40,0,75,0,150,0,36,0,167,0,12,0,67,0,0,0,76,0,105,0,105,0,19,0,84,0,81,0,30,0,62,0,0,0,198,0,18,0,57,0,20,0,15,0,8,0,115,0,242,0,0,0,216,0,0,0,249,0,0,0,161,0,76,0,234,0,53,0,0,0,233,0,139,0,30,0,89,0,76,0,229,0,239,0,62,0,0,0,9,0,155,0,66,0,0,0,220,0,0,0,226,0,122,0,34,0,0,0,201,0,12,0,112,0,229,0,242,0,182,0,194,0,137,0,226,0,127,0,0,0,63,0,176,0,255,0,11,0,34,0,188,0,0,0,9,0,187,0,21,0,0,0,8,0,55,0,255,0,76,0,14,0,54,0,1,0,81,0,182,0,0,0,97,0,10,0,48,0,189,0,123,0,6,0,110,0,18,0,98,0,22,0,168,0,54,0,39,0,41,0,92,0,46,0,49,0,177,0,145,0,47,0,51,0,15,0,25,0,39,0,66,0,0,0,53,0,65,0,106,0,110,0,174,0,169,0,0,0,81,0,104,0,58,0,70,0,71,0,0,0,206,0,199,0,0,0,253,0,98,0,47,0,78,0,0,0,125,0,146,0,66,0,167,0,202,0,148,0,225,0,106,0,85,0,153,0,0,0,55,0,222,0,178,0,96,0,41,0,24,0,122,0,85,0,75,0,163,0,214,0,3,0,0,0,0,0,0,0,41,0,120,0,255,0,82,0,223,0,160,0,49,0,0,0,219,0,18,0,190,0,252,0,35,0,0,0,0,0,214,0,233,0,110,0,176,0,1,0,114,0,95,0,175,0,36,0,49,0,198,0,0,0,0,0,224,0,101,0,0,0,0,0,99,0,100,0,31,0,0,0,0,0,224,0,171,0,43,0,155,0,74,0,0,0,52,0,246,0,0,0,162,0,223,0,225,0,0,0,2,0,221,0,218,0,183,0,0,0,184,0,0,0,162,0,84,0,226,0,0,0,120,0,54,0,68,0,0,0,206,0,164,0,192,0,0,0,0,0,250,0,0,0,8,0,97,0,79,0,235,0,207,0,61,0,171,0,125,0,132,0,145,0,0,0,177,0,0,0,0,0,0,0,130,0,0,0,12,0,218,0,0,0,222,0,0,0,131,0,206,0,0,0,0,0,79,0,98,0,14,0,210,0,0,0,41,0,0,0,232,0,177,0,45,0,0,0,156,0,5,0,123,0,45,0,127,0,60,0,115,0,39,0,17,0,152,0,216,0,248,0,26,0,242,0,77,0,0,0,16,0,42,0,0,0,0,0,63,0,123,0,0,0,30,0,0,0,56,0,39,0,46,0,18,0,0,0,7,0,222,0,207,0,161,0,111,0,173,0,5,0,152,0,212,0,151,0,0,0,70,0,48,0,0,0,35,0,213,0,196,0,149,0,154,0,35,0,61,0,168,0,0,0,154,0,115,0,53,0,0,0,96,0,18,0,0,0,0,0,38,0,92,0,73,0,71,0,160,0,242,0,225,0,232,0,132,0,0,0,0,0,54,0,229,0,0,0,221,0,0,0,144,0,0,0,35,0,190,0,166,0,0,0,103,0,0,0,142,0,10,0,43,0,156,0,196,0,133,0,34,0,13,0,121,0,186,0,0,0,238,0,160,0,0,0,39,0,0,0,0,0,0,0,78,0,39,0,147,0,227,0,86,0,82,0,0,0,13,0,182,0,249,0,110,0,40,0,108,0,45,0,198,0,209,0,123,0,0,0,171,0,34,0,99,0,178,0,194,0,170,0,0,0,0,0,0,0,16,0,132,0,122,0,184,0,67,0,62,0,165,0,87,0,46,0,0,0,34,0,62,0,0,0,143,0,160,0,83,0,0,0,0,0,101,0,161,0,37,0,182,0,237,0,95,0,243,0,0,0,93,0,8,0,65,0,46,0,37,0,0,0,254,0,147,0,0,0,224,0,54,0,0,0,105,0,243,0,217,0,83,0,66,0,87,0,13,0,199,0,75,0,26,0,169,0,169,0,0,0,147,0,26,0,0,0,19,0,241,0,64,0,175,0,0,0,0,0,143,0,134,0,26,0,240,0,239,0,0,0,0,0,229,0,170,0,195,0,0,0,232,0,0,0,39,0,85,0,218,0,119,0,225,0,136,0,0,0,186,0,94,0,155,0,15,0,219,0,137,0,250,0,229,0,153,0,124,0,21,0,118,0,0,0,150,0,143,0,0,0,172,0,0,0,134,0,161,0,0,0,83,0,239,0,144,0,117,0,232,0,17,0,230,0,44,0,164,0,123,0,0,0,138,0,17,0,0,0,56,0,4,0,75,0,38,0,187,0,218,0,195,0,28,0,58,0,89,0,86,0,69,0,90,0,4,0,178,0,104,0,209,0,118,0,99,0,127,0,1,0,128,0,225,0,72,0,0,0,146,0,254,0,12,0,47,0,0,0,132,0,176,0,251,0,93,0,178,0,189,0,0,0,230,0,69,0,236,0,0,0,15,0,145,0,69,0,74,0,126,0,20,0,222,0,115,0,92,0,0,0,215,0,98,0,0,0,0,0,210,0,130,0,98,0);
signal scenario_full  : scenario_type := (169,31,192,31,192,30,192,29,23,31,139,31,46,31,42,31,103,31,220,31,221,31,44,31,44,30,91,31,91,30,31,31,31,30,168,31,220,31,251,31,126,31,103,31,74,31,74,30,63,31,63,30,246,31,61,31,61,30,162,31,162,30,162,29,101,31,97,31,195,31,121,31,80,31,154,31,154,30,154,29,154,28,191,31,41,31,27,31,27,30,25,31,171,31,237,31,84,31,214,31,252,31,110,31,240,31,195,31,20,31,251,31,189,31,189,30,64,31,129,31,129,30,60,31,57,31,78,31,78,30,255,31,255,30,118,31,210,31,113,31,113,30,6,31,30,31,172,31,208,31,211,31,15,31,76,31,76,30,76,29,58,31,86,31,22,31,22,30,122,31,223,31,45,31,238,31,134,31,114,31,9,31,225,31,5,31,110,31,151,31,11,31,11,30,11,29,86,31,165,31,217,31,96,31,41,31,41,30,204,31,97,31,145,31,81,31,242,31,196,31,152,31,89,31,103,31,136,31,221,31,251,31,76,31,136,31,163,31,154,31,234,31,85,31,196,31,196,30,3,31,182,31,156,31,146,31,222,31,16,31,193,31,215,31,134,31,191,31,235,31,235,30,222,31,80,31,44,31,145,31,94,31,226,31,178,31,229,31,28,31,79,31,240,31,149,31,181,31,181,30,173,31,173,30,14,31,64,31,184,31,241,31,156,31,156,30,252,31,114,31,175,31,144,31,141,31,141,30,48,31,93,31,75,31,3,31,179,31,6,31,253,31,34,31,136,31,148,31,148,30,121,31,1,31,90,31,20,31,235,31,134,31,16,31,16,30,181,31,181,30,120,31,120,30,120,29,120,28,94,31,108,31,108,30,144,31,183,31,243,31,202,31,163,31,37,31,82,31,120,31,155,31,126,31,207,31,207,30,65,31,53,31,243,31,243,30,123,31,241,31,95,31,86,31,51,31,154,31,154,31,59,31,93,31,47,31,234,31,234,30,149,31,162,31,162,30,162,29,117,31,130,31,170,31,159,31,63,31,46,31,54,31,2,31,2,30,205,31,83,31,61,31,209,31,52,31,23,31,241,31,58,31,125,31,125,30,125,29,43,31,107,31,252,31,94,31,137,31,137,31,134,31,164,31,161,31,199,31,199,30,199,29,242,31,27,31,206,31,206,30,27,31,54,31,57,31,220,31,44,31,44,30,130,31,239,31,176,31,139,31,139,30,111,31,78,31,203,31,203,30,171,31,148,31,11,31,161,31,119,31,119,30,85,31,95,31,218,31,218,30,151,31,133,31,182,31,116,31,38,31,38,30,165,31,73,31,8,31,146,31,3,31,3,30,251,31,104,31,104,30,107,31,66,31,216,31,40,31,107,31,217,31,184,31,189,31,234,31,234,30,204,31,106,31,179,31,13,31,13,30,253,31,12,31,36,31,52,31,226,31,82,31,247,31,44,31,44,30,161,31,248,31,76,31,176,31,12,31,12,30,12,29,128,31,162,31,131,31,2,31,97,31,97,30,97,29,23,31,138,31,131,31,131,30,131,29,27,31,51,31,134,31,122,31,207,31,34,31,34,30,252,31,169,31,169,30,221,31,208,31,95,31,64,31,139,31,218,31,127,31,51,31,51,30,241,31,241,30,156,31,84,31,84,30,21,31,21,30,51,31,128,31,112,31,65,31,75,31,96,31,96,30,96,29,241,31,71,31,136,31,75,31,75,30,26,31,51,31,105,31,105,30,75,31,19,31,17,31,229,31,100,31,151,31,88,31,99,31,190,31,190,30,190,29,75,31,15,31,215,31,167,31,72,31,130,31,130,30,171,31,52,31,158,31,158,30,179,31,252,31,37,31,128,31,204,31,230,31,230,30,230,29,230,28,225,31,70,31,64,31,79,31,165,31,165,30,165,29,165,28,229,31,187,31,155,31,246,31,68,31,40,31,75,31,150,31,36,31,167,31,12,31,67,31,67,30,76,31,105,31,105,31,19,31,84,31,81,31,30,31,62,31,62,30,198,31,18,31,57,31,20,31,15,31,8,31,115,31,242,31,242,30,216,31,216,30,249,31,249,30,161,31,76,31,234,31,53,31,53,30,233,31,139,31,30,31,89,31,76,31,229,31,239,31,62,31,62,30,9,31,155,31,66,31,66,30,220,31,220,30,226,31,122,31,34,31,34,30,201,31,12,31,112,31,229,31,242,31,182,31,194,31,137,31,226,31,127,31,127,30,63,31,176,31,255,31,11,31,34,31,188,31,188,30,9,31,187,31,21,31,21,30,8,31,55,31,255,31,76,31,14,31,54,31,1,31,81,31,182,31,182,30,97,31,10,31,48,31,189,31,123,31,6,31,110,31,18,31,98,31,22,31,168,31,54,31,39,31,41,31,92,31,46,31,49,31,177,31,145,31,47,31,51,31,15,31,25,31,39,31,66,31,66,30,53,31,65,31,106,31,110,31,174,31,169,31,169,30,81,31,104,31,58,31,70,31,71,31,71,30,206,31,199,31,199,30,253,31,98,31,47,31,78,31,78,30,125,31,146,31,66,31,167,31,202,31,148,31,225,31,106,31,85,31,153,31,153,30,55,31,222,31,178,31,96,31,41,31,24,31,122,31,85,31,75,31,163,31,214,31,3,31,3,30,3,29,3,28,41,31,120,31,255,31,82,31,223,31,160,31,49,31,49,30,219,31,18,31,190,31,252,31,35,31,35,30,35,29,214,31,233,31,110,31,176,31,1,31,114,31,95,31,175,31,36,31,49,31,198,31,198,30,198,29,224,31,101,31,101,30,101,29,99,31,100,31,31,31,31,30,31,29,224,31,171,31,43,31,155,31,74,31,74,30,52,31,246,31,246,30,162,31,223,31,225,31,225,30,2,31,221,31,218,31,183,31,183,30,184,31,184,30,162,31,84,31,226,31,226,30,120,31,54,31,68,31,68,30,206,31,164,31,192,31,192,30,192,29,250,31,250,30,8,31,97,31,79,31,235,31,207,31,61,31,171,31,125,31,132,31,145,31,145,30,177,31,177,30,177,29,177,28,130,31,130,30,12,31,218,31,218,30,222,31,222,30,131,31,206,31,206,30,206,29,79,31,98,31,14,31,210,31,210,30,41,31,41,30,232,31,177,31,45,31,45,30,156,31,5,31,123,31,45,31,127,31,60,31,115,31,39,31,17,31,152,31,216,31,248,31,26,31,242,31,77,31,77,30,16,31,42,31,42,30,42,29,63,31,123,31,123,30,30,31,30,30,56,31,39,31,46,31,18,31,18,30,7,31,222,31,207,31,161,31,111,31,173,31,5,31,152,31,212,31,151,31,151,30,70,31,48,31,48,30,35,31,213,31,196,31,149,31,154,31,35,31,61,31,168,31,168,30,154,31,115,31,53,31,53,30,96,31,18,31,18,30,18,29,38,31,92,31,73,31,71,31,160,31,242,31,225,31,232,31,132,31,132,30,132,29,54,31,229,31,229,30,221,31,221,30,144,31,144,30,35,31,190,31,166,31,166,30,103,31,103,30,142,31,10,31,43,31,156,31,196,31,133,31,34,31,13,31,121,31,186,31,186,30,238,31,160,31,160,30,39,31,39,30,39,29,39,28,78,31,39,31,147,31,227,31,86,31,82,31,82,30,13,31,182,31,249,31,110,31,40,31,108,31,45,31,198,31,209,31,123,31,123,30,171,31,34,31,99,31,178,31,194,31,170,31,170,30,170,29,170,28,16,31,132,31,122,31,184,31,67,31,62,31,165,31,87,31,46,31,46,30,34,31,62,31,62,30,143,31,160,31,83,31,83,30,83,29,101,31,161,31,37,31,182,31,237,31,95,31,243,31,243,30,93,31,8,31,65,31,46,31,37,31,37,30,254,31,147,31,147,30,224,31,54,31,54,30,105,31,243,31,217,31,83,31,66,31,87,31,13,31,199,31,75,31,26,31,169,31,169,31,169,30,147,31,26,31,26,30,19,31,241,31,64,31,175,31,175,30,175,29,143,31,134,31,26,31,240,31,239,31,239,30,239,29,229,31,170,31,195,31,195,30,232,31,232,30,39,31,85,31,218,31,119,31,225,31,136,31,136,30,186,31,94,31,155,31,15,31,219,31,137,31,250,31,229,31,153,31,124,31,21,31,118,31,118,30,150,31,143,31,143,30,172,31,172,30,134,31,161,31,161,30,83,31,239,31,144,31,117,31,232,31,17,31,230,31,44,31,164,31,123,31,123,30,138,31,17,31,17,30,56,31,4,31,75,31,38,31,187,31,218,31,195,31,28,31,58,31,89,31,86,31,69,31,90,31,4,31,178,31,104,31,209,31,118,31,99,31,127,31,1,31,128,31,225,31,72,31,72,30,146,31,254,31,12,31,47,31,47,30,132,31,176,31,251,31,93,31,178,31,189,31,189,30,230,31,69,31,236,31,236,30,15,31,145,31,69,31,74,31,126,31,20,31,222,31,115,31,92,31,92,30,215,31,98,31,98,30,98,29,210,31,130,31,98,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
