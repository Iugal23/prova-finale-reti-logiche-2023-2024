-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_782 is
end project_tb_782;

architecture project_tb_arch_782 of project_tb_782 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 276;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (153,0,156,0,7,0,223,0,153,0,64,0,212,0,3,0,211,0,188,0,0,0,103,0,0,0,102,0,107,0,212,0,179,0,151,0,0,0,0,0,236,0,0,0,34,0,44,0,0,0,0,0,136,0,0,0,52,0,211,0,235,0,164,0,0,0,27,0,164,0,135,0,237,0,0,0,72,0,0,0,7,0,249,0,75,0,62,0,28,0,240,0,127,0,87,0,238,0,164,0,225,0,21,0,151,0,173,0,205,0,0,0,148,0,0,0,17,0,153,0,112,0,246,0,87,0,38,0,110,0,40,0,0,0,218,0,0,0,44,0,110,0,124,0,241,0,162,0,0,0,251,0,0,0,77,0,0,0,225,0,29,0,251,0,26,0,199,0,158,0,58,0,183,0,130,0,124,0,0,0,132,0,0,0,183,0,160,0,9,0,0,0,183,0,6,0,102,0,183,0,187,0,112,0,21,0,0,0,0,0,210,0,19,0,0,0,66,0,0,0,0,0,112,0,72,0,109,0,145,0,231,0,0,0,40,0,202,0,14,0,4,0,133,0,143,0,12,0,86,0,242,0,69,0,201,0,13,0,80,0,0,0,0,0,69,0,255,0,183,0,10,0,0,0,122,0,162,0,241,0,227,0,155,0,163,0,0,0,0,0,120,0,161,0,94,0,87,0,48,0,134,0,0,0,6,0,0,0,0,0,0,0,232,0,48,0,187,0,77,0,96,0,38,0,83,0,38,0,229,0,190,0,0,0,96,0,90,0,0,0,0,0,140,0,13,0,254,0,0,0,221,0,114,0,159,0,156,0,0,0,148,0,111,0,79,0,181,0,191,0,243,0,104,0,224,0,149,0,203,0,243,0,241,0,28,0,128,0,71,0,126,0,191,0,98,0,207,0,232,0,0,0,1,0,0,0,44,0,160,0,169,0,191,0,78,0,174,0,132,0,59,0,0,0,159,0,73,0,0,0,195,0,255,0,17,0,33,0,178,0,106,0,100,0,0,0,0,0,251,0,226,0,0,0,181,0,29,0,208,0,0,0,200,0,0,0,195,0,19,0,0,0,0,0,113,0,17,0,131,0,64,0,94,0,0,0,193,0,249,0,96,0,112,0,0,0,27,0,251,0,141,0,78,0,21,0,186,0,0,0,217,0,223,0,217,0,159,0,111,0,0,0,0,0,83,0,0,0,122,0,51,0,0,0,45,0,123,0,133,0,0,0,197,0,31,0,137,0,79,0,178,0);
signal scenario_full  : scenario_type := (153,31,156,31,7,31,223,31,153,31,64,31,212,31,3,31,211,31,188,31,188,30,103,31,103,30,102,31,107,31,212,31,179,31,151,31,151,30,151,29,236,31,236,30,34,31,44,31,44,30,44,29,136,31,136,30,52,31,211,31,235,31,164,31,164,30,27,31,164,31,135,31,237,31,237,30,72,31,72,30,7,31,249,31,75,31,62,31,28,31,240,31,127,31,87,31,238,31,164,31,225,31,21,31,151,31,173,31,205,31,205,30,148,31,148,30,17,31,153,31,112,31,246,31,87,31,38,31,110,31,40,31,40,30,218,31,218,30,44,31,110,31,124,31,241,31,162,31,162,30,251,31,251,30,77,31,77,30,225,31,29,31,251,31,26,31,199,31,158,31,58,31,183,31,130,31,124,31,124,30,132,31,132,30,183,31,160,31,9,31,9,30,183,31,6,31,102,31,183,31,187,31,112,31,21,31,21,30,21,29,210,31,19,31,19,30,66,31,66,30,66,29,112,31,72,31,109,31,145,31,231,31,231,30,40,31,202,31,14,31,4,31,133,31,143,31,12,31,86,31,242,31,69,31,201,31,13,31,80,31,80,30,80,29,69,31,255,31,183,31,10,31,10,30,122,31,162,31,241,31,227,31,155,31,163,31,163,30,163,29,120,31,161,31,94,31,87,31,48,31,134,31,134,30,6,31,6,30,6,29,6,28,232,31,48,31,187,31,77,31,96,31,38,31,83,31,38,31,229,31,190,31,190,30,96,31,90,31,90,30,90,29,140,31,13,31,254,31,254,30,221,31,114,31,159,31,156,31,156,30,148,31,111,31,79,31,181,31,191,31,243,31,104,31,224,31,149,31,203,31,243,31,241,31,28,31,128,31,71,31,126,31,191,31,98,31,207,31,232,31,232,30,1,31,1,30,44,31,160,31,169,31,191,31,78,31,174,31,132,31,59,31,59,30,159,31,73,31,73,30,195,31,255,31,17,31,33,31,178,31,106,31,100,31,100,30,100,29,251,31,226,31,226,30,181,31,29,31,208,31,208,30,200,31,200,30,195,31,19,31,19,30,19,29,113,31,17,31,131,31,64,31,94,31,94,30,193,31,249,31,96,31,112,31,112,30,27,31,251,31,141,31,78,31,21,31,186,31,186,30,217,31,223,31,217,31,159,31,111,31,111,30,111,29,83,31,83,30,122,31,51,31,51,30,45,31,123,31,133,31,133,30,197,31,31,31,137,31,79,31,178,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
