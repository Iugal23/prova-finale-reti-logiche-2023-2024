-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 417;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,28,0,117,0,168,0,0,0,40,0,86,0,231,0,39,0,254,0,170,0,27,0,0,0,24,0,0,0,30,0,68,0,62,0,180,0,158,0,213,0,240,0,147,0,82,0,229,0,42,0,0,0,0,0,84,0,144,0,187,0,0,0,222,0,195,0,154,0,204,0,0,0,73,0,172,0,0,0,20,0,26,0,159,0,139,0,0,0,97,0,0,0,69,0,137,0,71,0,210,0,217,0,97,0,101,0,66,0,228,0,56,0,101,0,48,0,0,0,0,0,229,0,254,0,121,0,180,0,0,0,52,0,222,0,169,0,214,0,95,0,175,0,147,0,65,0,207,0,108,0,207,0,226,0,0,0,0,0,0,0,60,0,0,0,12,0,119,0,0,0,191,0,197,0,200,0,122,0,0,0,0,0,172,0,130,0,88,0,149,0,12,0,59,0,85,0,216,0,121,0,29,0,0,0,156,0,254,0,185,0,160,0,78,0,158,0,0,0,0,0,239,0,113,0,171,0,22,0,75,0,0,0,193,0,0,0,143,0,90,0,62,0,8,0,105,0,206,0,109,0,113,0,74,0,86,0,0,0,0,0,247,0,25,0,0,0,212,0,172,0,218,0,173,0,190,0,204,0,0,0,224,0,160,0,166,0,7,0,0,0,144,0,204,0,101,0,169,0,70,0,211,0,123,0,191,0,251,0,62,0,90,0,57,0,103,0,13,0,104,0,59,0,0,0,51,0,11,0,0,0,251,0,137,0,99,0,82,0,217,0,70,0,166,0,227,0,145,0,137,0,0,0,25,0,0,0,5,0,244,0,137,0,246,0,255,0,168,0,247,0,130,0,0,0,4,0,220,0,28,0,248,0,199,0,95,0,0,0,50,0,36,0,0,0,157,0,0,0,103,0,0,0,22,0,149,0,0,0,0,0,179,0,126,0,88,0,16,0,0,0,247,0,202,0,168,0,236,0,195,0,0,0,162,0,11,0,0,0,0,0,220,0,70,0,186,0,70,0,156,0,115,0,17,0,0,0,123,0,213,0,205,0,20,0,0,0,58,0,0,0,0,0,163,0,76,0,254,0,221,0,22,0,247,0,0,0,132,0,22,0,22,0,62,0,66,0,8,0,201,0,211,0,254,0,198,0,0,0,0,0,108,0,11,0,167,0,248,0,146,0,228,0,0,0,115,0,0,0,69,0,0,0,0,0,0,0,79,0,16,0,0,0,239,0,30,0,21,0,88,0,154,0,26,0,84,0,4,0,106,0,208,0,0,0,20,0,239,0,48,0,234,0,162,0,115,0,0,0,1,0,0,0,122,0,1,0,29,0,154,0,69,0,36,0,0,0,0,0,244,0,68,0,0,0,85,0,104,0,85,0,0,0,122,0,0,0,0,0,0,0,197,0,129,0,18,0,0,0,169,0,181,0,97,0,85,0,50,0,199,0,194,0,0,0,102,0,31,0,195,0,41,0,172,0,0,0,29,0,69,0,0,0,0,0,28,0,0,0,245,0,96,0,239,0,244,0,0,0,229,0,83,0,230,0,63,0,49,0,177,0,49,0,0,0,18,0,123,0,210,0,233,0,37,0,117,0,238,0,51,0,20,0,87,0,50,0,23,0,0,0,17,0,109,0,57,0,0,0,44,0,90,0,0,0,0,0,116,0,208,0,167,0,0,0,0,0,0,0,0,0,77,0,179,0,109,0,131,0,0,0,167,0,130,0,21,0,0,0,38,0,147,0,164,0,16,0,198,0,191,0,167,0,126,0,43,0,0,0,132,0,0,0,154,0,60,0,180,0,111,0,151,0,252,0,212,0,127,0,211,0,0,0,189,0,161,0,60,0,57,0,160,0,0,0,111,0,213,0,14,0,0,0);
signal scenario_full  : scenario_type := (149,31,28,31,117,31,168,31,168,30,40,31,86,31,231,31,39,31,254,31,170,31,27,31,27,30,24,31,24,30,30,31,68,31,62,31,180,31,158,31,213,31,240,31,147,31,82,31,229,31,42,31,42,30,42,29,84,31,144,31,187,31,187,30,222,31,195,31,154,31,204,31,204,30,73,31,172,31,172,30,20,31,26,31,159,31,139,31,139,30,97,31,97,30,69,31,137,31,71,31,210,31,217,31,97,31,101,31,66,31,228,31,56,31,101,31,48,31,48,30,48,29,229,31,254,31,121,31,180,31,180,30,52,31,222,31,169,31,214,31,95,31,175,31,147,31,65,31,207,31,108,31,207,31,226,31,226,30,226,29,226,28,60,31,60,30,12,31,119,31,119,30,191,31,197,31,200,31,122,31,122,30,122,29,172,31,130,31,88,31,149,31,12,31,59,31,85,31,216,31,121,31,29,31,29,30,156,31,254,31,185,31,160,31,78,31,158,31,158,30,158,29,239,31,113,31,171,31,22,31,75,31,75,30,193,31,193,30,143,31,90,31,62,31,8,31,105,31,206,31,109,31,113,31,74,31,86,31,86,30,86,29,247,31,25,31,25,30,212,31,172,31,218,31,173,31,190,31,204,31,204,30,224,31,160,31,166,31,7,31,7,30,144,31,204,31,101,31,169,31,70,31,211,31,123,31,191,31,251,31,62,31,90,31,57,31,103,31,13,31,104,31,59,31,59,30,51,31,11,31,11,30,251,31,137,31,99,31,82,31,217,31,70,31,166,31,227,31,145,31,137,31,137,30,25,31,25,30,5,31,244,31,137,31,246,31,255,31,168,31,247,31,130,31,130,30,4,31,220,31,28,31,248,31,199,31,95,31,95,30,50,31,36,31,36,30,157,31,157,30,103,31,103,30,22,31,149,31,149,30,149,29,179,31,126,31,88,31,16,31,16,30,247,31,202,31,168,31,236,31,195,31,195,30,162,31,11,31,11,30,11,29,220,31,70,31,186,31,70,31,156,31,115,31,17,31,17,30,123,31,213,31,205,31,20,31,20,30,58,31,58,30,58,29,163,31,76,31,254,31,221,31,22,31,247,31,247,30,132,31,22,31,22,31,62,31,66,31,8,31,201,31,211,31,254,31,198,31,198,30,198,29,108,31,11,31,167,31,248,31,146,31,228,31,228,30,115,31,115,30,69,31,69,30,69,29,69,28,79,31,16,31,16,30,239,31,30,31,21,31,88,31,154,31,26,31,84,31,4,31,106,31,208,31,208,30,20,31,239,31,48,31,234,31,162,31,115,31,115,30,1,31,1,30,122,31,1,31,29,31,154,31,69,31,36,31,36,30,36,29,244,31,68,31,68,30,85,31,104,31,85,31,85,30,122,31,122,30,122,29,122,28,197,31,129,31,18,31,18,30,169,31,181,31,97,31,85,31,50,31,199,31,194,31,194,30,102,31,31,31,195,31,41,31,172,31,172,30,29,31,69,31,69,30,69,29,28,31,28,30,245,31,96,31,239,31,244,31,244,30,229,31,83,31,230,31,63,31,49,31,177,31,49,31,49,30,18,31,123,31,210,31,233,31,37,31,117,31,238,31,51,31,20,31,87,31,50,31,23,31,23,30,17,31,109,31,57,31,57,30,44,31,90,31,90,30,90,29,116,31,208,31,167,31,167,30,167,29,167,28,167,27,77,31,179,31,109,31,131,31,131,30,167,31,130,31,21,31,21,30,38,31,147,31,164,31,16,31,198,31,191,31,167,31,126,31,43,31,43,30,132,31,132,30,154,31,60,31,180,31,111,31,151,31,252,31,212,31,127,31,211,31,211,30,189,31,161,31,60,31,57,31,160,31,160,30,111,31,213,31,14,31,14,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
