-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 933;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,234,0,0,0,41,0,186,0,238,0,168,0,248,0,217,0,40,0,226,0,169,0,17,0,17,0,8,0,0,0,234,0,46,0,237,0,0,0,60,0,126,0,161,0,0,0,35,0,176,0,3,0,0,0,0,0,38,0,255,0,70,0,242,0,249,0,141,0,49,0,161,0,86,0,21,0,62,0,246,0,205,0,213,0,0,0,129,0,187,0,226,0,236,0,92,0,127,0,0,0,17,0,231,0,105,0,117,0,213,0,208,0,0,0,127,0,79,0,160,0,212,0,68,0,149,0,0,0,147,0,233,0,243,0,0,0,34,0,142,0,116,0,21,0,12,0,23,0,233,0,241,0,203,0,24,0,108,0,78,0,0,0,146,0,26,0,66,0,98,0,221,0,106,0,0,0,0,0,0,0,0,0,0,0,122,0,213,0,234,0,163,0,164,0,248,0,173,0,61,0,163,0,56,0,177,0,4,0,0,0,35,0,0,0,204,0,71,0,168,0,0,0,98,0,145,0,0,0,50,0,206,0,231,0,5,0,58,0,163,0,102,0,170,0,133,0,0,0,30,0,253,0,238,0,220,0,198,0,184,0,153,0,86,0,212,0,0,0,219,0,0,0,52,0,223,0,0,0,236,0,0,0,28,0,187,0,0,0,247,0,88,0,89,0,215,0,205,0,240,0,62,0,23,0,67,0,0,0,125,0,105,0,145,0,239,0,52,0,218,0,0,0,12,0,47,0,0,0,165,0,23,0,212,0,72,0,99,0,148,0,96,0,0,0,90,0,0,0,65,0,136,0,204,0,10,0,136,0,171,0,62,0,0,0,17,0,107,0,240,0,231,0,12,0,157,0,170,0,251,0,197,0,0,0,0,0,0,0,252,0,218,0,117,0,163,0,1,0,127,0,10,0,7,0,10,0,70,0,0,0,12,0,10,0,109,0,37,0,214,0,90,0,124,0,191,0,0,0,134,0,206,0,239,0,209,0,0,0,0,0,229,0,201,0,113,0,0,0,32,0,0,0,0,0,99,0,0,0,221,0,184,0,1,0,96,0,128,0,3,0,132,0,0,0,0,0,217,0,246,0,169,0,232,0,255,0,32,0,157,0,196,0,207,0,72,0,0,0,94,0,252,0,0,0,163,0,10,0,18,0,155,0,0,0,83,0,145,0,2,0,80,0,62,0,182,0,135,0,133,0,3,0,63,0,218,0,0,0,159,0,112,0,109,0,64,0,147,0,41,0,201,0,183,0,0,0,198,0,4,0,4,0,180,0,5,0,215,0,56,0,12,0,211,0,120,0,129,0,45,0,94,0,137,0,0,0,187,0,76,0,98,0,27,0,194,0,165,0,136,0,107,0,0,0,201,0,204,0,209,0,52,0,6,0,133,0,141,0,0,0,197,0,154,0,0,0,86,0,71,0,195,0,35,0,158,0,185,0,22,0,191,0,0,0,2,0,183,0,0,0,62,0,93,0,83,0,0,0,167,0,0,0,224,0,96,0,212,0,144,0,123,0,124,0,67,0,70,0,171,0,164,0,102,0,81,0,165,0,111,0,0,0,185,0,211,0,77,0,67,0,218,0,44,0,27,0,0,0,174,0,82,0,0,0,0,0,203,0,208,0,13,0,91,0,101,0,59,0,58,0,235,0,144,0,50,0,98,0,18,0,177,0,92,0,0,0,150,0,196,0,21,0,98,0,83,0,173,0,0,0,21,0,58,0,190,0,140,0,213,0,0,0,0,0,22,0,31,0,173,0,95,0,0,0,133,0,109,0,75,0,249,0,240,0,91,0,244,0,0,0,235,0,42,0,218,0,0,0,156,0,111,0,250,0,235,0,0,0,141,0,207,0,135,0,31,0,53,0,3,0,47,0,92,0,0,0,240,0,45,0,0,0,71,0,0,0,213,0,0,0,73,0,53,0,204,0,168,0,207,0,132,0,4,0,131,0,1,0,179,0,230,0,196,0,79,0,109,0,17,0,23,0,31,0,54,0,226,0,0,0,0,0,184,0,95,0,177,0,6,0,196,0,187,0,183,0,0,0,158,0,0,0,134,0,232,0,143,0,179,0,233,0,244,0,26,0,85,0,198,0,0,0,0,0,252,0,247,0,43,0,194,0,1,0,21,0,153,0,127,0,182,0,39,0,133,0,15,0,0,0,92,0,236,0,170,0,241,0,153,0,161,0,187,0,0,0,0,0,179,0,5,0,94,0,0,0,209,0,65,0,79,0,161,0,237,0,207,0,27,0,48,0,0,0,0,0,0,0,92,0,244,0,195,0,42,0,125,0,160,0,105,0,148,0,0,0,163,0,45,0,114,0,0,0,95,0,0,0,53,0,79,0,0,0,144,0,0,0,245,0,0,0,17,0,0,0,184,0,19,0,172,0,9,0,0,0,0,0,213,0,173,0,0,0,58,0,19,0,183,0,0,0,86,0,199,0,52,0,83,0,0,0,247,0,222,0,223,0,194,0,190,0,76,0,143,0,209,0,183,0,24,0,175,0,45,0,139,0,0,0,169,0,35,0,0,0,125,0,220,0,66,0,40,0,147,0,0,0,127,0,0,0,0,0,119,0,0,0,42,0,0,0,57,0,196,0,136,0,86,0,171,0,3,0,0,0,110,0,94,0,185,0,6,0,91,0,206,0,83,0,0,0,0,0,185,0,192,0,68,0,31,0,216,0,80,0,204,0,20,0,70,0,159,0,68,0,0,0,223,0,23,0,229,0,163,0,232,0,187,0,0,0,205,0,119,0,0,0,164,0,13,0,0,0,76,0,168,0,105,0,211,0,135,0,68,0,158,0,83,0,96,0,0,0,137,0,227,0,19,0,140,0,85,0,42,0,134,0,0,0,229,0,107,0,27,0,41,0,229,0,69,0,0,0,31,0,90,0,0,0,134,0,152,0,1,0,236,0,106,0,24,0,0,0,54,0,0,0,220,0,41,0,95,0,154,0,122,0,44,0,132,0,56,0,97,0,0,0,169,0,92,0,185,0,2,0,62,0,120,0,70,0,77,0,0,0,244,0,0,0,66,0,0,0,0,0,90,0,0,0,227,0,43,0,235,0,167,0,22,0,51,0,106,0,15,0,102,0,0,0,0,0,66,0,39,0,0,0,0,0,0,0,0,0,81,0,146,0,228,0,0,0,68,0,65,0,41,0,211,0,132,0,0,0,60,0,161,0,4,0,176,0,116,0,233,0,0,0,2,0,87,0,35,0,201,0,68,0,0,0,153,0,215,0,216,0,175,0,3,0,173,0,0,0,0,0,129,0,11,0,168,0,0,0,124,0,200,0,216,0,0,0,175,0,120,0,129,0,68,0,0,0,17,0,202,0,48,0,204,0,26,0,82,0,38,0,69,0,228,0,216,0,70,0,98,0,139,0,177,0,0,0,226,0,95,0,230,0,15,0,218,0,156,0,144,0,0,0,74,0,175,0,0,0,43,0,102,0,5,0,11,0,126,0,180,0,48,0,0,0,200,0,238,0,109,0,145,0,211,0,211,0,0,0,144,0,58,0,180,0,0,0,46,0,175,0,188,0,76,0,0,0,101,0,0,0,230,0,147,0,90,0,184,0,0,0,0,0,172,0,59,0,231,0,57,0,0,0,43,0,100,0,30,0,200,0,211,0,0,0,231,0,255,0,82,0,147,0,146,0,166,0,0,0,57,0,16,0,250,0,29,0,156,0,0,0,36,0,0,0,0,0,130,0,0,0,111,0,17,0,0,0,51,0,122,0,54,0,134,0,24,0,26,0,125,0,0,0,83,0,38,0,246,0,170,0,128,0,103,0,183,0,45,0,210,0,34,0,224,0,9,0,139,0,92,0,209,0,215,0,164,0,187,0,244,0,0,0,110,0,0,0,37,0,114,0,82,0,0,0,30,0,81,0,67,0,156,0,237,0,139,0,179,0,119,0,88,0,0,0,64,0,107,0,78,0,101,0,130,0,0,0,0,0,212,0,5,0,104,0,0,0,111,0,192,0,12,0,0,0,0,0,132,0,201,0,36,0,30,0,0,0,97,0,59,0,0,0,119,0,254,0,171,0,147,0,0,0,121,0,99,0,5,0,185,0,253,0,214,0,140,0,0,0,235,0,0,0,228,0,140,0,176,0,9,0,193,0,244,0,82,0,17,0,59,0,9,0,219,0,184,0,39,0,163,0,116,0,0,0,182,0,71,0);
signal scenario_full  : scenario_type := (181,31,234,31,234,30,41,31,186,31,238,31,168,31,248,31,217,31,40,31,226,31,169,31,17,31,17,31,8,31,8,30,234,31,46,31,237,31,237,30,60,31,126,31,161,31,161,30,35,31,176,31,3,31,3,30,3,29,38,31,255,31,70,31,242,31,249,31,141,31,49,31,161,31,86,31,21,31,62,31,246,31,205,31,213,31,213,30,129,31,187,31,226,31,236,31,92,31,127,31,127,30,17,31,231,31,105,31,117,31,213,31,208,31,208,30,127,31,79,31,160,31,212,31,68,31,149,31,149,30,147,31,233,31,243,31,243,30,34,31,142,31,116,31,21,31,12,31,23,31,233,31,241,31,203,31,24,31,108,31,78,31,78,30,146,31,26,31,66,31,98,31,221,31,106,31,106,30,106,29,106,28,106,27,106,26,122,31,213,31,234,31,163,31,164,31,248,31,173,31,61,31,163,31,56,31,177,31,4,31,4,30,35,31,35,30,204,31,71,31,168,31,168,30,98,31,145,31,145,30,50,31,206,31,231,31,5,31,58,31,163,31,102,31,170,31,133,31,133,30,30,31,253,31,238,31,220,31,198,31,184,31,153,31,86,31,212,31,212,30,219,31,219,30,52,31,223,31,223,30,236,31,236,30,28,31,187,31,187,30,247,31,88,31,89,31,215,31,205,31,240,31,62,31,23,31,67,31,67,30,125,31,105,31,145,31,239,31,52,31,218,31,218,30,12,31,47,31,47,30,165,31,23,31,212,31,72,31,99,31,148,31,96,31,96,30,90,31,90,30,65,31,136,31,204,31,10,31,136,31,171,31,62,31,62,30,17,31,107,31,240,31,231,31,12,31,157,31,170,31,251,31,197,31,197,30,197,29,197,28,252,31,218,31,117,31,163,31,1,31,127,31,10,31,7,31,10,31,70,31,70,30,12,31,10,31,109,31,37,31,214,31,90,31,124,31,191,31,191,30,134,31,206,31,239,31,209,31,209,30,209,29,229,31,201,31,113,31,113,30,32,31,32,30,32,29,99,31,99,30,221,31,184,31,1,31,96,31,128,31,3,31,132,31,132,30,132,29,217,31,246,31,169,31,232,31,255,31,32,31,157,31,196,31,207,31,72,31,72,30,94,31,252,31,252,30,163,31,10,31,18,31,155,31,155,30,83,31,145,31,2,31,80,31,62,31,182,31,135,31,133,31,3,31,63,31,218,31,218,30,159,31,112,31,109,31,64,31,147,31,41,31,201,31,183,31,183,30,198,31,4,31,4,31,180,31,5,31,215,31,56,31,12,31,211,31,120,31,129,31,45,31,94,31,137,31,137,30,187,31,76,31,98,31,27,31,194,31,165,31,136,31,107,31,107,30,201,31,204,31,209,31,52,31,6,31,133,31,141,31,141,30,197,31,154,31,154,30,86,31,71,31,195,31,35,31,158,31,185,31,22,31,191,31,191,30,2,31,183,31,183,30,62,31,93,31,83,31,83,30,167,31,167,30,224,31,96,31,212,31,144,31,123,31,124,31,67,31,70,31,171,31,164,31,102,31,81,31,165,31,111,31,111,30,185,31,211,31,77,31,67,31,218,31,44,31,27,31,27,30,174,31,82,31,82,30,82,29,203,31,208,31,13,31,91,31,101,31,59,31,58,31,235,31,144,31,50,31,98,31,18,31,177,31,92,31,92,30,150,31,196,31,21,31,98,31,83,31,173,31,173,30,21,31,58,31,190,31,140,31,213,31,213,30,213,29,22,31,31,31,173,31,95,31,95,30,133,31,109,31,75,31,249,31,240,31,91,31,244,31,244,30,235,31,42,31,218,31,218,30,156,31,111,31,250,31,235,31,235,30,141,31,207,31,135,31,31,31,53,31,3,31,47,31,92,31,92,30,240,31,45,31,45,30,71,31,71,30,213,31,213,30,73,31,53,31,204,31,168,31,207,31,132,31,4,31,131,31,1,31,179,31,230,31,196,31,79,31,109,31,17,31,23,31,31,31,54,31,226,31,226,30,226,29,184,31,95,31,177,31,6,31,196,31,187,31,183,31,183,30,158,31,158,30,134,31,232,31,143,31,179,31,233,31,244,31,26,31,85,31,198,31,198,30,198,29,252,31,247,31,43,31,194,31,1,31,21,31,153,31,127,31,182,31,39,31,133,31,15,31,15,30,92,31,236,31,170,31,241,31,153,31,161,31,187,31,187,30,187,29,179,31,5,31,94,31,94,30,209,31,65,31,79,31,161,31,237,31,207,31,27,31,48,31,48,30,48,29,48,28,92,31,244,31,195,31,42,31,125,31,160,31,105,31,148,31,148,30,163,31,45,31,114,31,114,30,95,31,95,30,53,31,79,31,79,30,144,31,144,30,245,31,245,30,17,31,17,30,184,31,19,31,172,31,9,31,9,30,9,29,213,31,173,31,173,30,58,31,19,31,183,31,183,30,86,31,199,31,52,31,83,31,83,30,247,31,222,31,223,31,194,31,190,31,76,31,143,31,209,31,183,31,24,31,175,31,45,31,139,31,139,30,169,31,35,31,35,30,125,31,220,31,66,31,40,31,147,31,147,30,127,31,127,30,127,29,119,31,119,30,42,31,42,30,57,31,196,31,136,31,86,31,171,31,3,31,3,30,110,31,94,31,185,31,6,31,91,31,206,31,83,31,83,30,83,29,185,31,192,31,68,31,31,31,216,31,80,31,204,31,20,31,70,31,159,31,68,31,68,30,223,31,23,31,229,31,163,31,232,31,187,31,187,30,205,31,119,31,119,30,164,31,13,31,13,30,76,31,168,31,105,31,211,31,135,31,68,31,158,31,83,31,96,31,96,30,137,31,227,31,19,31,140,31,85,31,42,31,134,31,134,30,229,31,107,31,27,31,41,31,229,31,69,31,69,30,31,31,90,31,90,30,134,31,152,31,1,31,236,31,106,31,24,31,24,30,54,31,54,30,220,31,41,31,95,31,154,31,122,31,44,31,132,31,56,31,97,31,97,30,169,31,92,31,185,31,2,31,62,31,120,31,70,31,77,31,77,30,244,31,244,30,66,31,66,30,66,29,90,31,90,30,227,31,43,31,235,31,167,31,22,31,51,31,106,31,15,31,102,31,102,30,102,29,66,31,39,31,39,30,39,29,39,28,39,27,81,31,146,31,228,31,228,30,68,31,65,31,41,31,211,31,132,31,132,30,60,31,161,31,4,31,176,31,116,31,233,31,233,30,2,31,87,31,35,31,201,31,68,31,68,30,153,31,215,31,216,31,175,31,3,31,173,31,173,30,173,29,129,31,11,31,168,31,168,30,124,31,200,31,216,31,216,30,175,31,120,31,129,31,68,31,68,30,17,31,202,31,48,31,204,31,26,31,82,31,38,31,69,31,228,31,216,31,70,31,98,31,139,31,177,31,177,30,226,31,95,31,230,31,15,31,218,31,156,31,144,31,144,30,74,31,175,31,175,30,43,31,102,31,5,31,11,31,126,31,180,31,48,31,48,30,200,31,238,31,109,31,145,31,211,31,211,31,211,30,144,31,58,31,180,31,180,30,46,31,175,31,188,31,76,31,76,30,101,31,101,30,230,31,147,31,90,31,184,31,184,30,184,29,172,31,59,31,231,31,57,31,57,30,43,31,100,31,30,31,200,31,211,31,211,30,231,31,255,31,82,31,147,31,146,31,166,31,166,30,57,31,16,31,250,31,29,31,156,31,156,30,36,31,36,30,36,29,130,31,130,30,111,31,17,31,17,30,51,31,122,31,54,31,134,31,24,31,26,31,125,31,125,30,83,31,38,31,246,31,170,31,128,31,103,31,183,31,45,31,210,31,34,31,224,31,9,31,139,31,92,31,209,31,215,31,164,31,187,31,244,31,244,30,110,31,110,30,37,31,114,31,82,31,82,30,30,31,81,31,67,31,156,31,237,31,139,31,179,31,119,31,88,31,88,30,64,31,107,31,78,31,101,31,130,31,130,30,130,29,212,31,5,31,104,31,104,30,111,31,192,31,12,31,12,30,12,29,132,31,201,31,36,31,30,31,30,30,97,31,59,31,59,30,119,31,254,31,171,31,147,31,147,30,121,31,99,31,5,31,185,31,253,31,214,31,140,31,140,30,235,31,235,30,228,31,140,31,176,31,9,31,193,31,244,31,82,31,17,31,59,31,9,31,219,31,184,31,39,31,163,31,116,31,116,30,182,31,71,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
