-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_971 is
end project_tb_971;

architecture project_tb_arch_971 of project_tb_971 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 182;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,172,0,245,0,242,0,122,0,192,0,99,0,0,0,156,0,234,0,5,0,0,0,0,0,0,0,104,0,46,0,0,0,208,0,0,0,227,0,220,0,190,0,230,0,0,0,190,0,80,0,0,0,26,0,216,0,0,0,144,0,24,0,26,0,132,0,171,0,177,0,208,0,98,0,240,0,124,0,96,0,142,0,71,0,164,0,199,0,0,0,14,0,68,0,0,0,3,0,3,0,0,0,204,0,0,0,146,0,105,0,0,0,82,0,49,0,0,0,140,0,255,0,70,0,181,0,249,0,0,0,0,0,137,0,89,0,11,0,207,0,0,0,147,0,89,0,184,0,0,0,248,0,207,0,135,0,179,0,51,0,58,0,196,0,126,0,190,0,65,0,246,0,229,0,166,0,28,0,55,0,206,0,209,0,213,0,151,0,0,0,135,0,176,0,21,0,59,0,61,0,175,0,95,0,191,0,0,0,154,0,0,0,140,0,241,0,0,0,241,0,242,0,66,0,150,0,44,0,205,0,0,0,132,0,242,0,54,0,121,0,17,0,119,0,247,0,63,0,243,0,52,0,235,0,0,0,0,0,218,0,240,0,145,0,16,0,0,0,233,0,189,0,17,0,41,0,213,0,213,0,112,0,75,0,0,0,98,0,103,0,106,0,173,0,108,0,143,0,205,0,98,0,93,0,132,0,0,0,54,0,144,0,102,0,16,0,97,0,4,0,106,0,146,0,100,0,0,0,72,0,72,0,186,0,181,0,202,0,0,0,75,0,40,0,225,0,207,0,177,0,30,0,0,0,116,0,183,0,76,0,234,0);
signal scenario_full  : scenario_type := (134,31,172,31,245,31,242,31,122,31,192,31,99,31,99,30,156,31,234,31,5,31,5,30,5,29,5,28,104,31,46,31,46,30,208,31,208,30,227,31,220,31,190,31,230,31,230,30,190,31,80,31,80,30,26,31,216,31,216,30,144,31,24,31,26,31,132,31,171,31,177,31,208,31,98,31,240,31,124,31,96,31,142,31,71,31,164,31,199,31,199,30,14,31,68,31,68,30,3,31,3,31,3,30,204,31,204,30,146,31,105,31,105,30,82,31,49,31,49,30,140,31,255,31,70,31,181,31,249,31,249,30,249,29,137,31,89,31,11,31,207,31,207,30,147,31,89,31,184,31,184,30,248,31,207,31,135,31,179,31,51,31,58,31,196,31,126,31,190,31,65,31,246,31,229,31,166,31,28,31,55,31,206,31,209,31,213,31,151,31,151,30,135,31,176,31,21,31,59,31,61,31,175,31,95,31,191,31,191,30,154,31,154,30,140,31,241,31,241,30,241,31,242,31,66,31,150,31,44,31,205,31,205,30,132,31,242,31,54,31,121,31,17,31,119,31,247,31,63,31,243,31,52,31,235,31,235,30,235,29,218,31,240,31,145,31,16,31,16,30,233,31,189,31,17,31,41,31,213,31,213,31,112,31,75,31,75,30,98,31,103,31,106,31,173,31,108,31,143,31,205,31,98,31,93,31,132,31,132,30,54,31,144,31,102,31,16,31,97,31,4,31,106,31,146,31,100,31,100,30,72,31,72,31,186,31,181,31,202,31,202,30,75,31,40,31,225,31,207,31,177,31,30,31,30,30,116,31,183,31,76,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
