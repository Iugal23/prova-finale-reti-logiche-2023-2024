-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 379;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,111,0,0,0,142,0,102,0,140,0,196,0,138,0,87,0,0,0,231,0,208,0,172,0,122,0,0,0,0,0,244,0,0,0,110,0,0,0,18,0,245,0,156,0,166,0,114,0,145,0,0,0,170,0,134,0,28,0,0,0,0,0,201,0,239,0,135,0,38,0,62,0,125,0,16,0,182,0,176,0,22,0,0,0,239,0,255,0,0,0,0,0,4,0,0,0,243,0,247,0,80,0,245,0,86,0,197,0,206,0,20,0,51,0,151,0,223,0,0,0,0,0,80,0,104,0,229,0,61,0,0,0,94,0,0,0,190,0,249,0,23,0,162,0,187,0,120,0,0,0,247,0,0,0,159,0,109,0,80,0,166,0,54,0,152,0,0,0,59,0,181,0,146,0,190,0,99,0,69,0,48,0,160,0,13,0,72,0,58,0,0,0,41,0,77,0,243,0,0,0,244,0,131,0,61,0,137,0,62,0,163,0,49,0,8,0,69,0,4,0,86,0,173,0,250,0,45,0,0,0,195,0,143,0,0,0,148,0,235,0,38,0,90,0,0,0,0,0,249,0,251,0,194,0,0,0,80,0,9,0,119,0,204,0,0,0,54,0,206,0,205,0,70,0,29,0,10,0,126,0,144,0,41,0,161,0,0,0,103,0,30,0,47,0,1,0,243,0,0,0,0,0,227,0,20,0,67,0,143,0,38,0,14,0,169,0,2,0,101,0,47,0,0,0,7,0,18,0,0,0,50,0,131,0,101,0,59,0,213,0,0,0,195,0,91,0,237,0,0,0,88,0,0,0,0,0,108,0,52,0,98,0,0,0,171,0,0,0,0,0,42,0,0,0,50,0,230,0,131,0,238,0,133,0,0,0,0,0,145,0,153,0,92,0,0,0,147,0,166,0,0,0,0,0,226,0,0,0,62,0,89,0,82,0,142,0,0,0,201,0,0,0,12,0,66,0,5,0,3,0,0,0,6,0,0,0,186,0,0,0,101,0,0,0,0,0,0,0,254,0,154,0,241,0,232,0,213,0,108,0,147,0,47,0,163,0,68,0,104,0,198,0,90,0,0,0,30,0,0,0,83,0,17,0,103,0,55,0,34,0,9,0,63,0,102,0,93,0,224,0,148,0,232,0,0,0,100,0,69,0,0,0,39,0,0,0,194,0,0,0,63,0,203,0,39,0,44,0,200,0,208,0,201,0,166,0,231,0,21,0,48,0,0,0,17,0,64,0,129,0,255,0,211,0,68,0,224,0,173,0,162,0,220,0,118,0,29,0,148,0,43,0,163,0,130,0,221,0,139,0,0,0,0,0,237,0,106,0,0,0,0,0,71,0,147,0,231,0,74,0,38,0,181,0,0,0,208,0,0,0,243,0,0,0,190,0,156,0,254,0,0,0,213,0,30,0,0,0,143,0,24,0,165,0,12,0,100,0,198,0,0,0,0,0,0,0,148,0,94,0,0,0,190,0,76,0,35,0,0,0,235,0,226,0,217,0,107,0,234,0,159,0,191,0,195,0,87,0,126,0,226,0,231,0,43,0,35,0,163,0,173,0,162,0,122,0,86,0,0,0,13,0,137,0,146,0,174,0,214,0,75,0,106,0,0,0,205,0,144,0,172,0,0,0,158,0,0,0,7,0,0,0,0,0,96,0,205,0,156,0,48,0,0,0,2,0,0,0,0,0,0,0,26,0,253,0);
signal scenario_full  : scenario_type := (0,0,111,31,111,30,142,31,102,31,140,31,196,31,138,31,87,31,87,30,231,31,208,31,172,31,122,31,122,30,122,29,244,31,244,30,110,31,110,30,18,31,245,31,156,31,166,31,114,31,145,31,145,30,170,31,134,31,28,31,28,30,28,29,201,31,239,31,135,31,38,31,62,31,125,31,16,31,182,31,176,31,22,31,22,30,239,31,255,31,255,30,255,29,4,31,4,30,243,31,247,31,80,31,245,31,86,31,197,31,206,31,20,31,51,31,151,31,223,31,223,30,223,29,80,31,104,31,229,31,61,31,61,30,94,31,94,30,190,31,249,31,23,31,162,31,187,31,120,31,120,30,247,31,247,30,159,31,109,31,80,31,166,31,54,31,152,31,152,30,59,31,181,31,146,31,190,31,99,31,69,31,48,31,160,31,13,31,72,31,58,31,58,30,41,31,77,31,243,31,243,30,244,31,131,31,61,31,137,31,62,31,163,31,49,31,8,31,69,31,4,31,86,31,173,31,250,31,45,31,45,30,195,31,143,31,143,30,148,31,235,31,38,31,90,31,90,30,90,29,249,31,251,31,194,31,194,30,80,31,9,31,119,31,204,31,204,30,54,31,206,31,205,31,70,31,29,31,10,31,126,31,144,31,41,31,161,31,161,30,103,31,30,31,47,31,1,31,243,31,243,30,243,29,227,31,20,31,67,31,143,31,38,31,14,31,169,31,2,31,101,31,47,31,47,30,7,31,18,31,18,30,50,31,131,31,101,31,59,31,213,31,213,30,195,31,91,31,237,31,237,30,88,31,88,30,88,29,108,31,52,31,98,31,98,30,171,31,171,30,171,29,42,31,42,30,50,31,230,31,131,31,238,31,133,31,133,30,133,29,145,31,153,31,92,31,92,30,147,31,166,31,166,30,166,29,226,31,226,30,62,31,89,31,82,31,142,31,142,30,201,31,201,30,12,31,66,31,5,31,3,31,3,30,6,31,6,30,186,31,186,30,101,31,101,30,101,29,101,28,254,31,154,31,241,31,232,31,213,31,108,31,147,31,47,31,163,31,68,31,104,31,198,31,90,31,90,30,30,31,30,30,83,31,17,31,103,31,55,31,34,31,9,31,63,31,102,31,93,31,224,31,148,31,232,31,232,30,100,31,69,31,69,30,39,31,39,30,194,31,194,30,63,31,203,31,39,31,44,31,200,31,208,31,201,31,166,31,231,31,21,31,48,31,48,30,17,31,64,31,129,31,255,31,211,31,68,31,224,31,173,31,162,31,220,31,118,31,29,31,148,31,43,31,163,31,130,31,221,31,139,31,139,30,139,29,237,31,106,31,106,30,106,29,71,31,147,31,231,31,74,31,38,31,181,31,181,30,208,31,208,30,243,31,243,30,190,31,156,31,254,31,254,30,213,31,30,31,30,30,143,31,24,31,165,31,12,31,100,31,198,31,198,30,198,29,198,28,148,31,94,31,94,30,190,31,76,31,35,31,35,30,235,31,226,31,217,31,107,31,234,31,159,31,191,31,195,31,87,31,126,31,226,31,231,31,43,31,35,31,163,31,173,31,162,31,122,31,86,31,86,30,13,31,137,31,146,31,174,31,214,31,75,31,106,31,106,30,205,31,144,31,172,31,172,30,158,31,158,30,7,31,7,30,7,29,96,31,205,31,156,31,48,31,48,30,2,31,2,30,2,29,2,28,26,31,253,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
