-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 175;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (51,0,140,0,82,0,124,0,81,0,135,0,200,0,0,0,145,0,0,0,62,0,70,0,0,0,0,0,255,0,140,0,98,0,103,0,181,0,44,0,102,0,187,0,0,0,52,0,206,0,47,0,0,0,130,0,38,0,15,0,0,0,0,0,55,0,0,0,55,0,28,0,182,0,219,0,23,0,213,0,0,0,42,0,180,0,84,0,60,0,110,0,0,0,47,0,100,0,0,0,76,0,237,0,0,0,150,0,2,0,50,0,127,0,170,0,41,0,66,0,48,0,224,0,0,0,93,0,12,0,0,0,89,0,94,0,129,0,230,0,58,0,184,0,0,0,124,0,0,0,122,0,3,0,138,0,129,0,83,0,167,0,205,0,254,0,19,0,0,0,25,0,0,0,50,0,151,0,100,0,0,0,4,0,0,0,0,0,235,0,57,0,120,0,1,0,159,0,5,0,0,0,0,0,163,0,46,0,0,0,54,0,147,0,0,0,234,0,0,0,4,0,134,0,226,0,50,0,187,0,0,0,201,0,97,0,98,0,154,0,246,0,143,0,92,0,8,0,11,0,247,0,177,0,89,0,206,0,88,0,98,0,0,0,89,0,110,0,249,0,119,0,10,0,0,0,193,0,79,0,98,0,0,0,0,0,83,0,0,0,217,0,181,0,192,0,139,0,200,0,5,0,0,0,146,0,136,0,79,0,195,0,192,0,211,0,242,0,203,0,0,0,197,0,161,0,5,0,34,0,173,0,182,0,136,0,254,0,0,0,166,0,78,0,111,0,0,0,177,0);
signal scenario_full  : scenario_type := (51,31,140,31,82,31,124,31,81,31,135,31,200,31,200,30,145,31,145,30,62,31,70,31,70,30,70,29,255,31,140,31,98,31,103,31,181,31,44,31,102,31,187,31,187,30,52,31,206,31,47,31,47,30,130,31,38,31,15,31,15,30,15,29,55,31,55,30,55,31,28,31,182,31,219,31,23,31,213,31,213,30,42,31,180,31,84,31,60,31,110,31,110,30,47,31,100,31,100,30,76,31,237,31,237,30,150,31,2,31,50,31,127,31,170,31,41,31,66,31,48,31,224,31,224,30,93,31,12,31,12,30,89,31,94,31,129,31,230,31,58,31,184,31,184,30,124,31,124,30,122,31,3,31,138,31,129,31,83,31,167,31,205,31,254,31,19,31,19,30,25,31,25,30,50,31,151,31,100,31,100,30,4,31,4,30,4,29,235,31,57,31,120,31,1,31,159,31,5,31,5,30,5,29,163,31,46,31,46,30,54,31,147,31,147,30,234,31,234,30,4,31,134,31,226,31,50,31,187,31,187,30,201,31,97,31,98,31,154,31,246,31,143,31,92,31,8,31,11,31,247,31,177,31,89,31,206,31,88,31,98,31,98,30,89,31,110,31,249,31,119,31,10,31,10,30,193,31,79,31,98,31,98,30,98,29,83,31,83,30,217,31,181,31,192,31,139,31,200,31,5,31,5,30,146,31,136,31,79,31,195,31,192,31,211,31,242,31,203,31,203,30,197,31,161,31,5,31,34,31,173,31,182,31,136,31,254,31,254,30,166,31,78,31,111,31,111,30,177,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
