-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 192;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,183,0,10,0,107,0,0,0,2,0,17,0,217,0,164,0,0,0,220,0,156,0,47,0,168,0,0,0,98,0,157,0,154,0,198,0,52,0,33,0,0,0,97,0,42,0,233,0,173,0,97,0,84,0,56,0,146,0,0,0,64,0,121,0,59,0,0,0,62,0,192,0,28,0,46,0,170,0,87,0,126,0,160,0,0,0,101,0,34,0,0,0,0,0,243,0,0,0,206,0,19,0,0,0,50,0,0,0,235,0,196,0,74,0,171,0,0,0,237,0,119,0,117,0,116,0,246,0,52,0,164,0,86,0,107,0,175,0,187,0,0,0,9,0,202,0,211,0,0,0,145,0,253,0,225,0,1,0,122,0,35,0,67,0,157,0,122,0,0,0,105,0,182,0,137,0,0,0,167,0,115,0,201,0,85,0,0,0,93,0,0,0,115,0,233,0,231,0,0,0,156,0,0,0,196,0,211,0,228,0,92,0,227,0,248,0,81,0,81,0,64,0,0,0,22,0,175,0,49,0,122,0,27,0,168,0,9,0,171,0,0,0,63,0,0,0,188,0,227,0,120,0,46,0,0,0,130,0,219,0,78,0,210,0,211,0,148,0,50,0,235,0,255,0,96,0,8,0,224,0,0,0,39,0,254,0,155,0,0,0,203,0,0,0,216,0,0,0,0,0,148,0,76,0,0,0,0,0,176,0,0,0,0,0,117,0,122,0,119,0,139,0,104,0,0,0,67,0,176,0,184,0,189,0,118,0,0,0,0,0,188,0,33,0,242,0,0,0,76,0,0,0,111,0,103,0,178,0,70,0,25,0,0,0,247,0,156,0,222,0,0,0,177,0,165,0,144,0,0,0,229,0);
signal scenario_full  : scenario_type := (147,31,183,31,10,31,107,31,107,30,2,31,17,31,217,31,164,31,164,30,220,31,156,31,47,31,168,31,168,30,98,31,157,31,154,31,198,31,52,31,33,31,33,30,97,31,42,31,233,31,173,31,97,31,84,31,56,31,146,31,146,30,64,31,121,31,59,31,59,30,62,31,192,31,28,31,46,31,170,31,87,31,126,31,160,31,160,30,101,31,34,31,34,30,34,29,243,31,243,30,206,31,19,31,19,30,50,31,50,30,235,31,196,31,74,31,171,31,171,30,237,31,119,31,117,31,116,31,246,31,52,31,164,31,86,31,107,31,175,31,187,31,187,30,9,31,202,31,211,31,211,30,145,31,253,31,225,31,1,31,122,31,35,31,67,31,157,31,122,31,122,30,105,31,182,31,137,31,137,30,167,31,115,31,201,31,85,31,85,30,93,31,93,30,115,31,233,31,231,31,231,30,156,31,156,30,196,31,211,31,228,31,92,31,227,31,248,31,81,31,81,31,64,31,64,30,22,31,175,31,49,31,122,31,27,31,168,31,9,31,171,31,171,30,63,31,63,30,188,31,227,31,120,31,46,31,46,30,130,31,219,31,78,31,210,31,211,31,148,31,50,31,235,31,255,31,96,31,8,31,224,31,224,30,39,31,254,31,155,31,155,30,203,31,203,30,216,31,216,30,216,29,148,31,76,31,76,30,76,29,176,31,176,30,176,29,117,31,122,31,119,31,139,31,104,31,104,30,67,31,176,31,184,31,189,31,118,31,118,30,118,29,188,31,33,31,242,31,242,30,76,31,76,30,111,31,103,31,178,31,70,31,25,31,25,30,247,31,156,31,222,31,222,30,177,31,165,31,144,31,144,30,229,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
