-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 567;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (91,0,49,0,181,0,99,0,249,0,18,0,58,0,38,0,57,0,15,0,229,0,85,0,0,0,36,0,0,0,218,0,2,0,0,0,84,0,63,0,0,0,17,0,0,0,0,0,0,0,145,0,0,0,204,0,208,0,122,0,0,0,214,0,231,0,63,0,134,0,6,0,252,0,16,0,111,0,236,0,108,0,3,0,0,0,210,0,146,0,184,0,111,0,166,0,151,0,226,0,74,0,99,0,33,0,128,0,0,0,0,0,111,0,121,0,115,0,48,0,114,0,0,0,158,0,45,0,236,0,0,0,170,0,120,0,0,0,0,0,123,0,239,0,99,0,10,0,0,0,200,0,33,0,252,0,0,0,145,0,191,0,0,0,24,0,26,0,0,0,133,0,190,0,67,0,150,0,214,0,34,0,241,0,98,0,0,0,244,0,90,0,95,0,183,0,0,0,55,0,103,0,167,0,122,0,22,0,212,0,123,0,0,0,111,0,83,0,225,0,97,0,219,0,101,0,103,0,135,0,210,0,98,0,0,0,206,0,13,0,36,0,0,0,197,0,68,0,10,0,109,0,55,0,93,0,179,0,255,0,0,0,91,0,0,0,189,0,92,0,44,0,53,0,38,0,76,0,0,0,180,0,185,0,238,0,160,0,0,0,122,0,66,0,0,0,121,0,23,0,167,0,0,0,0,0,177,0,0,0,225,0,202,0,101,0,151,0,55,0,122,0,169,0,233,0,0,0,85,0,198,0,0,0,41,0,0,0,220,0,70,0,180,0,78,0,135,0,41,0,146,0,15,0,0,0,43,0,37,0,144,0,130,0,205,0,0,0,215,0,117,0,44,0,154,0,203,0,77,0,0,0,8,0,0,0,109,0,91,0,255,0,98,0,175,0,0,0,6,0,190,0,41,0,172,0,0,0,124,0,208,0,29,0,85,0,187,0,0,0,226,0,0,0,0,0,98,0,170,0,124,0,0,0,252,0,187,0,174,0,225,0,192,0,185,0,35,0,224,0,56,0,157,0,154,0,238,0,51,0,0,0,0,0,243,0,234,0,0,0,117,0,111,0,71,0,164,0,96,0,182,0,187,0,0,0,83,0,14,0,0,0,95,0,0,0,0,0,0,0,0,0,74,0,61,0,206,0,0,0,254,0,167,0,0,0,208,0,116,0,118,0,213,0,136,0,0,0,0,0,247,0,131,0,60,0,15,0,181,0,0,0,185,0,229,0,104,0,226,0,0,0,176,0,185,0,147,0,57,0,21,0,253,0,120,0,162,0,7,0,191,0,173,0,0,0,187,0,20,0,20,0,176,0,144,0,48,0,111,0,3,0,64,0,158,0,214,0,0,0,150,0,116,0,67,0,0,0,0,0,56,0,119,0,48,0,0,0,224,0,199,0,184,0,181,0,36,0,0,0,179,0,173,0,92,0,189,0,113,0,0,0,193,0,0,0,77,0,243,0,0,0,85,0,205,0,136,0,43,0,190,0,173,0,74,0,180,0,229,0,198,0,185,0,59,0,137,0,0,0,178,0,106,0,70,0,0,0,190,0,67,0,37,0,216,0,164,0,0,0,252,0,130,0,209,0,232,0,0,0,0,0,3,0,0,0,0,0,0,0,225,0,21,0,108,0,66,0,0,0,110,0,211,0,167,0,50,0,0,0,10,0,204,0,64,0,0,0,178,0,194,0,0,0,99,0,177,0,255,0,151,0,0,0,0,0,106,0,211,0,251,0,32,0,159,0,224,0,0,0,148,0,78,0,70,0,41,0,0,0,216,0,145,0,0,0,0,0,0,0,25,0,0,0,0,0,71,0,233,0,5,0,0,0,31,0,0,0,72,0,0,0,226,0,22,0,28,0,86,0,75,0,189,0,223,0,122,0,152,0,3,0,84,0,246,0,254,0,129,0,226,0,201,0,198,0,231,0,156,0,0,0,127,0,83,0,247,0,0,0,27,0,0,0,94,0,0,0,242,0,0,0,0,0,26,0,248,0,0,0,0,0,201,0,0,0,91,0,0,0,0,0,194,0,63,0,149,0,168,0,174,0,93,0,193,0,246,0,125,0,0,0,0,0,15,0,92,0,244,0,245,0,15,0,0,0,117,0,119,0,0,0,146,0,0,0,96,0,0,0,170,0,20,0,0,0,0,0,111,0,141,0,81,0,189,0,228,0,238,0,148,0,117,0,96,0,179,0,68,0,26,0,126,0,214,0,174,0,52,0,32,0,0,0,168,0,37,0,192,0,107,0,0,0,43,0,251,0,0,0,202,0,242,0,164,0,0,0,0,0,200,0,195,0,0,0,34,0,60,0,222,0,55,0,75,0,53,0,0,0,0,0,99,0,0,0,102,0,0,0,131,0,0,0,0,0,146,0,55,0,130,0,226,0,0,0,0,0,84,0,199,0,40,0,119,0,0,0,36,0,248,0,154,0,0,0,197,0,0,0,0,0,37,0,199,0,0,0,67,0,254,0,165,0,182,0,0,0,66,0,0,0,89,0,236,0,102,0,29,0,206,0,0,0,144,0,178,0,78,0,128,0,119,0);
signal scenario_full  : scenario_type := (91,31,49,31,181,31,99,31,249,31,18,31,58,31,38,31,57,31,15,31,229,31,85,31,85,30,36,31,36,30,218,31,2,31,2,30,84,31,63,31,63,30,17,31,17,30,17,29,17,28,145,31,145,30,204,31,208,31,122,31,122,30,214,31,231,31,63,31,134,31,6,31,252,31,16,31,111,31,236,31,108,31,3,31,3,30,210,31,146,31,184,31,111,31,166,31,151,31,226,31,74,31,99,31,33,31,128,31,128,30,128,29,111,31,121,31,115,31,48,31,114,31,114,30,158,31,45,31,236,31,236,30,170,31,120,31,120,30,120,29,123,31,239,31,99,31,10,31,10,30,200,31,33,31,252,31,252,30,145,31,191,31,191,30,24,31,26,31,26,30,133,31,190,31,67,31,150,31,214,31,34,31,241,31,98,31,98,30,244,31,90,31,95,31,183,31,183,30,55,31,103,31,167,31,122,31,22,31,212,31,123,31,123,30,111,31,83,31,225,31,97,31,219,31,101,31,103,31,135,31,210,31,98,31,98,30,206,31,13,31,36,31,36,30,197,31,68,31,10,31,109,31,55,31,93,31,179,31,255,31,255,30,91,31,91,30,189,31,92,31,44,31,53,31,38,31,76,31,76,30,180,31,185,31,238,31,160,31,160,30,122,31,66,31,66,30,121,31,23,31,167,31,167,30,167,29,177,31,177,30,225,31,202,31,101,31,151,31,55,31,122,31,169,31,233,31,233,30,85,31,198,31,198,30,41,31,41,30,220,31,70,31,180,31,78,31,135,31,41,31,146,31,15,31,15,30,43,31,37,31,144,31,130,31,205,31,205,30,215,31,117,31,44,31,154,31,203,31,77,31,77,30,8,31,8,30,109,31,91,31,255,31,98,31,175,31,175,30,6,31,190,31,41,31,172,31,172,30,124,31,208,31,29,31,85,31,187,31,187,30,226,31,226,30,226,29,98,31,170,31,124,31,124,30,252,31,187,31,174,31,225,31,192,31,185,31,35,31,224,31,56,31,157,31,154,31,238,31,51,31,51,30,51,29,243,31,234,31,234,30,117,31,111,31,71,31,164,31,96,31,182,31,187,31,187,30,83,31,14,31,14,30,95,31,95,30,95,29,95,28,95,27,74,31,61,31,206,31,206,30,254,31,167,31,167,30,208,31,116,31,118,31,213,31,136,31,136,30,136,29,247,31,131,31,60,31,15,31,181,31,181,30,185,31,229,31,104,31,226,31,226,30,176,31,185,31,147,31,57,31,21,31,253,31,120,31,162,31,7,31,191,31,173,31,173,30,187,31,20,31,20,31,176,31,144,31,48,31,111,31,3,31,64,31,158,31,214,31,214,30,150,31,116,31,67,31,67,30,67,29,56,31,119,31,48,31,48,30,224,31,199,31,184,31,181,31,36,31,36,30,179,31,173,31,92,31,189,31,113,31,113,30,193,31,193,30,77,31,243,31,243,30,85,31,205,31,136,31,43,31,190,31,173,31,74,31,180,31,229,31,198,31,185,31,59,31,137,31,137,30,178,31,106,31,70,31,70,30,190,31,67,31,37,31,216,31,164,31,164,30,252,31,130,31,209,31,232,31,232,30,232,29,3,31,3,30,3,29,3,28,225,31,21,31,108,31,66,31,66,30,110,31,211,31,167,31,50,31,50,30,10,31,204,31,64,31,64,30,178,31,194,31,194,30,99,31,177,31,255,31,151,31,151,30,151,29,106,31,211,31,251,31,32,31,159,31,224,31,224,30,148,31,78,31,70,31,41,31,41,30,216,31,145,31,145,30,145,29,145,28,25,31,25,30,25,29,71,31,233,31,5,31,5,30,31,31,31,30,72,31,72,30,226,31,22,31,28,31,86,31,75,31,189,31,223,31,122,31,152,31,3,31,84,31,246,31,254,31,129,31,226,31,201,31,198,31,231,31,156,31,156,30,127,31,83,31,247,31,247,30,27,31,27,30,94,31,94,30,242,31,242,30,242,29,26,31,248,31,248,30,248,29,201,31,201,30,91,31,91,30,91,29,194,31,63,31,149,31,168,31,174,31,93,31,193,31,246,31,125,31,125,30,125,29,15,31,92,31,244,31,245,31,15,31,15,30,117,31,119,31,119,30,146,31,146,30,96,31,96,30,170,31,20,31,20,30,20,29,111,31,141,31,81,31,189,31,228,31,238,31,148,31,117,31,96,31,179,31,68,31,26,31,126,31,214,31,174,31,52,31,32,31,32,30,168,31,37,31,192,31,107,31,107,30,43,31,251,31,251,30,202,31,242,31,164,31,164,30,164,29,200,31,195,31,195,30,34,31,60,31,222,31,55,31,75,31,53,31,53,30,53,29,99,31,99,30,102,31,102,30,131,31,131,30,131,29,146,31,55,31,130,31,226,31,226,30,226,29,84,31,199,31,40,31,119,31,119,30,36,31,248,31,154,31,154,30,197,31,197,30,197,29,37,31,199,31,199,30,67,31,254,31,165,31,182,31,182,30,66,31,66,30,89,31,236,31,102,31,29,31,206,31,206,30,144,31,178,31,78,31,128,31,119,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
