-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 784;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,114,0,61,0,0,0,0,0,209,0,0,0,153,0,145,0,48,0,171,0,63,0,125,0,234,0,218,0,189,0,0,0,65,0,47,0,5,0,93,0,214,0,0,0,218,0,31,0,31,0,0,0,0,0,197,0,61,0,171,0,93,0,135,0,183,0,96,0,188,0,15,0,186,0,0,0,195,0,229,0,226,0,187,0,246,0,165,0,0,0,188,0,176,0,252,0,32,0,0,0,167,0,119,0,0,0,58,0,251,0,134,0,8,0,224,0,0,0,5,0,0,0,67,0,0,0,235,0,0,0,138,0,19,0,116,0,253,0,210,0,56,0,133,0,253,0,1,0,0,0,230,0,128,0,209,0,0,0,143,0,136,0,183,0,226,0,56,0,93,0,136,0,86,0,227,0,255,0,166,0,223,0,105,0,88,0,115,0,40,0,177,0,254,0,0,0,167,0,17,0,132,0,18,0,219,0,0,0,43,0,29,0,71,0,116,0,31,0,38,0,243,0,0,0,157,0,37,0,0,0,177,0,10,0,27,0,168,0,162,0,188,0,159,0,64,0,141,0,0,0,200,0,158,0,164,0,12,0,219,0,0,0,0,0,8,0,138,0,174,0,0,0,88,0,0,0,236,0,96,0,115,0,0,0,155,0,107,0,103,0,244,0,0,0,107,0,143,0,178,0,96,0,98,0,124,0,161,0,241,0,0,0,9,0,0,0,70,0,110,0,153,0,81,0,41,0,73,0,79,0,126,0,94,0,0,0,56,0,109,0,150,0,165,0,0,0,176,0,116,0,87,0,12,0,119,0,218,0,150,0,134,0,61,0,106,0,25,0,0,0,0,0,104,0,0,0,118,0,157,0,233,0,4,0,33,0,118,0,211,0,125,0,181,0,0,0,194,0,175,0,0,0,168,0,0,0,0,0,40,0,228,0,201,0,184,0,0,0,200,0,73,0,25,0,137,0,0,0,153,0,235,0,83,0,0,0,71,0,229,0,91,0,218,0,0,0,0,0,91,0,111,0,45,0,131,0,91,0,55,0,94,0,191,0,144,0,176,0,253,0,14,0,101,0,48,0,23,0,215,0,190,0,202,0,164,0,110,0,0,0,0,0,128,0,60,0,192,0,73,0,138,0,171,0,34,0,129,0,0,0,18,0,34,0,0,0,194,0,48,0,31,0,219,0,196,0,0,0,2,0,137,0,5,0,199,0,113,0,197,0,101,0,8,0,212,0,44,0,182,0,111,0,241,0,39,0,242,0,207,0,252,0,128,0,0,0,154,0,0,0,164,0,167,0,194,0,97,0,31,0,7,0,246,0,216,0,153,0,17,0,136,0,152,0,0,0,185,0,87,0,25,0,67,0,252,0,134,0,0,0,0,0,17,0,0,0,70,0,124,0,0,0,150,0,92,0,18,0,131,0,160,0,165,0,156,0,242,0,0,0,223,0,135,0,167,0,175,0,72,0,0,0,220,0,0,0,45,0,67,0,100,0,192,0,156,0,189,0,201,0,0,0,0,0,38,0,60,0,106,0,137,0,83,0,101,0,123,0,0,0,0,0,56,0,0,0,175,0,186,0,226,0,30,0,217,0,0,0,17,0,27,0,0,0,212,0,100,0,145,0,45,0,199,0,76,0,7,0,34,0,0,0,0,0,68,0,187,0,66,0,23,0,150,0,0,0,10,0,119,0,0,0,204,0,249,0,0,0,163,0,141,0,186,0,58,0,222,0,14,0,221,0,227,0,175,0,0,0,0,0,18,0,51,0,41,0,142,0,125,0,235,0,243,0,192,0,235,0,126,0,11,0,5,0,0,0,239,0,53,0,0,0,128,0,0,0,177,0,135,0,0,0,0,0,120,0,50,0,168,0,0,0,0,0,185,0,0,0,0,0,99,0,239,0,0,0,153,0,235,0,151,0,37,0,196,0,125,0,98,0,24,0,193,0,129,0,51,0,0,0,55,0,117,0,55,0,85,0,55,0,0,0,0,0,111,0,0,0,19,0,196,0,133,0,219,0,0,0,158,0,0,0,0,0,151,0,185,0,230,0,106,0,60,0,142,0,0,0,0,0,72,0,195,0,81,0,115,0,0,0,153,0,0,0,221,0,90,0,161,0,36,0,10,0,118,0,0,0,46,0,2,0,225,0,218,0,20,0,217,0,140,0,197,0,222,0,127,0,103,0,162,0,0,0,180,0,89,0,67,0,243,0,0,0,237,0,0,0,80,0,0,0,103,0,59,0,222,0,29,0,0,0,142,0,0,0,152,0,175,0,0,0,0,0,144,0,109,0,97,0,234,0,20,0,99,0,0,0,5,0,250,0,134,0,119,0,228,0,101,0,171,0,227,0,206,0,0,0,243,0,127,0,45,0,32,0,19,0,145,0,112,0,69,0,218,0,237,0,241,0,57,0,134,0,36,0,0,0,0,0,93,0,81,0,123,0,0,0,121,0,84,0,161,0,142,0,61,0,188,0,0,0,0,0,126,0,2,0,199,0,103,0,247,0,57,0,131,0,107,0,146,0,26,0,0,0,199,0,132,0,0,0,0,0,19,0,254,0,92,0,83,0,115,0,124,0,160,0,0,0,156,0,251,0,0,0,158,0,0,0,172,0,0,0,115,0,195,0,105,0,140,0,241,0,137,0,89,0,157,0,32,0,238,0,193,0,0,0,0,0,187,0,43,0,152,0,85,0,32,0,38,0,0,0,0,0,0,0,153,0,83,0,0,0,76,0,100,0,50,0,0,0,186,0,209,0,202,0,0,0,11,0,30,0,221,0,0,0,0,0,183,0,33,0,226,0,130,0,94,0,33,0,28,0,158,0,0,0,64,0,80,0,187,0,0,0,188,0,74,0,181,0,129,0,133,0,162,0,186,0,25,0,244,0,0,0,0,0,0,0,31,0,72,0,51,0,0,0,251,0,201,0,0,0,236,0,50,0,155,0,217,0,116,0,129,0,130,0,237,0,242,0,136,0,0,0,0,0,13,0,0,0,0,0,67,0,36,0,100,0,0,0,222,0,155,0,192,0,192,0,216,0,169,0,39,0,198,0,193,0,149,0,171,0,223,0,14,0,0,0,243,0,0,0,192,0,179,0,247,0,2,0,0,0,234,0,116,0,102,0,226,0,213,0,238,0,68,0,129,0,0,0,0,0,92,0,166,0,200,0,34,0,98,0,129,0,56,0,238,0,243,0,177,0,12,0,116,0,244,0,170,0,144,0,0,0,0,0,94,0,154,0,3,0,214,0,135,0,114,0,80,0,202,0,153,0,211,0,0,0,142,0,92,0,35,0,0,0,100,0,0,0,11,0,208,0,0,0,54,0,38,0,189,0,164,0,0,0,0,0,0,0,177,0,5,0,140,0,79,0,168,0,198,0,128,0,190,0,207,0,196,0,33,0,22,0,0,0,82,0,212,0,121,0,234,0,162,0,30,0,214,0,254,0,236,0,252,0,0,0,0,0,48,0,80,0,28,0,13,0,173,0,188,0,7,0,0,0,22,0,154,0,0,0,54,0);
signal scenario_full  : scenario_type := (197,31,114,31,61,31,61,30,61,29,209,31,209,30,153,31,145,31,48,31,171,31,63,31,125,31,234,31,218,31,189,31,189,30,65,31,47,31,5,31,93,31,214,31,214,30,218,31,31,31,31,31,31,30,31,29,197,31,61,31,171,31,93,31,135,31,183,31,96,31,188,31,15,31,186,31,186,30,195,31,229,31,226,31,187,31,246,31,165,31,165,30,188,31,176,31,252,31,32,31,32,30,167,31,119,31,119,30,58,31,251,31,134,31,8,31,224,31,224,30,5,31,5,30,67,31,67,30,235,31,235,30,138,31,19,31,116,31,253,31,210,31,56,31,133,31,253,31,1,31,1,30,230,31,128,31,209,31,209,30,143,31,136,31,183,31,226,31,56,31,93,31,136,31,86,31,227,31,255,31,166,31,223,31,105,31,88,31,115,31,40,31,177,31,254,31,254,30,167,31,17,31,132,31,18,31,219,31,219,30,43,31,29,31,71,31,116,31,31,31,38,31,243,31,243,30,157,31,37,31,37,30,177,31,10,31,27,31,168,31,162,31,188,31,159,31,64,31,141,31,141,30,200,31,158,31,164,31,12,31,219,31,219,30,219,29,8,31,138,31,174,31,174,30,88,31,88,30,236,31,96,31,115,31,115,30,155,31,107,31,103,31,244,31,244,30,107,31,143,31,178,31,96,31,98,31,124,31,161,31,241,31,241,30,9,31,9,30,70,31,110,31,153,31,81,31,41,31,73,31,79,31,126,31,94,31,94,30,56,31,109,31,150,31,165,31,165,30,176,31,116,31,87,31,12,31,119,31,218,31,150,31,134,31,61,31,106,31,25,31,25,30,25,29,104,31,104,30,118,31,157,31,233,31,4,31,33,31,118,31,211,31,125,31,181,31,181,30,194,31,175,31,175,30,168,31,168,30,168,29,40,31,228,31,201,31,184,31,184,30,200,31,73,31,25,31,137,31,137,30,153,31,235,31,83,31,83,30,71,31,229,31,91,31,218,31,218,30,218,29,91,31,111,31,45,31,131,31,91,31,55,31,94,31,191,31,144,31,176,31,253,31,14,31,101,31,48,31,23,31,215,31,190,31,202,31,164,31,110,31,110,30,110,29,128,31,60,31,192,31,73,31,138,31,171,31,34,31,129,31,129,30,18,31,34,31,34,30,194,31,48,31,31,31,219,31,196,31,196,30,2,31,137,31,5,31,199,31,113,31,197,31,101,31,8,31,212,31,44,31,182,31,111,31,241,31,39,31,242,31,207,31,252,31,128,31,128,30,154,31,154,30,164,31,167,31,194,31,97,31,31,31,7,31,246,31,216,31,153,31,17,31,136,31,152,31,152,30,185,31,87,31,25,31,67,31,252,31,134,31,134,30,134,29,17,31,17,30,70,31,124,31,124,30,150,31,92,31,18,31,131,31,160,31,165,31,156,31,242,31,242,30,223,31,135,31,167,31,175,31,72,31,72,30,220,31,220,30,45,31,67,31,100,31,192,31,156,31,189,31,201,31,201,30,201,29,38,31,60,31,106,31,137,31,83,31,101,31,123,31,123,30,123,29,56,31,56,30,175,31,186,31,226,31,30,31,217,31,217,30,17,31,27,31,27,30,212,31,100,31,145,31,45,31,199,31,76,31,7,31,34,31,34,30,34,29,68,31,187,31,66,31,23,31,150,31,150,30,10,31,119,31,119,30,204,31,249,31,249,30,163,31,141,31,186,31,58,31,222,31,14,31,221,31,227,31,175,31,175,30,175,29,18,31,51,31,41,31,142,31,125,31,235,31,243,31,192,31,235,31,126,31,11,31,5,31,5,30,239,31,53,31,53,30,128,31,128,30,177,31,135,31,135,30,135,29,120,31,50,31,168,31,168,30,168,29,185,31,185,30,185,29,99,31,239,31,239,30,153,31,235,31,151,31,37,31,196,31,125,31,98,31,24,31,193,31,129,31,51,31,51,30,55,31,117,31,55,31,85,31,55,31,55,30,55,29,111,31,111,30,19,31,196,31,133,31,219,31,219,30,158,31,158,30,158,29,151,31,185,31,230,31,106,31,60,31,142,31,142,30,142,29,72,31,195,31,81,31,115,31,115,30,153,31,153,30,221,31,90,31,161,31,36,31,10,31,118,31,118,30,46,31,2,31,225,31,218,31,20,31,217,31,140,31,197,31,222,31,127,31,103,31,162,31,162,30,180,31,89,31,67,31,243,31,243,30,237,31,237,30,80,31,80,30,103,31,59,31,222,31,29,31,29,30,142,31,142,30,152,31,175,31,175,30,175,29,144,31,109,31,97,31,234,31,20,31,99,31,99,30,5,31,250,31,134,31,119,31,228,31,101,31,171,31,227,31,206,31,206,30,243,31,127,31,45,31,32,31,19,31,145,31,112,31,69,31,218,31,237,31,241,31,57,31,134,31,36,31,36,30,36,29,93,31,81,31,123,31,123,30,121,31,84,31,161,31,142,31,61,31,188,31,188,30,188,29,126,31,2,31,199,31,103,31,247,31,57,31,131,31,107,31,146,31,26,31,26,30,199,31,132,31,132,30,132,29,19,31,254,31,92,31,83,31,115,31,124,31,160,31,160,30,156,31,251,31,251,30,158,31,158,30,172,31,172,30,115,31,195,31,105,31,140,31,241,31,137,31,89,31,157,31,32,31,238,31,193,31,193,30,193,29,187,31,43,31,152,31,85,31,32,31,38,31,38,30,38,29,38,28,153,31,83,31,83,30,76,31,100,31,50,31,50,30,186,31,209,31,202,31,202,30,11,31,30,31,221,31,221,30,221,29,183,31,33,31,226,31,130,31,94,31,33,31,28,31,158,31,158,30,64,31,80,31,187,31,187,30,188,31,74,31,181,31,129,31,133,31,162,31,186,31,25,31,244,31,244,30,244,29,244,28,31,31,72,31,51,31,51,30,251,31,201,31,201,30,236,31,50,31,155,31,217,31,116,31,129,31,130,31,237,31,242,31,136,31,136,30,136,29,13,31,13,30,13,29,67,31,36,31,100,31,100,30,222,31,155,31,192,31,192,31,216,31,169,31,39,31,198,31,193,31,149,31,171,31,223,31,14,31,14,30,243,31,243,30,192,31,179,31,247,31,2,31,2,30,234,31,116,31,102,31,226,31,213,31,238,31,68,31,129,31,129,30,129,29,92,31,166,31,200,31,34,31,98,31,129,31,56,31,238,31,243,31,177,31,12,31,116,31,244,31,170,31,144,31,144,30,144,29,94,31,154,31,3,31,214,31,135,31,114,31,80,31,202,31,153,31,211,31,211,30,142,31,92,31,35,31,35,30,100,31,100,30,11,31,208,31,208,30,54,31,38,31,189,31,164,31,164,30,164,29,164,28,177,31,5,31,140,31,79,31,168,31,198,31,128,31,190,31,207,31,196,31,33,31,22,31,22,30,82,31,212,31,121,31,234,31,162,31,30,31,214,31,254,31,236,31,252,31,252,30,252,29,48,31,80,31,28,31,13,31,173,31,188,31,7,31,7,30,22,31,154,31,154,30,54,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
