-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_601 is
end project_tb_601;

architecture project_tb_arch_601 of project_tb_601 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 897;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,243,0,0,0,165,0,8,0,79,0,119,0,250,0,0,0,0,0,0,0,221,0,229,0,0,0,101,0,82,0,23,0,128,0,107,0,10,0,133,0,182,0,0,0,86,0,57,0,0,0,32,0,1,0,0,0,130,0,0,0,0,0,252,0,192,0,161,0,134,0,117,0,202,0,83,0,48,0,0,0,172,0,70,0,31,0,23,0,113,0,121,0,0,0,127,0,177,0,11,0,14,0,87,0,134,0,60,0,161,0,0,0,169,0,28,0,89,0,145,0,203,0,75,0,183,0,0,0,226,0,221,0,39,0,0,0,55,0,133,0,217,0,251,0,225,0,117,0,189,0,167,0,241,0,179,0,35,0,168,0,66,0,17,0,167,0,1,0,163,0,0,0,1,0,36,0,82,0,253,0,81,0,162,0,43,0,0,0,0,0,68,0,44,0,0,0,160,0,229,0,110,0,117,0,0,0,203,0,170,0,0,0,23,0,141,0,0,0,14,0,210,0,202,0,113,0,133,0,0,0,233,0,186,0,0,0,0,0,0,0,0,0,0,0,143,0,84,0,228,0,165,0,84,0,134,0,0,0,79,0,247,0,27,0,158,0,121,0,0,0,0,0,236,0,225,0,0,0,106,0,156,0,86,0,0,0,254,0,79,0,38,0,121,0,0,0,191,0,20,0,24,0,249,0,36,0,200,0,0,0,184,0,109,0,73,0,228,0,140,0,14,0,90,0,0,0,141,0,245,0,5,0,124,0,58,0,132,0,113,0,52,0,85,0,38,0,71,0,44,0,33,0,122,0,251,0,41,0,191,0,145,0,7,0,113,0,0,0,170,0,119,0,64,0,18,0,143,0,0,0,0,0,0,0,207,0,140,0,8,0,0,0,196,0,147,0,0,0,202,0,0,0,180,0,101,0,119,0,0,0,184,0,192,0,188,0,69,0,129,0,104,0,116,0,0,0,0,0,139,0,55,0,0,0,193,0,92,0,0,0,0,0,160,0,168,0,226,0,123,0,51,0,26,0,64,0,131,0,0,0,74,0,255,0,9,0,56,0,64,0,254,0,0,0,239,0,86,0,124,0,113,0,146,0,142,0,133,0,0,0,203,0,188,0,232,0,59,0,167,0,0,0,0,0,187,0,0,0,11,0,193,0,13,0,195,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,57,0,0,0,177,0,174,0,246,0,0,0,8,0,223,0,99,0,19,0,30,0,0,0,0,0,18,0,0,0,20,0,110,0,125,0,54,0,237,0,178,0,24,0,129,0,70,0,10,0,65,0,151,0,56,0,185,0,175,0,202,0,138,0,165,0,40,0,100,0,106,0,122,0,248,0,116,0,118,0,201,0,151,0,188,0,250,0,0,0,0,0,0,0,127,0,0,0,99,0,202,0,0,0,88,0,124,0,23,0,57,0,206,0,7,0,161,0,141,0,11,0,0,0,228,0,196,0,231,0,238,0,34,0,117,0,141,0,0,0,167,0,155,0,0,0,182,0,105,0,231,0,0,0,202,0,208,0,180,0,208,0,240,0,252,0,169,0,0,0,98,0,0,0,0,0,13,0,0,0,0,0,135,0,133,0,86,0,89,0,0,0,0,0,44,0,247,0,154,0,36,0,57,0,0,0,81,0,120,0,255,0,181,0,175,0,0,0,27,0,75,0,10,0,155,0,168,0,32,0,81,0,252,0,124,0,0,0,169,0,248,0,88,0,198,0,0,0,38,0,157,0,131,0,146,0,70,0,0,0,136,0,0,0,103,0,111,0,169,0,0,0,161,0,153,0,120,0,197,0,44,0,0,0,0,0,61,0,218,0,41,0,46,0,0,0,108,0,28,0,0,0,121,0,184,0,0,0,174,0,229,0,0,0,154,0,70,0,80,0,144,0,180,0,50,0,203,0,0,0,186,0,88,0,147,0,0,0,64,0,76,0,64,0,156,0,234,0,0,0,32,0,8,0,0,0,237,0,0,0,86,0,128,0,59,0,0,0,170,0,196,0,0,0,75,0,30,0,192,0,223,0,61,0,0,0,228,0,91,0,0,0,56,0,137,0,226,0,202,0,161,0,157,0,0,0,169,0,187,0,98,0,0,0,173,0,99,0,127,0,0,0,182,0,0,0,15,0,252,0,107,0,0,0,231,0,16,0,0,0,0,0,20,0,186,0,0,0,63,0,250,0,197,0,137,0,204,0,195,0,135,0,213,0,247,0,142,0,32,0,155,0,72,0,172,0,95,0,170,0,0,0,204,0,14,0,213,0,0,0,149,0,153,0,111,0,248,0,206,0,103,0,197,0,244,0,0,0,218,0,119,0,202,0,0,0,0,0,224,0,46,0,198,0,0,0,242,0,222,0,180,0,0,0,83,0,140,0,140,0,0,0,218,0,226,0,177,0,67,0,96,0,0,0,52,0,0,0,175,0,44,0,242,0,0,0,0,0,83,0,17,0,49,0,222,0,87,0,98,0,234,0,38,0,178,0,230,0,215,0,175,0,221,0,181,0,252,0,0,0,0,0,84,0,8,0,240,0,60,0,64,0,0,0,156,0,0,0,95,0,203,0,94,0,116,0,167,0,187,0,0,0,220,0,0,0,0,0,46,0,50,0,118,0,0,0,0,0,196,0,108,0,145,0,35,0,10,0,192,0,0,0,24,0,45,0,12,0,0,0,155,0,185,0,85,0,166,0,0,0,0,0,252,0,66,0,57,0,0,0,80,0,196,0,31,0,0,0,56,0,0,0,169,0,0,0,99,0,12,0,175,0,50,0,0,0,38,0,253,0,119,0,47,0,7,0,0,0,0,0,200,0,245,0,175,0,0,0,10,0,250,0,0,0,151,0,92,0,177,0,222,0,196,0,206,0,36,0,0,0,0,0,75,0,0,0,0,0,10,0,74,0,58,0,145,0,165,0,0,0,203,0,117,0,45,0,0,0,131,0,140,0,140,0,0,0,111,0,15,0,94,0,46,0,59,0,22,0,238,0,2,0,181,0,56,0,155,0,255,0,115,0,250,0,164,0,177,0,213,0,91,0,200,0,127,0,0,0,0,0,140,0,157,0,102,0,0,0,48,0,199,0,208,0,145,0,149,0,197,0,17,0,69,0,202,0,73,0,68,0,194,0,240,0,1,0,100,0,215,0,0,0,0,0,28,0,127,0,0,0,213,0,241,0,98,0,131,0,161,0,51,0,22,0,0,0,0,0,80,0,20,0,19,0,126,0,92,0,0,0,80,0,67,0,0,0,28,0,219,0,0,0,17,0,73,0,0,0,246,0,250,0,194,0,254,0,99,0,24,0,141,0,249,0,0,0,146,0,0,0,0,0,187,0,0,0,0,0,0,0,24,0,173,0,80,0,90,0,0,0,66,0,145,0,210,0,76,0,249,0,45,0,130,0,75,0,236,0,9,0,0,0,185,0,131,0,198,0,182,0,0,0,185,0,86,0,179,0,244,0,16,0,103,0,231,0,176,0,61,0,251,0,0,0,0,0,28,0,0,0,140,0,26,0,172,0,24,0,247,0,117,0,0,0,80,0,0,0,132,0,16,0,232,0,246,0,203,0,0,0,0,0,72,0,30,0,230,0,117,0,231,0,253,0,218,0,0,0,16,0,146,0,0,0,108,0,244,0,159,0,46,0,125,0,173,0,96,0,0,0,0,0,16,0,34,0,70,0,205,0,109,0,105,0,189,0,70,0,123,0,0,0,191,0,181,0,175,0,179,0,0,0,0,0,57,0,211,0,1,0,59,0,51,0,0,0,106,0,206,0,54,0,62,0,34,0,243,0,85,0,0,0,0,0,207,0,61,0,85,0,0,0,96,0,11,0,8,0,100,0,237,0,0,0,227,0,0,0,130,0,156,0,0,0,16,0,0,0,73,0,225,0,40,0,0,0,116,0,0,0,178,0,242,0,137,0,136,0,26,0,116,0,28,0,0,0,150,0,177,0,227,0,0,0,84,0,6,0,243,0,115,0,92,0,11,0,173,0,211,0,92,0);
signal scenario_full  : scenario_type := (0,0,243,31,243,30,165,31,8,31,79,31,119,31,250,31,250,30,250,29,250,28,221,31,229,31,229,30,101,31,82,31,23,31,128,31,107,31,10,31,133,31,182,31,182,30,86,31,57,31,57,30,32,31,1,31,1,30,130,31,130,30,130,29,252,31,192,31,161,31,134,31,117,31,202,31,83,31,48,31,48,30,172,31,70,31,31,31,23,31,113,31,121,31,121,30,127,31,177,31,11,31,14,31,87,31,134,31,60,31,161,31,161,30,169,31,28,31,89,31,145,31,203,31,75,31,183,31,183,30,226,31,221,31,39,31,39,30,55,31,133,31,217,31,251,31,225,31,117,31,189,31,167,31,241,31,179,31,35,31,168,31,66,31,17,31,167,31,1,31,163,31,163,30,1,31,36,31,82,31,253,31,81,31,162,31,43,31,43,30,43,29,68,31,44,31,44,30,160,31,229,31,110,31,117,31,117,30,203,31,170,31,170,30,23,31,141,31,141,30,14,31,210,31,202,31,113,31,133,31,133,30,233,31,186,31,186,30,186,29,186,28,186,27,186,26,143,31,84,31,228,31,165,31,84,31,134,31,134,30,79,31,247,31,27,31,158,31,121,31,121,30,121,29,236,31,225,31,225,30,106,31,156,31,86,31,86,30,254,31,79,31,38,31,121,31,121,30,191,31,20,31,24,31,249,31,36,31,200,31,200,30,184,31,109,31,73,31,228,31,140,31,14,31,90,31,90,30,141,31,245,31,5,31,124,31,58,31,132,31,113,31,52,31,85,31,38,31,71,31,44,31,33,31,122,31,251,31,41,31,191,31,145,31,7,31,113,31,113,30,170,31,119,31,64,31,18,31,143,31,143,30,143,29,143,28,207,31,140,31,8,31,8,30,196,31,147,31,147,30,202,31,202,30,180,31,101,31,119,31,119,30,184,31,192,31,188,31,69,31,129,31,104,31,116,31,116,30,116,29,139,31,55,31,55,30,193,31,92,31,92,30,92,29,160,31,168,31,226,31,123,31,51,31,26,31,64,31,131,31,131,30,74,31,255,31,9,31,56,31,64,31,254,31,254,30,239,31,86,31,124,31,113,31,146,31,142,31,133,31,133,30,203,31,188,31,232,31,59,31,167,31,167,30,167,29,187,31,187,30,11,31,193,31,13,31,195,31,195,30,195,29,195,28,195,27,195,26,195,25,195,24,57,31,57,30,177,31,174,31,246,31,246,30,8,31,223,31,99,31,19,31,30,31,30,30,30,29,18,31,18,30,20,31,110,31,125,31,54,31,237,31,178,31,24,31,129,31,70,31,10,31,65,31,151,31,56,31,185,31,175,31,202,31,138,31,165,31,40,31,100,31,106,31,122,31,248,31,116,31,118,31,201,31,151,31,188,31,250,31,250,30,250,29,250,28,127,31,127,30,99,31,202,31,202,30,88,31,124,31,23,31,57,31,206,31,7,31,161,31,141,31,11,31,11,30,228,31,196,31,231,31,238,31,34,31,117,31,141,31,141,30,167,31,155,31,155,30,182,31,105,31,231,31,231,30,202,31,208,31,180,31,208,31,240,31,252,31,169,31,169,30,98,31,98,30,98,29,13,31,13,30,13,29,135,31,133,31,86,31,89,31,89,30,89,29,44,31,247,31,154,31,36,31,57,31,57,30,81,31,120,31,255,31,181,31,175,31,175,30,27,31,75,31,10,31,155,31,168,31,32,31,81,31,252,31,124,31,124,30,169,31,248,31,88,31,198,31,198,30,38,31,157,31,131,31,146,31,70,31,70,30,136,31,136,30,103,31,111,31,169,31,169,30,161,31,153,31,120,31,197,31,44,31,44,30,44,29,61,31,218,31,41,31,46,31,46,30,108,31,28,31,28,30,121,31,184,31,184,30,174,31,229,31,229,30,154,31,70,31,80,31,144,31,180,31,50,31,203,31,203,30,186,31,88,31,147,31,147,30,64,31,76,31,64,31,156,31,234,31,234,30,32,31,8,31,8,30,237,31,237,30,86,31,128,31,59,31,59,30,170,31,196,31,196,30,75,31,30,31,192,31,223,31,61,31,61,30,228,31,91,31,91,30,56,31,137,31,226,31,202,31,161,31,157,31,157,30,169,31,187,31,98,31,98,30,173,31,99,31,127,31,127,30,182,31,182,30,15,31,252,31,107,31,107,30,231,31,16,31,16,30,16,29,20,31,186,31,186,30,63,31,250,31,197,31,137,31,204,31,195,31,135,31,213,31,247,31,142,31,32,31,155,31,72,31,172,31,95,31,170,31,170,30,204,31,14,31,213,31,213,30,149,31,153,31,111,31,248,31,206,31,103,31,197,31,244,31,244,30,218,31,119,31,202,31,202,30,202,29,224,31,46,31,198,31,198,30,242,31,222,31,180,31,180,30,83,31,140,31,140,31,140,30,218,31,226,31,177,31,67,31,96,31,96,30,52,31,52,30,175,31,44,31,242,31,242,30,242,29,83,31,17,31,49,31,222,31,87,31,98,31,234,31,38,31,178,31,230,31,215,31,175,31,221,31,181,31,252,31,252,30,252,29,84,31,8,31,240,31,60,31,64,31,64,30,156,31,156,30,95,31,203,31,94,31,116,31,167,31,187,31,187,30,220,31,220,30,220,29,46,31,50,31,118,31,118,30,118,29,196,31,108,31,145,31,35,31,10,31,192,31,192,30,24,31,45,31,12,31,12,30,155,31,185,31,85,31,166,31,166,30,166,29,252,31,66,31,57,31,57,30,80,31,196,31,31,31,31,30,56,31,56,30,169,31,169,30,99,31,12,31,175,31,50,31,50,30,38,31,253,31,119,31,47,31,7,31,7,30,7,29,200,31,245,31,175,31,175,30,10,31,250,31,250,30,151,31,92,31,177,31,222,31,196,31,206,31,36,31,36,30,36,29,75,31,75,30,75,29,10,31,74,31,58,31,145,31,165,31,165,30,203,31,117,31,45,31,45,30,131,31,140,31,140,31,140,30,111,31,15,31,94,31,46,31,59,31,22,31,238,31,2,31,181,31,56,31,155,31,255,31,115,31,250,31,164,31,177,31,213,31,91,31,200,31,127,31,127,30,127,29,140,31,157,31,102,31,102,30,48,31,199,31,208,31,145,31,149,31,197,31,17,31,69,31,202,31,73,31,68,31,194,31,240,31,1,31,100,31,215,31,215,30,215,29,28,31,127,31,127,30,213,31,241,31,98,31,131,31,161,31,51,31,22,31,22,30,22,29,80,31,20,31,19,31,126,31,92,31,92,30,80,31,67,31,67,30,28,31,219,31,219,30,17,31,73,31,73,30,246,31,250,31,194,31,254,31,99,31,24,31,141,31,249,31,249,30,146,31,146,30,146,29,187,31,187,30,187,29,187,28,24,31,173,31,80,31,90,31,90,30,66,31,145,31,210,31,76,31,249,31,45,31,130,31,75,31,236,31,9,31,9,30,185,31,131,31,198,31,182,31,182,30,185,31,86,31,179,31,244,31,16,31,103,31,231,31,176,31,61,31,251,31,251,30,251,29,28,31,28,30,140,31,26,31,172,31,24,31,247,31,117,31,117,30,80,31,80,30,132,31,16,31,232,31,246,31,203,31,203,30,203,29,72,31,30,31,230,31,117,31,231,31,253,31,218,31,218,30,16,31,146,31,146,30,108,31,244,31,159,31,46,31,125,31,173,31,96,31,96,30,96,29,16,31,34,31,70,31,205,31,109,31,105,31,189,31,70,31,123,31,123,30,191,31,181,31,175,31,179,31,179,30,179,29,57,31,211,31,1,31,59,31,51,31,51,30,106,31,206,31,54,31,62,31,34,31,243,31,85,31,85,30,85,29,207,31,61,31,85,31,85,30,96,31,11,31,8,31,100,31,237,31,237,30,227,31,227,30,130,31,156,31,156,30,16,31,16,30,73,31,225,31,40,31,40,30,116,31,116,30,178,31,242,31,137,31,136,31,26,31,116,31,28,31,28,30,150,31,177,31,227,31,227,30,84,31,6,31,243,31,115,31,92,31,11,31,173,31,211,31,92,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
