-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 983;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (85,0,199,0,255,0,27,0,101,0,95,0,148,0,118,0,158,0,88,0,206,0,102,0,0,0,237,0,65,0,0,0,181,0,91,0,13,0,20,0,0,0,13,0,0,0,17,0,0,0,54,0,0,0,249,0,188,0,88,0,72,0,23,0,232,0,0,0,0,0,11,0,180,0,127,0,42,0,216,0,90,0,232,0,175,0,63,0,157,0,0,0,0,0,179,0,72,0,185,0,63,0,238,0,0,0,35,0,117,0,74,0,0,0,159,0,84,0,59,0,142,0,0,0,38,0,208,0,255,0,51,0,227,0,93,0,55,0,117,0,206,0,97,0,80,0,212,0,121,0,0,0,0,0,247,0,0,0,0,0,0,0,189,0,36,0,36,0,175,0,215,0,122,0,207,0,244,0,237,0,163,0,153,0,176,0,102,0,93,0,251,0,83,0,0,0,136,0,110,0,214,0,0,0,106,0,0,0,4,0,216,0,0,0,113,0,43,0,0,0,103,0,118,0,12,0,199,0,197,0,195,0,186,0,225,0,114,0,235,0,241,0,41,0,0,0,113,0,126,0,8,0,196,0,0,0,0,0,218,0,0,0,49,0,0,0,171,0,220,0,11,0,0,0,144,0,0,0,0,0,0,0,164,0,147,0,177,0,85,0,0,0,222,0,0,0,57,0,106,0,0,0,0,0,26,0,143,0,246,0,0,0,216,0,149,0,164,0,0,0,213,0,0,0,189,0,0,0,127,0,111,0,223,0,199,0,239,0,135,0,189,0,170,0,237,0,102,0,147,0,48,0,137,0,198,0,224,0,48,0,246,0,52,0,207,0,188,0,80,0,0,0,0,0,58,0,0,0,0,0,129,0,49,0,42,0,26,0,206,0,238,0,166,0,85,0,236,0,172,0,166,0,0,0,14,0,170,0,172,0,228,0,0,0,46,0,145,0,151,0,0,0,64,0,51,0,0,0,144,0,0,0,254,0,0,0,213,0,0,0,187,0,0,0,0,0,137,0,225,0,179,0,70,0,77,0,112,0,60,0,0,0,5,0,117,0,0,0,0,0,60,0,43,0,0,0,23,0,101,0,0,0,10,0,242,0,0,0,174,0,227,0,80,0,90,0,110,0,34,0,208,0,20,0,72,0,250,0,0,0,37,0,237,0,61,0,163,0,22,0,26,0,0,0,0,0,115,0,170,0,125,0,0,0,169,0,203,0,34,0,239,0,185,0,0,0,138,0,13,0,0,0,12,0,237,0,73,0,121,0,0,0,235,0,87,0,199,0,222,0,120,0,198,0,212,0,95,0,152,0,175,0,131,0,204,0,0,0,142,0,26,0,217,0,0,0,0,0,238,0,0,0,0,0,246,0,193,0,0,0,126,0,57,0,0,0,248,0,0,0,93,0,173,0,182,0,65,0,4,0,41,0,186,0,92,0,151,0,46,0,125,0,113,0,168,0,170,0,222,0,0,0,190,0,0,0,166,0,174,0,0,0,138,0,193,0,141,0,0,0,220,0,0,0,162,0,168,0,180,0,217,0,0,0,45,0,155,0,0,0,105,0,174,0,38,0,219,0,215,0,23,0,0,0,0,0,176,0,0,0,48,0,233,0,20,0,155,0,177,0,227,0,3,0,128,0,87,0,133,0,234,0,130,0,0,0,15,0,0,0,95,0,254,0,226,0,0,0,253,0,200,0,47,0,68,0,244,0,6,0,54,0,0,0,191,0,0,0,177,0,100,0,3,0,215,0,229,0,0,0,78,0,0,0,109,0,189,0,251,0,240,0,187,0,158,0,43,0,24,0,0,0,125,0,109,0,33,0,83,0,134,0,0,0,255,0,0,0,138,0,107,0,213,0,5,0,75,0,197,0,189,0,148,0,92,0,27,0,113,0,16,0,196,0,28,0,21,0,86,0,132,0,204,0,228,0,69,0,19,0,151,0,0,0,157,0,254,0,200,0,18,0,10,0,65,0,132,0,0,0,0,0,230,0,0,0,0,0,204,0,0,0,103,0,220,0,232,0,233,0,31,0,61,0,199,0,0,0,143,0,195,0,0,0,242,0,43,0,179,0,195,0,168,0,40,0,219,0,83,0,114,0,62,0,220,0,98,0,0,0,93,0,250,0,204,0,68,0,48,0,75,0,26,0,145,0,247,0,0,0,85,0,0,0,81,0,57,0,89,0,156,0,255,0,33,0,168,0,0,0,142,0,174,0,74,0,71,0,170,0,150,0,28,0,204,0,0,0,0,0,235,0,112,0,0,0,33,0,254,0,98,0,126,0,0,0,0,0,58,0,80,0,13,0,0,0,223,0,9,0,152,0,0,0,114,0,130,0,0,0,0,0,187,0,0,0,34,0,136,0,218,0,228,0,171,0,102,0,232,0,0,0,188,0,144,0,98,0,140,0,235,0,17,0,16,0,126,0,119,0,80,0,72,0,175,0,108,0,0,0,41,0,101,0,172,0,28,0,18,0,223,0,0,0,206,0,192,0,7,0,0,0,63,0,253,0,221,0,132,0,0,0,198,0,168,0,246,0,225,0,86,0,15,0,161,0,40,0,127,0,31,0,120,0,117,0,0,0,227,0,99,0,200,0,46,0,133,0,63,0,10,0,104,0,36,0,240,0,124,0,58,0,152,0,248,0,103,0,207,0,0,0,128,0,81,0,138,0,160,0,85,0,45,0,0,0,74,0,161,0,0,0,79,0,105,0,0,0,159,0,113,0,0,0,152,0,0,0,102,0,148,0,215,0,127,0,232,0,81,0,142,0,248,0,137,0,114,0,231,0,153,0,0,0,8,0,50,0,221,0,66,0,108,0,248,0,71,0,0,0,176,0,243,0,88,0,0,0,189,0,69,0,13,0,9,0,72,0,254,0,74,0,25,0,66,0,78,0,141,0,252,0,160,0,164,0,54,0,3,0,0,0,62,0,0,0,40,0,92,0,0,0,212,0,4,0,232,0,0,0,217,0,76,0,171,0,73,0,0,0,42,0,40,0,101,0,117,0,0,0,188,0,165,0,226,0,155,0,49,0,244,0,155,0,190,0,7,0,0,0,96,0,234,0,142,0,141,0,244,0,0,0,0,0,110,0,128,0,168,0,154,0,0,0,69,0,0,0,69,0,0,0,0,0,0,0,197,0,0,0,160,0,0,0,97,0,0,0,117,0,106,0,22,0,182,0,188,0,0,0,255,0,210,0,58,0,192,0,0,0,142,0,50,0,0,0,173,0,0,0,126,0,174,0,171,0,0,0,0,0,24,0,37,0,154,0,0,0,0,0,64,0,205,0,35,0,203,0,0,0,9,0,160,0,116,0,129,0,175,0,233,0,152,0,0,0,147,0,55,0,241,0,99,0,78,0,224,0,106,0,113,0,239,0,115,0,84,0,87,0,162,0,59,0,0,0,63,0,83,0,110,0,162,0,226,0,94,0,0,0,35,0,128,0,231,0,0,0,197,0,201,0,3,0,73,0,0,0,208,0,0,0,0,0,225,0,33,0,238,0,0,0,79,0,19,0,177,0,174,0,51,0,53,0,189,0,178,0,219,0,122,0,255,0,79,0,0,0,180,0,0,0,45,0,152,0,188,0,160,0,200,0,0,0,0,0,172,0,27,0,0,0,60,0,39,0,194,0,34,0,212,0,209,0,0,0,190,0,158,0,0,0,38,0,197,0,199,0,245,0,239,0,172,0,166,0,188,0,0,0,179,0,81,0,85,0,244,0,0,0,140,0,64,0,67,0,114,0,208,0,183,0,221,0,83,0,0,0,160,0,193,0,189,0,114,0,149,0,19,0,22,0,184,0,253,0,0,0,142,0,43,0,60,0,202,0,94,0,56,0,0,0,28,0,76,0,115,0,0,0,37,0,232,0,235,0,179,0,169,0,162,0,61,0,69,0,192,0,208,0,133,0,0,0,72,0,223,0,0,0,167,0,180,0,234,0,30,0,0,0,51,0,238,0,178,0,223,0,0,0,43,0,0,0,196,0,25,0,179,0,145,0,145,0,120,0,0,0,39,0,134,0,235,0,0,0,0,0,212,0,31,0,243,0,0,0,238,0,56,0,78,0,49,0,140,0,228,0,68,0,147,0,252,0,101,0,0,0,164,0,0,0,0,0,176,0,0,0,143,0,206,0,164,0,0,0,215,0,121,0,34,0,152,0,0,0,115,0,0,0,86,0,6,0,24,0,174,0,118,0,5,0,72,0,178,0,200,0,0,0,151,0,70,0,0,0,0,0,0,0,0,0,0,0,50,0,235,0,0,0,170,0,218,0,0,0,202,0,115,0,38,0,0,0,0,0,117,0,178,0,176,0,110,0,221,0,114,0,19,0,151,0,143,0,157,0,190,0,53,0,0,0,23,0,0,0,0,0,148,0,218,0,243,0,0,0,0,0,56,0,237,0,160,0,0,0);
signal scenario_full  : scenario_type := (85,31,199,31,255,31,27,31,101,31,95,31,148,31,118,31,158,31,88,31,206,31,102,31,102,30,237,31,65,31,65,30,181,31,91,31,13,31,20,31,20,30,13,31,13,30,17,31,17,30,54,31,54,30,249,31,188,31,88,31,72,31,23,31,232,31,232,30,232,29,11,31,180,31,127,31,42,31,216,31,90,31,232,31,175,31,63,31,157,31,157,30,157,29,179,31,72,31,185,31,63,31,238,31,238,30,35,31,117,31,74,31,74,30,159,31,84,31,59,31,142,31,142,30,38,31,208,31,255,31,51,31,227,31,93,31,55,31,117,31,206,31,97,31,80,31,212,31,121,31,121,30,121,29,247,31,247,30,247,29,247,28,189,31,36,31,36,31,175,31,215,31,122,31,207,31,244,31,237,31,163,31,153,31,176,31,102,31,93,31,251,31,83,31,83,30,136,31,110,31,214,31,214,30,106,31,106,30,4,31,216,31,216,30,113,31,43,31,43,30,103,31,118,31,12,31,199,31,197,31,195,31,186,31,225,31,114,31,235,31,241,31,41,31,41,30,113,31,126,31,8,31,196,31,196,30,196,29,218,31,218,30,49,31,49,30,171,31,220,31,11,31,11,30,144,31,144,30,144,29,144,28,164,31,147,31,177,31,85,31,85,30,222,31,222,30,57,31,106,31,106,30,106,29,26,31,143,31,246,31,246,30,216,31,149,31,164,31,164,30,213,31,213,30,189,31,189,30,127,31,111,31,223,31,199,31,239,31,135,31,189,31,170,31,237,31,102,31,147,31,48,31,137,31,198,31,224,31,48,31,246,31,52,31,207,31,188,31,80,31,80,30,80,29,58,31,58,30,58,29,129,31,49,31,42,31,26,31,206,31,238,31,166,31,85,31,236,31,172,31,166,31,166,30,14,31,170,31,172,31,228,31,228,30,46,31,145,31,151,31,151,30,64,31,51,31,51,30,144,31,144,30,254,31,254,30,213,31,213,30,187,31,187,30,187,29,137,31,225,31,179,31,70,31,77,31,112,31,60,31,60,30,5,31,117,31,117,30,117,29,60,31,43,31,43,30,23,31,101,31,101,30,10,31,242,31,242,30,174,31,227,31,80,31,90,31,110,31,34,31,208,31,20,31,72,31,250,31,250,30,37,31,237,31,61,31,163,31,22,31,26,31,26,30,26,29,115,31,170,31,125,31,125,30,169,31,203,31,34,31,239,31,185,31,185,30,138,31,13,31,13,30,12,31,237,31,73,31,121,31,121,30,235,31,87,31,199,31,222,31,120,31,198,31,212,31,95,31,152,31,175,31,131,31,204,31,204,30,142,31,26,31,217,31,217,30,217,29,238,31,238,30,238,29,246,31,193,31,193,30,126,31,57,31,57,30,248,31,248,30,93,31,173,31,182,31,65,31,4,31,41,31,186,31,92,31,151,31,46,31,125,31,113,31,168,31,170,31,222,31,222,30,190,31,190,30,166,31,174,31,174,30,138,31,193,31,141,31,141,30,220,31,220,30,162,31,168,31,180,31,217,31,217,30,45,31,155,31,155,30,105,31,174,31,38,31,219,31,215,31,23,31,23,30,23,29,176,31,176,30,48,31,233,31,20,31,155,31,177,31,227,31,3,31,128,31,87,31,133,31,234,31,130,31,130,30,15,31,15,30,95,31,254,31,226,31,226,30,253,31,200,31,47,31,68,31,244,31,6,31,54,31,54,30,191,31,191,30,177,31,100,31,3,31,215,31,229,31,229,30,78,31,78,30,109,31,189,31,251,31,240,31,187,31,158,31,43,31,24,31,24,30,125,31,109,31,33,31,83,31,134,31,134,30,255,31,255,30,138,31,107,31,213,31,5,31,75,31,197,31,189,31,148,31,92,31,27,31,113,31,16,31,196,31,28,31,21,31,86,31,132,31,204,31,228,31,69,31,19,31,151,31,151,30,157,31,254,31,200,31,18,31,10,31,65,31,132,31,132,30,132,29,230,31,230,30,230,29,204,31,204,30,103,31,220,31,232,31,233,31,31,31,61,31,199,31,199,30,143,31,195,31,195,30,242,31,43,31,179,31,195,31,168,31,40,31,219,31,83,31,114,31,62,31,220,31,98,31,98,30,93,31,250,31,204,31,68,31,48,31,75,31,26,31,145,31,247,31,247,30,85,31,85,30,81,31,57,31,89,31,156,31,255,31,33,31,168,31,168,30,142,31,174,31,74,31,71,31,170,31,150,31,28,31,204,31,204,30,204,29,235,31,112,31,112,30,33,31,254,31,98,31,126,31,126,30,126,29,58,31,80,31,13,31,13,30,223,31,9,31,152,31,152,30,114,31,130,31,130,30,130,29,187,31,187,30,34,31,136,31,218,31,228,31,171,31,102,31,232,31,232,30,188,31,144,31,98,31,140,31,235,31,17,31,16,31,126,31,119,31,80,31,72,31,175,31,108,31,108,30,41,31,101,31,172,31,28,31,18,31,223,31,223,30,206,31,192,31,7,31,7,30,63,31,253,31,221,31,132,31,132,30,198,31,168,31,246,31,225,31,86,31,15,31,161,31,40,31,127,31,31,31,120,31,117,31,117,30,227,31,99,31,200,31,46,31,133,31,63,31,10,31,104,31,36,31,240,31,124,31,58,31,152,31,248,31,103,31,207,31,207,30,128,31,81,31,138,31,160,31,85,31,45,31,45,30,74,31,161,31,161,30,79,31,105,31,105,30,159,31,113,31,113,30,152,31,152,30,102,31,148,31,215,31,127,31,232,31,81,31,142,31,248,31,137,31,114,31,231,31,153,31,153,30,8,31,50,31,221,31,66,31,108,31,248,31,71,31,71,30,176,31,243,31,88,31,88,30,189,31,69,31,13,31,9,31,72,31,254,31,74,31,25,31,66,31,78,31,141,31,252,31,160,31,164,31,54,31,3,31,3,30,62,31,62,30,40,31,92,31,92,30,212,31,4,31,232,31,232,30,217,31,76,31,171,31,73,31,73,30,42,31,40,31,101,31,117,31,117,30,188,31,165,31,226,31,155,31,49,31,244,31,155,31,190,31,7,31,7,30,96,31,234,31,142,31,141,31,244,31,244,30,244,29,110,31,128,31,168,31,154,31,154,30,69,31,69,30,69,31,69,30,69,29,69,28,197,31,197,30,160,31,160,30,97,31,97,30,117,31,106,31,22,31,182,31,188,31,188,30,255,31,210,31,58,31,192,31,192,30,142,31,50,31,50,30,173,31,173,30,126,31,174,31,171,31,171,30,171,29,24,31,37,31,154,31,154,30,154,29,64,31,205,31,35,31,203,31,203,30,9,31,160,31,116,31,129,31,175,31,233,31,152,31,152,30,147,31,55,31,241,31,99,31,78,31,224,31,106,31,113,31,239,31,115,31,84,31,87,31,162,31,59,31,59,30,63,31,83,31,110,31,162,31,226,31,94,31,94,30,35,31,128,31,231,31,231,30,197,31,201,31,3,31,73,31,73,30,208,31,208,30,208,29,225,31,33,31,238,31,238,30,79,31,19,31,177,31,174,31,51,31,53,31,189,31,178,31,219,31,122,31,255,31,79,31,79,30,180,31,180,30,45,31,152,31,188,31,160,31,200,31,200,30,200,29,172,31,27,31,27,30,60,31,39,31,194,31,34,31,212,31,209,31,209,30,190,31,158,31,158,30,38,31,197,31,199,31,245,31,239,31,172,31,166,31,188,31,188,30,179,31,81,31,85,31,244,31,244,30,140,31,64,31,67,31,114,31,208,31,183,31,221,31,83,31,83,30,160,31,193,31,189,31,114,31,149,31,19,31,22,31,184,31,253,31,253,30,142,31,43,31,60,31,202,31,94,31,56,31,56,30,28,31,76,31,115,31,115,30,37,31,232,31,235,31,179,31,169,31,162,31,61,31,69,31,192,31,208,31,133,31,133,30,72,31,223,31,223,30,167,31,180,31,234,31,30,31,30,30,51,31,238,31,178,31,223,31,223,30,43,31,43,30,196,31,25,31,179,31,145,31,145,31,120,31,120,30,39,31,134,31,235,31,235,30,235,29,212,31,31,31,243,31,243,30,238,31,56,31,78,31,49,31,140,31,228,31,68,31,147,31,252,31,101,31,101,30,164,31,164,30,164,29,176,31,176,30,143,31,206,31,164,31,164,30,215,31,121,31,34,31,152,31,152,30,115,31,115,30,86,31,6,31,24,31,174,31,118,31,5,31,72,31,178,31,200,31,200,30,151,31,70,31,70,30,70,29,70,28,70,27,70,26,50,31,235,31,235,30,170,31,218,31,218,30,202,31,115,31,38,31,38,30,38,29,117,31,178,31,176,31,110,31,221,31,114,31,19,31,151,31,143,31,157,31,190,31,53,31,53,30,23,31,23,30,23,29,148,31,218,31,243,31,243,30,243,29,56,31,237,31,160,31,160,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
