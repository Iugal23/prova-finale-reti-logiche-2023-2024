-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 444;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (177,0,46,0,69,0,222,0,159,0,35,0,89,0,121,0,233,0,190,0,209,0,0,0,0,0,55,0,248,0,87,0,200,0,149,0,215,0,107,0,241,0,228,0,123,0,57,0,4,0,101,0,0,0,102,0,72,0,113,0,60,0,108,0,150,0,54,0,121,0,177,0,212,0,242,0,130,0,34,0,165,0,219,0,198,0,8,0,0,0,47,0,0,0,5,0,237,0,234,0,0,0,25,0,3,0,0,0,39,0,146,0,0,0,0,0,0,0,47,0,99,0,93,0,178,0,0,0,194,0,96,0,0,0,84,0,252,0,93,0,0,0,119,0,246,0,203,0,136,0,12,0,248,0,113,0,188,0,37,0,96,0,151,0,213,0,0,0,179,0,10,0,163,0,177,0,10,0,71,0,64,0,176,0,0,0,10,0,31,0,83,0,95,0,52,0,110,0,69,0,178,0,124,0,246,0,225,0,0,0,0,0,20,0,1,0,244,0,0,0,208,0,102,0,39,0,149,0,84,0,80,0,40,0,102,0,109,0,37,0,18,0,186,0,0,0,0,0,0,0,93,0,0,0,125,0,104,0,76,0,82,0,21,0,0,0,151,0,0,0,4,0,144,0,129,0,88,0,219,0,244,0,141,0,0,0,125,0,0,0,61,0,207,0,40,0,156,0,170,0,40,0,236,0,191,0,17,0,148,0,172,0,141,0,0,0,250,0,128,0,242,0,154,0,43,0,248,0,149,0,255,0,203,0,242,0,170,0,55,0,132,0,135,0,8,0,229,0,211,0,0,0,3,0,13,0,166,0,0,0,64,0,155,0,92,0,91,0,210,0,48,0,141,0,11,0,0,0,0,0,215,0,75,0,198,0,24,0,109,0,0,0,71,0,0,0,18,0,17,0,226,0,232,0,0,0,225,0,171,0,229,0,74,0,106,0,199,0,192,0,0,0,207,0,148,0,147,0,237,0,0,0,245,0,85,0,245,0,0,0,200,0,0,0,0,0,233,0,111,0,58,0,121,0,196,0,63,0,0,0,0,0,0,0,143,0,115,0,17,0,66,0,30,0,36,0,250,0,183,0,58,0,183,0,195,0,236,0,38,0,0,0,227,0,138,0,178,0,252,0,33,0,167,0,0,0,184,0,158,0,176,0,41,0,0,0,105,0,214,0,218,0,0,0,252,0,9,0,223,0,0,0,255,0,247,0,45,0,0,0,52,0,74,0,55,0,0,0,121,0,119,0,0,0,43,0,0,0,0,0,0,0,0,0,0,0,22,0,30,0,0,0,0,0,166,0,96,0,108,0,255,0,137,0,173,0,248,0,90,0,0,0,0,0,32,0,4,0,0,0,0,0,78,0,90,0,108,0,160,0,53,0,0,0,0,0,133,0,37,0,61,0,0,0,82,0,237,0,0,0,4,0,117,0,0,0,107,0,11,0,69,0,94,0,113,0,21,0,98,0,0,0,242,0,127,0,74,0,66,0,209,0,0,0,189,0,0,0,18,0,174,0,189,0,215,0,166,0,4,0,0,0,155,0,220,0,147,0,133,0,39,0,170,0,154,0,231,0,221,0,243,0,42,0,248,0,226,0,34,0,144,0,233,0,158,0,5,0,40,0,0,0,242,0,0,0,70,0,0,0,73,0,138,0,183,0,0,0,173,0,0,0,90,0,0,0,40,0,104,0,0,0,6,0,227,0,214,0,95,0,0,0,95,0,192,0,0,0,0,0,0,0,229,0,0,0,213,0,72,0,0,0,82,0,34,0,0,0,162,0,0,0,211,0,81,0,202,0,179,0,68,0,81,0,171,0,29,0,240,0,249,0,0,0,0,0,163,0,46,0,40,0,24,0,199,0,0,0,27,0,29,0,28,0,189,0,46,0,244,0,0,0,65,0,220,0,249,0,239,0,187,0,48,0,47,0,206,0,0,0,118,0,158,0,96,0,135,0,70,0,246,0,136,0,128,0,246,0,40,0,0,0,115,0,73,0,104,0);
signal scenario_full  : scenario_type := (177,31,46,31,69,31,222,31,159,31,35,31,89,31,121,31,233,31,190,31,209,31,209,30,209,29,55,31,248,31,87,31,200,31,149,31,215,31,107,31,241,31,228,31,123,31,57,31,4,31,101,31,101,30,102,31,72,31,113,31,60,31,108,31,150,31,54,31,121,31,177,31,212,31,242,31,130,31,34,31,165,31,219,31,198,31,8,31,8,30,47,31,47,30,5,31,237,31,234,31,234,30,25,31,3,31,3,30,39,31,146,31,146,30,146,29,146,28,47,31,99,31,93,31,178,31,178,30,194,31,96,31,96,30,84,31,252,31,93,31,93,30,119,31,246,31,203,31,136,31,12,31,248,31,113,31,188,31,37,31,96,31,151,31,213,31,213,30,179,31,10,31,163,31,177,31,10,31,71,31,64,31,176,31,176,30,10,31,31,31,83,31,95,31,52,31,110,31,69,31,178,31,124,31,246,31,225,31,225,30,225,29,20,31,1,31,244,31,244,30,208,31,102,31,39,31,149,31,84,31,80,31,40,31,102,31,109,31,37,31,18,31,186,31,186,30,186,29,186,28,93,31,93,30,125,31,104,31,76,31,82,31,21,31,21,30,151,31,151,30,4,31,144,31,129,31,88,31,219,31,244,31,141,31,141,30,125,31,125,30,61,31,207,31,40,31,156,31,170,31,40,31,236,31,191,31,17,31,148,31,172,31,141,31,141,30,250,31,128,31,242,31,154,31,43,31,248,31,149,31,255,31,203,31,242,31,170,31,55,31,132,31,135,31,8,31,229,31,211,31,211,30,3,31,13,31,166,31,166,30,64,31,155,31,92,31,91,31,210,31,48,31,141,31,11,31,11,30,11,29,215,31,75,31,198,31,24,31,109,31,109,30,71,31,71,30,18,31,17,31,226,31,232,31,232,30,225,31,171,31,229,31,74,31,106,31,199,31,192,31,192,30,207,31,148,31,147,31,237,31,237,30,245,31,85,31,245,31,245,30,200,31,200,30,200,29,233,31,111,31,58,31,121,31,196,31,63,31,63,30,63,29,63,28,143,31,115,31,17,31,66,31,30,31,36,31,250,31,183,31,58,31,183,31,195,31,236,31,38,31,38,30,227,31,138,31,178,31,252,31,33,31,167,31,167,30,184,31,158,31,176,31,41,31,41,30,105,31,214,31,218,31,218,30,252,31,9,31,223,31,223,30,255,31,247,31,45,31,45,30,52,31,74,31,55,31,55,30,121,31,119,31,119,30,43,31,43,30,43,29,43,28,43,27,43,26,22,31,30,31,30,30,30,29,166,31,96,31,108,31,255,31,137,31,173,31,248,31,90,31,90,30,90,29,32,31,4,31,4,30,4,29,78,31,90,31,108,31,160,31,53,31,53,30,53,29,133,31,37,31,61,31,61,30,82,31,237,31,237,30,4,31,117,31,117,30,107,31,11,31,69,31,94,31,113,31,21,31,98,31,98,30,242,31,127,31,74,31,66,31,209,31,209,30,189,31,189,30,18,31,174,31,189,31,215,31,166,31,4,31,4,30,155,31,220,31,147,31,133,31,39,31,170,31,154,31,231,31,221,31,243,31,42,31,248,31,226,31,34,31,144,31,233,31,158,31,5,31,40,31,40,30,242,31,242,30,70,31,70,30,73,31,138,31,183,31,183,30,173,31,173,30,90,31,90,30,40,31,104,31,104,30,6,31,227,31,214,31,95,31,95,30,95,31,192,31,192,30,192,29,192,28,229,31,229,30,213,31,72,31,72,30,82,31,34,31,34,30,162,31,162,30,211,31,81,31,202,31,179,31,68,31,81,31,171,31,29,31,240,31,249,31,249,30,249,29,163,31,46,31,40,31,24,31,199,31,199,30,27,31,29,31,28,31,189,31,46,31,244,31,244,30,65,31,220,31,249,31,239,31,187,31,48,31,47,31,206,31,206,30,118,31,158,31,96,31,135,31,70,31,246,31,136,31,128,31,246,31,40,31,40,30,115,31,73,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
