-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_644 is
end project_tb_644;

architecture project_tb_arch_644 of project_tb_644 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 944;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,0,0,0,0,10,0,116,0,242,0,208,0,134,0,131,0,0,0,214,0,129,0,83,0,247,0,233,0,130,0,216,0,166,0,0,0,0,0,0,0,73,0,200,0,0,0,183,0,0,0,0,0,0,0,170,0,217,0,22,0,6,0,134,0,30,0,165,0,0,0,246,0,23,0,182,0,0,0,212,0,0,0,221,0,248,0,201,0,149,0,202,0,0,0,183,0,33,0,114,0,0,0,54,0,0,0,174,0,58,0,0,0,138,0,162,0,195,0,175,0,121,0,0,0,181,0,30,0,127,0,32,0,0,0,126,0,40,0,76,0,0,0,75,0,163,0,237,0,0,0,62,0,38,0,162,0,94,0,96,0,203,0,0,0,123,0,201,0,68,0,7,0,8,0,165,0,19,0,114,0,0,0,90,0,68,0,138,0,152,0,208,0,236,0,0,0,0,0,249,0,0,0,108,0,33,0,229,0,57,0,136,0,170,0,12,0,73,0,235,0,142,0,129,0,173,0,0,0,0,0,103,0,25,0,62,0,0,0,16,0,33,0,202,0,57,0,0,0,40,0,189,0,42,0,78,0,192,0,79,0,0,0,160,0,194,0,90,0,152,0,99,0,46,0,104,0,0,0,200,0,152,0,0,0,54,0,0,0,0,0,0,0,82,0,0,0,75,0,0,0,8,0,142,0,10,0,86,0,91,0,160,0,241,0,222,0,0,0,90,0,245,0,0,0,198,0,89,0,192,0,67,0,0,0,241,0,20,0,120,0,54,0,3,0,204,0,15,0,201,0,150,0,52,0,0,0,0,0,196,0,109,0,238,0,0,0,64,0,214,0,105,0,57,0,226,0,154,0,166,0,185,0,39,0,16,0,0,0,216,0,185,0,197,0,34,0,100,0,72,0,0,0,196,0,177,0,136,0,31,0,12,0,208,0,171,0,145,0,228,0,0,0,214,0,0,0,61,0,190,0,144,0,182,0,193,0,1,0,171,0,65,0,0,0,239,0,74,0,126,0,250,0,44,0,59,0,74,0,161,0,0,0,211,0,21,0,0,0,163,0,0,0,44,0,216,0,119,0,156,0,0,0,37,0,60,0,116,0,186,0,0,0,0,0,57,0,173,0,93,0,24,0,218,0,0,0,120,0,0,0,0,0,128,0,0,0,241,0,59,0,0,0,233,0,165,0,16,0,0,0,196,0,61,0,0,0,226,0,253,0,89,0,156,0,15,0,0,0,100,0,164,0,186,0,0,0,118,0,118,0,114,0,157,0,21,0,244,0,0,0,81,0,31,0,196,0,213,0,0,0,158,0,0,0,176,0,0,0,206,0,18,0,0,0,0,0,24,0,174,0,210,0,132,0,0,0,0,0,35,0,144,0,0,0,232,0,0,0,82,0,55,0,119,0,161,0,254,0,69,0,184,0,36,0,114,0,88,0,55,0,227,0,117,0,0,0,112,0,160,0,124,0,0,0,230,0,0,0,0,0,0,0,76,0,106,0,0,0,0,0,40,0,200,0,0,0,0,0,124,0,64,0,62,0,0,0,79,0,0,0,245,0,252,0,156,0,39,0,70,0,228,0,219,0,242,0,189,0,242,0,47,0,122,0,183,0,0,0,57,0,99,0,194,0,23,0,87,0,79,0,72,0,79,0,16,0,255,0,74,0,213,0,0,0,46,0,111,0,0,0,52,0,0,0,253,0,213,0,124,0,0,0,194,0,195,0,2,0,131,0,100,0,134,0,66,0,68,0,68,0,0,0,117,0,239,0,144,0,165,0,120,0,0,0,76,0,141,0,139,0,66,0,236,0,100,0,0,0,82,0,145,0,0,0,0,0,0,0,35,0,205,0,186,0,115,0,0,0,147,0,138,0,229,0,0,0,191,0,48,0,121,0,138,0,32,0,0,0,48,0,160,0,141,0,148,0,0,0,0,0,182,0,43,0,131,0,129,0,163,0,62,0,0,0,50,0,140,0,238,0,240,0,121,0,228,0,218,0,130,0,192,0,0,0,236,0,0,0,0,0,70,0,185,0,0,0,34,0,0,0,129,0,141,0,0,0,164,0,0,0,38,0,240,0,0,0,0,0,26,0,160,0,4,0,115,0,88,0,240,0,0,0,196,0,52,0,95,0,36,0,250,0,49,0,81,0,13,0,250,0,91,0,81,0,0,0,0,0,0,0,157,0,225,0,51,0,0,0,122,0,10,0,200,0,24,0,0,0,251,0,68,0,64,0,75,0,72,0,0,0,0,0,198,0,179,0,28,0,0,0,43,0,123,0,0,0,0,0,38,0,172,0,69,0,18,0,99,0,32,0,63,0,139,0,95,0,177,0,79,0,166,0,202,0,120,0,121,0,72,0,158,0,90,0,70,0,0,0,218,0,0,0,0,0,235,0,132,0,26,0,0,0,142,0,80,0,68,0,163,0,82,0,131,0,43,0,238,0,0,0,103,0,117,0,69,0,87,0,150,0,0,0,26,0,131,0,200,0,0,0,196,0,0,0,165,0,209,0,48,0,0,0,127,0,104,0,0,0,17,0,218,0,243,0,0,0,183,0,7,0,73,0,175,0,152,0,139,0,238,0,9,0,230,0,158,0,123,0,80,0,0,0,0,0,113,0,190,0,3,0,184,0,159,0,27,0,84,0,52,0,246,0,125,0,0,0,136,0,234,0,166,0,229,0,61,0,90,0,0,0,215,0,99,0,0,0,247,0,0,0,9,0,136,0,88,0,196,0,0,0,184,0,0,0,155,0,177,0,196,0,123,0,1,0,208,0,129,0,50,0,176,0,139,0,95,0,245,0,0,0,0,0,32,0,147,0,79,0,218,0,220,0,106,0,0,0,0,0,65,0,48,0,0,0,51,0,0,0,203,0,64,0,240,0,183,0,139,0,128,0,255,0,0,0,156,0,0,0,0,0,144,0,0,0,122,0,127,0,157,0,0,0,0,0,0,0,0,0,244,0,23,0,0,0,38,0,43,0,216,0,58,0,219,0,179,0,102,0,85,0,64,0,173,0,0,0,0,0,55,0,24,0,12,0,73,0,0,0,106,0,214,0,0,0,103,0,0,0,93,0,42,0,143,0,85,0,102,0,132,0,105,0,244,0,57,0,30,0,173,0,0,0,192,0,180,0,7,0,191,0,145,0,98,0,180,0,14,0,19,0,35,0,69,0,207,0,240,0,34,0,0,0,127,0,85,0,200,0,178,0,2,0,122,0,128,0,61,0,143,0,32,0,167,0,157,0,231,0,136,0,2,0,9,0,73,0,11,0,0,0,174,0,214,0,97,0,88,0,62,0,177,0,0,0,159,0,237,0,17,0,108,0,174,0,235,0,0,0,255,0,240,0,57,0,105,0,0,0,244,0,73,0,138,0,0,0,53,0,0,0,165,0,201,0,222,0,0,0,1,0,24,0,0,0,159,0,143,0,80,0,204,0,65,0,132,0,148,0,108,0,0,0,69,0,36,0,4,0,205,0,167,0,70,0,0,0,0,0,0,0,142,0,108,0,216,0,31,0,106,0,0,0,172,0,215,0,193,0,251,0,234,0,131,0,88,0,102,0,248,0,28,0,105,0,152,0,0,0,135,0,36,0,175,0,213,0,225,0,122,0,195,0,241,0,242,0,223,0,0,0,5,0,0,0,52,0,77,0,0,0,85,0,242,0,0,0,0,0,135,0,146,0,19,0,142,0,140,0,119,0,0,0,0,0,252,0,0,0,150,0,189,0,135,0,50,0,248,0,251,0,43,0,91,0,111,0,113,0,50,0,56,0,250,0,225,0,0,0,34,0,108,0,12,0,222,0,230,0,228,0,180,0,22,0,36,0,124,0,0,0,14,0,189,0,78,0,0,0,90,0,0,0,0,0,205,0,247,0,173,0,66,0,0,0,8,0,190,0,254,0,221,0,0,0,0,0,195,0,95,0,158,0,138,0,196,0,39,0,28,0,252,0,45,0,76,0,146,0,4,0,49,0,20,0,106,0,218,0,154,0,211,0,146,0,228,0,2,0,82,0,156,0,0,0,82,0,1,0,50,0,52,0,161,0,42,0,104,0,207,0,77,0,153,0,246,0,25,0,126,0,0,0,66,0,145,0,49,0,190,0,160,0,238,0,94,0,122,0,74,0,66,0,128,0,6,0,60,0,244,0,190,0,240,0,62,0,20,0,58,0,242,0,159,0,230,0,159,0,163,0,192,0,163,0,40,0,180,0,0,0,0,0,1,0,40,0);
signal scenario_full  : scenario_type := (135,31,135,30,135,29,10,31,116,31,242,31,208,31,134,31,131,31,131,30,214,31,129,31,83,31,247,31,233,31,130,31,216,31,166,31,166,30,166,29,166,28,73,31,200,31,200,30,183,31,183,30,183,29,183,28,170,31,217,31,22,31,6,31,134,31,30,31,165,31,165,30,246,31,23,31,182,31,182,30,212,31,212,30,221,31,248,31,201,31,149,31,202,31,202,30,183,31,33,31,114,31,114,30,54,31,54,30,174,31,58,31,58,30,138,31,162,31,195,31,175,31,121,31,121,30,181,31,30,31,127,31,32,31,32,30,126,31,40,31,76,31,76,30,75,31,163,31,237,31,237,30,62,31,38,31,162,31,94,31,96,31,203,31,203,30,123,31,201,31,68,31,7,31,8,31,165,31,19,31,114,31,114,30,90,31,68,31,138,31,152,31,208,31,236,31,236,30,236,29,249,31,249,30,108,31,33,31,229,31,57,31,136,31,170,31,12,31,73,31,235,31,142,31,129,31,173,31,173,30,173,29,103,31,25,31,62,31,62,30,16,31,33,31,202,31,57,31,57,30,40,31,189,31,42,31,78,31,192,31,79,31,79,30,160,31,194,31,90,31,152,31,99,31,46,31,104,31,104,30,200,31,152,31,152,30,54,31,54,30,54,29,54,28,82,31,82,30,75,31,75,30,8,31,142,31,10,31,86,31,91,31,160,31,241,31,222,31,222,30,90,31,245,31,245,30,198,31,89,31,192,31,67,31,67,30,241,31,20,31,120,31,54,31,3,31,204,31,15,31,201,31,150,31,52,31,52,30,52,29,196,31,109,31,238,31,238,30,64,31,214,31,105,31,57,31,226,31,154,31,166,31,185,31,39,31,16,31,16,30,216,31,185,31,197,31,34,31,100,31,72,31,72,30,196,31,177,31,136,31,31,31,12,31,208,31,171,31,145,31,228,31,228,30,214,31,214,30,61,31,190,31,144,31,182,31,193,31,1,31,171,31,65,31,65,30,239,31,74,31,126,31,250,31,44,31,59,31,74,31,161,31,161,30,211,31,21,31,21,30,163,31,163,30,44,31,216,31,119,31,156,31,156,30,37,31,60,31,116,31,186,31,186,30,186,29,57,31,173,31,93,31,24,31,218,31,218,30,120,31,120,30,120,29,128,31,128,30,241,31,59,31,59,30,233,31,165,31,16,31,16,30,196,31,61,31,61,30,226,31,253,31,89,31,156,31,15,31,15,30,100,31,164,31,186,31,186,30,118,31,118,31,114,31,157,31,21,31,244,31,244,30,81,31,31,31,196,31,213,31,213,30,158,31,158,30,176,31,176,30,206,31,18,31,18,30,18,29,24,31,174,31,210,31,132,31,132,30,132,29,35,31,144,31,144,30,232,31,232,30,82,31,55,31,119,31,161,31,254,31,69,31,184,31,36,31,114,31,88,31,55,31,227,31,117,31,117,30,112,31,160,31,124,31,124,30,230,31,230,30,230,29,230,28,76,31,106,31,106,30,106,29,40,31,200,31,200,30,200,29,124,31,64,31,62,31,62,30,79,31,79,30,245,31,252,31,156,31,39,31,70,31,228,31,219,31,242,31,189,31,242,31,47,31,122,31,183,31,183,30,57,31,99,31,194,31,23,31,87,31,79,31,72,31,79,31,16,31,255,31,74,31,213,31,213,30,46,31,111,31,111,30,52,31,52,30,253,31,213,31,124,31,124,30,194,31,195,31,2,31,131,31,100,31,134,31,66,31,68,31,68,31,68,30,117,31,239,31,144,31,165,31,120,31,120,30,76,31,141,31,139,31,66,31,236,31,100,31,100,30,82,31,145,31,145,30,145,29,145,28,35,31,205,31,186,31,115,31,115,30,147,31,138,31,229,31,229,30,191,31,48,31,121,31,138,31,32,31,32,30,48,31,160,31,141,31,148,31,148,30,148,29,182,31,43,31,131,31,129,31,163,31,62,31,62,30,50,31,140,31,238,31,240,31,121,31,228,31,218,31,130,31,192,31,192,30,236,31,236,30,236,29,70,31,185,31,185,30,34,31,34,30,129,31,141,31,141,30,164,31,164,30,38,31,240,31,240,30,240,29,26,31,160,31,4,31,115,31,88,31,240,31,240,30,196,31,52,31,95,31,36,31,250,31,49,31,81,31,13,31,250,31,91,31,81,31,81,30,81,29,81,28,157,31,225,31,51,31,51,30,122,31,10,31,200,31,24,31,24,30,251,31,68,31,64,31,75,31,72,31,72,30,72,29,198,31,179,31,28,31,28,30,43,31,123,31,123,30,123,29,38,31,172,31,69,31,18,31,99,31,32,31,63,31,139,31,95,31,177,31,79,31,166,31,202,31,120,31,121,31,72,31,158,31,90,31,70,31,70,30,218,31,218,30,218,29,235,31,132,31,26,31,26,30,142,31,80,31,68,31,163,31,82,31,131,31,43,31,238,31,238,30,103,31,117,31,69,31,87,31,150,31,150,30,26,31,131,31,200,31,200,30,196,31,196,30,165,31,209,31,48,31,48,30,127,31,104,31,104,30,17,31,218,31,243,31,243,30,183,31,7,31,73,31,175,31,152,31,139,31,238,31,9,31,230,31,158,31,123,31,80,31,80,30,80,29,113,31,190,31,3,31,184,31,159,31,27,31,84,31,52,31,246,31,125,31,125,30,136,31,234,31,166,31,229,31,61,31,90,31,90,30,215,31,99,31,99,30,247,31,247,30,9,31,136,31,88,31,196,31,196,30,184,31,184,30,155,31,177,31,196,31,123,31,1,31,208,31,129,31,50,31,176,31,139,31,95,31,245,31,245,30,245,29,32,31,147,31,79,31,218,31,220,31,106,31,106,30,106,29,65,31,48,31,48,30,51,31,51,30,203,31,64,31,240,31,183,31,139,31,128,31,255,31,255,30,156,31,156,30,156,29,144,31,144,30,122,31,127,31,157,31,157,30,157,29,157,28,157,27,244,31,23,31,23,30,38,31,43,31,216,31,58,31,219,31,179,31,102,31,85,31,64,31,173,31,173,30,173,29,55,31,24,31,12,31,73,31,73,30,106,31,214,31,214,30,103,31,103,30,93,31,42,31,143,31,85,31,102,31,132,31,105,31,244,31,57,31,30,31,173,31,173,30,192,31,180,31,7,31,191,31,145,31,98,31,180,31,14,31,19,31,35,31,69,31,207,31,240,31,34,31,34,30,127,31,85,31,200,31,178,31,2,31,122,31,128,31,61,31,143,31,32,31,167,31,157,31,231,31,136,31,2,31,9,31,73,31,11,31,11,30,174,31,214,31,97,31,88,31,62,31,177,31,177,30,159,31,237,31,17,31,108,31,174,31,235,31,235,30,255,31,240,31,57,31,105,31,105,30,244,31,73,31,138,31,138,30,53,31,53,30,165,31,201,31,222,31,222,30,1,31,24,31,24,30,159,31,143,31,80,31,204,31,65,31,132,31,148,31,108,31,108,30,69,31,36,31,4,31,205,31,167,31,70,31,70,30,70,29,70,28,142,31,108,31,216,31,31,31,106,31,106,30,172,31,215,31,193,31,251,31,234,31,131,31,88,31,102,31,248,31,28,31,105,31,152,31,152,30,135,31,36,31,175,31,213,31,225,31,122,31,195,31,241,31,242,31,223,31,223,30,5,31,5,30,52,31,77,31,77,30,85,31,242,31,242,30,242,29,135,31,146,31,19,31,142,31,140,31,119,31,119,30,119,29,252,31,252,30,150,31,189,31,135,31,50,31,248,31,251,31,43,31,91,31,111,31,113,31,50,31,56,31,250,31,225,31,225,30,34,31,108,31,12,31,222,31,230,31,228,31,180,31,22,31,36,31,124,31,124,30,14,31,189,31,78,31,78,30,90,31,90,30,90,29,205,31,247,31,173,31,66,31,66,30,8,31,190,31,254,31,221,31,221,30,221,29,195,31,95,31,158,31,138,31,196,31,39,31,28,31,252,31,45,31,76,31,146,31,4,31,49,31,20,31,106,31,218,31,154,31,211,31,146,31,228,31,2,31,82,31,156,31,156,30,82,31,1,31,50,31,52,31,161,31,42,31,104,31,207,31,77,31,153,31,246,31,25,31,126,31,126,30,66,31,145,31,49,31,190,31,160,31,238,31,94,31,122,31,74,31,66,31,128,31,6,31,60,31,244,31,190,31,240,31,62,31,20,31,58,31,242,31,159,31,230,31,159,31,163,31,192,31,163,31,40,31,180,31,180,30,180,29,1,31,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
