-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 890;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (81,0,0,0,242,0,57,0,0,0,81,0,229,0,45,0,254,0,53,0,227,0,246,0,203,0,75,0,0,0,47,0,143,0,103,0,191,0,152,0,179,0,73,0,45,0,0,0,0,0,10,0,54,0,149,0,45,0,0,0,93,0,51,0,32,0,8,0,103,0,49,0,167,0,247,0,92,0,144,0,0,0,159,0,231,0,6,0,43,0,35,0,34,0,66,0,253,0,0,0,0,0,49,0,134,0,0,0,185,0,232,0,146,0,0,0,232,0,187,0,136,0,36,0,0,0,0,0,69,0,36,0,0,0,8,0,154,0,0,0,0,0,96,0,238,0,0,0,12,0,0,0,0,0,62,0,95,0,147,0,213,0,92,0,158,0,11,0,0,0,43,0,17,0,0,0,0,0,0,0,238,0,226,0,0,0,37,0,21,0,154,0,248,0,147,0,0,0,166,0,0,0,116,0,4,0,247,0,0,0,24,0,0,0,51,0,240,0,158,0,124,0,141,0,165,0,0,0,194,0,228,0,145,0,188,0,120,0,21,0,156,0,246,0,64,0,63,0,41,0,0,0,73,0,133,0,156,0,63,0,208,0,172,0,0,0,46,0,158,0,207,0,14,0,233,0,218,0,160,0,226,0,198,0,6,0,143,0,85,0,197,0,210,0,0,0,159,0,8,0,0,0,254,0,245,0,228,0,33,0,131,0,111,0,0,0,253,0,159,0,227,0,8,0,187,0,68,0,94,0,213,0,0,0,129,0,114,0,179,0,152,0,0,0,0,0,0,0,218,0,0,0,207,0,0,0,93,0,219,0,142,0,14,0,221,0,194,0,231,0,31,0,63,0,206,0,190,0,46,0,0,0,0,0,192,0,0,0,56,0,0,0,179,0,163,0,199,0,151,0,0,0,59,0,39,0,118,0,49,0,0,0,194,0,0,0,0,0,191,0,86,0,19,0,97,0,0,0,67,0,125,0,38,0,110,0,153,0,145,0,136,0,0,0,123,0,220,0,252,0,53,0,92,0,215,0,225,0,254,0,178,0,197,0,143,0,109,0,143,0,229,0,167,0,195,0,216,0,88,0,241,0,44,0,16,0,96,0,236,0,206,0,151,0,57,0,219,0,41,0,108,0,216,0,223,0,0,0,53,0,253,0,0,0,112,0,0,0,155,0,77,0,17,0,8,0,209,0,0,0,48,0,176,0,237,0,65,0,98,0,0,0,136,0,81,0,0,0,217,0,60,0,214,0,94,0,0,0,163,0,0,0,84,0,239,0,211,0,171,0,6,0,69,0,98,0,226,0,124,0,140,0,237,0,29,0,224,0,145,0,247,0,61,0,45,0,211,0,176,0,12,0,83,0,156,0,192,0,0,0,42,0,0,0,133,0,73,0,0,0,255,0,214,0,0,0,0,0,157,0,141,0,141,0,0,0,250,0,0,0,77,0,168,0,0,0,0,0,103,0,105,0,63,0,186,0,24,0,216,0,223,0,67,0,79,0,113,0,67,0,194,0,160,0,41,0,195,0,22,0,84,0,0,0,0,0,193,0,3,0,88,0,13,0,0,0,197,0,7,0,204,0,138,0,70,0,53,0,92,0,100,0,220,0,124,0,227,0,77,0,185,0,166,0,0,0,113,0,58,0,183,0,167,0,0,0,188,0,199,0,0,0,29,0,162,0,150,0,142,0,0,0,35,0,23,0,110,0,59,0,190,0,22,0,34,0,63,0,26,0,21,0,246,0,26,0,174,0,109,0,105,0,0,0,106,0,0,0,204,0,71,0,60,0,0,0,239,0,225,0,84,0,169,0,107,0,179,0,81,0,120,0,0,0,0,0,89,0,217,0,125,0,192,0,195,0,185,0,159,0,181,0,97,0,0,0,72,0,65,0,57,0,0,0,198,0,47,0,0,0,235,0,194,0,198,0,142,0,75,0,77,0,81,0,64,0,52,0,0,0,161,0,0,0,91,0,169,0,219,0,248,0,159,0,93,0,168,0,78,0,72,0,212,0,151,0,61,0,29,0,0,0,0,0,41,0,168,0,196,0,45,0,180,0,108,0,253,0,128,0,78,0,85,0,63,0,126,0,149,0,234,0,60,0,66,0,58,0,0,0,28,0,250,0,182,0,64,0,192,0,10,0,238,0,0,0,135,0,64,0,0,0,216,0,129,0,163,0,70,0,25,0,200,0,74,0,106,0,0,0,178,0,224,0,18,0,94,0,0,0,83,0,78,0,0,0,64,0,217,0,184,0,253,0,182,0,165,0,52,0,127,0,121,0,126,0,124,0,181,0,218,0,82,0,27,0,114,0,228,0,68,0,77,0,0,0,60,0,0,0,0,0,0,0,243,0,0,0,77,0,71,0,2,0,111,0,239,0,0,0,178,0,89,0,145,0,39,0,127,0,247,0,150,0,0,0,211,0,28,0,145,0,228,0,80,0,22,0,247,0,94,0,229,0,0,0,28,0,174,0,0,0,0,0,0,0,120,0,0,0,47,0,205,0,37,0,0,0,4,0,129,0,0,0,119,0,0,0,254,0,0,0,24,0,134,0,180,0,188,0,85,0,199,0,196,0,0,0,173,0,117,0,134,0,5,0,0,0,0,0,97,0,191,0,143,0,108,0,247,0,223,0,0,0,144,0,244,0,11,0,0,0,100,0,69,0,205,0,187,0,0,0,44,0,174,0,69,0,227,0,66,0,0,0,0,0,95,0,71,0,46,0,0,0,9,0,110,0,236,0,82,0,125,0,0,0,112,0,0,0,0,0,16,0,191,0,30,0,0,0,163,0,109,0,62,0,161,0,51,0,119,0,169,0,115,0,198,0,25,0,210,0,24,0,0,0,239,0,224,0,59,0,121,0,200,0,0,0,54,0,67,0,54,0,119,0,29,0,172,0,208,0,181,0,160,0,108,0,154,0,0,0,80,0,0,0,0,0,0,0,158,0,0,0,143,0,195,0,206,0,0,0,0,0,193,0,58,0,156,0,154,0,202,0,0,0,53,0,39,0,48,0,23,0,0,0,21,0,0,0,116,0,237,0,213,0,75,0,9,0,93,0,163,0,18,0,148,0,0,0,148,0,58,0,0,0,174,0,0,0,0,0,63,0,252,0,231,0,76,0,140,0,199,0,137,0,203,0,144,0,165,0,0,0,78,0,62,0,220,0,187,0,188,0,0,0,103,0,0,0,0,0,29,0,0,0,122,0,161,0,26,0,0,0,153,0,25,0,91,0,0,0,83,0,86,0,146,0,50,0,233,0,101,0,5,0,208,0,208,0,83,0,201,0,103,0,28,0,187,0,110,0,0,0,234,0,191,0,210,0,0,0,203,0,107,0,0,0,0,0,205,0,252,0,225,0,124,0,65,0,36,0,75,0,193,0,240,0,3,0,29,0,173,0,90,0,0,0,63,0,44,0,0,0,127,0,48,0,117,0,0,0,158,0,27,0,0,0,0,0,14,0,141,0,237,0,78,0,176,0,231,0,89,0,28,0,114,0,71,0,232,0,15,0,179,0,185,0,202,0,187,0,135,0,0,0,5,0,162,0,242,0,102,0,0,0,249,0,155,0,140,0,79,0,87,0,144,0,207,0,45,0,151,0,27,0,130,0,44,0,33,0,168,0,0,0,193,0,248,0,108,0,107,0,58,0,135,0,0,0,106,0,36,0,0,0,210,0,65,0,0,0,30,0,208,0,20,0,247,0,0,0,230,0,0,0,205,0,139,0,41,0,42,0,157,0,0,0,0,0,101,0,0,0,70,0,135,0,187,0,70,0,106,0,0,0,114,0,100,0,66,0,229,0,141,0,219,0,190,0,0,0,0,0,239,0,0,0,100,0,92,0,200,0,145,0,218,0,0,0,162,0,0,0,158,0,101,0,0,0,141,0,240,0,16,0,232,0,233,0,232,0,117,0,181,0,141,0,62,0,61,0,68,0,233,0,114,0,0,0,157,0,237,0,0,0,0,0,106,0,239,0,0,0,28,0,46,0,226,0);
signal scenario_full  : scenario_type := (81,31,81,30,242,31,57,31,57,30,81,31,229,31,45,31,254,31,53,31,227,31,246,31,203,31,75,31,75,30,47,31,143,31,103,31,191,31,152,31,179,31,73,31,45,31,45,30,45,29,10,31,54,31,149,31,45,31,45,30,93,31,51,31,32,31,8,31,103,31,49,31,167,31,247,31,92,31,144,31,144,30,159,31,231,31,6,31,43,31,35,31,34,31,66,31,253,31,253,30,253,29,49,31,134,31,134,30,185,31,232,31,146,31,146,30,232,31,187,31,136,31,36,31,36,30,36,29,69,31,36,31,36,30,8,31,154,31,154,30,154,29,96,31,238,31,238,30,12,31,12,30,12,29,62,31,95,31,147,31,213,31,92,31,158,31,11,31,11,30,43,31,17,31,17,30,17,29,17,28,238,31,226,31,226,30,37,31,21,31,154,31,248,31,147,31,147,30,166,31,166,30,116,31,4,31,247,31,247,30,24,31,24,30,51,31,240,31,158,31,124,31,141,31,165,31,165,30,194,31,228,31,145,31,188,31,120,31,21,31,156,31,246,31,64,31,63,31,41,31,41,30,73,31,133,31,156,31,63,31,208,31,172,31,172,30,46,31,158,31,207,31,14,31,233,31,218,31,160,31,226,31,198,31,6,31,143,31,85,31,197,31,210,31,210,30,159,31,8,31,8,30,254,31,245,31,228,31,33,31,131,31,111,31,111,30,253,31,159,31,227,31,8,31,187,31,68,31,94,31,213,31,213,30,129,31,114,31,179,31,152,31,152,30,152,29,152,28,218,31,218,30,207,31,207,30,93,31,219,31,142,31,14,31,221,31,194,31,231,31,31,31,63,31,206,31,190,31,46,31,46,30,46,29,192,31,192,30,56,31,56,30,179,31,163,31,199,31,151,31,151,30,59,31,39,31,118,31,49,31,49,30,194,31,194,30,194,29,191,31,86,31,19,31,97,31,97,30,67,31,125,31,38,31,110,31,153,31,145,31,136,31,136,30,123,31,220,31,252,31,53,31,92,31,215,31,225,31,254,31,178,31,197,31,143,31,109,31,143,31,229,31,167,31,195,31,216,31,88,31,241,31,44,31,16,31,96,31,236,31,206,31,151,31,57,31,219,31,41,31,108,31,216,31,223,31,223,30,53,31,253,31,253,30,112,31,112,30,155,31,77,31,17,31,8,31,209,31,209,30,48,31,176,31,237,31,65,31,98,31,98,30,136,31,81,31,81,30,217,31,60,31,214,31,94,31,94,30,163,31,163,30,84,31,239,31,211,31,171,31,6,31,69,31,98,31,226,31,124,31,140,31,237,31,29,31,224,31,145,31,247,31,61,31,45,31,211,31,176,31,12,31,83,31,156,31,192,31,192,30,42,31,42,30,133,31,73,31,73,30,255,31,214,31,214,30,214,29,157,31,141,31,141,31,141,30,250,31,250,30,77,31,168,31,168,30,168,29,103,31,105,31,63,31,186,31,24,31,216,31,223,31,67,31,79,31,113,31,67,31,194,31,160,31,41,31,195,31,22,31,84,31,84,30,84,29,193,31,3,31,88,31,13,31,13,30,197,31,7,31,204,31,138,31,70,31,53,31,92,31,100,31,220,31,124,31,227,31,77,31,185,31,166,31,166,30,113,31,58,31,183,31,167,31,167,30,188,31,199,31,199,30,29,31,162,31,150,31,142,31,142,30,35,31,23,31,110,31,59,31,190,31,22,31,34,31,63,31,26,31,21,31,246,31,26,31,174,31,109,31,105,31,105,30,106,31,106,30,204,31,71,31,60,31,60,30,239,31,225,31,84,31,169,31,107,31,179,31,81,31,120,31,120,30,120,29,89,31,217,31,125,31,192,31,195,31,185,31,159,31,181,31,97,31,97,30,72,31,65,31,57,31,57,30,198,31,47,31,47,30,235,31,194,31,198,31,142,31,75,31,77,31,81,31,64,31,52,31,52,30,161,31,161,30,91,31,169,31,219,31,248,31,159,31,93,31,168,31,78,31,72,31,212,31,151,31,61,31,29,31,29,30,29,29,41,31,168,31,196,31,45,31,180,31,108,31,253,31,128,31,78,31,85,31,63,31,126,31,149,31,234,31,60,31,66,31,58,31,58,30,28,31,250,31,182,31,64,31,192,31,10,31,238,31,238,30,135,31,64,31,64,30,216,31,129,31,163,31,70,31,25,31,200,31,74,31,106,31,106,30,178,31,224,31,18,31,94,31,94,30,83,31,78,31,78,30,64,31,217,31,184,31,253,31,182,31,165,31,52,31,127,31,121,31,126,31,124,31,181,31,218,31,82,31,27,31,114,31,228,31,68,31,77,31,77,30,60,31,60,30,60,29,60,28,243,31,243,30,77,31,71,31,2,31,111,31,239,31,239,30,178,31,89,31,145,31,39,31,127,31,247,31,150,31,150,30,211,31,28,31,145,31,228,31,80,31,22,31,247,31,94,31,229,31,229,30,28,31,174,31,174,30,174,29,174,28,120,31,120,30,47,31,205,31,37,31,37,30,4,31,129,31,129,30,119,31,119,30,254,31,254,30,24,31,134,31,180,31,188,31,85,31,199,31,196,31,196,30,173,31,117,31,134,31,5,31,5,30,5,29,97,31,191,31,143,31,108,31,247,31,223,31,223,30,144,31,244,31,11,31,11,30,100,31,69,31,205,31,187,31,187,30,44,31,174,31,69,31,227,31,66,31,66,30,66,29,95,31,71,31,46,31,46,30,9,31,110,31,236,31,82,31,125,31,125,30,112,31,112,30,112,29,16,31,191,31,30,31,30,30,163,31,109,31,62,31,161,31,51,31,119,31,169,31,115,31,198,31,25,31,210,31,24,31,24,30,239,31,224,31,59,31,121,31,200,31,200,30,54,31,67,31,54,31,119,31,29,31,172,31,208,31,181,31,160,31,108,31,154,31,154,30,80,31,80,30,80,29,80,28,158,31,158,30,143,31,195,31,206,31,206,30,206,29,193,31,58,31,156,31,154,31,202,31,202,30,53,31,39,31,48,31,23,31,23,30,21,31,21,30,116,31,237,31,213,31,75,31,9,31,93,31,163,31,18,31,148,31,148,30,148,31,58,31,58,30,174,31,174,30,174,29,63,31,252,31,231,31,76,31,140,31,199,31,137,31,203,31,144,31,165,31,165,30,78,31,62,31,220,31,187,31,188,31,188,30,103,31,103,30,103,29,29,31,29,30,122,31,161,31,26,31,26,30,153,31,25,31,91,31,91,30,83,31,86,31,146,31,50,31,233,31,101,31,5,31,208,31,208,31,83,31,201,31,103,31,28,31,187,31,110,31,110,30,234,31,191,31,210,31,210,30,203,31,107,31,107,30,107,29,205,31,252,31,225,31,124,31,65,31,36,31,75,31,193,31,240,31,3,31,29,31,173,31,90,31,90,30,63,31,44,31,44,30,127,31,48,31,117,31,117,30,158,31,27,31,27,30,27,29,14,31,141,31,237,31,78,31,176,31,231,31,89,31,28,31,114,31,71,31,232,31,15,31,179,31,185,31,202,31,187,31,135,31,135,30,5,31,162,31,242,31,102,31,102,30,249,31,155,31,140,31,79,31,87,31,144,31,207,31,45,31,151,31,27,31,130,31,44,31,33,31,168,31,168,30,193,31,248,31,108,31,107,31,58,31,135,31,135,30,106,31,36,31,36,30,210,31,65,31,65,30,30,31,208,31,20,31,247,31,247,30,230,31,230,30,205,31,139,31,41,31,42,31,157,31,157,30,157,29,101,31,101,30,70,31,135,31,187,31,70,31,106,31,106,30,114,31,100,31,66,31,229,31,141,31,219,31,190,31,190,30,190,29,239,31,239,30,100,31,92,31,200,31,145,31,218,31,218,30,162,31,162,30,158,31,101,31,101,30,141,31,240,31,16,31,232,31,233,31,232,31,117,31,181,31,141,31,62,31,61,31,68,31,233,31,114,31,114,30,157,31,237,31,237,30,237,29,106,31,239,31,239,30,28,31,46,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
