-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 811;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (240,0,126,0,93,0,0,0,182,0,28,0,0,0,0,0,104,0,0,0,192,0,115,0,236,0,187,0,78,0,0,0,172,0,141,0,162,0,11,0,246,0,0,0,217,0,141,0,100,0,203,0,88,0,180,0,187,0,5,0,0,0,54,0,205,0,216,0,129,0,221,0,189,0,174,0,138,0,60,0,180,0,0,0,189,0,0,0,176,0,0,0,145,0,180,0,0,0,15,0,133,0,58,0,43,0,193,0,0,0,1,0,0,0,120,0,161,0,138,0,233,0,38,0,155,0,80,0,198,0,71,0,7,0,0,0,4,0,42,0,198,0,177,0,223,0,0,0,220,0,254,0,39,0,213,0,150,0,0,0,8,0,166,0,125,0,219,0,121,0,34,0,240,0,0,0,176,0,156,0,80,0,0,0,0,0,250,0,36,0,195,0,124,0,0,0,55,0,192,0,173,0,36,0,162,0,0,0,167,0,82,0,128,0,83,0,239,0,254,0,164,0,156,0,180,0,199,0,93,0,107,0,190,0,91,0,139,0,0,0,146,0,209,0,212,0,0,0,21,0,249,0,241,0,90,0,68,0,149,0,0,0,125,0,136,0,43,0,223,0,67,0,48,0,0,0,2,0,0,0,30,0,42,0,207,0,160,0,232,0,255,0,77,0,129,0,0,0,74,0,247,0,0,0,108,0,202,0,53,0,68,0,234,0,0,0,190,0,199,0,198,0,0,0,71,0,7,0,0,0,24,0,211,0,0,0,239,0,67,0,205,0,88,0,102,0,153,0,81,0,0,0,0,0,119,0,57,0,226,0,201,0,132,0,119,0,63,0,214,0,0,0,45,0,28,0,0,0,142,0,134,0,185,0,245,0,157,0,94,0,50,0,225,0,239,0,232,0,5,0,116,0,181,0,221,0,17,0,0,0,4,0,243,0,45,0,0,0,141,0,146,0,119,0,133,0,171,0,187,0,150,0,24,0,180,0,0,0,146,0,77,0,57,0,42,0,113,0,84,0,0,0,158,0,0,0,219,0,186,0,74,0,0,0,206,0,231,0,201,0,12,0,0,0,48,0,34,0,83,0,2,0,232,0,0,0,168,0,217,0,246,0,105,0,91,0,204,0,99,0,9,0,135,0,0,0,240,0,84,0,81,0,59,0,202,0,93,0,44,0,214,0,0,0,171,0,57,0,0,0,230,0,132,0,24,0,254,0,219,0,89,0,233,0,0,0,226,0,222,0,217,0,0,0,250,0,30,0,45,0,58,0,92,0,140,0,11,0,143,0,0,0,116,0,208,0,156,0,139,0,65,0,248,0,178,0,21,0,61,0,0,0,28,0,228,0,59,0,205,0,147,0,0,0,131,0,185,0,243,0,15,0,0,0,30,0,0,0,0,0,80,0,107,0,0,0,112,0,0,0,0,0,0,0,191,0,82,0,86,0,166,0,0,0,39,0,115,0,224,0,77,0,32,0,28,0,196,0,241,0,163,0,83,0,108,0,128,0,180,0,112,0,219,0,0,0,50,0,22,0,161,0,6,0,183,0,163,0,116,0,243,0,224,0,160,0,194,0,88,0,0,0,103,0,230,0,223,0,223,0,70,0,179,0,142,0,54,0,44,0,133,0,129,0,180,0,95,0,158,0,129,0,149,0,44,0,156,0,188,0,96,0,0,0,237,0,230,0,198,0,0,0,216,0,248,0,208,0,156,0,126,0,0,0,195,0,26,0,88,0,33,0,0,0,0,0,149,0,50,0,0,0,0,0,0,0,91,0,231,0,0,0,9,0,0,0,222,0,152,0,33,0,17,0,0,0,61,0,201,0,40,0,161,0,0,0,129,0,3,0,95,0,209,0,0,0,180,0,230,0,0,0,0,0,0,0,9,0,138,0,0,0,0,0,0,0,87,0,10,0,100,0,0,0,53,0,88,0,77,0,0,0,212,0,0,0,68,0,118,0,0,0,175,0,184,0,0,0,184,0,201,0,145,0,143,0,164,0,0,0,0,0,242,0,228,0,0,0,29,0,233,0,145,0,227,0,19,0,164,0,215,0,44,0,21,0,0,0,117,0,0,0,221,0,48,0,64,0,4,0,176,0,0,0,68,0,254,0,3,0,35,0,0,0,216,0,3,0,9,0,132,0,1,0,111,0,130,0,186,0,155,0,234,0,233,0,52,0,0,0,0,0,29,0,157,0,144,0,232,0,146,0,212,0,248,0,0,0,253,0,178,0,21,0,0,0,2,0,64,0,243,0,236,0,51,0,157,0,13,0,67,0,106,0,31,0,235,0,106,0,70,0,22,0,169,0,12,0,151,0,161,0,0,0,48,0,132,0,0,0,153,0,163,0,18,0,116,0,71,0,0,0,0,0,48,0,224,0,0,0,238,0,0,0,46,0,0,0,190,0,217,0,62,0,153,0,0,0,139,0,164,0,72,0,44,0,34,0,84,0,116,0,179,0,38,0,34,0,0,0,0,0,197,0,114,0,0,0,91,0,0,0,212,0,44,0,65,0,53,0,174,0,117,0,169,0,81,0,56,0,90,0,2,0,248,0,234,0,137,0,56,0,157,0,148,0,117,0,155,0,212,0,54,0,0,0,0,0,157,0,0,0,0,0,185,0,130,0,0,0,42,0,145,0,0,0,175,0,0,0,129,0,61,0,179,0,120,0,252,0,195,0,113,0,153,0,189,0,0,0,52,0,0,0,233,0,0,0,247,0,33,0,65,0,160,0,234,0,162,0,81,0,0,0,0,0,159,0,254,0,15,0,24,0,167,0,0,0,196,0,163,0,142,0,150,0,0,0,15,0,44,0,46,0,1,0,242,0,138,0,15,0,79,0,192,0,141,0,201,0,81,0,81,0,87,0,40,0,0,0,181,0,0,0,52,0,107,0,11,0,194,0,97,0,191,0,45,0,124,0,188,0,46,0,111,0,142,0,241,0,123,0,0,0,43,0,0,0,192,0,0,0,46,0,232,0,72,0,164,0,47,0,142,0,63,0,60,0,212,0,179,0,106,0,73,0,8,0,0,0,116,0,219,0,88,0,151,0,231,0,155,0,174,0,153,0,79,0,0,0,136,0,0,0,230,0,221,0,124,0,253,0,125,0,0,0,156,0,88,0,210,0,0,0,53,0,0,0,125,0,38,0,50,0,22,0,142,0,109,0,87,0,223,0,229,0,0,0,51,0,77,0,53,0,55,0,75,0,30,0,83,0,0,0,133,0,0,0,243,0,173,0,106,0,240,0,228,0,74,0,0,0,147,0,121,0,100,0,105,0,52,0,255,0,60,0,99,0,12,0,242,0,127,0,122,0,239,0,79,0,92,0,201,0,157,0,0,0,28,0,218,0,188,0,50,0,0,0,0,0,0,0,140,0,175,0,203,0,162,0,0,0,63,0,161,0,155,0,216,0,0,0,172,0,128,0,30,0,0,0,49,0,11,0,100,0,77,0,72,0,0,0,221,0,178,0,33,0,113,0,185,0,191,0,2,0,115,0,0,0,9,0,248,0,0,0,8,0,94,0,186,0,169,0,0,0,70,0,106,0,0,0,178,0,166,0,156,0,216,0,105,0,21,0,160,0,0,0,96,0,177,0,109,0,64,0,252,0,9,0,0,0,36,0,0,0,21,0,0,0,200,0);
signal scenario_full  : scenario_type := (240,31,126,31,93,31,93,30,182,31,28,31,28,30,28,29,104,31,104,30,192,31,115,31,236,31,187,31,78,31,78,30,172,31,141,31,162,31,11,31,246,31,246,30,217,31,141,31,100,31,203,31,88,31,180,31,187,31,5,31,5,30,54,31,205,31,216,31,129,31,221,31,189,31,174,31,138,31,60,31,180,31,180,30,189,31,189,30,176,31,176,30,145,31,180,31,180,30,15,31,133,31,58,31,43,31,193,31,193,30,1,31,1,30,120,31,161,31,138,31,233,31,38,31,155,31,80,31,198,31,71,31,7,31,7,30,4,31,42,31,198,31,177,31,223,31,223,30,220,31,254,31,39,31,213,31,150,31,150,30,8,31,166,31,125,31,219,31,121,31,34,31,240,31,240,30,176,31,156,31,80,31,80,30,80,29,250,31,36,31,195,31,124,31,124,30,55,31,192,31,173,31,36,31,162,31,162,30,167,31,82,31,128,31,83,31,239,31,254,31,164,31,156,31,180,31,199,31,93,31,107,31,190,31,91,31,139,31,139,30,146,31,209,31,212,31,212,30,21,31,249,31,241,31,90,31,68,31,149,31,149,30,125,31,136,31,43,31,223,31,67,31,48,31,48,30,2,31,2,30,30,31,42,31,207,31,160,31,232,31,255,31,77,31,129,31,129,30,74,31,247,31,247,30,108,31,202,31,53,31,68,31,234,31,234,30,190,31,199,31,198,31,198,30,71,31,7,31,7,30,24,31,211,31,211,30,239,31,67,31,205,31,88,31,102,31,153,31,81,31,81,30,81,29,119,31,57,31,226,31,201,31,132,31,119,31,63,31,214,31,214,30,45,31,28,31,28,30,142,31,134,31,185,31,245,31,157,31,94,31,50,31,225,31,239,31,232,31,5,31,116,31,181,31,221,31,17,31,17,30,4,31,243,31,45,31,45,30,141,31,146,31,119,31,133,31,171,31,187,31,150,31,24,31,180,31,180,30,146,31,77,31,57,31,42,31,113,31,84,31,84,30,158,31,158,30,219,31,186,31,74,31,74,30,206,31,231,31,201,31,12,31,12,30,48,31,34,31,83,31,2,31,232,31,232,30,168,31,217,31,246,31,105,31,91,31,204,31,99,31,9,31,135,31,135,30,240,31,84,31,81,31,59,31,202,31,93,31,44,31,214,31,214,30,171,31,57,31,57,30,230,31,132,31,24,31,254,31,219,31,89,31,233,31,233,30,226,31,222,31,217,31,217,30,250,31,30,31,45,31,58,31,92,31,140,31,11,31,143,31,143,30,116,31,208,31,156,31,139,31,65,31,248,31,178,31,21,31,61,31,61,30,28,31,228,31,59,31,205,31,147,31,147,30,131,31,185,31,243,31,15,31,15,30,30,31,30,30,30,29,80,31,107,31,107,30,112,31,112,30,112,29,112,28,191,31,82,31,86,31,166,31,166,30,39,31,115,31,224,31,77,31,32,31,28,31,196,31,241,31,163,31,83,31,108,31,128,31,180,31,112,31,219,31,219,30,50,31,22,31,161,31,6,31,183,31,163,31,116,31,243,31,224,31,160,31,194,31,88,31,88,30,103,31,230,31,223,31,223,31,70,31,179,31,142,31,54,31,44,31,133,31,129,31,180,31,95,31,158,31,129,31,149,31,44,31,156,31,188,31,96,31,96,30,237,31,230,31,198,31,198,30,216,31,248,31,208,31,156,31,126,31,126,30,195,31,26,31,88,31,33,31,33,30,33,29,149,31,50,31,50,30,50,29,50,28,91,31,231,31,231,30,9,31,9,30,222,31,152,31,33,31,17,31,17,30,61,31,201,31,40,31,161,31,161,30,129,31,3,31,95,31,209,31,209,30,180,31,230,31,230,30,230,29,230,28,9,31,138,31,138,30,138,29,138,28,87,31,10,31,100,31,100,30,53,31,88,31,77,31,77,30,212,31,212,30,68,31,118,31,118,30,175,31,184,31,184,30,184,31,201,31,145,31,143,31,164,31,164,30,164,29,242,31,228,31,228,30,29,31,233,31,145,31,227,31,19,31,164,31,215,31,44,31,21,31,21,30,117,31,117,30,221,31,48,31,64,31,4,31,176,31,176,30,68,31,254,31,3,31,35,31,35,30,216,31,3,31,9,31,132,31,1,31,111,31,130,31,186,31,155,31,234,31,233,31,52,31,52,30,52,29,29,31,157,31,144,31,232,31,146,31,212,31,248,31,248,30,253,31,178,31,21,31,21,30,2,31,64,31,243,31,236,31,51,31,157,31,13,31,67,31,106,31,31,31,235,31,106,31,70,31,22,31,169,31,12,31,151,31,161,31,161,30,48,31,132,31,132,30,153,31,163,31,18,31,116,31,71,31,71,30,71,29,48,31,224,31,224,30,238,31,238,30,46,31,46,30,190,31,217,31,62,31,153,31,153,30,139,31,164,31,72,31,44,31,34,31,84,31,116,31,179,31,38,31,34,31,34,30,34,29,197,31,114,31,114,30,91,31,91,30,212,31,44,31,65,31,53,31,174,31,117,31,169,31,81,31,56,31,90,31,2,31,248,31,234,31,137,31,56,31,157,31,148,31,117,31,155,31,212,31,54,31,54,30,54,29,157,31,157,30,157,29,185,31,130,31,130,30,42,31,145,31,145,30,175,31,175,30,129,31,61,31,179,31,120,31,252,31,195,31,113,31,153,31,189,31,189,30,52,31,52,30,233,31,233,30,247,31,33,31,65,31,160,31,234,31,162,31,81,31,81,30,81,29,159,31,254,31,15,31,24,31,167,31,167,30,196,31,163,31,142,31,150,31,150,30,15,31,44,31,46,31,1,31,242,31,138,31,15,31,79,31,192,31,141,31,201,31,81,31,81,31,87,31,40,31,40,30,181,31,181,30,52,31,107,31,11,31,194,31,97,31,191,31,45,31,124,31,188,31,46,31,111,31,142,31,241,31,123,31,123,30,43,31,43,30,192,31,192,30,46,31,232,31,72,31,164,31,47,31,142,31,63,31,60,31,212,31,179,31,106,31,73,31,8,31,8,30,116,31,219,31,88,31,151,31,231,31,155,31,174,31,153,31,79,31,79,30,136,31,136,30,230,31,221,31,124,31,253,31,125,31,125,30,156,31,88,31,210,31,210,30,53,31,53,30,125,31,38,31,50,31,22,31,142,31,109,31,87,31,223,31,229,31,229,30,51,31,77,31,53,31,55,31,75,31,30,31,83,31,83,30,133,31,133,30,243,31,173,31,106,31,240,31,228,31,74,31,74,30,147,31,121,31,100,31,105,31,52,31,255,31,60,31,99,31,12,31,242,31,127,31,122,31,239,31,79,31,92,31,201,31,157,31,157,30,28,31,218,31,188,31,50,31,50,30,50,29,50,28,140,31,175,31,203,31,162,31,162,30,63,31,161,31,155,31,216,31,216,30,172,31,128,31,30,31,30,30,49,31,11,31,100,31,77,31,72,31,72,30,221,31,178,31,33,31,113,31,185,31,191,31,2,31,115,31,115,30,9,31,248,31,248,30,8,31,94,31,186,31,169,31,169,30,70,31,106,31,106,30,178,31,166,31,156,31,216,31,105,31,21,31,160,31,160,30,96,31,177,31,109,31,64,31,252,31,9,31,9,30,36,31,36,30,21,31,21,30,200,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
