-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_389 is
end project_tb_389;

architecture project_tb_arch_389 of project_tb_389 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 953;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (81,0,82,0,43,0,214,0,21,0,51,0,0,0,218,0,5,0,7,0,0,0,176,0,179,0,87,0,0,0,0,0,0,0,70,0,230,0,187,0,186,0,26,0,95,0,28,0,161,0,41,0,156,0,0,0,175,0,0,0,52,0,82,0,65,0,206,0,231,0,0,0,245,0,245,0,97,0,0,0,92,0,0,0,28,0,172,0,96,0,113,0,25,0,95,0,168,0,26,0,223,0,97,0,240,0,0,0,126,0,157,0,0,0,30,0,194,0,148,0,174,0,25,0,212,0,0,0,181,0,0,0,0,0,66,0,149,0,162,0,0,0,0,0,85,0,34,0,0,0,59,0,215,0,247,0,95,0,0,0,23,0,217,0,0,0,0,0,62,0,19,0,48,0,243,0,191,0,165,0,0,0,41,0,0,0,210,0,199,0,54,0,197,0,0,0,72,0,173,0,70,0,175,0,117,0,0,0,23,0,179,0,73,0,21,0,204,0,18,0,0,0,27,0,183,0,119,0,230,0,56,0,38,0,70,0,119,0,196,0,0,0,204,0,99,0,208,0,224,0,225,0,46,0,0,0,241,0,0,0,53,0,231,0,0,0,100,0,177,0,55,0,86,0,168,0,128,0,9,0,212,0,118,0,253,0,132,0,241,0,248,0,39,0,0,0,188,0,86,0,168,0,39,0,17,0,202,0,149,0,184,0,87,0,175,0,0,0,198,0,177,0,128,0,0,0,102,0,141,0,81,0,24,0,27,0,25,0,0,0,0,0,131,0,0,0,156,0,186,0,41,0,224,0,0,0,178,0,245,0,0,0,124,0,17,0,0,0,0,0,0,0,91,0,170,0,148,0,141,0,0,0,0,0,0,0,0,0,139,0,101,0,185,0,9,0,0,0,0,0,207,0,211,0,162,0,217,0,171,0,231,0,0,0,159,0,20,0,0,0,20,0,170,0,0,0,218,0,32,0,236,0,74,0,2,0,0,0,114,0,128,0,162,0,236,0,221,0,101,0,0,0,0,0,240,0,174,0,182,0,246,0,237,0,115,0,65,0,189,0,166,0,201,0,29,0,12,0,190,0,6,0,161,0,42,0,165,0,229,0,91,0,9,0,56,0,184,0,122,0,196,0,64,0,0,0,237,0,13,0,44,0,225,0,223,0,86,0,74,0,155,0,124,0,226,0,247,0,93,0,21,0,85,0,106,0,133,0,143,0,34,0,82,0,61,0,53,0,0,0,177,0,194,0,219,0,21,0,236,0,0,0,119,0,229,0,0,0,3,0,202,0,0,0,113,0,156,0,35,0,230,0,0,0,25,0,0,0,31,0,67,0,196,0,103,0,0,0,162,0,134,0,243,0,209,0,64,0,43,0,0,0,184,0,235,0,212,0,0,0,10,0,0,0,191,0,161,0,50,0,133,0,244,0,26,0,105,0,150,0,0,0,4,0,64,0,0,0,202,0,163,0,115,0,0,0,156,0,49,0,219,0,10,0,128,0,140,0,23,0,219,0,0,0,206,0,124,0,6,0,50,0,0,0,45,0,0,0,252,0,0,0,134,0,108,0,189,0,240,0,178,0,249,0,253,0,137,0,233,0,91,0,193,0,0,0,183,0,0,0,100,0,0,0,158,0,0,0,157,0,35,0,151,0,0,0,131,0,0,0,94,0,0,0,41,0,0,0,238,0,3,0,10,0,163,0,3,0,0,0,0,0,107,0,105,0,138,0,160,0,0,0,128,0,243,0,112,0,0,0,56,0,38,0,212,0,0,0,0,0,38,0,86,0,88,0,0,0,234,0,50,0,231,0,0,0,238,0,213,0,73,0,182,0,157,0,7,0,0,0,113,0,64,0,0,0,0,0,122,0,162,0,162,0,65,0,0,0,0,0,42,0,143,0,12,0,136,0,244,0,217,0,224,0,0,0,0,0,34,0,217,0,89,0,3,0,186,0,147,0,116,0,135,0,178,0,25,0,0,0,45,0,9,0,208,0,193,0,185,0,206,0,22,0,19,0,18,0,211,0,163,0,16,0,98,0,197,0,18,0,200,0,247,0,208,0,245,0,234,0,31,0,24,0,0,0,117,0,70,0,210,0,240,0,165,0,240,0,244,0,138,0,0,0,233,0,116,0,32,0,130,0,154,0,248,0,86,0,166,0,35,0,250,0,246,0,154,0,20,0,7,0,222,0,0,0,0,0,6,0,10,0,149,0,112,0,0,0,122,0,113,0,174,0,180,0,87,0,17,0,185,0,184,0,35,0,0,0,41,0,127,0,0,0,48,0,0,0,49,0,253,0,236,0,0,0,252,0,110,0,9,0,228,0,0,0,0,0,159,0,250,0,105,0,77,0,228,0,166,0,103,0,111,0,76,0,52,0,120,0,246,0,0,0,136,0,187,0,253,0,78,0,0,0,244,0,123,0,173,0,185,0,0,0,0,0,119,0,157,0,85,0,0,0,60,0,217,0,199,0,120,0,230,0,78,0,172,0,151,0,61,0,204,0,0,0,79,0,27,0,162,0,197,0,220,0,100,0,0,0,231,0,93,0,179,0,179,0,0,0,6,0,35,0,0,0,190,0,236,0,9,0,221,0,34,0,10,0,131,0,92,0,243,0,130,0,54,0,49,0,42,0,112,0,133,0,142,0,243,0,109,0,196,0,112,0,158,0,0,0,232,0,34,0,181,0,128,0,9,0,124,0,100,0,97,0,192,0,226,0,0,0,136,0,131,0,1,0,76,0,244,0,187,0,168,0,30,0,0,0,196,0,0,0,255,0,177,0,75,0,0,0,116,0,217,0,243,0,71,0,120,0,71,0,89,0,217,0,194,0,154,0,53,0,8,0,26,0,190,0,0,0,130,0,170,0,17,0,77,0,84,0,0,0,92,0,205,0,232,0,207,0,108,0,126,0,183,0,82,0,29,0,222,0,48,0,0,0,10,0,26,0,184,0,40,0,0,0,249,0,39,0,0,0,38,0,0,0,242,0,62,0,38,0,70,0,197,0,0,0,125,0,0,0,150,0,0,0,93,0,99,0,95,0,14,0,207,0,27,0,121,0,166,0,192,0,229,0,12,0,108,0,207,0,247,0,169,0,0,0,217,0,0,0,134,0,169,0,29,0,0,0,27,0,206,0,12,0,0,0,255,0,0,0,8,0,53,0,0,0,0,0,159,0,74,0,69,0,138,0,107,0,116,0,175,0,124,0,203,0,74,0,22,0,109,0,186,0,84,0,105,0,0,0,220,0,0,0,58,0,0,0,0,0,172,0,0,0,167,0,221,0,90,0,0,0,251,0,71,0,225,0,204,0,188,0,252,0,130,0,147,0,130,0,3,0,242,0,5,0,223,0,20,0,103,0,40,0,148,0,68,0,101,0,212,0,251,0,62,0,53,0,138,0,199,0,105,0,219,0,64,0,57,0,166,0,31,0,0,0,0,0,214,0,4,0,0,0,198,0,150,0,40,0,251,0,33,0,243,0,109,0,213,0,0,0,48,0,125,0,79,0,253,0,158,0,4,0,190,0,215,0,50,0,234,0,207,0,178,0,0,0,0,0,251,0,167,0,15,0,190,0,107,0,64,0,179,0,91,0,0,0,132,0,218,0,32,0,25,0,88,0,44,0,78,0,0,0,88,0,180,0,0,0,79,0,123,0,27,0,31,0,150,0,67,0,151,0,0,0,98,0,34,0,132,0,215,0,120,0,97,0,39,0,216,0,174,0,0,0,133,0,168,0,211,0,33,0,189,0,173,0,91,0,0,0,120,0,86,0,0,0,0,0,205,0,118,0,191,0,241,0,0,0,183,0,192,0,37,0,132,0,0,0,0,0,7,0,227,0,245,0,22,0,66,0,65,0,200,0,157,0,98,0,18,0,50,0,169,0,192,0,0,0,97,0,0,0,221,0,120,0,0,0,113,0,252,0,158,0,60,0,141,0,164,0,223,0,76,0,44,0,0,0,182,0,32,0,227,0,9,0,86,0,105,0,148,0,60,0,166,0,169,0,175,0,34,0,0,0,29,0,219,0,238,0,145,0,177,0,0,0,0,0,0,0,0,0,28,0,209,0,124,0,49,0,223,0,162,0,175,0,36,0,0,0,0,0,2,0,56,0,120,0,75,0,202,0,47,0,253,0,0,0,119,0,181,0,165,0,83,0,69,0,79,0,228,0,189,0,254,0,88,0,62,0,129,0,14,0,108,0,247,0,194,0,220,0,151,0,54,0,179,0,105,0,0,0,0,0,92,0,57,0,116,0,36,0,22,0,57,0,11,0,0,0);
signal scenario_full  : scenario_type := (81,31,82,31,43,31,214,31,21,31,51,31,51,30,218,31,5,31,7,31,7,30,176,31,179,31,87,31,87,30,87,29,87,28,70,31,230,31,187,31,186,31,26,31,95,31,28,31,161,31,41,31,156,31,156,30,175,31,175,30,52,31,82,31,65,31,206,31,231,31,231,30,245,31,245,31,97,31,97,30,92,31,92,30,28,31,172,31,96,31,113,31,25,31,95,31,168,31,26,31,223,31,97,31,240,31,240,30,126,31,157,31,157,30,30,31,194,31,148,31,174,31,25,31,212,31,212,30,181,31,181,30,181,29,66,31,149,31,162,31,162,30,162,29,85,31,34,31,34,30,59,31,215,31,247,31,95,31,95,30,23,31,217,31,217,30,217,29,62,31,19,31,48,31,243,31,191,31,165,31,165,30,41,31,41,30,210,31,199,31,54,31,197,31,197,30,72,31,173,31,70,31,175,31,117,31,117,30,23,31,179,31,73,31,21,31,204,31,18,31,18,30,27,31,183,31,119,31,230,31,56,31,38,31,70,31,119,31,196,31,196,30,204,31,99,31,208,31,224,31,225,31,46,31,46,30,241,31,241,30,53,31,231,31,231,30,100,31,177,31,55,31,86,31,168,31,128,31,9,31,212,31,118,31,253,31,132,31,241,31,248,31,39,31,39,30,188,31,86,31,168,31,39,31,17,31,202,31,149,31,184,31,87,31,175,31,175,30,198,31,177,31,128,31,128,30,102,31,141,31,81,31,24,31,27,31,25,31,25,30,25,29,131,31,131,30,156,31,186,31,41,31,224,31,224,30,178,31,245,31,245,30,124,31,17,31,17,30,17,29,17,28,91,31,170,31,148,31,141,31,141,30,141,29,141,28,141,27,139,31,101,31,185,31,9,31,9,30,9,29,207,31,211,31,162,31,217,31,171,31,231,31,231,30,159,31,20,31,20,30,20,31,170,31,170,30,218,31,32,31,236,31,74,31,2,31,2,30,114,31,128,31,162,31,236,31,221,31,101,31,101,30,101,29,240,31,174,31,182,31,246,31,237,31,115,31,65,31,189,31,166,31,201,31,29,31,12,31,190,31,6,31,161,31,42,31,165,31,229,31,91,31,9,31,56,31,184,31,122,31,196,31,64,31,64,30,237,31,13,31,44,31,225,31,223,31,86,31,74,31,155,31,124,31,226,31,247,31,93,31,21,31,85,31,106,31,133,31,143,31,34,31,82,31,61,31,53,31,53,30,177,31,194,31,219,31,21,31,236,31,236,30,119,31,229,31,229,30,3,31,202,31,202,30,113,31,156,31,35,31,230,31,230,30,25,31,25,30,31,31,67,31,196,31,103,31,103,30,162,31,134,31,243,31,209,31,64,31,43,31,43,30,184,31,235,31,212,31,212,30,10,31,10,30,191,31,161,31,50,31,133,31,244,31,26,31,105,31,150,31,150,30,4,31,64,31,64,30,202,31,163,31,115,31,115,30,156,31,49,31,219,31,10,31,128,31,140,31,23,31,219,31,219,30,206,31,124,31,6,31,50,31,50,30,45,31,45,30,252,31,252,30,134,31,108,31,189,31,240,31,178,31,249,31,253,31,137,31,233,31,91,31,193,31,193,30,183,31,183,30,100,31,100,30,158,31,158,30,157,31,35,31,151,31,151,30,131,31,131,30,94,31,94,30,41,31,41,30,238,31,3,31,10,31,163,31,3,31,3,30,3,29,107,31,105,31,138,31,160,31,160,30,128,31,243,31,112,31,112,30,56,31,38,31,212,31,212,30,212,29,38,31,86,31,88,31,88,30,234,31,50,31,231,31,231,30,238,31,213,31,73,31,182,31,157,31,7,31,7,30,113,31,64,31,64,30,64,29,122,31,162,31,162,31,65,31,65,30,65,29,42,31,143,31,12,31,136,31,244,31,217,31,224,31,224,30,224,29,34,31,217,31,89,31,3,31,186,31,147,31,116,31,135,31,178,31,25,31,25,30,45,31,9,31,208,31,193,31,185,31,206,31,22,31,19,31,18,31,211,31,163,31,16,31,98,31,197,31,18,31,200,31,247,31,208,31,245,31,234,31,31,31,24,31,24,30,117,31,70,31,210,31,240,31,165,31,240,31,244,31,138,31,138,30,233,31,116,31,32,31,130,31,154,31,248,31,86,31,166,31,35,31,250,31,246,31,154,31,20,31,7,31,222,31,222,30,222,29,6,31,10,31,149,31,112,31,112,30,122,31,113,31,174,31,180,31,87,31,17,31,185,31,184,31,35,31,35,30,41,31,127,31,127,30,48,31,48,30,49,31,253,31,236,31,236,30,252,31,110,31,9,31,228,31,228,30,228,29,159,31,250,31,105,31,77,31,228,31,166,31,103,31,111,31,76,31,52,31,120,31,246,31,246,30,136,31,187,31,253,31,78,31,78,30,244,31,123,31,173,31,185,31,185,30,185,29,119,31,157,31,85,31,85,30,60,31,217,31,199,31,120,31,230,31,78,31,172,31,151,31,61,31,204,31,204,30,79,31,27,31,162,31,197,31,220,31,100,31,100,30,231,31,93,31,179,31,179,31,179,30,6,31,35,31,35,30,190,31,236,31,9,31,221,31,34,31,10,31,131,31,92,31,243,31,130,31,54,31,49,31,42,31,112,31,133,31,142,31,243,31,109,31,196,31,112,31,158,31,158,30,232,31,34,31,181,31,128,31,9,31,124,31,100,31,97,31,192,31,226,31,226,30,136,31,131,31,1,31,76,31,244,31,187,31,168,31,30,31,30,30,196,31,196,30,255,31,177,31,75,31,75,30,116,31,217,31,243,31,71,31,120,31,71,31,89,31,217,31,194,31,154,31,53,31,8,31,26,31,190,31,190,30,130,31,170,31,17,31,77,31,84,31,84,30,92,31,205,31,232,31,207,31,108,31,126,31,183,31,82,31,29,31,222,31,48,31,48,30,10,31,26,31,184,31,40,31,40,30,249,31,39,31,39,30,38,31,38,30,242,31,62,31,38,31,70,31,197,31,197,30,125,31,125,30,150,31,150,30,93,31,99,31,95,31,14,31,207,31,27,31,121,31,166,31,192,31,229,31,12,31,108,31,207,31,247,31,169,31,169,30,217,31,217,30,134,31,169,31,29,31,29,30,27,31,206,31,12,31,12,30,255,31,255,30,8,31,53,31,53,30,53,29,159,31,74,31,69,31,138,31,107,31,116,31,175,31,124,31,203,31,74,31,22,31,109,31,186,31,84,31,105,31,105,30,220,31,220,30,58,31,58,30,58,29,172,31,172,30,167,31,221,31,90,31,90,30,251,31,71,31,225,31,204,31,188,31,252,31,130,31,147,31,130,31,3,31,242,31,5,31,223,31,20,31,103,31,40,31,148,31,68,31,101,31,212,31,251,31,62,31,53,31,138,31,199,31,105,31,219,31,64,31,57,31,166,31,31,31,31,30,31,29,214,31,4,31,4,30,198,31,150,31,40,31,251,31,33,31,243,31,109,31,213,31,213,30,48,31,125,31,79,31,253,31,158,31,4,31,190,31,215,31,50,31,234,31,207,31,178,31,178,30,178,29,251,31,167,31,15,31,190,31,107,31,64,31,179,31,91,31,91,30,132,31,218,31,32,31,25,31,88,31,44,31,78,31,78,30,88,31,180,31,180,30,79,31,123,31,27,31,31,31,150,31,67,31,151,31,151,30,98,31,34,31,132,31,215,31,120,31,97,31,39,31,216,31,174,31,174,30,133,31,168,31,211,31,33,31,189,31,173,31,91,31,91,30,120,31,86,31,86,30,86,29,205,31,118,31,191,31,241,31,241,30,183,31,192,31,37,31,132,31,132,30,132,29,7,31,227,31,245,31,22,31,66,31,65,31,200,31,157,31,98,31,18,31,50,31,169,31,192,31,192,30,97,31,97,30,221,31,120,31,120,30,113,31,252,31,158,31,60,31,141,31,164,31,223,31,76,31,44,31,44,30,182,31,32,31,227,31,9,31,86,31,105,31,148,31,60,31,166,31,169,31,175,31,34,31,34,30,29,31,219,31,238,31,145,31,177,31,177,30,177,29,177,28,177,27,28,31,209,31,124,31,49,31,223,31,162,31,175,31,36,31,36,30,36,29,2,31,56,31,120,31,75,31,202,31,47,31,253,31,253,30,119,31,181,31,165,31,83,31,69,31,79,31,228,31,189,31,254,31,88,31,62,31,129,31,14,31,108,31,247,31,194,31,220,31,151,31,54,31,179,31,105,31,105,30,105,29,92,31,57,31,116,31,36,31,22,31,57,31,11,31,11,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
