-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1001;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,229,0,0,0,197,0,8,0,159,0,54,0,99,0,161,0,181,0,15,0,161,0,0,0,200,0,95,0,243,0,226,0,225,0,0,0,77,0,56,0,92,0,185,0,0,0,229,0,127,0,14,0,104,0,19,0,0,0,30,0,203,0,167,0,98,0,250,0,185,0,0,0,241,0,140,0,228,0,0,0,0,0,223,0,6,0,42,0,0,0,157,0,3,0,0,0,183,0,48,0,34,0,37,0,127,0,48,0,42,0,182,0,153,0,216,0,200,0,29,0,171,0,61,0,20,0,199,0,134,0,20,0,162,0,40,0,194,0,22,0,186,0,0,0,83,0,0,0,229,0,70,0,212,0,249,0,0,0,125,0,15,0,251,0,98,0,105,0,226,0,108,0,143,0,0,0,0,0,127,0,157,0,0,0,90,0,183,0,225,0,108,0,0,0,213,0,214,0,94,0,205,0,164,0,167,0,184,0,44,0,0,0,140,0,196,0,88,0,208,0,235,0,16,0,0,0,116,0,142,0,32,0,1,0,0,0,41,0,158,0,220,0,49,0,169,0,253,0,164,0,122,0,31,0,203,0,71,0,204,0,0,0,58,0,23,0,247,0,174,0,82,0,196,0,79,0,87,0,0,0,121,0,0,0,133,0,23,0,26,0,126,0,186,0,213,0,193,0,245,0,232,0,0,0,136,0,31,0,81,0,0,0,177,0,54,0,28,0,0,0,170,0,12,0,0,0,232,0,242,0,240,0,0,0,235,0,13,0,62,0,10,0,177,0,129,0,176,0,191,0,0,0,0,0,0,0,0,0,201,0,65,0,36,0,134,0,0,0,6,0,109,0,35,0,0,0,153,0,179,0,211,0,180,0,167,0,177,0,149,0,152,0,145,0,44,0,20,0,88,0,129,0,144,0,13,0,37,0,5,0,153,0,4,0,213,0,113,0,0,0,151,0,174,0,209,0,212,0,194,0,229,0,32,0,80,0,216,0,102,0,0,0,65,0,62,0,0,0,229,0,50,0,149,0,215,0,21,0,61,0,0,0,235,0,90,0,116,0,110,0,103,0,242,0,197,0,97,0,241,0,107,0,246,0,0,0,162,0,0,0,51,0,205,0,46,0,133,0,60,0,153,0,241,0,186,0,161,0,30,0,139,0,0,0,219,0,163,0,51,0,115,0,217,0,80,0,213,0,0,0,219,0,25,0,31,0,0,0,219,0,45,0,170,0,126,0,8,0,88,0,75,0,146,0,210,0,136,0,0,0,4,0,0,0,122,0,241,0,210,0,1,0,175,0,107,0,0,0,0,0,155,0,226,0,141,0,90,0,132,0,0,0,77,0,74,0,225,0,0,0,0,0,81,0,0,0,5,0,0,0,0,0,2,0,93,0,189,0,162,0,252,0,0,0,48,0,12,0,116,0,0,0,73,0,0,0,114,0,110,0,65,0,0,0,202,0,0,0,206,0,0,0,20,0,243,0,61,0,226,0,0,0,0,0,0,0,142,0,112,0,231,0,79,0,129,0,146,0,180,0,241,0,217,0,169,0,85,0,136,0,165,0,26,0,0,0,211,0,0,0,207,0,0,0,238,0,97,0,219,0,88,0,25,0,70,0,212,0,0,0,228,0,0,0,0,0,116,0,22,0,44,0,135,0,75,0,180,0,103,0,0,0,17,0,173,0,195,0,0,0,238,0,44,0,0,0,30,0,0,0,131,0,166,0,207,0,0,0,127,0,204,0,97,0,0,0,99,0,237,0,201,0,254,0,128,0,83,0,37,0,77,0,110,0,0,0,0,0,188,0,6,0,255,0,168,0,100,0,0,0,114,0,14,0,161,0,0,0,108,0,113,0,196,0,198,0,150,0,0,0,56,0,138,0,93,0,95,0,166,0,0,0,207,0,195,0,94,0,0,0,0,0,48,0,215,0,160,0,0,0,57,0,188,0,84,0,0,0,233,0,76,0,157,0,0,0,112,0,0,0,242,0,32,0,118,0,167,0,74,0,60,0,17,0,29,0,102,0,70,0,143,0,207,0,149,0,214,0,168,0,80,0,80,0,148,0,0,0,50,0,71,0,73,0,23,0,12,0,0,0,0,0,133,0,220,0,127,0,184,0,5,0,118,0,210,0,32,0,107,0,136,0,143,0,49,0,87,0,219,0,99,0,187,0,166,0,112,0,99,0,230,0,215,0,241,0,125,0,99,0,68,0,147,0,2,0,0,0,177,0,84,0,64,0,145,0,167,0,137,0,45,0,129,0,224,0,163,0,96,0,165,0,67,0,151,0,125,0,255,0,253,0,0,0,26,0,0,0,0,0,237,0,205,0,0,0,238,0,120,0,200,0,10,0,187,0,18,0,82,0,0,0,71,0,81,0,0,0,51,0,92,0,235,0,106,0,155,0,0,0,0,0,135,0,0,0,0,0,0,0,16,0,11,0,124,0,85,0,43,0,209,0,65,0,32,0,0,0,41,0,197,0,44,0,128,0,118,0,87,0,159,0,200,0,92,0,193,0,114,0,212,0,120,0,149,0,38,0,149,0,66,0,207,0,1,0,219,0,0,0,201,0,150,0,162,0,87,0,0,0,190,0,15,0,0,0,227,0,34,0,226,0,174,0,151,0,67,0,206,0,237,0,142,0,47,0,199,0,178,0,31,0,176,0,61,0,66,0,130,0,69,0,222,0,231,0,199,0,24,0,201,0,208,0,215,0,0,0,192,0,162,0,43,0,100,0,35,0,192,0,208,0,205,0,126,0,231,0,0,0,0,0,50,0,146,0,0,0,9,0,244,0,21,0,213,0,27,0,236,0,250,0,161,0,165,0,128,0,101,0,204,0,21,0,147,0,92,0,129,0,0,0,0,0,128,0,0,0,201,0,167,0,2,0,78,0,11,0,70,0,14,0,232,0,213,0,0,0,240,0,110,0,149,0,114,0,31,0,14,0,0,0,209,0,239,0,191,0,199,0,53,0,0,0,0,0,227,0,152,0,32,0,106,0,242,0,195,0,54,0,151,0,27,0,0,0,228,0,0,0,246,0,231,0,95,0,238,0,31,0,162,0,0,0,63,0,180,0,120,0,172,0,32,0,159,0,134,0,0,0,93,0,65,0,173,0,178,0,58,0,112,0,0,0,183,0,151,0,55,0,0,0,117,0,64,0,0,0,161,0,0,0,128,0,0,0,170,0,111,0,15,0,0,0,213,0,39,0,71,0,89,0,60,0,0,0,0,0,241,0,106,0,34,0,17,0,0,0,0,0,29,0,56,0,0,0,0,0,46,0,0,0,18,0,102,0,86,0,30,0,134,0,48,0,227,0,234,0,0,0,146,0,71,0,99,0,0,0,0,0,101,0,208,0,12,0,112,0,160,0,241,0,145,0,186,0,0,0,202,0,150,0,161,0,0,0,146,0,0,0,135,0,186,0,89,0,0,0,226,0,41,0,142,0,146,0,75,0,7,0,96,0,5,0,188,0,208,0,242,0,0,0,90,0,240,0,231,0,170,0,16,0,0,0,0,0,98,0,221,0,0,0,160,0,223,0,0,0,194,0,155,0,14,0,0,0,153,0,88,0,51,0,124,0,68,0,250,0,128,0,61,0,0,0,245,0,248,0,62,0,119,0,65,0,51,0,194,0,0,0,129,0,0,0,53,0,174,0,63,0,98,0,170,0,209,0,138,0,62,0,107,0,128,0,166,0,202,0,111,0,0,0,119,0,96,0,73,0,0,0,147,0,30,0,180,0,1,0,128,0,0,0,139,0,144,0,0,0,240,0,201,0,172,0,90,0,0,0,214,0,175,0,66,0,0,0,53,0,237,0,77,0,41,0,59,0,0,0,238,0,25,0,12,0,191,0,245,0,169,0,0,0,0,0,0,0,177,0,0,0,225,0,171,0,198,0,203,0,145,0,22,0,221,0,177,0,62,0,86,0,139,0,139,0,146,0,5,0,117,0,130,0,46,0,197,0,20,0,86,0,99,0,0,0,0,0,0,0,0,0,0,0,70,0,48,0,213,0,233,0,202,0,112,0,70,0,0,0,63,0,181,0,204,0,218,0,0,0,0,0,209,0,0,0,211,0,0,0,161,0,104,0,251,0,0,0,81,0,194,0,85,0,125,0,0,0,225,0,0,0,118,0,80,0,241,0,0,0,107,0,0,0,196,0,189,0,129,0,0,0,110,0,240,0,5,0,112,0,0,0,221,0,72,0,93,0,73,0,187,0,27,0,142,0,212,0,155,0,197,0,153,0,167,0,163,0,53,0,31,0,135,0,0,0,194,0,104,0,41,0,122,0,31,0,93,0,190,0,0,0,163,0,82,0,162,0,188,0,59,0,230,0,133,0,155,0,124,0,48,0,0,0,45,0,26,0,59,0,152,0,229,0,22,0,0,0,234,0,148,0,126,0,206,0,248,0,154,0,236,0,1,0,23,0,51,0,151,0,40,0,252,0,177,0,140,0,72,0,133,0,0,0,0,0,147,0,34,0,246,0);
signal scenario_full  : scenario_type := (0,0,229,31,229,30,197,31,8,31,159,31,54,31,99,31,161,31,181,31,15,31,161,31,161,30,200,31,95,31,243,31,226,31,225,31,225,30,77,31,56,31,92,31,185,31,185,30,229,31,127,31,14,31,104,31,19,31,19,30,30,31,203,31,167,31,98,31,250,31,185,31,185,30,241,31,140,31,228,31,228,30,228,29,223,31,6,31,42,31,42,30,157,31,3,31,3,30,183,31,48,31,34,31,37,31,127,31,48,31,42,31,182,31,153,31,216,31,200,31,29,31,171,31,61,31,20,31,199,31,134,31,20,31,162,31,40,31,194,31,22,31,186,31,186,30,83,31,83,30,229,31,70,31,212,31,249,31,249,30,125,31,15,31,251,31,98,31,105,31,226,31,108,31,143,31,143,30,143,29,127,31,157,31,157,30,90,31,183,31,225,31,108,31,108,30,213,31,214,31,94,31,205,31,164,31,167,31,184,31,44,31,44,30,140,31,196,31,88,31,208,31,235,31,16,31,16,30,116,31,142,31,32,31,1,31,1,30,41,31,158,31,220,31,49,31,169,31,253,31,164,31,122,31,31,31,203,31,71,31,204,31,204,30,58,31,23,31,247,31,174,31,82,31,196,31,79,31,87,31,87,30,121,31,121,30,133,31,23,31,26,31,126,31,186,31,213,31,193,31,245,31,232,31,232,30,136,31,31,31,81,31,81,30,177,31,54,31,28,31,28,30,170,31,12,31,12,30,232,31,242,31,240,31,240,30,235,31,13,31,62,31,10,31,177,31,129,31,176,31,191,31,191,30,191,29,191,28,191,27,201,31,65,31,36,31,134,31,134,30,6,31,109,31,35,31,35,30,153,31,179,31,211,31,180,31,167,31,177,31,149,31,152,31,145,31,44,31,20,31,88,31,129,31,144,31,13,31,37,31,5,31,153,31,4,31,213,31,113,31,113,30,151,31,174,31,209,31,212,31,194,31,229,31,32,31,80,31,216,31,102,31,102,30,65,31,62,31,62,30,229,31,50,31,149,31,215,31,21,31,61,31,61,30,235,31,90,31,116,31,110,31,103,31,242,31,197,31,97,31,241,31,107,31,246,31,246,30,162,31,162,30,51,31,205,31,46,31,133,31,60,31,153,31,241,31,186,31,161,31,30,31,139,31,139,30,219,31,163,31,51,31,115,31,217,31,80,31,213,31,213,30,219,31,25,31,31,31,31,30,219,31,45,31,170,31,126,31,8,31,88,31,75,31,146,31,210,31,136,31,136,30,4,31,4,30,122,31,241,31,210,31,1,31,175,31,107,31,107,30,107,29,155,31,226,31,141,31,90,31,132,31,132,30,77,31,74,31,225,31,225,30,225,29,81,31,81,30,5,31,5,30,5,29,2,31,93,31,189,31,162,31,252,31,252,30,48,31,12,31,116,31,116,30,73,31,73,30,114,31,110,31,65,31,65,30,202,31,202,30,206,31,206,30,20,31,243,31,61,31,226,31,226,30,226,29,226,28,142,31,112,31,231,31,79,31,129,31,146,31,180,31,241,31,217,31,169,31,85,31,136,31,165,31,26,31,26,30,211,31,211,30,207,31,207,30,238,31,97,31,219,31,88,31,25,31,70,31,212,31,212,30,228,31,228,30,228,29,116,31,22,31,44,31,135,31,75,31,180,31,103,31,103,30,17,31,173,31,195,31,195,30,238,31,44,31,44,30,30,31,30,30,131,31,166,31,207,31,207,30,127,31,204,31,97,31,97,30,99,31,237,31,201,31,254,31,128,31,83,31,37,31,77,31,110,31,110,30,110,29,188,31,6,31,255,31,168,31,100,31,100,30,114,31,14,31,161,31,161,30,108,31,113,31,196,31,198,31,150,31,150,30,56,31,138,31,93,31,95,31,166,31,166,30,207,31,195,31,94,31,94,30,94,29,48,31,215,31,160,31,160,30,57,31,188,31,84,31,84,30,233,31,76,31,157,31,157,30,112,31,112,30,242,31,32,31,118,31,167,31,74,31,60,31,17,31,29,31,102,31,70,31,143,31,207,31,149,31,214,31,168,31,80,31,80,31,148,31,148,30,50,31,71,31,73,31,23,31,12,31,12,30,12,29,133,31,220,31,127,31,184,31,5,31,118,31,210,31,32,31,107,31,136,31,143,31,49,31,87,31,219,31,99,31,187,31,166,31,112,31,99,31,230,31,215,31,241,31,125,31,99,31,68,31,147,31,2,31,2,30,177,31,84,31,64,31,145,31,167,31,137,31,45,31,129,31,224,31,163,31,96,31,165,31,67,31,151,31,125,31,255,31,253,31,253,30,26,31,26,30,26,29,237,31,205,31,205,30,238,31,120,31,200,31,10,31,187,31,18,31,82,31,82,30,71,31,81,31,81,30,51,31,92,31,235,31,106,31,155,31,155,30,155,29,135,31,135,30,135,29,135,28,16,31,11,31,124,31,85,31,43,31,209,31,65,31,32,31,32,30,41,31,197,31,44,31,128,31,118,31,87,31,159,31,200,31,92,31,193,31,114,31,212,31,120,31,149,31,38,31,149,31,66,31,207,31,1,31,219,31,219,30,201,31,150,31,162,31,87,31,87,30,190,31,15,31,15,30,227,31,34,31,226,31,174,31,151,31,67,31,206,31,237,31,142,31,47,31,199,31,178,31,31,31,176,31,61,31,66,31,130,31,69,31,222,31,231,31,199,31,24,31,201,31,208,31,215,31,215,30,192,31,162,31,43,31,100,31,35,31,192,31,208,31,205,31,126,31,231,31,231,30,231,29,50,31,146,31,146,30,9,31,244,31,21,31,213,31,27,31,236,31,250,31,161,31,165,31,128,31,101,31,204,31,21,31,147,31,92,31,129,31,129,30,129,29,128,31,128,30,201,31,167,31,2,31,78,31,11,31,70,31,14,31,232,31,213,31,213,30,240,31,110,31,149,31,114,31,31,31,14,31,14,30,209,31,239,31,191,31,199,31,53,31,53,30,53,29,227,31,152,31,32,31,106,31,242,31,195,31,54,31,151,31,27,31,27,30,228,31,228,30,246,31,231,31,95,31,238,31,31,31,162,31,162,30,63,31,180,31,120,31,172,31,32,31,159,31,134,31,134,30,93,31,65,31,173,31,178,31,58,31,112,31,112,30,183,31,151,31,55,31,55,30,117,31,64,31,64,30,161,31,161,30,128,31,128,30,170,31,111,31,15,31,15,30,213,31,39,31,71,31,89,31,60,31,60,30,60,29,241,31,106,31,34,31,17,31,17,30,17,29,29,31,56,31,56,30,56,29,46,31,46,30,18,31,102,31,86,31,30,31,134,31,48,31,227,31,234,31,234,30,146,31,71,31,99,31,99,30,99,29,101,31,208,31,12,31,112,31,160,31,241,31,145,31,186,31,186,30,202,31,150,31,161,31,161,30,146,31,146,30,135,31,186,31,89,31,89,30,226,31,41,31,142,31,146,31,75,31,7,31,96,31,5,31,188,31,208,31,242,31,242,30,90,31,240,31,231,31,170,31,16,31,16,30,16,29,98,31,221,31,221,30,160,31,223,31,223,30,194,31,155,31,14,31,14,30,153,31,88,31,51,31,124,31,68,31,250,31,128,31,61,31,61,30,245,31,248,31,62,31,119,31,65,31,51,31,194,31,194,30,129,31,129,30,53,31,174,31,63,31,98,31,170,31,209,31,138,31,62,31,107,31,128,31,166,31,202,31,111,31,111,30,119,31,96,31,73,31,73,30,147,31,30,31,180,31,1,31,128,31,128,30,139,31,144,31,144,30,240,31,201,31,172,31,90,31,90,30,214,31,175,31,66,31,66,30,53,31,237,31,77,31,41,31,59,31,59,30,238,31,25,31,12,31,191,31,245,31,169,31,169,30,169,29,169,28,177,31,177,30,225,31,171,31,198,31,203,31,145,31,22,31,221,31,177,31,62,31,86,31,139,31,139,31,146,31,5,31,117,31,130,31,46,31,197,31,20,31,86,31,99,31,99,30,99,29,99,28,99,27,99,26,70,31,48,31,213,31,233,31,202,31,112,31,70,31,70,30,63,31,181,31,204,31,218,31,218,30,218,29,209,31,209,30,211,31,211,30,161,31,104,31,251,31,251,30,81,31,194,31,85,31,125,31,125,30,225,31,225,30,118,31,80,31,241,31,241,30,107,31,107,30,196,31,189,31,129,31,129,30,110,31,240,31,5,31,112,31,112,30,221,31,72,31,93,31,73,31,187,31,27,31,142,31,212,31,155,31,197,31,153,31,167,31,163,31,53,31,31,31,135,31,135,30,194,31,104,31,41,31,122,31,31,31,93,31,190,31,190,30,163,31,82,31,162,31,188,31,59,31,230,31,133,31,155,31,124,31,48,31,48,30,45,31,26,31,59,31,152,31,229,31,22,31,22,30,234,31,148,31,126,31,206,31,248,31,154,31,236,31,1,31,23,31,51,31,151,31,40,31,252,31,177,31,140,31,72,31,133,31,133,30,133,29,147,31,34,31,246,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
