-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_750 is
end project_tb_750;

architecture project_tb_arch_750 of project_tb_750 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 976;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,38,0,247,0,101,0,217,0,31,0,237,0,30,0,201,0,86,0,103,0,21,0,0,0,11,0,233,0,181,0,83,0,208,0,0,0,213,0,244,0,0,0,210,0,154,0,194,0,1,0,134,0,0,0,33,0,34,0,207,0,48,0,205,0,64,0,171,0,201,0,160,0,130,0,0,0,138,0,0,0,153,0,209,0,83,0,0,0,0,0,204,0,243,0,172,0,0,0,185,0,48,0,19,0,170,0,19,0,0,0,103,0,0,0,136,0,55,0,0,0,129,0,80,0,6,0,0,0,7,0,86,0,141,0,95,0,122,0,22,0,29,0,169,0,190,0,12,0,33,0,9,0,197,0,71,0,197,0,30,0,184,0,63,0,118,0,199,0,159,0,0,0,170,0,0,0,155,0,231,0,179,0,0,0,193,0,144,0,34,0,194,0,105,0,53,0,133,0,46,0,0,0,9,0,0,0,0,0,205,0,12,0,231,0,0,0,24,0,124,0,171,0,0,0,18,0,255,0,14,0,127,0,0,0,196,0,172,0,210,0,247,0,0,0,0,0,212,0,35,0,0,0,224,0,235,0,111,0,232,0,238,0,0,0,52,0,0,0,255,0,0,0,0,0,74,0,109,0,17,0,181,0,105,0,156,0,22,0,0,0,165,0,111,0,126,0,239,0,223,0,196,0,0,0,208,0,229,0,64,0,23,0,201,0,69,0,60,0,148,0,199,0,0,0,0,0,103,0,216,0,25,0,179,0,0,0,74,0,27,0,45,0,221,0,162,0,42,0,220,0,158,0,227,0,23,0,102,0,169,0,161,0,0,0,0,0,230,0,226,0,48,0,61,0,249,0,4,0,103,0,0,0,92,0,0,0,47,0,172,0,110,0,101,0,0,0,71,0,35,0,239,0,194,0,113,0,0,0,77,0,0,0,64,0,254,0,30,0,123,0,48,0,29,0,43,0,59,0,0,0,71,0,8,0,166,0,192,0,0,0,120,0,151,0,80,0,0,0,157,0,33,0,144,0,42,0,0,0,105,0,154,0,110,0,101,0,21,0,157,0,0,0,81,0,45,0,0,0,188,0,49,0,244,0,239,0,17,0,150,0,237,0,40,0,96,0,47,0,161,0,31,0,0,0,67,0,211,0,88,0,0,0,252,0,142,0,240,0,0,0,0,0,0,0,155,0,8,0,0,0,250,0,0,0,0,0,0,0,114,0,107,0,232,0,79,0,38,0,36,0,46,0,6,0,216,0,115,0,0,0,22,0,146,0,147,0,240,0,0,0,126,0,217,0,122,0,140,0,208,0,219,0,91,0,220,0,0,0,181,0,151,0,200,0,85,0,165,0,0,0,72,0,233,0,0,0,251,0,128,0,156,0,59,0,32,0,235,0,112,0,126,0,24,0,45,0,78,0,145,0,91,0,193,0,0,0,242,0,70,0,0,0,44,0,210,0,93,0,0,0,47,0,7,0,55,0,244,0,89,0,0,0,156,0,0,0,0,0,107,0,1,0,202,0,22,0,98,0,0,0,9,0,127,0,0,0,237,0,192,0,131,0,196,0,42,0,37,0,60,0,90,0,165,0,0,0,178,0,201,0,0,0,87,0,44,0,0,0,54,0,241,0,93,0,0,0,30,0,144,0,135,0,0,0,254,0,114,0,214,0,168,0,70,0,56,0,60,0,77,0,235,0,146,0,130,0,218,0,0,0,36,0,0,0,0,0,80,0,0,0,158,0,82,0,234,0,7,0,177,0,141,0,0,0,203,0,2,0,60,0,0,0,108,0,0,0,82,0,75,0,56,0,211,0,172,0,95,0,68,0,155,0,181,0,93,0,205,0,47,0,0,0,0,0,247,0,119,0,185,0,167,0,101,0,0,0,61,0,168,0,0,0,174,0,45,0,0,0,0,0,0,0,28,0,71,0,4,0,160,0,0,0,120,0,155,0,231,0,251,0,77,0,95,0,161,0,49,0,9,0,156,0,48,0,39,0,131,0,68,0,197,0,158,0,127,0,177,0,209,0,103,0,159,0,229,0,148,0,0,0,190,0,177,0,51,0,0,0,218,0,240,0,16,0,0,0,0,0,236,0,0,0,113,0,209,0,0,0,0,0,0,0,0,0,78,0,75,0,246,0,124,0,202,0,248,0,201,0,0,0,0,0,248,0,152,0,29,0,202,0,54,0,0,0,222,0,48,0,7,0,144,0,108,0,45,0,75,0,194,0,85,0,220,0,94,0,74,0,205,0,53,0,213,0,172,0,162,0,51,0,171,0,208,0,4,0,13,0,0,0,33,0,40,0,91,0,136,0,89,0,45,0,253,0,197,0,230,0,5,0,0,0,0,0,209,0,242,0,0,0,83,0,99,0,0,0,37,0,191,0,0,0,185,0,0,0,0,0,167,0,235,0,34,0,84,0,48,0,25,0,0,0,21,0,218,0,209,0,19,0,79,0,109,0,240,0,70,0,57,0,44,0,11,0,195,0,0,0,0,0,131,0,0,0,0,0,123,0,0,0,0,0,172,0,230,0,248,0,36,0,245,0,0,0,60,0,46,0,19,0,28,0,154,0,0,0,225,0,0,0,167,0,0,0,236,0,49,0,0,0,207,0,0,0,0,0,78,0,189,0,25,0,140,0,167,0,213,0,119,0,146,0,228,0,152,0,0,0,122,0,12,0,223,0,0,0,0,0,0,0,0,0,208,0,0,0,0,0,71,0,0,0,92,0,0,0,0,0,161,0,67,0,63,0,70,0,0,0,79,0,180,0,0,0,178,0,59,0,49,0,136,0,34,0,81,0,51,0,217,0,219,0,51,0,0,0,79,0,191,0,0,0,0,0,72,0,67,0,85,0,105,0,253,0,121,0,78,0,0,0,66,0,253,0,106,0,0,0,157,0,192,0,0,0,0,0,40,0,0,0,0,0,173,0,175,0,221,0,0,0,138,0,177,0,204,0,60,0,237,0,138,0,153,0,108,0,97,0,142,0,89,0,101,0,212,0,126,0,185,0,133,0,117,0,66,0,25,0,11,0,0,0,223,0,165,0,0,0,0,0,78,0,111,0,0,0,85,0,224,0,8,0,60,0,0,0,226,0,45,0,0,0,233,0,36,0,58,0,234,0,233,0,0,0,151,0,131,0,191,0,0,0,0,0,0,0,230,0,86,0,0,0,107,0,0,0,0,0,58,0,234,0,93,0,145,0,152,0,115,0,224,0,200,0,202,0,0,0,113,0,243,0,192,0,0,0,96,0,143,0,0,0,184,0,200,0,0,0,242,0,167,0,77,0,40,0,0,0,187,0,109,0,125,0,83,0,100,0,4,0,211,0,42,0,0,0,173,0,0,0,6,0,68,0,1,0,78,0,246,0,0,0,140,0,0,0,25,0,0,0,9,0,37,0,175,0,141,0,164,0,0,0,193,0,132,0,0,0,0,0,207,0,83,0,0,0,76,0,0,0,220,0,0,0,168,0,0,0,242,0,15,0,202,0,50,0,226,0,38,0,126,0,202,0,90,0,25,0,182,0,149,0,0,0,47,0,153,0,186,0,252,0,30,0,214,0,0,0,198,0,42,0,0,0,177,0,235,0,116,0,0,0,144,0,98,0,0,0,167,0,0,0,33,0,159,0,119,0,176,0,182,0,0,0,0,0,0,0,0,0,186,0,0,0,60,0,67,0,189,0,148,0,5,0,186,0,237,0,238,0,0,0,154,0,135,0,212,0,142,0,129,0,203,0,160,0,0,0,59,0,203,0,51,0,73,0,46,0,218,0,225,0,181,0,239,0,45,0,37,0,124,0,0,0,180,0,196,0,233,0,11,0,197,0,199,0,100,0,100,0,17,0,43,0,134,0,253,0,49,0,136,0,174,0,208,0,119,0,0,0,0,0,86,0,129,0,175,0,103,0,90,0,0,0,232,0,0,0,244,0,133,0,42,0,64,0,232,0,93,0,3,0,155,0,101,0,13,0,98,0,0,0,131,0,29,0,8,0,0,0,66,0,99,0,189,0,44,0,74,0,230,0,184,0,198,0,145,0,143,0,103,0,235,0,191,0,188,0,99,0,75,0,0,0,83,0,0,0,109,0,254,0,112,0,145,0,0,0,233,0,172,0,92,0,7,0,205,0,0,0,0,0,246,0,59,0,90,0,87,0,251,0,156,0,59,0,208,0,0,0,106,0,100,0,24,0,254,0,223,0,76,0,3,0,203,0,154,0,12,0,209,0,238,0,96,0,0,0,192,0,23,0,0,0,53,0,0,0,140,0,30,0,9,0,183,0,29,0,231,0,72,0,133,0,186,0,190,0,0,0,220,0,0,0,0,0,172,0,140,0,246,0,99,0,151,0,247,0,0,0,212,0,167,0,192,0,120,0,64,0);
signal scenario_full  : scenario_type := (0,0,38,31,247,31,101,31,217,31,31,31,237,31,30,31,201,31,86,31,103,31,21,31,21,30,11,31,233,31,181,31,83,31,208,31,208,30,213,31,244,31,244,30,210,31,154,31,194,31,1,31,134,31,134,30,33,31,34,31,207,31,48,31,205,31,64,31,171,31,201,31,160,31,130,31,130,30,138,31,138,30,153,31,209,31,83,31,83,30,83,29,204,31,243,31,172,31,172,30,185,31,48,31,19,31,170,31,19,31,19,30,103,31,103,30,136,31,55,31,55,30,129,31,80,31,6,31,6,30,7,31,86,31,141,31,95,31,122,31,22,31,29,31,169,31,190,31,12,31,33,31,9,31,197,31,71,31,197,31,30,31,184,31,63,31,118,31,199,31,159,31,159,30,170,31,170,30,155,31,231,31,179,31,179,30,193,31,144,31,34,31,194,31,105,31,53,31,133,31,46,31,46,30,9,31,9,30,9,29,205,31,12,31,231,31,231,30,24,31,124,31,171,31,171,30,18,31,255,31,14,31,127,31,127,30,196,31,172,31,210,31,247,31,247,30,247,29,212,31,35,31,35,30,224,31,235,31,111,31,232,31,238,31,238,30,52,31,52,30,255,31,255,30,255,29,74,31,109,31,17,31,181,31,105,31,156,31,22,31,22,30,165,31,111,31,126,31,239,31,223,31,196,31,196,30,208,31,229,31,64,31,23,31,201,31,69,31,60,31,148,31,199,31,199,30,199,29,103,31,216,31,25,31,179,31,179,30,74,31,27,31,45,31,221,31,162,31,42,31,220,31,158,31,227,31,23,31,102,31,169,31,161,31,161,30,161,29,230,31,226,31,48,31,61,31,249,31,4,31,103,31,103,30,92,31,92,30,47,31,172,31,110,31,101,31,101,30,71,31,35,31,239,31,194,31,113,31,113,30,77,31,77,30,64,31,254,31,30,31,123,31,48,31,29,31,43,31,59,31,59,30,71,31,8,31,166,31,192,31,192,30,120,31,151,31,80,31,80,30,157,31,33,31,144,31,42,31,42,30,105,31,154,31,110,31,101,31,21,31,157,31,157,30,81,31,45,31,45,30,188,31,49,31,244,31,239,31,17,31,150,31,237,31,40,31,96,31,47,31,161,31,31,31,31,30,67,31,211,31,88,31,88,30,252,31,142,31,240,31,240,30,240,29,240,28,155,31,8,31,8,30,250,31,250,30,250,29,250,28,114,31,107,31,232,31,79,31,38,31,36,31,46,31,6,31,216,31,115,31,115,30,22,31,146,31,147,31,240,31,240,30,126,31,217,31,122,31,140,31,208,31,219,31,91,31,220,31,220,30,181,31,151,31,200,31,85,31,165,31,165,30,72,31,233,31,233,30,251,31,128,31,156,31,59,31,32,31,235,31,112,31,126,31,24,31,45,31,78,31,145,31,91,31,193,31,193,30,242,31,70,31,70,30,44,31,210,31,93,31,93,30,47,31,7,31,55,31,244,31,89,31,89,30,156,31,156,30,156,29,107,31,1,31,202,31,22,31,98,31,98,30,9,31,127,31,127,30,237,31,192,31,131,31,196,31,42,31,37,31,60,31,90,31,165,31,165,30,178,31,201,31,201,30,87,31,44,31,44,30,54,31,241,31,93,31,93,30,30,31,144,31,135,31,135,30,254,31,114,31,214,31,168,31,70,31,56,31,60,31,77,31,235,31,146,31,130,31,218,31,218,30,36,31,36,30,36,29,80,31,80,30,158,31,82,31,234,31,7,31,177,31,141,31,141,30,203,31,2,31,60,31,60,30,108,31,108,30,82,31,75,31,56,31,211,31,172,31,95,31,68,31,155,31,181,31,93,31,205,31,47,31,47,30,47,29,247,31,119,31,185,31,167,31,101,31,101,30,61,31,168,31,168,30,174,31,45,31,45,30,45,29,45,28,28,31,71,31,4,31,160,31,160,30,120,31,155,31,231,31,251,31,77,31,95,31,161,31,49,31,9,31,156,31,48,31,39,31,131,31,68,31,197,31,158,31,127,31,177,31,209,31,103,31,159,31,229,31,148,31,148,30,190,31,177,31,51,31,51,30,218,31,240,31,16,31,16,30,16,29,236,31,236,30,113,31,209,31,209,30,209,29,209,28,209,27,78,31,75,31,246,31,124,31,202,31,248,31,201,31,201,30,201,29,248,31,152,31,29,31,202,31,54,31,54,30,222,31,48,31,7,31,144,31,108,31,45,31,75,31,194,31,85,31,220,31,94,31,74,31,205,31,53,31,213,31,172,31,162,31,51,31,171,31,208,31,4,31,13,31,13,30,33,31,40,31,91,31,136,31,89,31,45,31,253,31,197,31,230,31,5,31,5,30,5,29,209,31,242,31,242,30,83,31,99,31,99,30,37,31,191,31,191,30,185,31,185,30,185,29,167,31,235,31,34,31,84,31,48,31,25,31,25,30,21,31,218,31,209,31,19,31,79,31,109,31,240,31,70,31,57,31,44,31,11,31,195,31,195,30,195,29,131,31,131,30,131,29,123,31,123,30,123,29,172,31,230,31,248,31,36,31,245,31,245,30,60,31,46,31,19,31,28,31,154,31,154,30,225,31,225,30,167,31,167,30,236,31,49,31,49,30,207,31,207,30,207,29,78,31,189,31,25,31,140,31,167,31,213,31,119,31,146,31,228,31,152,31,152,30,122,31,12,31,223,31,223,30,223,29,223,28,223,27,208,31,208,30,208,29,71,31,71,30,92,31,92,30,92,29,161,31,67,31,63,31,70,31,70,30,79,31,180,31,180,30,178,31,59,31,49,31,136,31,34,31,81,31,51,31,217,31,219,31,51,31,51,30,79,31,191,31,191,30,191,29,72,31,67,31,85,31,105,31,253,31,121,31,78,31,78,30,66,31,253,31,106,31,106,30,157,31,192,31,192,30,192,29,40,31,40,30,40,29,173,31,175,31,221,31,221,30,138,31,177,31,204,31,60,31,237,31,138,31,153,31,108,31,97,31,142,31,89,31,101,31,212,31,126,31,185,31,133,31,117,31,66,31,25,31,11,31,11,30,223,31,165,31,165,30,165,29,78,31,111,31,111,30,85,31,224,31,8,31,60,31,60,30,226,31,45,31,45,30,233,31,36,31,58,31,234,31,233,31,233,30,151,31,131,31,191,31,191,30,191,29,191,28,230,31,86,31,86,30,107,31,107,30,107,29,58,31,234,31,93,31,145,31,152,31,115,31,224,31,200,31,202,31,202,30,113,31,243,31,192,31,192,30,96,31,143,31,143,30,184,31,200,31,200,30,242,31,167,31,77,31,40,31,40,30,187,31,109,31,125,31,83,31,100,31,4,31,211,31,42,31,42,30,173,31,173,30,6,31,68,31,1,31,78,31,246,31,246,30,140,31,140,30,25,31,25,30,9,31,37,31,175,31,141,31,164,31,164,30,193,31,132,31,132,30,132,29,207,31,83,31,83,30,76,31,76,30,220,31,220,30,168,31,168,30,242,31,15,31,202,31,50,31,226,31,38,31,126,31,202,31,90,31,25,31,182,31,149,31,149,30,47,31,153,31,186,31,252,31,30,31,214,31,214,30,198,31,42,31,42,30,177,31,235,31,116,31,116,30,144,31,98,31,98,30,167,31,167,30,33,31,159,31,119,31,176,31,182,31,182,30,182,29,182,28,182,27,186,31,186,30,60,31,67,31,189,31,148,31,5,31,186,31,237,31,238,31,238,30,154,31,135,31,212,31,142,31,129,31,203,31,160,31,160,30,59,31,203,31,51,31,73,31,46,31,218,31,225,31,181,31,239,31,45,31,37,31,124,31,124,30,180,31,196,31,233,31,11,31,197,31,199,31,100,31,100,31,17,31,43,31,134,31,253,31,49,31,136,31,174,31,208,31,119,31,119,30,119,29,86,31,129,31,175,31,103,31,90,31,90,30,232,31,232,30,244,31,133,31,42,31,64,31,232,31,93,31,3,31,155,31,101,31,13,31,98,31,98,30,131,31,29,31,8,31,8,30,66,31,99,31,189,31,44,31,74,31,230,31,184,31,198,31,145,31,143,31,103,31,235,31,191,31,188,31,99,31,75,31,75,30,83,31,83,30,109,31,254,31,112,31,145,31,145,30,233,31,172,31,92,31,7,31,205,31,205,30,205,29,246,31,59,31,90,31,87,31,251,31,156,31,59,31,208,31,208,30,106,31,100,31,24,31,254,31,223,31,76,31,3,31,203,31,154,31,12,31,209,31,238,31,96,31,96,30,192,31,23,31,23,30,53,31,53,30,140,31,30,31,9,31,183,31,29,31,231,31,72,31,133,31,186,31,190,31,190,30,220,31,220,30,220,29,172,31,140,31,246,31,99,31,151,31,247,31,247,30,212,31,167,31,192,31,120,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
