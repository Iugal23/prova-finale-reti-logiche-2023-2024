-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_104 is
end project_tb_104;

architecture project_tb_arch_104 of project_tb_104 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 611;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (247,0,0,0,0,0,81,0,50,0,46,0,201,0,61,0,0,0,226,0,118,0,198,0,147,0,0,0,0,0,98,0,173,0,157,0,160,0,200,0,241,0,0,0,0,0,0,0,212,0,129,0,78,0,62,0,153,0,52,0,0,0,53,0,132,0,1,0,226,0,155,0,137,0,15,0,0,0,63,0,161,0,60,0,95,0,235,0,215,0,205,0,39,0,0,0,89,0,36,0,149,0,17,0,154,0,193,0,33,0,118,0,0,0,41,0,254,0,0,0,54,0,219,0,114,0,244,0,3,0,153,0,253,0,25,0,200,0,102,0,0,0,109,0,32,0,162,0,228,0,18,0,214,0,116,0,192,0,214,0,57,0,0,0,63,0,0,0,21,0,0,0,109,0,30,0,245,0,0,0,159,0,49,0,247,0,152,0,65,0,245,0,0,0,242,0,96,0,42,0,189,0,114,0,0,0,222,0,247,0,0,0,143,0,159,0,22,0,114,0,0,0,100,0,84,0,22,0,0,0,131,0,189,0,137,0,56,0,251,0,3,0,223,0,176,0,21,0,185,0,0,0,187,0,141,0,167,0,128,0,249,0,0,0,199,0,162,0,191,0,131,0,38,0,116,0,0,0,0,0,253,0,108,0,13,0,90,0,92,0,198,0,0,0,217,0,100,0,174,0,0,0,11,0,217,0,130,0,244,0,172,0,0,0,0,0,191,0,0,0,26,0,201,0,116,0,0,0,150,0,253,0,204,0,232,0,0,0,142,0,97,0,160,0,98,0,6,0,237,0,0,0,221,0,0,0,172,0,60,0,66,0,146,0,0,0,0,0,115,0,247,0,0,0,0,0,98,0,185,0,117,0,58,0,0,0,177,0,185,0,179,0,170,0,254,0,254,0,0,0,96,0,89,0,0,0,67,0,216,0,73,0,251,0,34,0,76,0,226,0,76,0,210,0,0,0,128,0,12,0,63,0,0,0,78,0,227,0,87,0,1,0,99,0,174,0,30,0,0,0,255,0,194,0,18,0,134,0,101,0,132,0,251,0,253,0,223,0,232,0,65,0,138,0,30,0,230,0,0,0,130,0,180,0,69,0,255,0,66,0,185,0,180,0,226,0,0,0,0,0,0,0,0,0,101,0,0,0,165,0,74,0,219,0,21,0,38,0,234,0,213,0,24,0,244,0,188,0,63,0,0,0,0,0,70,0,0,0,0,0,161,0,28,0,107,0,103,0,0,0,118,0,0,0,50,0,56,0,171,0,48,0,0,0,228,0,113,0,142,0,252,0,76,0,163,0,203,0,141,0,92,0,130,0,59,0,242,0,138,0,22,0,155,0,0,0,229,0,60,0,0,0,69,0,197,0,58,0,221,0,0,0,183,0,79,0,189,0,238,0,131,0,127,0,108,0,244,0,214,0,99,0,169,0,129,0,10,0,251,0,38,0,0,0,69,0,0,0,0,0,0,0,198,0,83,0,57,0,77,0,75,0,224,0,0,0,0,0,133,0,0,0,225,0,0,0,208,0,53,0,115,0,111,0,68,0,99,0,215,0,123,0,234,0,0,0,201,0,234,0,0,0,171,0,186,0,122,0,0,0,117,0,101,0,204,0,29,0,31,0,210,0,39,0,137,0,47,0,8,0,123,0,190,0,155,0,41,0,213,0,87,0,0,0,99,0,0,0,0,0,90,0,74,0,253,0,217,0,0,0,199,0,244,0,194,0,148,0,197,0,5,0,0,0,110,0,23,0,89,0,0,0,79,0,222,0,148,0,72,0,12,0,6,0,0,0,246,0,0,0,115,0,242,0,12,0,241,0,108,0,49,0,103,0,169,0,93,0,207,0,39,0,226,0,0,0,59,0,143,0,172,0,28,0,0,0,171,0,63,0,225,0,0,0,204,0,72,0,202,0,54,0,71,0,131,0,238,0,0,0,122,0,157,0,239,0,16,0,100,0,0,0,30,0,174,0,2,0,164,0,175,0,191,0,0,0,143,0,244,0,118,0,253,0,209,0,76,0,182,0,222,0,219,0,72,0,45,0,0,0,217,0,2,0,213,0,0,0,52,0,0,0,16,0,0,0,117,0,154,0,0,0,169,0,13,0,220,0,143,0,186,0,43,0,12,0,104,0,0,0,0,0,35,0,0,0,78,0,70,0,100,0,0,0,7,0,89,0,0,0,226,0,62,0,0,0,243,0,0,0,218,0,112,0,0,0,116,0,124,0,229,0,64,0,0,0,248,0,0,0,185,0,0,0,0,0,0,0,84,0,238,0,187,0,127,0,0,0,244,0,98,0,221,0,158,0,197,0,0,0,0,0,132,0,0,0,120,0,0,0,0,0,0,0,4,0,182,0,13,0,2,0,0,0,15,0,0,0,33,0,24,0,74,0,233,0,114,0,55,0,46,0,108,0,189,0,128,0,0,0,132,0,116,0,96,0,0,0,80,0,250,0,244,0,17,0,243,0,106,0,0,0,0,0,102,0,186,0,0,0,0,0,158,0,25,0,204,0,106,0,0,0,222,0,8,0,20,0,81,0,8,0,0,0,183,0,40,0,170,0,49,0,0,0,207,0,0,0,31,0,149,0,202,0,92,0,0,0,99,0,76,0,21,0,197,0,0,0,0,0,0,0,209,0,103,0,120,0,108,0,87,0,0,0,159,0,20,0,0,0,13,0,198,0,166,0,216,0,92,0,49,0,0,0,0,0,31,0,143,0,0,0,0,0,119,0,170,0,220,0,112,0);
signal scenario_full  : scenario_type := (247,31,247,30,247,29,81,31,50,31,46,31,201,31,61,31,61,30,226,31,118,31,198,31,147,31,147,30,147,29,98,31,173,31,157,31,160,31,200,31,241,31,241,30,241,29,241,28,212,31,129,31,78,31,62,31,153,31,52,31,52,30,53,31,132,31,1,31,226,31,155,31,137,31,15,31,15,30,63,31,161,31,60,31,95,31,235,31,215,31,205,31,39,31,39,30,89,31,36,31,149,31,17,31,154,31,193,31,33,31,118,31,118,30,41,31,254,31,254,30,54,31,219,31,114,31,244,31,3,31,153,31,253,31,25,31,200,31,102,31,102,30,109,31,32,31,162,31,228,31,18,31,214,31,116,31,192,31,214,31,57,31,57,30,63,31,63,30,21,31,21,30,109,31,30,31,245,31,245,30,159,31,49,31,247,31,152,31,65,31,245,31,245,30,242,31,96,31,42,31,189,31,114,31,114,30,222,31,247,31,247,30,143,31,159,31,22,31,114,31,114,30,100,31,84,31,22,31,22,30,131,31,189,31,137,31,56,31,251,31,3,31,223,31,176,31,21,31,185,31,185,30,187,31,141,31,167,31,128,31,249,31,249,30,199,31,162,31,191,31,131,31,38,31,116,31,116,30,116,29,253,31,108,31,13,31,90,31,92,31,198,31,198,30,217,31,100,31,174,31,174,30,11,31,217,31,130,31,244,31,172,31,172,30,172,29,191,31,191,30,26,31,201,31,116,31,116,30,150,31,253,31,204,31,232,31,232,30,142,31,97,31,160,31,98,31,6,31,237,31,237,30,221,31,221,30,172,31,60,31,66,31,146,31,146,30,146,29,115,31,247,31,247,30,247,29,98,31,185,31,117,31,58,31,58,30,177,31,185,31,179,31,170,31,254,31,254,31,254,30,96,31,89,31,89,30,67,31,216,31,73,31,251,31,34,31,76,31,226,31,76,31,210,31,210,30,128,31,12,31,63,31,63,30,78,31,227,31,87,31,1,31,99,31,174,31,30,31,30,30,255,31,194,31,18,31,134,31,101,31,132,31,251,31,253,31,223,31,232,31,65,31,138,31,30,31,230,31,230,30,130,31,180,31,69,31,255,31,66,31,185,31,180,31,226,31,226,30,226,29,226,28,226,27,101,31,101,30,165,31,74,31,219,31,21,31,38,31,234,31,213,31,24,31,244,31,188,31,63,31,63,30,63,29,70,31,70,30,70,29,161,31,28,31,107,31,103,31,103,30,118,31,118,30,50,31,56,31,171,31,48,31,48,30,228,31,113,31,142,31,252,31,76,31,163,31,203,31,141,31,92,31,130,31,59,31,242,31,138,31,22,31,155,31,155,30,229,31,60,31,60,30,69,31,197,31,58,31,221,31,221,30,183,31,79,31,189,31,238,31,131,31,127,31,108,31,244,31,214,31,99,31,169,31,129,31,10,31,251,31,38,31,38,30,69,31,69,30,69,29,69,28,198,31,83,31,57,31,77,31,75,31,224,31,224,30,224,29,133,31,133,30,225,31,225,30,208,31,53,31,115,31,111,31,68,31,99,31,215,31,123,31,234,31,234,30,201,31,234,31,234,30,171,31,186,31,122,31,122,30,117,31,101,31,204,31,29,31,31,31,210,31,39,31,137,31,47,31,8,31,123,31,190,31,155,31,41,31,213,31,87,31,87,30,99,31,99,30,99,29,90,31,74,31,253,31,217,31,217,30,199,31,244,31,194,31,148,31,197,31,5,31,5,30,110,31,23,31,89,31,89,30,79,31,222,31,148,31,72,31,12,31,6,31,6,30,246,31,246,30,115,31,242,31,12,31,241,31,108,31,49,31,103,31,169,31,93,31,207,31,39,31,226,31,226,30,59,31,143,31,172,31,28,31,28,30,171,31,63,31,225,31,225,30,204,31,72,31,202,31,54,31,71,31,131,31,238,31,238,30,122,31,157,31,239,31,16,31,100,31,100,30,30,31,174,31,2,31,164,31,175,31,191,31,191,30,143,31,244,31,118,31,253,31,209,31,76,31,182,31,222,31,219,31,72,31,45,31,45,30,217,31,2,31,213,31,213,30,52,31,52,30,16,31,16,30,117,31,154,31,154,30,169,31,13,31,220,31,143,31,186,31,43,31,12,31,104,31,104,30,104,29,35,31,35,30,78,31,70,31,100,31,100,30,7,31,89,31,89,30,226,31,62,31,62,30,243,31,243,30,218,31,112,31,112,30,116,31,124,31,229,31,64,31,64,30,248,31,248,30,185,31,185,30,185,29,185,28,84,31,238,31,187,31,127,31,127,30,244,31,98,31,221,31,158,31,197,31,197,30,197,29,132,31,132,30,120,31,120,30,120,29,120,28,4,31,182,31,13,31,2,31,2,30,15,31,15,30,33,31,24,31,74,31,233,31,114,31,55,31,46,31,108,31,189,31,128,31,128,30,132,31,116,31,96,31,96,30,80,31,250,31,244,31,17,31,243,31,106,31,106,30,106,29,102,31,186,31,186,30,186,29,158,31,25,31,204,31,106,31,106,30,222,31,8,31,20,31,81,31,8,31,8,30,183,31,40,31,170,31,49,31,49,30,207,31,207,30,31,31,149,31,202,31,92,31,92,30,99,31,76,31,21,31,197,31,197,30,197,29,197,28,209,31,103,31,120,31,108,31,87,31,87,30,159,31,20,31,20,30,13,31,198,31,166,31,216,31,92,31,49,31,49,30,49,29,31,31,143,31,143,30,143,29,119,31,170,31,220,31,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
