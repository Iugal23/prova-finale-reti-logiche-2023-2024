-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_59 is
end project_tb_59;

architecture project_tb_arch_59 of project_tb_59 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 657;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,70,0,76,0,113,0,190,0,0,0,69,0,142,0,13,0,0,0,20,0,204,0,149,0,0,0,71,0,9,0,0,0,89,0,0,0,109,0,38,0,41,0,87,0,164,0,32,0,100,0,240,0,128,0,203,0,134,0,107,0,30,0,117,0,167,0,63,0,226,0,190,0,43,0,0,0,146,0,115,0,129,0,148,0,85,0,0,0,0,0,108,0,0,0,171,0,148,0,184,0,0,0,96,0,69,0,7,0,0,0,23,0,122,0,0,0,56,0,165,0,0,0,169,0,191,0,143,0,203,0,221,0,8,0,239,0,141,0,85,0,130,0,77,0,0,0,45,0,107,0,97,0,55,0,214,0,164,0,12,0,233,0,17,0,205,0,103,0,52,0,242,0,136,0,17,0,164,0,111,0,97,0,160,0,20,0,53,0,0,0,85,0,115,0,71,0,43,0,232,0,212,0,0,0,79,0,159,0,8,0,235,0,0,0,228,0,58,0,25,0,95,0,191,0,72,0,87,0,118,0,0,0,51,0,133,0,127,0,0,0,0,0,41,0,0,0,46,0,74,0,162,0,0,0,32,0,53,0,0,0,109,0,80,0,32,0,228,0,141,0,121,0,222,0,0,0,183,0,219,0,197,0,78,0,35,0,0,0,0,0,113,0,0,0,0,0,140,0,244,0,42,0,0,0,0,0,231,0,243,0,65,0,203,0,199,0,151,0,18,0,121,0,215,0,0,0,143,0,0,0,119,0,10,0,0,0,189,0,0,0,18,0,44,0,153,0,0,0,113,0,48,0,167,0,203,0,0,0,12,0,227,0,208,0,250,0,20,0,167,0,45,0,64,0,125,0,11,0,23,0,0,0,180,0,0,0,203,0,44,0,111,0,244,0,125,0,17,0,145,0,92,0,1,0,207,0,48,0,0,0,52,0,207,0,99,0,40,0,35,0,184,0,0,0,51,0,0,0,154,0,78,0,246,0,0,0,245,0,23,0,135,0,185,0,125,0,68,0,0,0,106,0,191,0,0,0,242,0,0,0,0,0,164,0,0,0,221,0,225,0,53,0,0,0,0,0,81,0,99,0,71,0,86,0,0,0,59,0,0,0,16,0,104,0,52,0,0,0,254,0,63,0,83,0,207,0,116,0,0,0,0,0,21,0,0,0,3,0,9,0,64,0,0,0,74,0,238,0,0,0,68,0,6,0,31,0,41,0,139,0,0,0,241,0,44,0,110,0,133,0,0,0,184,0,72,0,121,0,103,0,250,0,0,0,0,0,92,0,71,0,82,0,254,0,0,0,192,0,252,0,217,0,138,0,0,0,142,0,120,0,49,0,105,0,0,0,120,0,192,0,0,0,179,0,111,0,195,0,125,0,86,0,0,0,213,0,228,0,235,0,50,0,0,0,23,0,64,0,186,0,219,0,152,0,237,0,120,0,31,0,120,0,0,0,154,0,254,0,0,0,220,0,113,0,0,0,163,0,85,0,56,0,102,0,93,0,109,0,75,0,247,0,97,0,0,0,56,0,94,0,133,0,0,0,162,0,0,0,23,0,0,0,56,0,195,0,152,0,207,0,31,0,0,0,157,0,50,0,130,0,205,0,247,0,99,0,2,0,215,0,0,0,0,0,138,0,126,0,0,0,0,0,77,0,247,0,100,0,53,0,0,0,15,0,98,0,72,0,189,0,212,0,226,0,0,0,137,0,31,0,178,0,195,0,16,0,45,0,0,0,192,0,83,0,144,0,232,0,71,0,84,0,140,0,79,0,0,0,68,0,0,0,14,0,40,0,94,0,93,0,0,0,240,0,199,0,112,0,165,0,176,0,80,0,180,0,0,0,0,0,0,0,215,0,0,0,188,0,93,0,131,0,156,0,105,0,0,0,67,0,183,0,94,0,175,0,0,0,0,0,0,0,216,0,145,0,0,0,47,0,53,0,0,0,0,0,198,0,0,0,10,0,69,0,51,0,223,0,73,0,195,0,93,0,60,0,168,0,124,0,84,0,0,0,0,0,251,0,0,0,115,0,34,0,54,0,50,0,88,0,1,0,159,0,143,0,145,0,49,0,121,0,187,0,174,0,80,0,0,0,52,0,97,0,129,0,0,0,37,0,184,0,0,0,0,0,21,0,223,0,186,0,90,0,0,0,0,0,122,0,15,0,118,0,15,0,218,0,0,0,125,0,151,0,146,0,132,0,89,0,78,0,0,0,153,0,122,0,151,0,0,0,185,0,181,0,141,0,144,0,63,0,0,0,200,0,0,0,41,0,134,0,0,0,191,0,236,0,188,0,44,0,224,0,113,0,227,0,0,0,93,0,98,0,34,0,0,0,100,0,98,0,0,0,0,0,36,0,155,0,48,0,234,0,141,0,0,0,247,0,251,0,0,0,117,0,135,0,94,0,192,0,36,0,0,0,0,0,174,0,15,0,190,0,0,0,91,0,0,0,1,0,0,0,197,0,102,0,94,0,156,0,165,0,76,0,126,0,59,0,47,0,72,0,158,0,175,0,112,0,228,0,133,0,0,0,36,0,142,0,155,0,158,0,197,0,207,0,103,0,191,0,125,0,0,0,179,0,0,0,79,0,77,0,53,0,38,0,234,0,155,0,56,0,78,0,49,0,23,0,93,0,77,0,164,0,118,0,240,0,153,0,0,0,0,0,27,0,243,0,0,0,147,0,200,0,34,0,254,0,127,0,58,0,0,0,177,0,1,0,224,0,239,0,37,0,0,0,0,0,75,0,83,0,242,0,186,0,86,0,220,0,92,0,151,0,222,0,0,0,223,0,26,0,231,0,137,0,26,0,107,0,0,0,10,0,54,0,161,0,236,0,13,0,70,0,47,0,142,0,36,0,122,0,0,0,0,0,122,0,161,0,57,0,213,0,128,0,216,0,30,0,87,0,227,0,0,0,0,0,16,0,42,0,92,0,64,0,245,0,16,0);
signal scenario_full  : scenario_type := (0,0,70,31,76,31,113,31,190,31,190,30,69,31,142,31,13,31,13,30,20,31,204,31,149,31,149,30,71,31,9,31,9,30,89,31,89,30,109,31,38,31,41,31,87,31,164,31,32,31,100,31,240,31,128,31,203,31,134,31,107,31,30,31,117,31,167,31,63,31,226,31,190,31,43,31,43,30,146,31,115,31,129,31,148,31,85,31,85,30,85,29,108,31,108,30,171,31,148,31,184,31,184,30,96,31,69,31,7,31,7,30,23,31,122,31,122,30,56,31,165,31,165,30,169,31,191,31,143,31,203,31,221,31,8,31,239,31,141,31,85,31,130,31,77,31,77,30,45,31,107,31,97,31,55,31,214,31,164,31,12,31,233,31,17,31,205,31,103,31,52,31,242,31,136,31,17,31,164,31,111,31,97,31,160,31,20,31,53,31,53,30,85,31,115,31,71,31,43,31,232,31,212,31,212,30,79,31,159,31,8,31,235,31,235,30,228,31,58,31,25,31,95,31,191,31,72,31,87,31,118,31,118,30,51,31,133,31,127,31,127,30,127,29,41,31,41,30,46,31,74,31,162,31,162,30,32,31,53,31,53,30,109,31,80,31,32,31,228,31,141,31,121,31,222,31,222,30,183,31,219,31,197,31,78,31,35,31,35,30,35,29,113,31,113,30,113,29,140,31,244,31,42,31,42,30,42,29,231,31,243,31,65,31,203,31,199,31,151,31,18,31,121,31,215,31,215,30,143,31,143,30,119,31,10,31,10,30,189,31,189,30,18,31,44,31,153,31,153,30,113,31,48,31,167,31,203,31,203,30,12,31,227,31,208,31,250,31,20,31,167,31,45,31,64,31,125,31,11,31,23,31,23,30,180,31,180,30,203,31,44,31,111,31,244,31,125,31,17,31,145,31,92,31,1,31,207,31,48,31,48,30,52,31,207,31,99,31,40,31,35,31,184,31,184,30,51,31,51,30,154,31,78,31,246,31,246,30,245,31,23,31,135,31,185,31,125,31,68,31,68,30,106,31,191,31,191,30,242,31,242,30,242,29,164,31,164,30,221,31,225,31,53,31,53,30,53,29,81,31,99,31,71,31,86,31,86,30,59,31,59,30,16,31,104,31,52,31,52,30,254,31,63,31,83,31,207,31,116,31,116,30,116,29,21,31,21,30,3,31,9,31,64,31,64,30,74,31,238,31,238,30,68,31,6,31,31,31,41,31,139,31,139,30,241,31,44,31,110,31,133,31,133,30,184,31,72,31,121,31,103,31,250,31,250,30,250,29,92,31,71,31,82,31,254,31,254,30,192,31,252,31,217,31,138,31,138,30,142,31,120,31,49,31,105,31,105,30,120,31,192,31,192,30,179,31,111,31,195,31,125,31,86,31,86,30,213,31,228,31,235,31,50,31,50,30,23,31,64,31,186,31,219,31,152,31,237,31,120,31,31,31,120,31,120,30,154,31,254,31,254,30,220,31,113,31,113,30,163,31,85,31,56,31,102,31,93,31,109,31,75,31,247,31,97,31,97,30,56,31,94,31,133,31,133,30,162,31,162,30,23,31,23,30,56,31,195,31,152,31,207,31,31,31,31,30,157,31,50,31,130,31,205,31,247,31,99,31,2,31,215,31,215,30,215,29,138,31,126,31,126,30,126,29,77,31,247,31,100,31,53,31,53,30,15,31,98,31,72,31,189,31,212,31,226,31,226,30,137,31,31,31,178,31,195,31,16,31,45,31,45,30,192,31,83,31,144,31,232,31,71,31,84,31,140,31,79,31,79,30,68,31,68,30,14,31,40,31,94,31,93,31,93,30,240,31,199,31,112,31,165,31,176,31,80,31,180,31,180,30,180,29,180,28,215,31,215,30,188,31,93,31,131,31,156,31,105,31,105,30,67,31,183,31,94,31,175,31,175,30,175,29,175,28,216,31,145,31,145,30,47,31,53,31,53,30,53,29,198,31,198,30,10,31,69,31,51,31,223,31,73,31,195,31,93,31,60,31,168,31,124,31,84,31,84,30,84,29,251,31,251,30,115,31,34,31,54,31,50,31,88,31,1,31,159,31,143,31,145,31,49,31,121,31,187,31,174,31,80,31,80,30,52,31,97,31,129,31,129,30,37,31,184,31,184,30,184,29,21,31,223,31,186,31,90,31,90,30,90,29,122,31,15,31,118,31,15,31,218,31,218,30,125,31,151,31,146,31,132,31,89,31,78,31,78,30,153,31,122,31,151,31,151,30,185,31,181,31,141,31,144,31,63,31,63,30,200,31,200,30,41,31,134,31,134,30,191,31,236,31,188,31,44,31,224,31,113,31,227,31,227,30,93,31,98,31,34,31,34,30,100,31,98,31,98,30,98,29,36,31,155,31,48,31,234,31,141,31,141,30,247,31,251,31,251,30,117,31,135,31,94,31,192,31,36,31,36,30,36,29,174,31,15,31,190,31,190,30,91,31,91,30,1,31,1,30,197,31,102,31,94,31,156,31,165,31,76,31,126,31,59,31,47,31,72,31,158,31,175,31,112,31,228,31,133,31,133,30,36,31,142,31,155,31,158,31,197,31,207,31,103,31,191,31,125,31,125,30,179,31,179,30,79,31,77,31,53,31,38,31,234,31,155,31,56,31,78,31,49,31,23,31,93,31,77,31,164,31,118,31,240,31,153,31,153,30,153,29,27,31,243,31,243,30,147,31,200,31,34,31,254,31,127,31,58,31,58,30,177,31,1,31,224,31,239,31,37,31,37,30,37,29,75,31,83,31,242,31,186,31,86,31,220,31,92,31,151,31,222,31,222,30,223,31,26,31,231,31,137,31,26,31,107,31,107,30,10,31,54,31,161,31,236,31,13,31,70,31,47,31,142,31,36,31,122,31,122,30,122,29,122,31,161,31,57,31,213,31,128,31,216,31,30,31,87,31,227,31,227,30,227,29,16,31,42,31,92,31,64,31,245,31,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
