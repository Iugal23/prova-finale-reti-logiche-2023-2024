-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 466;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (110,0,69,0,0,0,19,0,179,0,0,0,135,0,0,0,97,0,0,0,17,0,32,0,101,0,222,0,0,0,72,0,61,0,0,0,88,0,0,0,138,0,106,0,115,0,0,0,0,0,189,0,38,0,214,0,92,0,113,0,0,0,13,0,213,0,80,0,255,0,243,0,20,0,46,0,0,0,46,0,232,0,0,0,184,0,32,0,110,0,0,0,193,0,255,0,0,0,0,0,60,0,75,0,191,0,73,0,0,0,88,0,9,0,43,0,126,0,206,0,63,0,188,0,0,0,0,0,0,0,217,0,145,0,0,0,236,0,11,0,141,0,232,0,0,0,8,0,210,0,181,0,110,0,232,0,147,0,0,0,85,0,37,0,0,0,0,0,18,0,7,0,26,0,82,0,125,0,205,0,18,0,164,0,74,0,51,0,59,0,0,0,113,0,0,0,110,0,208,0,0,0,217,0,84,0,34,0,139,0,59,0,0,0,87,0,0,0,13,0,0,0,0,0,234,0,38,0,90,0,0,0,7,0,0,0,0,0,104,0,0,0,214,0,183,0,0,0,119,0,86,0,0,0,252,0,236,0,78,0,168,0,249,0,55,0,0,0,234,0,218,0,167,0,246,0,187,0,161,0,94,0,194,0,244,0,0,0,220,0,0,0,116,0,25,0,102,0,194,0,162,0,84,0,208,0,192,0,0,0,0,0,158,0,80,0,244,0,210,0,121,0,149,0,36,0,32,0,21,0,0,0,179,0,0,0,0,0,0,0,15,0,0,0,155,0,0,0,223,0,139,0,230,0,81,0,197,0,114,0,17,0,3,0,151,0,105,0,5,0,97,0,43,0,111,0,71,0,189,0,2,0,188,0,56,0,155,0,194,0,76,0,150,0,22,0,226,0,0,0,212,0,10,0,69,0,0,0,142,0,245,0,177,0,189,0,29,0,132,0,103,0,204,0,30,0,27,0,227,0,0,0,70,0,0,0,181,0,103,0,190,0,0,0,168,0,0,0,0,0,92,0,28,0,7,0,188,0,102,0,239,0,188,0,0,0,73,0,0,0,105,0,129,0,67,0,70,0,11,0,200,0,170,0,169,0,23,0,0,0,183,0,86,0,86,0,147,0,0,0,165,0,209,0,0,0,96,0,55,0,117,0,120,0,0,0,83,0,237,0,187,0,239,0,71,0,216,0,207,0,0,0,99,0,242,0,156,0,156,0,120,0,90,0,253,0,0,0,0,0,223,0,211,0,0,0,193,0,244,0,182,0,5,0,255,0,187,0,246,0,255,0,20,0,0,0,37,0,225,0,250,0,141,0,207,0,248,0,0,0,0,0,207,0,230,0,172,0,44,0,68,0,62,0,63,0,194,0,2,0,34,0,38,0,254,0,82,0,23,0,148,0,140,0,211,0,225,0,0,0,55,0,220,0,191,0,102,0,0,0,0,0,0,0,168,0,67,0,67,0,87,0,73,0,188,0,228,0,180,0,192,0,5,0,44,0,0,0,211,0,127,0,80,0,191,0,202,0,239,0,214,0,73,0,0,0,130,0,0,0,229,0,121,0,89,0,131,0,0,0,170,0,0,0,84,0,219,0,7,0,143,0,216,0,57,0,167,0,198,0,77,0,18,0,77,0,255,0,93,0,109,0,76,0,0,0,226,0,44,0,238,0,0,0,60,0,253,0,104,0,0,0,2,0,110,0,0,0,236,0,228,0,43,0,0,0,148,0,70,0,0,0,126,0,169,0,50,0,51,0,98,0,220,0,95,0,57,0,75,0,10,0,123,0,0,0,79,0,210,0,213,0,48,0,131,0,0,0,55,0,44,0,96,0,0,0,141,0,40,0,69,0,25,0,195,0,44,0,84,0,158,0,231,0,0,0,6,0,0,0,8,0,121,0,239,0,99,0,235,0,242,0,209,0,220,0,141,0,0,0,109,0,83,0,102,0,201,0,107,0,1,0,108,0,165,0,183,0,253,0,0,0,0,0,78,0,123,0,140,0,121,0,212,0,55,0,0,0,0,0,197,0,142,0,181,0,137,0,212,0,253,0,173,0,249,0,251,0,0,0,245,0,58,0,0,0,225,0,237,0,0,0);
signal scenario_full  : scenario_type := (110,31,69,31,69,30,19,31,179,31,179,30,135,31,135,30,97,31,97,30,17,31,32,31,101,31,222,31,222,30,72,31,61,31,61,30,88,31,88,30,138,31,106,31,115,31,115,30,115,29,189,31,38,31,214,31,92,31,113,31,113,30,13,31,213,31,80,31,255,31,243,31,20,31,46,31,46,30,46,31,232,31,232,30,184,31,32,31,110,31,110,30,193,31,255,31,255,30,255,29,60,31,75,31,191,31,73,31,73,30,88,31,9,31,43,31,126,31,206,31,63,31,188,31,188,30,188,29,188,28,217,31,145,31,145,30,236,31,11,31,141,31,232,31,232,30,8,31,210,31,181,31,110,31,232,31,147,31,147,30,85,31,37,31,37,30,37,29,18,31,7,31,26,31,82,31,125,31,205,31,18,31,164,31,74,31,51,31,59,31,59,30,113,31,113,30,110,31,208,31,208,30,217,31,84,31,34,31,139,31,59,31,59,30,87,31,87,30,13,31,13,30,13,29,234,31,38,31,90,31,90,30,7,31,7,30,7,29,104,31,104,30,214,31,183,31,183,30,119,31,86,31,86,30,252,31,236,31,78,31,168,31,249,31,55,31,55,30,234,31,218,31,167,31,246,31,187,31,161,31,94,31,194,31,244,31,244,30,220,31,220,30,116,31,25,31,102,31,194,31,162,31,84,31,208,31,192,31,192,30,192,29,158,31,80,31,244,31,210,31,121,31,149,31,36,31,32,31,21,31,21,30,179,31,179,30,179,29,179,28,15,31,15,30,155,31,155,30,223,31,139,31,230,31,81,31,197,31,114,31,17,31,3,31,151,31,105,31,5,31,97,31,43,31,111,31,71,31,189,31,2,31,188,31,56,31,155,31,194,31,76,31,150,31,22,31,226,31,226,30,212,31,10,31,69,31,69,30,142,31,245,31,177,31,189,31,29,31,132,31,103,31,204,31,30,31,27,31,227,31,227,30,70,31,70,30,181,31,103,31,190,31,190,30,168,31,168,30,168,29,92,31,28,31,7,31,188,31,102,31,239,31,188,31,188,30,73,31,73,30,105,31,129,31,67,31,70,31,11,31,200,31,170,31,169,31,23,31,23,30,183,31,86,31,86,31,147,31,147,30,165,31,209,31,209,30,96,31,55,31,117,31,120,31,120,30,83,31,237,31,187,31,239,31,71,31,216,31,207,31,207,30,99,31,242,31,156,31,156,31,120,31,90,31,253,31,253,30,253,29,223,31,211,31,211,30,193,31,244,31,182,31,5,31,255,31,187,31,246,31,255,31,20,31,20,30,37,31,225,31,250,31,141,31,207,31,248,31,248,30,248,29,207,31,230,31,172,31,44,31,68,31,62,31,63,31,194,31,2,31,34,31,38,31,254,31,82,31,23,31,148,31,140,31,211,31,225,31,225,30,55,31,220,31,191,31,102,31,102,30,102,29,102,28,168,31,67,31,67,31,87,31,73,31,188,31,228,31,180,31,192,31,5,31,44,31,44,30,211,31,127,31,80,31,191,31,202,31,239,31,214,31,73,31,73,30,130,31,130,30,229,31,121,31,89,31,131,31,131,30,170,31,170,30,84,31,219,31,7,31,143,31,216,31,57,31,167,31,198,31,77,31,18,31,77,31,255,31,93,31,109,31,76,31,76,30,226,31,44,31,238,31,238,30,60,31,253,31,104,31,104,30,2,31,110,31,110,30,236,31,228,31,43,31,43,30,148,31,70,31,70,30,126,31,169,31,50,31,51,31,98,31,220,31,95,31,57,31,75,31,10,31,123,31,123,30,79,31,210,31,213,31,48,31,131,31,131,30,55,31,44,31,96,31,96,30,141,31,40,31,69,31,25,31,195,31,44,31,84,31,158,31,231,31,231,30,6,31,6,30,8,31,121,31,239,31,99,31,235,31,242,31,209,31,220,31,141,31,141,30,109,31,83,31,102,31,201,31,107,31,1,31,108,31,165,31,183,31,253,31,253,30,253,29,78,31,123,31,140,31,121,31,212,31,55,31,55,30,55,29,197,31,142,31,181,31,137,31,212,31,253,31,173,31,249,31,251,31,251,30,245,31,58,31,58,30,225,31,237,31,237,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
