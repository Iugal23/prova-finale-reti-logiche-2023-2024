-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_394 is
end project_tb_394;

architecture project_tb_arch_394 of project_tb_394 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 332;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,2,0,83,0,134,0,152,0,0,0,12,0,45,0,5,0,161,0,181,0,25,0,186,0,100,0,55,0,250,0,12,0,129,0,0,0,11,0,82,0,1,0,245,0,29,0,202,0,162,0,119,0,34,0,78,0,151,0,57,0,0,0,149,0,77,0,0,0,0,0,145,0,149,0,203,0,0,0,154,0,183,0,250,0,49,0,85,0,221,0,6,0,160,0,0,0,171,0,0,0,29,0,0,0,85,0,33,0,156,0,0,0,57,0,227,0,92,0,41,0,2,0,31,0,242,0,71,0,0,0,14,0,88,0,16,0,255,0,236,0,50,0,78,0,153,0,209,0,166,0,1,0,16,0,60,0,73,0,29,0,27,0,173,0,0,0,183,0,96,0,12,0,131,0,52,0,0,0,226,0,2,0,0,0,0,0,0,0,64,0,55,0,2,0,0,0,0,0,187,0,0,0,65,0,151,0,200,0,107,0,98,0,0,0,129,0,193,0,206,0,2,0,82,0,79,0,152,0,225,0,111,0,120,0,130,0,75,0,140,0,107,0,89,0,167,0,49,0,0,0,93,0,151,0,196,0,1,0,237,0,57,0,128,0,226,0,0,0,33,0,0,0,7,0,178,0,115,0,38,0,0,0,188,0,249,0,185,0,75,0,216,0,161,0,93,0,178,0,56,0,102,0,7,0,217,0,42,0,175,0,232,0,149,0,162,0,40,0,213,0,106,0,215,0,143,0,0,0,226,0,36,0,116,0,102,0,136,0,242,0,18,0,241,0,153,0,87,0,255,0,0,0,32,0,205,0,0,0,187,0,110,0,254,0,0,0,0,0,0,0,4,0,238,0,65,0,88,0,0,0,0,0,183,0,35,0,90,0,0,0,109,0,154,0,196,0,154,0,0,0,0,0,208,0,220,0,212,0,147,0,153,0,9,0,131,0,28,0,181,0,247,0,50,0,0,0,0,0,118,0,69,0,64,0,181,0,110,0,34,0,91,0,0,0,76,0,151,0,0,0,179,0,13,0,5,0,0,0,46,0,0,0,103,0,197,0,0,0,207,0,80,0,0,0,144,0,113,0,15,0,7,0,77,0,210,0,0,0,182,0,245,0,0,0,0,0,24,0,0,0,0,0,48,0,184,0,188,0,148,0,0,0,249,0,95,0,113,0,153,0,0,0,81,0,53,0,214,0,0,0,110,0,0,0,0,0,37,0,216,0,142,0,223,0,0,0,123,0,114,0,114,0,213,0,81,0,190,0,0,0,231,0,147,0,240,0,157,0,0,0,255,0,0,0,127,0,18,0,209,0,165,0,252,0,149,0,0,0,49,0,0,0,177,0,11,0,199,0,59,0,246,0,159,0,0,0,147,0,96,0,34,0,0,0,34,0,109,0,121,0,150,0,135,0,2,0,136,0,27,0,184,0,54,0,123,0,36,0,0,0,172,0,101,0,148,0,231,0,129,0,125,0,108,0,186,0,7,0,46,0,123,0);
signal scenario_full  : scenario_type := (0,0,2,31,83,31,134,31,152,31,152,30,12,31,45,31,5,31,161,31,181,31,25,31,186,31,100,31,55,31,250,31,12,31,129,31,129,30,11,31,82,31,1,31,245,31,29,31,202,31,162,31,119,31,34,31,78,31,151,31,57,31,57,30,149,31,77,31,77,30,77,29,145,31,149,31,203,31,203,30,154,31,183,31,250,31,49,31,85,31,221,31,6,31,160,31,160,30,171,31,171,30,29,31,29,30,85,31,33,31,156,31,156,30,57,31,227,31,92,31,41,31,2,31,31,31,242,31,71,31,71,30,14,31,88,31,16,31,255,31,236,31,50,31,78,31,153,31,209,31,166,31,1,31,16,31,60,31,73,31,29,31,27,31,173,31,173,30,183,31,96,31,12,31,131,31,52,31,52,30,226,31,2,31,2,30,2,29,2,28,64,31,55,31,2,31,2,30,2,29,187,31,187,30,65,31,151,31,200,31,107,31,98,31,98,30,129,31,193,31,206,31,2,31,82,31,79,31,152,31,225,31,111,31,120,31,130,31,75,31,140,31,107,31,89,31,167,31,49,31,49,30,93,31,151,31,196,31,1,31,237,31,57,31,128,31,226,31,226,30,33,31,33,30,7,31,178,31,115,31,38,31,38,30,188,31,249,31,185,31,75,31,216,31,161,31,93,31,178,31,56,31,102,31,7,31,217,31,42,31,175,31,232,31,149,31,162,31,40,31,213,31,106,31,215,31,143,31,143,30,226,31,36,31,116,31,102,31,136,31,242,31,18,31,241,31,153,31,87,31,255,31,255,30,32,31,205,31,205,30,187,31,110,31,254,31,254,30,254,29,254,28,4,31,238,31,65,31,88,31,88,30,88,29,183,31,35,31,90,31,90,30,109,31,154,31,196,31,154,31,154,30,154,29,208,31,220,31,212,31,147,31,153,31,9,31,131,31,28,31,181,31,247,31,50,31,50,30,50,29,118,31,69,31,64,31,181,31,110,31,34,31,91,31,91,30,76,31,151,31,151,30,179,31,13,31,5,31,5,30,46,31,46,30,103,31,197,31,197,30,207,31,80,31,80,30,144,31,113,31,15,31,7,31,77,31,210,31,210,30,182,31,245,31,245,30,245,29,24,31,24,30,24,29,48,31,184,31,188,31,148,31,148,30,249,31,95,31,113,31,153,31,153,30,81,31,53,31,214,31,214,30,110,31,110,30,110,29,37,31,216,31,142,31,223,31,223,30,123,31,114,31,114,31,213,31,81,31,190,31,190,30,231,31,147,31,240,31,157,31,157,30,255,31,255,30,127,31,18,31,209,31,165,31,252,31,149,31,149,30,49,31,49,30,177,31,11,31,199,31,59,31,246,31,159,31,159,30,147,31,96,31,34,31,34,30,34,31,109,31,121,31,150,31,135,31,2,31,136,31,27,31,184,31,54,31,123,31,36,31,36,30,172,31,101,31,148,31,231,31,129,31,125,31,108,31,186,31,7,31,46,31,123,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
