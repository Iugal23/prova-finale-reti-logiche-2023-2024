-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_542 is
end project_tb_542;

architecture project_tb_arch_542 of project_tb_542 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 326;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (41,0,39,0,0,0,129,0,109,0,124,0,33,0,22,0,92,0,0,0,106,0,102,0,81,0,84,0,65,0,76,0,31,0,0,0,199,0,53,0,0,0,32,0,17,0,197,0,245,0,119,0,142,0,72,0,196,0,160,0,181,0,0,0,87,0,129,0,178,0,178,0,3,0,107,0,7,0,0,0,228,0,138,0,148,0,252,0,45,0,232,0,28,0,52,0,69,0,146,0,147,0,120,0,144,0,240,0,14,0,200,0,35,0,189,0,0,0,244,0,0,0,240,0,127,0,195,0,176,0,0,0,183,0,245,0,32,0,173,0,0,0,246,0,115,0,203,0,0,0,0,0,221,0,0,0,203,0,163,0,20,0,110,0,204,0,82,0,136,0,0,0,111,0,0,0,119,0,160,0,114,0,236,0,211,0,45,0,225,0,0,0,232,0,135,0,160,0,80,0,218,0,65,0,0,0,121,0,148,0,0,0,4,0,37,0,31,0,55,0,218,0,115,0,230,0,99,0,0,0,139,0,95,0,206,0,0,0,45,0,69,0,0,0,225,0,211,0,193,0,0,0,210,0,4,0,40,0,207,0,61,0,142,0,151,0,142,0,99,0,213,0,8,0,219,0,101,0,0,0,129,0,101,0,0,0,124,0,208,0,142,0,89,0,0,0,130,0,165,0,0,0,135,0,241,0,0,0,26,0,219,0,65,0,8,0,0,0,0,0,34,0,34,0,26,0,151,0,213,0,170,0,103,0,34,0,202,0,137,0,9,0,201,0,170,0,244,0,6,0,0,0,40,0,181,0,78,0,31,0,0,0,223,0,71,0,0,0,50,0,253,0,59,0,186,0,9,0,221,0,64,0,0,0,0,0,36,0,0,0,194,0,208,0,155,0,0,0,1,0,127,0,69,0,50,0,106,0,24,0,0,0,234,0,13,0,27,0,234,0,56,0,0,0,44,0,66,0,228,0,8,0,210,0,190,0,0,0,212,0,81,0,3,0,94,0,220,0,0,0,1,0,150,0,0,0,206,0,59,0,217,0,55,0,0,0,253,0,32,0,38,0,0,0,170,0,150,0,57,0,237,0,69,0,0,0,47,0,0,0,215,0,0,0,174,0,137,0,20,0,200,0,100,0,0,0,172,0,52,0,195,0,0,0,0,0,0,0,112,0,217,0,62,0,86,0,125,0,0,0,0,0,240,0,146,0,196,0,130,0,110,0,0,0,100,0,72,0,148,0,230,0,9,0,226,0,112,0,13,0,35,0,71,0,65,0,97,0,0,0,83,0,0,0,57,0,0,0,0,0,175,0,63,0,238,0,113,0,223,0,234,0,234,0,36,0,160,0,239,0,218,0,114,0,21,0,124,0,0,0,32,0,58,0,205,0,241,0,218,0,46,0,202,0,0,0,0,0,67,0,187,0,128,0,52,0,217,0,13,0,183,0,218,0,224,0,41,0,111,0,18,0);
signal scenario_full  : scenario_type := (41,31,39,31,39,30,129,31,109,31,124,31,33,31,22,31,92,31,92,30,106,31,102,31,81,31,84,31,65,31,76,31,31,31,31,30,199,31,53,31,53,30,32,31,17,31,197,31,245,31,119,31,142,31,72,31,196,31,160,31,181,31,181,30,87,31,129,31,178,31,178,31,3,31,107,31,7,31,7,30,228,31,138,31,148,31,252,31,45,31,232,31,28,31,52,31,69,31,146,31,147,31,120,31,144,31,240,31,14,31,200,31,35,31,189,31,189,30,244,31,244,30,240,31,127,31,195,31,176,31,176,30,183,31,245,31,32,31,173,31,173,30,246,31,115,31,203,31,203,30,203,29,221,31,221,30,203,31,163,31,20,31,110,31,204,31,82,31,136,31,136,30,111,31,111,30,119,31,160,31,114,31,236,31,211,31,45,31,225,31,225,30,232,31,135,31,160,31,80,31,218,31,65,31,65,30,121,31,148,31,148,30,4,31,37,31,31,31,55,31,218,31,115,31,230,31,99,31,99,30,139,31,95,31,206,31,206,30,45,31,69,31,69,30,225,31,211,31,193,31,193,30,210,31,4,31,40,31,207,31,61,31,142,31,151,31,142,31,99,31,213,31,8,31,219,31,101,31,101,30,129,31,101,31,101,30,124,31,208,31,142,31,89,31,89,30,130,31,165,31,165,30,135,31,241,31,241,30,26,31,219,31,65,31,8,31,8,30,8,29,34,31,34,31,26,31,151,31,213,31,170,31,103,31,34,31,202,31,137,31,9,31,201,31,170,31,244,31,6,31,6,30,40,31,181,31,78,31,31,31,31,30,223,31,71,31,71,30,50,31,253,31,59,31,186,31,9,31,221,31,64,31,64,30,64,29,36,31,36,30,194,31,208,31,155,31,155,30,1,31,127,31,69,31,50,31,106,31,24,31,24,30,234,31,13,31,27,31,234,31,56,31,56,30,44,31,66,31,228,31,8,31,210,31,190,31,190,30,212,31,81,31,3,31,94,31,220,31,220,30,1,31,150,31,150,30,206,31,59,31,217,31,55,31,55,30,253,31,32,31,38,31,38,30,170,31,150,31,57,31,237,31,69,31,69,30,47,31,47,30,215,31,215,30,174,31,137,31,20,31,200,31,100,31,100,30,172,31,52,31,195,31,195,30,195,29,195,28,112,31,217,31,62,31,86,31,125,31,125,30,125,29,240,31,146,31,196,31,130,31,110,31,110,30,100,31,72,31,148,31,230,31,9,31,226,31,112,31,13,31,35,31,71,31,65,31,97,31,97,30,83,31,83,30,57,31,57,30,57,29,175,31,63,31,238,31,113,31,223,31,234,31,234,31,36,31,160,31,239,31,218,31,114,31,21,31,124,31,124,30,32,31,58,31,205,31,241,31,218,31,46,31,202,31,202,30,202,29,67,31,187,31,128,31,52,31,217,31,13,31,183,31,218,31,224,31,41,31,111,31,18,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
