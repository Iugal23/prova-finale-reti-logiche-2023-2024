-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 933;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (60,0,114,0,101,0,217,0,0,0,0,0,233,0,176,0,0,0,251,0,83,0,95,0,0,0,241,0,159,0,20,0,0,0,202,0,102,0,110,0,97,0,59,0,147,0,226,0,166,0,245,0,217,0,147,0,243,0,130,0,226,0,159,0,2,0,184,0,72,0,19,0,207,0,0,0,209,0,204,0,0,0,207,0,101,0,237,0,32,0,116,0,246,0,144,0,71,0,0,0,193,0,0,0,168,0,0,0,201,0,9,0,238,0,0,0,145,0,121,0,150,0,68,0,152,0,210,0,0,0,0,0,153,0,223,0,10,0,176,0,243,0,126,0,134,0,145,0,70,0,130,0,0,0,192,0,117,0,0,0,83,0,232,0,0,0,98,0,195,0,63,0,219,0,251,0,0,0,120,0,217,0,227,0,177,0,0,0,138,0,0,0,0,0,20,0,227,0,0,0,156,0,172,0,175,0,0,0,126,0,146,0,0,0,208,0,33,0,154,0,228,0,133,0,0,0,0,0,10,0,0,0,164,0,81,0,217,0,77,0,205,0,76,0,247,0,3,0,146,0,170,0,67,0,118,0,202,0,164,0,0,0,0,0,0,0,117,0,74,0,92,0,128,0,197,0,16,0,44,0,192,0,18,0,237,0,114,0,47,0,40,0,17,0,0,0,52,0,120,0,81,0,0,0,63,0,166,0,0,0,143,0,99,0,22,0,0,0,21,0,15,0,170,0,87,0,0,0,175,0,217,0,146,0,0,0,241,0,140,0,246,0,243,0,242,0,141,0,135,0,0,0,228,0,0,0,205,0,139,0,130,0,73,0,0,0,131,0,98,0,230,0,47,0,0,0,162,0,119,0,71,0,130,0,203,0,26,0,179,0,148,0,171,0,0,0,37,0,103,0,0,0,219,0,0,0,0,0,47,0,182,0,45,0,0,0,0,0,72,0,223,0,232,0,136,0,247,0,10,0,16,0,203,0,0,0,158,0,52,0,0,0,28,0,0,0,149,0,93,0,30,0,171,0,197,0,156,0,0,0,0,0,137,0,50,0,0,0,202,0,0,0,228,0,13,0,40,0,91,0,253,0,5,0,100,0,14,0,173,0,116,0,220,0,231,0,41,0,122,0,152,0,54,0,176,0,0,0,67,0,0,0,132,0,124,0,97,0,191,0,72,0,0,0,200,0,177,0,0,0,238,0,0,0,96,0,200,0,154,0,165,0,122,0,194,0,57,0,0,0,161,0,9,0,93,0,216,0,0,0,177,0,30,0,115,0,131,0,254,0,217,0,0,0,151,0,28,0,225,0,179,0,200,0,0,0,168,0,0,0,0,0,197,0,228,0,0,0,72,0,58,0,90,0,119,0,48,0,141,0,0,0,0,0,33,0,0,0,78,0,255,0,220,0,0,0,0,0,128,0,21,0,245,0,0,0,224,0,252,0,102,0,0,0,178,0,83,0,0,0,235,0,109,0,32,0,110,0,126,0,0,0,95,0,0,0,232,0,16,0,56,0,0,0,215,0,0,0,221,0,230,0,206,0,156,0,236,0,0,0,224,0,38,0,175,0,209,0,25,0,68,0,164,0,215,0,0,0,0,0,0,0,0,0,126,0,0,0,63,0,0,0,228,0,60,0,24,0,134,0,3,0,117,0,27,0,199,0,224,0,41,0,0,0,0,0,0,0,94,0,82,0,0,0,92,0,201,0,151,0,0,0,244,0,238,0,53,0,241,0,0,0,0,0,77,0,170,0,12,0,44,0,88,0,220,0,0,0,0,0,76,0,233,0,5,0,0,0,210,0,228,0,186,0,161,0,126,0,7,0,16,0,0,0,200,0,56,0,205,0,129,0,0,0,31,0,66,0,253,0,151,0,49,0,192,0,133,0,20,0,140,0,226,0,182,0,120,0,120,0,82,0,226,0,140,0,222,0,176,0,240,0,7,0,97,0,0,0,0,0,183,0,0,0,44,0,34,0,178,0,0,0,137,0,0,0,96,0,219,0,126,0,198,0,0,0,177,0,236,0,171,0,67,0,202,0,198,0,227,0,0,0,166,0,246,0,14,0,27,0,241,0,0,0,85,0,180,0,121,0,115,0,0,0,211,0,174,0,48,0,0,0,222,0,178,0,139,0,37,0,113,0,221,0,139,0,0,0,212,0,110,0,240,0,205,0,0,0,163,0,79,0,84,0,42,0,160,0,68,0,233,0,118,0,55,0,38,0,51,0,94,0,31,0,84,0,0,0,196,0,32,0,0,0,102,0,101,0,102,0,179,0,0,0,140,0,218,0,178,0,249,0,0,0,74,0,0,0,45,0,74,0,87,0,30,0,5,0,124,0,92,0,0,0,179,0,98,0,0,0,55,0,196,0,218,0,0,0,233,0,206,0,8,0,62,0,142,0,111,0,183,0,119,0,173,0,42,0,204,0,0,0,244,0,171,0,187,0,142,0,209,0,160,0,84,0,0,0,85,0,0,0,136,0,157,0,90,0,0,0,176,0,89,0,114,0,189,0,226,0,232,0,241,0,135,0,36,0,0,0,71,0,64,0,192,0,204,0,189,0,111,0,121,0,146,0,0,0,18,0,167,0,45,0,0,0,235,0,236,0,169,0,124,0,175,0,88,0,0,0,190,0,71,0,130,0,66,0,13,0,121,0,204,0,0,0,0,0,117,0,19,0,120,0,166,0,101,0,182,0,193,0,33,0,148,0,37,0,172,0,0,0,168,0,30,0,226,0,193,0,219,0,3,0,208,0,71,0,217,0,0,0,181,0,0,0,118,0,0,0,0,0,78,0,211,0,22,0,251,0,255,0,107,0,159,0,197,0,222,0,148,0,148,0,134,0,229,0,78,0,228,0,229,0,34,0,41,0,66,0,210,0,133,0,182,0,189,0,110,0,182,0,246,0,163,0,0,0,47,0,73,0,63,0,0,0,57,0,155,0,193,0,28,0,149,0,104,0,0,0,110,0,0,0,179,0,251,0,0,0,0,0,226,0,37,0,254,0,70,0,199,0,54,0,126,0,229,0,92,0,31,0,51,0,179,0,124,0,75,0,237,0,142,0,254,0,226,0,201,0,196,0,0,0,0,0,206,0,222,0,143,0,121,0,68,0,147,0,249,0,92,0,170,0,55,0,85,0,52,0,63,0,190,0,0,0,30,0,0,0,107,0,232,0,162,0,0,0,0,0,119,0,77,0,58,0,0,0,255,0,0,0,232,0,47,0,0,0,56,0,0,0,234,0,0,0,50,0,0,0,25,0,0,0,121,0,67,0,227,0,186,0,185,0,225,0,196,0,51,0,181,0,0,0,0,0,159,0,202,0,248,0,0,0,26,0,3,0,58,0,0,0,245,0,95,0,223,0,187,0,53,0,70,0,132,0,0,0,80,0,250,0,219,0,255,0,45,0,86,0,117,0,109,0,121,0,0,0,6,0,10,0,207,0,5,0,95,0,188,0,162,0,0,0,127,0,98,0,116,0,0,0,151,0,59,0,254,0,175,0,0,0,15,0,85,0,0,0,153,0,26,0,234,0,34,0,0,0,17,0,59,0,0,0,129,0,253,0,180,0,102,0,174,0,54,0,52,0,39,0,244,0,119,0,231,0,0,0,173,0,26,0,226,0,209,0,220,0,0,0,40,0,42,0,164,0,0,0,15,0,54,0,125,0,44,0,101,0,173,0,0,0,44,0,252,0,113,0,66,0,182,0,68,0,0,0,165,0,40,0,201,0,42,0,174,0,202,0,117,0,0,0,0,0,125,0,103,0,81,0,128,0,0,0,0,0,66,0,200,0,0,0,10,0,121,0,0,0,26,0,39,0,174,0,0,0,14,0,197,0,0,0,45,0,0,0,0,0,0,0,54,0,146,0,0,0,106,0,219,0,174,0,0,0,209,0,216,0,0,0,59,0,231,0,0,0,233,0,207,0,48,0,50,0,236,0,203,0,164,0,89,0,156,0,230,0,0,0,129,0,0,0,237,0,254,0,80,0,20,0,120,0,0,0,43,0,80,0,0,0,203,0,0,0,61,0,237,0,142,0,90,0,123,0,189,0,0,0,172,0,91,0,5,0,55,0,152,0,0,0,27,0,102,0,5,0,155,0,137,0,65,0,0,0,206,0,0,0,146,0,83,0,204,0,0,0,109,0,0,0,138,0,0,0,23,0,133,0,249,0,112,0,183,0,0,0);
signal scenario_full  : scenario_type := (60,31,114,31,101,31,217,31,217,30,217,29,233,31,176,31,176,30,251,31,83,31,95,31,95,30,241,31,159,31,20,31,20,30,202,31,102,31,110,31,97,31,59,31,147,31,226,31,166,31,245,31,217,31,147,31,243,31,130,31,226,31,159,31,2,31,184,31,72,31,19,31,207,31,207,30,209,31,204,31,204,30,207,31,101,31,237,31,32,31,116,31,246,31,144,31,71,31,71,30,193,31,193,30,168,31,168,30,201,31,9,31,238,31,238,30,145,31,121,31,150,31,68,31,152,31,210,31,210,30,210,29,153,31,223,31,10,31,176,31,243,31,126,31,134,31,145,31,70,31,130,31,130,30,192,31,117,31,117,30,83,31,232,31,232,30,98,31,195,31,63,31,219,31,251,31,251,30,120,31,217,31,227,31,177,31,177,30,138,31,138,30,138,29,20,31,227,31,227,30,156,31,172,31,175,31,175,30,126,31,146,31,146,30,208,31,33,31,154,31,228,31,133,31,133,30,133,29,10,31,10,30,164,31,81,31,217,31,77,31,205,31,76,31,247,31,3,31,146,31,170,31,67,31,118,31,202,31,164,31,164,30,164,29,164,28,117,31,74,31,92,31,128,31,197,31,16,31,44,31,192,31,18,31,237,31,114,31,47,31,40,31,17,31,17,30,52,31,120,31,81,31,81,30,63,31,166,31,166,30,143,31,99,31,22,31,22,30,21,31,15,31,170,31,87,31,87,30,175,31,217,31,146,31,146,30,241,31,140,31,246,31,243,31,242,31,141,31,135,31,135,30,228,31,228,30,205,31,139,31,130,31,73,31,73,30,131,31,98,31,230,31,47,31,47,30,162,31,119,31,71,31,130,31,203,31,26,31,179,31,148,31,171,31,171,30,37,31,103,31,103,30,219,31,219,30,219,29,47,31,182,31,45,31,45,30,45,29,72,31,223,31,232,31,136,31,247,31,10,31,16,31,203,31,203,30,158,31,52,31,52,30,28,31,28,30,149,31,93,31,30,31,171,31,197,31,156,31,156,30,156,29,137,31,50,31,50,30,202,31,202,30,228,31,13,31,40,31,91,31,253,31,5,31,100,31,14,31,173,31,116,31,220,31,231,31,41,31,122,31,152,31,54,31,176,31,176,30,67,31,67,30,132,31,124,31,97,31,191,31,72,31,72,30,200,31,177,31,177,30,238,31,238,30,96,31,200,31,154,31,165,31,122,31,194,31,57,31,57,30,161,31,9,31,93,31,216,31,216,30,177,31,30,31,115,31,131,31,254,31,217,31,217,30,151,31,28,31,225,31,179,31,200,31,200,30,168,31,168,30,168,29,197,31,228,31,228,30,72,31,58,31,90,31,119,31,48,31,141,31,141,30,141,29,33,31,33,30,78,31,255,31,220,31,220,30,220,29,128,31,21,31,245,31,245,30,224,31,252,31,102,31,102,30,178,31,83,31,83,30,235,31,109,31,32,31,110,31,126,31,126,30,95,31,95,30,232,31,16,31,56,31,56,30,215,31,215,30,221,31,230,31,206,31,156,31,236,31,236,30,224,31,38,31,175,31,209,31,25,31,68,31,164,31,215,31,215,30,215,29,215,28,215,27,126,31,126,30,63,31,63,30,228,31,60,31,24,31,134,31,3,31,117,31,27,31,199,31,224,31,41,31,41,30,41,29,41,28,94,31,82,31,82,30,92,31,201,31,151,31,151,30,244,31,238,31,53,31,241,31,241,30,241,29,77,31,170,31,12,31,44,31,88,31,220,31,220,30,220,29,76,31,233,31,5,31,5,30,210,31,228,31,186,31,161,31,126,31,7,31,16,31,16,30,200,31,56,31,205,31,129,31,129,30,31,31,66,31,253,31,151,31,49,31,192,31,133,31,20,31,140,31,226,31,182,31,120,31,120,31,82,31,226,31,140,31,222,31,176,31,240,31,7,31,97,31,97,30,97,29,183,31,183,30,44,31,34,31,178,31,178,30,137,31,137,30,96,31,219,31,126,31,198,31,198,30,177,31,236,31,171,31,67,31,202,31,198,31,227,31,227,30,166,31,246,31,14,31,27,31,241,31,241,30,85,31,180,31,121,31,115,31,115,30,211,31,174,31,48,31,48,30,222,31,178,31,139,31,37,31,113,31,221,31,139,31,139,30,212,31,110,31,240,31,205,31,205,30,163,31,79,31,84,31,42,31,160,31,68,31,233,31,118,31,55,31,38,31,51,31,94,31,31,31,84,31,84,30,196,31,32,31,32,30,102,31,101,31,102,31,179,31,179,30,140,31,218,31,178,31,249,31,249,30,74,31,74,30,45,31,74,31,87,31,30,31,5,31,124,31,92,31,92,30,179,31,98,31,98,30,55,31,196,31,218,31,218,30,233,31,206,31,8,31,62,31,142,31,111,31,183,31,119,31,173,31,42,31,204,31,204,30,244,31,171,31,187,31,142,31,209,31,160,31,84,31,84,30,85,31,85,30,136,31,157,31,90,31,90,30,176,31,89,31,114,31,189,31,226,31,232,31,241,31,135,31,36,31,36,30,71,31,64,31,192,31,204,31,189,31,111,31,121,31,146,31,146,30,18,31,167,31,45,31,45,30,235,31,236,31,169,31,124,31,175,31,88,31,88,30,190,31,71,31,130,31,66,31,13,31,121,31,204,31,204,30,204,29,117,31,19,31,120,31,166,31,101,31,182,31,193,31,33,31,148,31,37,31,172,31,172,30,168,31,30,31,226,31,193,31,219,31,3,31,208,31,71,31,217,31,217,30,181,31,181,30,118,31,118,30,118,29,78,31,211,31,22,31,251,31,255,31,107,31,159,31,197,31,222,31,148,31,148,31,134,31,229,31,78,31,228,31,229,31,34,31,41,31,66,31,210,31,133,31,182,31,189,31,110,31,182,31,246,31,163,31,163,30,47,31,73,31,63,31,63,30,57,31,155,31,193,31,28,31,149,31,104,31,104,30,110,31,110,30,179,31,251,31,251,30,251,29,226,31,37,31,254,31,70,31,199,31,54,31,126,31,229,31,92,31,31,31,51,31,179,31,124,31,75,31,237,31,142,31,254,31,226,31,201,31,196,31,196,30,196,29,206,31,222,31,143,31,121,31,68,31,147,31,249,31,92,31,170,31,55,31,85,31,52,31,63,31,190,31,190,30,30,31,30,30,107,31,232,31,162,31,162,30,162,29,119,31,77,31,58,31,58,30,255,31,255,30,232,31,47,31,47,30,56,31,56,30,234,31,234,30,50,31,50,30,25,31,25,30,121,31,67,31,227,31,186,31,185,31,225,31,196,31,51,31,181,31,181,30,181,29,159,31,202,31,248,31,248,30,26,31,3,31,58,31,58,30,245,31,95,31,223,31,187,31,53,31,70,31,132,31,132,30,80,31,250,31,219,31,255,31,45,31,86,31,117,31,109,31,121,31,121,30,6,31,10,31,207,31,5,31,95,31,188,31,162,31,162,30,127,31,98,31,116,31,116,30,151,31,59,31,254,31,175,31,175,30,15,31,85,31,85,30,153,31,26,31,234,31,34,31,34,30,17,31,59,31,59,30,129,31,253,31,180,31,102,31,174,31,54,31,52,31,39,31,244,31,119,31,231,31,231,30,173,31,26,31,226,31,209,31,220,31,220,30,40,31,42,31,164,31,164,30,15,31,54,31,125,31,44,31,101,31,173,31,173,30,44,31,252,31,113,31,66,31,182,31,68,31,68,30,165,31,40,31,201,31,42,31,174,31,202,31,117,31,117,30,117,29,125,31,103,31,81,31,128,31,128,30,128,29,66,31,200,31,200,30,10,31,121,31,121,30,26,31,39,31,174,31,174,30,14,31,197,31,197,30,45,31,45,30,45,29,45,28,54,31,146,31,146,30,106,31,219,31,174,31,174,30,209,31,216,31,216,30,59,31,231,31,231,30,233,31,207,31,48,31,50,31,236,31,203,31,164,31,89,31,156,31,230,31,230,30,129,31,129,30,237,31,254,31,80,31,20,31,120,31,120,30,43,31,80,31,80,30,203,31,203,30,61,31,237,31,142,31,90,31,123,31,189,31,189,30,172,31,91,31,5,31,55,31,152,31,152,30,27,31,102,31,5,31,155,31,137,31,65,31,65,30,206,31,206,30,146,31,83,31,204,31,204,30,109,31,109,30,138,31,138,30,23,31,133,31,249,31,112,31,183,31,183,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
