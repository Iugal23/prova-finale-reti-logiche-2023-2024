-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_280 is
end project_tb_280;

architecture project_tb_arch_280 of project_tb_280 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 968;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,183,0,189,0,0,0,188,0,57,0,231,0,57,0,90,0,0,0,32,0,12,0,180,0,0,0,138,0,143,0,188,0,250,0,18,0,187,0,31,0,0,0,0,0,238,0,6,0,28,0,151,0,87,0,8,0,59,0,9,0,89,0,27,0,28,0,54,0,0,0,22,0,0,0,133,0,110,0,184,0,249,0,172,0,235,0,158,0,203,0,116,0,238,0,12,0,248,0,210,0,208,0,28,0,0,0,115,0,98,0,222,0,61,0,107,0,0,0,113,0,48,0,0,0,99,0,0,0,116,0,215,0,92,0,222,0,204,0,192,0,10,0,199,0,0,0,0,0,0,0,6,0,181,0,239,0,65,0,183,0,200,0,80,0,107,0,112,0,88,0,0,0,230,0,0,0,236,0,210,0,0,0,125,0,249,0,112,0,23,0,13,0,124,0,0,0,250,0,228,0,6,0,39,0,0,0,255,0,115,0,80,0,0,0,0,0,203,0,0,0,127,0,0,0,23,0,143,0,68,0,42,0,66,0,195,0,128,0,169,0,36,0,52,0,126,0,169,0,0,0,123,0,43,0,187,0,136,0,0,0,153,0,185,0,192,0,0,0,16,0,167,0,186,0,249,0,130,0,236,0,230,0,29,0,84,0,109,0,23,0,41,0,0,0,222,0,7,0,184,0,57,0,0,0,247,0,5,0,80,0,0,0,149,0,109,0,204,0,171,0,143,0,99,0,247,0,78,0,227,0,96,0,72,0,222,0,49,0,202,0,241,0,80,0,0,0,58,0,0,0,218,0,22,0,133,0,154,0,163,0,19,0,211,0,0,0,203,0,0,0,0,0,0,0,29,0,0,0,0,0,186,0,0,0,135,0,0,0,0,0,84,0,5,0,73,0,26,0,196,0,55,0,87,0,169,0,97,0,26,0,96,0,165,0,251,0,106,0,225,0,254,0,128,0,0,0,156,0,0,0,0,0,232,0,0,0,119,0,225,0,172,0,188,0,67,0,82,0,48,0,178,0,87,0,10,0,182,0,0,0,242,0,39,0,32,0,50,0,16,0,109,0,70,0,33,0,122,0,0,0,128,0,25,0,214,0,0,0,111,0,14,0,87,0,60,0,89,0,28,0,0,0,209,0,77,0,73,0,91,0,132,0,177,0,143,0,159,0,44,0,204,0,191,0,127,0,0,0,193,0,96,0,134,0,110,0,83,0,0,0,18,0,93,0,0,0,177,0,136,0,194,0,3,0,187,0,194,0,1,0,197,0,0,0,252,0,82,0,16,0,84,0,171,0,29,0,244,0,210,0,82,0,224,0,0,0,175,0,247,0,208,0,177,0,248,0,0,0,119,0,63,0,90,0,114,0,0,0,49,0,249,0,121,0,170,0,2,0,249,0,230,0,238,0,53,0,89,0,0,0,67,0,143,0,254,0,61,0,85,0,0,0,33,0,0,0,123,0,27,0,0,0,229,0,46,0,226,0,71,0,218,0,119,0,213,0,0,0,107,0,0,0,248,0,0,0,35,0,81,0,0,0,169,0,215,0,98,0,0,0,0,0,106,0,212,0,35,0,63,0,154,0,40,0,161,0,88,0,144,0,0,0,101,0,69,0,207,0,93,0,166,0,182,0,110,0,40,0,114,0,33,0,0,0,87,0,0,0,59,0,30,0,245,0,0,0,171,0,247,0,65,0,0,0,86,0,236,0,94,0,0,0,12,0,141,0,144,0,0,0,209,0,0,0,220,0,135,0,230,0,253,0,0,0,0,0,3,0,0,0,167,0,142,0,209,0,139,0,8,0,0,0,251,0,185,0,187,0,51,0,4,0,153,0,196,0,165,0,0,0,231,0,248,0,165,0,0,0,0,0,201,0,0,0,253,0,178,0,166,0,2,0,169,0,167,0,0,0,150,0,11,0,171,0,127,0,87,0,0,0,0,0,205,0,243,0,0,0,231,0,0,0,43,0,210,0,180,0,91,0,0,0,29,0,0,0,82,0,114,0,85,0,57,0,0,0,0,0,10,0,0,0,0,0,101,0,248,0,0,0,177,0,54,0,163,0,11,0,205,0,232,0,234,0,148,0,0,0,0,0,0,0,67,0,153,0,203,0,37,0,65,0,156,0,189,0,0,0,181,0,229,0,223,0,37,0,17,0,127,0,0,0,168,0,100,0,100,0,220,0,0,0,0,0,0,0,0,0,10,0,0,0,180,0,215,0,156,0,55,0,214,0,19,0,0,0,94,0,250,0,125,0,59,0,73,0,116,0,72,0,0,0,0,0,116,0,210,0,1,0,173,0,192,0,0,0,0,0,9,0,0,0,0,0,0,0,0,0,238,0,0,0,155,0,0,0,196,0,229,0,188,0,194,0,242,0,188,0,53,0,70,0,225,0,97,0,150,0,234,0,73,0,6,0,0,0,218,0,65,0,104,0,80,0,221,0,162,0,118,0,153,0,39,0,204,0,83,0,0,0,63,0,118,0,0,0,0,0,180,0,0,0,218,0,0,0,0,0,125,0,127,0,14,0,39,0,71,0,179,0,96,0,27,0,183,0,0,0,47,0,164,0,82,0,51,0,0,0,231,0,98,0,179,0,186,0,124,0,120,0,20,0,178,0,25,0,237,0,251,0,0,0,166,0,0,0,233,0,113,0,202,0,110,0,37,0,35,0,105,0,220,0,163,0,252,0,54,0,0,0,43,0,58,0,128,0,77,0,0,0,53,0,159,0,43,0,156,0,81,0,78,0,0,0,222,0,2,0,167,0,37,0,220,0,123,0,0,0,243,0,0,0,174,0,74,0,135,0,26,0,0,0,188,0,0,0,9,0,49,0,0,0,79,0,244,0,235,0,42,0,254,0,0,0,0,0,35,0,140,0,0,0,178,0,148,0,169,0,209,0,125,0,167,0,149,0,157,0,58,0,0,0,0,0,0,0,254,0,169,0,0,0,7,0,160,0,142,0,182,0,0,0,13,0,106,0,0,0,216,0,137,0,114,0,0,0,0,0,0,0,167,0,123,0,214,0,63,0,202,0,149,0,17,0,0,0,185,0,103,0,0,0,90,0,0,0,0,0,56,0,123,0,239,0,0,0,87,0,0,0,238,0,145,0,0,0,175,0,74,0,0,0,90,0,86,0,0,0,48,0,0,0,80,0,155,0,102,0,53,0,18,0,19,0,247,0,138,0,171,0,194,0,0,0,104,0,43,0,59,0,11,0,252,0,145,0,0,0,0,0,232,0,0,0,0,0,146,0,3,0,0,0,0,0,0,0,137,0,136,0,174,0,0,0,19,0,226,0,219,0,67,0,0,0,33,0,100,0,71,0,0,0,236,0,0,0,0,0,112,0,180,0,56,0,0,0,180,0,202,0,0,0,67,0,0,0,125,0,155,0,0,0,30,0,79,0,90,0,127,0,192,0,66,0,251,0,0,0,0,0,0,0,233,0,205,0,0,0,85,0,233,0,73,0,133,0,197,0,202,0,99,0,0,0,202,0,152,0,255,0,24,0,103,0,116,0,72,0,166,0,0,0,0,0,91,0,249,0,23,0,68,0,221,0,210,0,19,0,30,0,0,0,167,0,0,0,156,0,88,0,107,0,69,0,146,0,250,0,62,0,128,0,15,0,118,0,0,0,4,0,128,0,98,0,242,0,0,0,62,0,210,0,23,0,177,0,128,0,0,0,143,0,67,0,6,0,0,0,0,0,0,0,0,0,187,0,147,0,178,0,86,0,227,0,232,0,178,0,53,0,249,0,80,0,200,0,155,0,156,0,0,0,19,0,94,0,0,0,44,0,31,0,65,0,81,0,4,0,41,0,137,0,185,0,156,0,93,0,170,0,128,0,229,0,217,0,180,0,0,0,74,0,18,0,1,0,75,0,171,0,244,0,161,0,0,0,171,0,106,0,101,0,0,0,71,0,0,0,108,0,175,0,154,0,88,0,157,0,255,0,74,0,59,0,184,0,71,0,201,0,132,0,248,0,168,0,137,0,120,0,0,0,24,0,223,0,0,0,196,0,123,0,0,0,235,0,0,0,137,0,0,0,0,0,212,0,189,0,150,0,147,0,159,0,217,0,210,0,215,0,0,0,36,0,74,0,18,0,141,0,74,0,51,0,251,0,230,0,191,0,222,0,157,0,0,0,91,0,3,0,0,0,24,0,117,0,109,0,57,0,198,0,150,0,236,0,155,0,82,0,0,0,16,0,78,0,0,0,249,0,192,0,0,0,239,0,79,0,1,0,248,0,252,0,0,0,145,0,143,0,165,0,66,0,30,0,0,0,143,0,54,0,0,0,78,0,148,0,251,0,231,0,234,0,195,0,244,0,0,0,81,0,99,0);
signal scenario_full  : scenario_type := (16,31,183,31,189,31,189,30,188,31,57,31,231,31,57,31,90,31,90,30,32,31,12,31,180,31,180,30,138,31,143,31,188,31,250,31,18,31,187,31,31,31,31,30,31,29,238,31,6,31,28,31,151,31,87,31,8,31,59,31,9,31,89,31,27,31,28,31,54,31,54,30,22,31,22,30,133,31,110,31,184,31,249,31,172,31,235,31,158,31,203,31,116,31,238,31,12,31,248,31,210,31,208,31,28,31,28,30,115,31,98,31,222,31,61,31,107,31,107,30,113,31,48,31,48,30,99,31,99,30,116,31,215,31,92,31,222,31,204,31,192,31,10,31,199,31,199,30,199,29,199,28,6,31,181,31,239,31,65,31,183,31,200,31,80,31,107,31,112,31,88,31,88,30,230,31,230,30,236,31,210,31,210,30,125,31,249,31,112,31,23,31,13,31,124,31,124,30,250,31,228,31,6,31,39,31,39,30,255,31,115,31,80,31,80,30,80,29,203,31,203,30,127,31,127,30,23,31,143,31,68,31,42,31,66,31,195,31,128,31,169,31,36,31,52,31,126,31,169,31,169,30,123,31,43,31,187,31,136,31,136,30,153,31,185,31,192,31,192,30,16,31,167,31,186,31,249,31,130,31,236,31,230,31,29,31,84,31,109,31,23,31,41,31,41,30,222,31,7,31,184,31,57,31,57,30,247,31,5,31,80,31,80,30,149,31,109,31,204,31,171,31,143,31,99,31,247,31,78,31,227,31,96,31,72,31,222,31,49,31,202,31,241,31,80,31,80,30,58,31,58,30,218,31,22,31,133,31,154,31,163,31,19,31,211,31,211,30,203,31,203,30,203,29,203,28,29,31,29,30,29,29,186,31,186,30,135,31,135,30,135,29,84,31,5,31,73,31,26,31,196,31,55,31,87,31,169,31,97,31,26,31,96,31,165,31,251,31,106,31,225,31,254,31,128,31,128,30,156,31,156,30,156,29,232,31,232,30,119,31,225,31,172,31,188,31,67,31,82,31,48,31,178,31,87,31,10,31,182,31,182,30,242,31,39,31,32,31,50,31,16,31,109,31,70,31,33,31,122,31,122,30,128,31,25,31,214,31,214,30,111,31,14,31,87,31,60,31,89,31,28,31,28,30,209,31,77,31,73,31,91,31,132,31,177,31,143,31,159,31,44,31,204,31,191,31,127,31,127,30,193,31,96,31,134,31,110,31,83,31,83,30,18,31,93,31,93,30,177,31,136,31,194,31,3,31,187,31,194,31,1,31,197,31,197,30,252,31,82,31,16,31,84,31,171,31,29,31,244,31,210,31,82,31,224,31,224,30,175,31,247,31,208,31,177,31,248,31,248,30,119,31,63,31,90,31,114,31,114,30,49,31,249,31,121,31,170,31,2,31,249,31,230,31,238,31,53,31,89,31,89,30,67,31,143,31,254,31,61,31,85,31,85,30,33,31,33,30,123,31,27,31,27,30,229,31,46,31,226,31,71,31,218,31,119,31,213,31,213,30,107,31,107,30,248,31,248,30,35,31,81,31,81,30,169,31,215,31,98,31,98,30,98,29,106,31,212,31,35,31,63,31,154,31,40,31,161,31,88,31,144,31,144,30,101,31,69,31,207,31,93,31,166,31,182,31,110,31,40,31,114,31,33,31,33,30,87,31,87,30,59,31,30,31,245,31,245,30,171,31,247,31,65,31,65,30,86,31,236,31,94,31,94,30,12,31,141,31,144,31,144,30,209,31,209,30,220,31,135,31,230,31,253,31,253,30,253,29,3,31,3,30,167,31,142,31,209,31,139,31,8,31,8,30,251,31,185,31,187,31,51,31,4,31,153,31,196,31,165,31,165,30,231,31,248,31,165,31,165,30,165,29,201,31,201,30,253,31,178,31,166,31,2,31,169,31,167,31,167,30,150,31,11,31,171,31,127,31,87,31,87,30,87,29,205,31,243,31,243,30,231,31,231,30,43,31,210,31,180,31,91,31,91,30,29,31,29,30,82,31,114,31,85,31,57,31,57,30,57,29,10,31,10,30,10,29,101,31,248,31,248,30,177,31,54,31,163,31,11,31,205,31,232,31,234,31,148,31,148,30,148,29,148,28,67,31,153,31,203,31,37,31,65,31,156,31,189,31,189,30,181,31,229,31,223,31,37,31,17,31,127,31,127,30,168,31,100,31,100,31,220,31,220,30,220,29,220,28,220,27,10,31,10,30,180,31,215,31,156,31,55,31,214,31,19,31,19,30,94,31,250,31,125,31,59,31,73,31,116,31,72,31,72,30,72,29,116,31,210,31,1,31,173,31,192,31,192,30,192,29,9,31,9,30,9,29,9,28,9,27,238,31,238,30,155,31,155,30,196,31,229,31,188,31,194,31,242,31,188,31,53,31,70,31,225,31,97,31,150,31,234,31,73,31,6,31,6,30,218,31,65,31,104,31,80,31,221,31,162,31,118,31,153,31,39,31,204,31,83,31,83,30,63,31,118,31,118,30,118,29,180,31,180,30,218,31,218,30,218,29,125,31,127,31,14,31,39,31,71,31,179,31,96,31,27,31,183,31,183,30,47,31,164,31,82,31,51,31,51,30,231,31,98,31,179,31,186,31,124,31,120,31,20,31,178,31,25,31,237,31,251,31,251,30,166,31,166,30,233,31,113,31,202,31,110,31,37,31,35,31,105,31,220,31,163,31,252,31,54,31,54,30,43,31,58,31,128,31,77,31,77,30,53,31,159,31,43,31,156,31,81,31,78,31,78,30,222,31,2,31,167,31,37,31,220,31,123,31,123,30,243,31,243,30,174,31,74,31,135,31,26,31,26,30,188,31,188,30,9,31,49,31,49,30,79,31,244,31,235,31,42,31,254,31,254,30,254,29,35,31,140,31,140,30,178,31,148,31,169,31,209,31,125,31,167,31,149,31,157,31,58,31,58,30,58,29,58,28,254,31,169,31,169,30,7,31,160,31,142,31,182,31,182,30,13,31,106,31,106,30,216,31,137,31,114,31,114,30,114,29,114,28,167,31,123,31,214,31,63,31,202,31,149,31,17,31,17,30,185,31,103,31,103,30,90,31,90,30,90,29,56,31,123,31,239,31,239,30,87,31,87,30,238,31,145,31,145,30,175,31,74,31,74,30,90,31,86,31,86,30,48,31,48,30,80,31,155,31,102,31,53,31,18,31,19,31,247,31,138,31,171,31,194,31,194,30,104,31,43,31,59,31,11,31,252,31,145,31,145,30,145,29,232,31,232,30,232,29,146,31,3,31,3,30,3,29,3,28,137,31,136,31,174,31,174,30,19,31,226,31,219,31,67,31,67,30,33,31,100,31,71,31,71,30,236,31,236,30,236,29,112,31,180,31,56,31,56,30,180,31,202,31,202,30,67,31,67,30,125,31,155,31,155,30,30,31,79,31,90,31,127,31,192,31,66,31,251,31,251,30,251,29,251,28,233,31,205,31,205,30,85,31,233,31,73,31,133,31,197,31,202,31,99,31,99,30,202,31,152,31,255,31,24,31,103,31,116,31,72,31,166,31,166,30,166,29,91,31,249,31,23,31,68,31,221,31,210,31,19,31,30,31,30,30,167,31,167,30,156,31,88,31,107,31,69,31,146,31,250,31,62,31,128,31,15,31,118,31,118,30,4,31,128,31,98,31,242,31,242,30,62,31,210,31,23,31,177,31,128,31,128,30,143,31,67,31,6,31,6,30,6,29,6,28,6,27,187,31,147,31,178,31,86,31,227,31,232,31,178,31,53,31,249,31,80,31,200,31,155,31,156,31,156,30,19,31,94,31,94,30,44,31,31,31,65,31,81,31,4,31,41,31,137,31,185,31,156,31,93,31,170,31,128,31,229,31,217,31,180,31,180,30,74,31,18,31,1,31,75,31,171,31,244,31,161,31,161,30,171,31,106,31,101,31,101,30,71,31,71,30,108,31,175,31,154,31,88,31,157,31,255,31,74,31,59,31,184,31,71,31,201,31,132,31,248,31,168,31,137,31,120,31,120,30,24,31,223,31,223,30,196,31,123,31,123,30,235,31,235,30,137,31,137,30,137,29,212,31,189,31,150,31,147,31,159,31,217,31,210,31,215,31,215,30,36,31,74,31,18,31,141,31,74,31,51,31,251,31,230,31,191,31,222,31,157,31,157,30,91,31,3,31,3,30,24,31,117,31,109,31,57,31,198,31,150,31,236,31,155,31,82,31,82,30,16,31,78,31,78,30,249,31,192,31,192,30,239,31,79,31,1,31,248,31,252,31,252,30,145,31,143,31,165,31,66,31,30,31,30,30,143,31,54,31,54,30,78,31,148,31,251,31,231,31,234,31,195,31,244,31,244,30,81,31,99,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
