-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_52 is
end project_tb_52;

architecture project_tb_arch_52 of project_tb_52 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 573;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (161,0,70,0,9,0,136,0,233,0,106,0,237,0,40,0,239,0,142,0,19,0,221,0,0,0,97,0,234,0,103,0,0,0,0,0,44,0,41,0,133,0,0,0,216,0,184,0,145,0,204,0,229,0,68,0,0,0,234,0,49,0,149,0,0,0,166,0,3,0,107,0,0,0,127,0,0,0,164,0,0,0,143,0,90,0,0,0,69,0,194,0,19,0,160,0,141,0,60,0,76,0,2,0,0,0,0,0,6,0,0,0,196,0,133,0,5,0,92,0,121,0,114,0,74,0,194,0,226,0,65,0,9,0,100,0,154,0,199,0,0,0,118,0,43,0,0,0,27,0,148,0,227,0,25,0,42,0,203,0,72,0,179,0,0,0,93,0,41,0,61,0,0,0,123,0,0,0,0,0,40,0,72,0,0,0,79,0,115,0,62,0,57,0,72,0,0,0,214,0,83,0,41,0,127,0,130,0,0,0,152,0,1,0,115,0,17,0,0,0,15,0,0,0,228,0,61,0,191,0,245,0,203,0,145,0,92,0,206,0,201,0,0,0,150,0,87,0,137,0,221,0,0,0,200,0,8,0,6,0,234,0,210,0,59,0,71,0,10,0,0,0,148,0,37,0,0,0,31,0,0,0,136,0,0,0,35,0,107,0,0,0,234,0,16,0,0,0,242,0,84,0,251,0,150,0,112,0,178,0,232,0,27,0,145,0,234,0,139,0,0,0,25,0,181,0,91,0,81,0,174,0,241,0,162,0,35,0,107,0,0,0,236,0,0,0,27,0,131,0,66,0,140,0,152,0,19,0,80,0,0,0,21,0,0,0,191,0,53,0,232,0,198,0,17,0,0,0,149,0,28,0,91,0,90,0,3,0,124,0,0,0,163,0,88,0,40,0,146,0,123,0,191,0,165,0,168,0,88,0,224,0,209,0,0,0,190,0,92,0,99,0,108,0,100,0,33,0,147,0,123,0,69,0,0,0,187,0,64,0,3,0,9,0,53,0,172,0,149,0,0,0,233,0,69,0,69,0,208,0,61,0,29,0,169,0,0,0,100,0,36,0,198,0,246,0,6,0,187,0,251,0,0,0,4,0,35,0,146,0,125,0,82,0,0,0,180,0,0,0,91,0,214,0,176,0,64,0,0,0,121,0,212,0,66,0,249,0,161,0,91,0,98,0,0,0,0,0,0,0,135,0,16,0,58,0,0,0,91,0,0,0,0,0,0,0,109,0,46,0,114,0,0,0,157,0,249,0,0,0,51,0,7,0,61,0,97,0,188,0,0,0,131,0,158,0,105,0,224,0,136,0,61,0,115,0,0,0,19,0,0,0,0,0,195,0,0,0,0,0,0,0,136,0,0,0,169,0,197,0,203,0,0,0,0,0,232,0,3,0,89,0,91,0,156,0,40,0,115,0,22,0,126,0,0,0,153,0,54,0,0,0,1,0,0,0,0,0,28,0,61,0,85,0,85,0,162,0,94,0,81,0,115,0,148,0,206,0,68,0,45,0,0,0,35,0,122,0,0,0,40,0,114,0,0,0,0,0,224,0,103,0,33,0,97,0,248,0,22,0,250,0,22,0,136,0,40,0,186,0,13,0,112,0,127,0,130,0,0,0,214,0,0,0,175,0,147,0,0,0,92,0,222,0,0,0,20,0,89,0,76,0,116,0,115,0,243,0,7,0,25,0,76,0,202,0,0,0,171,0,231,0,132,0,153,0,135,0,0,0,122,0,244,0,130,0,161,0,4,0,110,0,13,0,121,0,251,0,179,0,151,0,162,0,255,0,14,0,243,0,82,0,0,0,44,0,182,0,41,0,0,0,29,0,25,0,69,0,92,0,115,0,219,0,100,0,1,0,219,0,140,0,82,0,171,0,36,0,227,0,181,0,215,0,18,0,215,0,186,0,70,0,89,0,0,0,84,0,0,0,48,0,165,0,18,0,1,0,0,0,92,0,199,0,90,0,87,0,119,0,54,0,115,0,77,0,181,0,40,0,193,0,117,0,71,0,0,0,98,0,255,0,61,0,93,0,58,0,234,0,17,0,68,0,199,0,215,0,0,0,194,0,44,0,0,0,68,0,129,0,164,0,150,0,57,0,185,0,7,0,185,0,197,0,157,0,189,0,126,0,0,0,217,0,138,0,0,0,187,0,127,0,0,0,174,0,63,0,0,0,0,0,0,0,87,0,172,0,147,0,130,0,0,0,115,0,192,0,101,0,162,0,139,0,83,0,134,0,184,0,187,0,125,0,3,0,16,0,214,0,43,0,108,0,0,0,0,0,141,0,221,0,165,0,254,0,54,0,0,0,0,0,33,0,0,0,182,0,0,0,123,0,217,0,39,0,0,0,250,0,40,0,97,0,155,0,0,0,0,0,0,0,128,0,0,0,10,0,102,0,0,0,177,0,100,0,0,0,0,0,207,0,50,0,37,0,202,0,133,0,0,0,214,0,57,0,1,0,64,0,102,0,16,0,237,0,63,0,60,0,28,0,240,0,91,0,105,0,220,0,168,0,172,0,227,0,174,0,206,0,251,0,247,0,246,0,169,0,35,0,250,0,252,0,240,0);
signal scenario_full  : scenario_type := (161,31,70,31,9,31,136,31,233,31,106,31,237,31,40,31,239,31,142,31,19,31,221,31,221,30,97,31,234,31,103,31,103,30,103,29,44,31,41,31,133,31,133,30,216,31,184,31,145,31,204,31,229,31,68,31,68,30,234,31,49,31,149,31,149,30,166,31,3,31,107,31,107,30,127,31,127,30,164,31,164,30,143,31,90,31,90,30,69,31,194,31,19,31,160,31,141,31,60,31,76,31,2,31,2,30,2,29,6,31,6,30,196,31,133,31,5,31,92,31,121,31,114,31,74,31,194,31,226,31,65,31,9,31,100,31,154,31,199,31,199,30,118,31,43,31,43,30,27,31,148,31,227,31,25,31,42,31,203,31,72,31,179,31,179,30,93,31,41,31,61,31,61,30,123,31,123,30,123,29,40,31,72,31,72,30,79,31,115,31,62,31,57,31,72,31,72,30,214,31,83,31,41,31,127,31,130,31,130,30,152,31,1,31,115,31,17,31,17,30,15,31,15,30,228,31,61,31,191,31,245,31,203,31,145,31,92,31,206,31,201,31,201,30,150,31,87,31,137,31,221,31,221,30,200,31,8,31,6,31,234,31,210,31,59,31,71,31,10,31,10,30,148,31,37,31,37,30,31,31,31,30,136,31,136,30,35,31,107,31,107,30,234,31,16,31,16,30,242,31,84,31,251,31,150,31,112,31,178,31,232,31,27,31,145,31,234,31,139,31,139,30,25,31,181,31,91,31,81,31,174,31,241,31,162,31,35,31,107,31,107,30,236,31,236,30,27,31,131,31,66,31,140,31,152,31,19,31,80,31,80,30,21,31,21,30,191,31,53,31,232,31,198,31,17,31,17,30,149,31,28,31,91,31,90,31,3,31,124,31,124,30,163,31,88,31,40,31,146,31,123,31,191,31,165,31,168,31,88,31,224,31,209,31,209,30,190,31,92,31,99,31,108,31,100,31,33,31,147,31,123,31,69,31,69,30,187,31,64,31,3,31,9,31,53,31,172,31,149,31,149,30,233,31,69,31,69,31,208,31,61,31,29,31,169,31,169,30,100,31,36,31,198,31,246,31,6,31,187,31,251,31,251,30,4,31,35,31,146,31,125,31,82,31,82,30,180,31,180,30,91,31,214,31,176,31,64,31,64,30,121,31,212,31,66,31,249,31,161,31,91,31,98,31,98,30,98,29,98,28,135,31,16,31,58,31,58,30,91,31,91,30,91,29,91,28,109,31,46,31,114,31,114,30,157,31,249,31,249,30,51,31,7,31,61,31,97,31,188,31,188,30,131,31,158,31,105,31,224,31,136,31,61,31,115,31,115,30,19,31,19,30,19,29,195,31,195,30,195,29,195,28,136,31,136,30,169,31,197,31,203,31,203,30,203,29,232,31,3,31,89,31,91,31,156,31,40,31,115,31,22,31,126,31,126,30,153,31,54,31,54,30,1,31,1,30,1,29,28,31,61,31,85,31,85,31,162,31,94,31,81,31,115,31,148,31,206,31,68,31,45,31,45,30,35,31,122,31,122,30,40,31,114,31,114,30,114,29,224,31,103,31,33,31,97,31,248,31,22,31,250,31,22,31,136,31,40,31,186,31,13,31,112,31,127,31,130,31,130,30,214,31,214,30,175,31,147,31,147,30,92,31,222,31,222,30,20,31,89,31,76,31,116,31,115,31,243,31,7,31,25,31,76,31,202,31,202,30,171,31,231,31,132,31,153,31,135,31,135,30,122,31,244,31,130,31,161,31,4,31,110,31,13,31,121,31,251,31,179,31,151,31,162,31,255,31,14,31,243,31,82,31,82,30,44,31,182,31,41,31,41,30,29,31,25,31,69,31,92,31,115,31,219,31,100,31,1,31,219,31,140,31,82,31,171,31,36,31,227,31,181,31,215,31,18,31,215,31,186,31,70,31,89,31,89,30,84,31,84,30,48,31,165,31,18,31,1,31,1,30,92,31,199,31,90,31,87,31,119,31,54,31,115,31,77,31,181,31,40,31,193,31,117,31,71,31,71,30,98,31,255,31,61,31,93,31,58,31,234,31,17,31,68,31,199,31,215,31,215,30,194,31,44,31,44,30,68,31,129,31,164,31,150,31,57,31,185,31,7,31,185,31,197,31,157,31,189,31,126,31,126,30,217,31,138,31,138,30,187,31,127,31,127,30,174,31,63,31,63,30,63,29,63,28,87,31,172,31,147,31,130,31,130,30,115,31,192,31,101,31,162,31,139,31,83,31,134,31,184,31,187,31,125,31,3,31,16,31,214,31,43,31,108,31,108,30,108,29,141,31,221,31,165,31,254,31,54,31,54,30,54,29,33,31,33,30,182,31,182,30,123,31,217,31,39,31,39,30,250,31,40,31,97,31,155,31,155,30,155,29,155,28,128,31,128,30,10,31,102,31,102,30,177,31,100,31,100,30,100,29,207,31,50,31,37,31,202,31,133,31,133,30,214,31,57,31,1,31,64,31,102,31,16,31,237,31,63,31,60,31,28,31,240,31,91,31,105,31,220,31,168,31,172,31,227,31,174,31,206,31,251,31,247,31,246,31,169,31,35,31,250,31,252,31,240,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
