-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 934;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (127,0,31,0,10,0,86,0,254,0,221,0,0,0,196,0,0,0,36,0,231,0,46,0,175,0,0,0,212,0,171,0,174,0,0,0,220,0,168,0,56,0,204,0,219,0,0,0,0,0,245,0,178,0,0,0,0,0,232,0,115,0,234,0,225,0,94,0,24,0,250,0,99,0,66,0,18,0,132,0,177,0,84,0,99,0,65,0,119,0,89,0,105,0,95,0,251,0,136,0,0,0,122,0,0,0,2,0,6,0,0,0,175,0,235,0,192,0,42,0,149,0,0,0,30,0,32,0,183,0,147,0,0,0,207,0,14,0,0,0,153,0,175,0,5,0,110,0,104,0,39,0,118,0,254,0,227,0,0,0,0,0,181,0,202,0,129,0,248,0,127,0,0,0,121,0,161,0,0,0,75,0,0,0,30,0,196,0,78,0,110,0,0,0,41,0,39,0,52,0,62,0,229,0,227,0,182,0,99,0,119,0,227,0,68,0,163,0,0,0,0,0,90,0,13,0,66,0,25,0,0,0,0,0,0,0,188,0,106,0,253,0,122,0,83,0,222,0,81,0,246,0,170,0,143,0,0,0,107,0,45,0,95,0,82,0,107,0,1,0,0,0,0,0,211,0,0,0,148,0,232,0,0,0,141,0,157,0,0,0,36,0,239,0,166,0,0,0,0,0,255,0,0,0,164,0,0,0,7,0,142,0,0,0,219,0,253,0,116,0,0,0,0,0,27,0,6,0,69,0,0,0,68,0,119,0,0,0,0,0,27,0,18,0,113,0,43,0,114,0,169,0,136,0,14,0,178,0,140,0,204,0,55,0,23,0,0,0,16,0,189,0,58,0,18,0,0,0,230,0,121,0,96,0,189,0,145,0,149,0,50,0,0,0,6,0,112,0,176,0,146,0,0,0,0,0,0,0,156,0,176,0,111,0,89,0,113,0,40,0,169,0,156,0,118,0,170,0,244,0,188,0,138,0,34,0,0,0,63,0,183,0,249,0,150,0,4,0,0,0,0,0,0,0,246,0,0,0,135,0,215,0,98,0,226,0,0,0,157,0,221,0,134,0,42,0,182,0,145,0,0,0,0,0,0,0,239,0,19,0,182,0,0,0,15,0,166,0,119,0,243,0,203,0,0,0,57,0,0,0,0,0,31,0,157,0,0,0,192,0,200,0,44,0,26,0,0,0,246,0,215,0,164,0,6,0,0,0,140,0,0,0,219,0,130,0,243,0,4,0,73,0,64,0,5,0,0,0,52,0,0,0,132,0,249,0,0,0,121,0,21,0,98,0,146,0,24,0,4,0,133,0,0,0,161,0,0,0,119,0,0,0,54,0,170,0,0,0,85,0,189,0,183,0,234,0,164,0,29,0,0,0,133,0,0,0,0,0,203,0,0,0,119,0,0,0,16,0,241,0,69,0,113,0,101,0,77,0,0,0,0,0,3,0,139,0,187,0,88,0,0,0,31,0,68,0,123,0,0,0,87,0,82,0,188,0,0,0,0,0,252,0,4,0,0,0,144,0,0,0,125,0,200,0,162,0,251,0,83,0,248,0,234,0,73,0,0,0,132,0,161,0,231,0,155,0,21,0,34,0,0,0,122,0,127,0,30,0,96,0,102,0,223,0,183,0,152,0,218,0,250,0,50,0,0,0,195,0,0,0,234,0,128,0,50,0,200,0,126,0,4,0,153,0,160,0,0,0,170,0,144,0,240,0,18,0,60,0,65,0,1,0,3,0,0,0,0,0,15,0,0,0,0,0,162,0,22,0,0,0,173,0,104,0,0,0,218,0,219,0,62,0,177,0,221,0,0,0,241,0,204,0,174,0,0,0,114,0,121,0,251,0,117,0,58,0,148,0,0,0,0,0,87,0,0,0,235,0,10,0,223,0,13,0,63,0,96,0,231,0,48,0,235,0,26,0,140,0,70,0,59,0,127,0,121,0,0,0,108,0,167,0,0,0,110,0,0,0,137,0,230,0,163,0,28,0,120,0,158,0,96,0,87,0,0,0,54,0,70,0,95,0,163,0,200,0,183,0,0,0,51,0,39,0,15,0,130,0,188,0,0,0,0,0,164,0,61,0,0,0,0,0,94,0,55,0,2,0,69,0,0,0,74,0,161,0,190,0,0,0,76,0,155,0,0,0,0,0,7,0,209,0,26,0,75,0,194,0,77,0,233,0,251,0,229,0,145,0,156,0,133,0,23,0,7,0,61,0,17,0,139,0,127,0,140,0,0,0,92,0,94,0,42,0,119,0,185,0,105,0,24,0,249,0,132,0,0,0,61,0,228,0,219,0,121,0,0,0,191,0,28,0,228,0,0,0,0,0,249,0,66,0,131,0,222,0,193,0,0,0,226,0,102,0,117,0,0,0,182,0,99,0,167,0,0,0,162,0,105,0,129,0,237,0,41,0,130,0,29,0,131,0,0,0,105,0,76,0,94,0,0,0,244,0,131,0,88,0,98,0,14,0,0,0,47,0,68,0,141,0,232,0,144,0,10,0,42,0,77,0,130,0,217,0,40,0,100,0,1,0,205,0,0,0,209,0,0,0,209,0,83,0,0,0,32,0,84,0,160,0,155,0,145,0,167,0,247,0,209,0,154,0,244,0,140,0,232,0,99,0,4,0,105,0,214,0,205,0,254,0,0,0,176,0,0,0,241,0,102,0,85,0,161,0,244,0,121,0,44,0,203,0,0,0,151,0,116,0,18,0,76,0,186,0,188,0,0,0,39,0,0,0,202,0,204,0,0,0,0,0,0,0,0,0,41,0,128,0,244,0,176,0,114,0,229,0,60,0,254,0,187,0,10,0,45,0,172,0,172,0,175,0,204,0,173,0,164,0,61,0,0,0,0,0,250,0,89,0,0,0,240,0,67,0,75,0,63,0,0,0,51,0,123,0,82,0,137,0,17,0,159,0,0,0,82,0,246,0,5,0,0,0,22,0,49,0,0,0,139,0,201,0,193,0,147,0,16,0,156,0,129,0,0,0,224,0,160,0,111,0,47,0,58,0,255,0,8,0,123,0,37,0,0,0,0,0,29,0,0,0,24,0,40,0,201,0,214,0,80,0,244,0,0,0,237,0,0,0,0,0,234,0,106,0,0,0,0,0,0,0,76,0,29,0,37,0,6,0,163,0,128,0,0,0,0,0,0,0,32,0,15,0,71,0,184,0,0,0,104,0,0,0,4,0,160,0,93,0,81,0,174,0,58,0,223,0,0,0,147,0,17,0,178,0,235,0,0,0,0,0,19,0,0,0,147,0,170,0,121,0,83,0,42,0,237,0,0,0,86,0,75,0,169,0,58,0,0,0,103,0,201,0,73,0,159,0,41,0,58,0,0,0,88,0,46,0,16,0,0,0,0,0,86,0,235,0,50,0,127,0,0,0,42,0,246,0,0,0,220,0,183,0,189,0,0,0,129,0,189,0,98,0,226,0,0,0,117,0,57,0,0,0,97,0,244,0,202,0,162,0,121,0,30,0,220,0,176,0,138,0,104,0,147,0,0,0,201,0,42,0,0,0,0,0,101,0,0,0,159,0,23,0,248,0,216,0,129,0,136,0,204,0,36,0,156,0,170,0,61,0,129,0,174,0,49,0,124,0,66,0,124,0,36,0,211,0,137,0,44,0,220,0,91,0,86,0,105,0,58,0,0,0,215,0,179,0,0,0,0,0,22,0,0,0,181,0,5,0,208,0,0,0,11,0,214,0,68,0,0,0,35,0,0,0,17,0,227,0,186,0,0,0,0,0,0,0,239,0,94,0,160,0,13,0,201,0,111,0,0,0,12,0,207,0,161,0,219,0,0,0,239,0,213,0,40,0,0,0,192,0,144,0,98,0,0,0,122,0,66,0,98,0,20,0,5,0,96,0,24,0,119,0,0,0,184,0,237,0,253,0,160,0,71,0,116,0,7,0,114,0,133,0,165,0,0,0,68,0,241,0,201,0,149,0,94,0,123,0,245,0,53,0,0,0,25,0,0,0,9,0,244,0,0,0,114,0,0,0,172,0,141,0,0,0,129,0,240,0,166,0,139,0,169,0,140,0,175,0,0,0,0,0,120,0,0,0,14,0,0,0,94,0,164,0,0,0,116,0,96,0,152,0,46,0,0,0,42,0,246,0,103,0,179,0,10,0,217,0,14,0,0,0,98,0,0,0,95,0,80,0,87,0,68,0,0,0,0,0);
signal scenario_full  : scenario_type := (127,31,31,31,10,31,86,31,254,31,221,31,221,30,196,31,196,30,36,31,231,31,46,31,175,31,175,30,212,31,171,31,174,31,174,30,220,31,168,31,56,31,204,31,219,31,219,30,219,29,245,31,178,31,178,30,178,29,232,31,115,31,234,31,225,31,94,31,24,31,250,31,99,31,66,31,18,31,132,31,177,31,84,31,99,31,65,31,119,31,89,31,105,31,95,31,251,31,136,31,136,30,122,31,122,30,2,31,6,31,6,30,175,31,235,31,192,31,42,31,149,31,149,30,30,31,32,31,183,31,147,31,147,30,207,31,14,31,14,30,153,31,175,31,5,31,110,31,104,31,39,31,118,31,254,31,227,31,227,30,227,29,181,31,202,31,129,31,248,31,127,31,127,30,121,31,161,31,161,30,75,31,75,30,30,31,196,31,78,31,110,31,110,30,41,31,39,31,52,31,62,31,229,31,227,31,182,31,99,31,119,31,227,31,68,31,163,31,163,30,163,29,90,31,13,31,66,31,25,31,25,30,25,29,25,28,188,31,106,31,253,31,122,31,83,31,222,31,81,31,246,31,170,31,143,31,143,30,107,31,45,31,95,31,82,31,107,31,1,31,1,30,1,29,211,31,211,30,148,31,232,31,232,30,141,31,157,31,157,30,36,31,239,31,166,31,166,30,166,29,255,31,255,30,164,31,164,30,7,31,142,31,142,30,219,31,253,31,116,31,116,30,116,29,27,31,6,31,69,31,69,30,68,31,119,31,119,30,119,29,27,31,18,31,113,31,43,31,114,31,169,31,136,31,14,31,178,31,140,31,204,31,55,31,23,31,23,30,16,31,189,31,58,31,18,31,18,30,230,31,121,31,96,31,189,31,145,31,149,31,50,31,50,30,6,31,112,31,176,31,146,31,146,30,146,29,146,28,156,31,176,31,111,31,89,31,113,31,40,31,169,31,156,31,118,31,170,31,244,31,188,31,138,31,34,31,34,30,63,31,183,31,249,31,150,31,4,31,4,30,4,29,4,28,246,31,246,30,135,31,215,31,98,31,226,31,226,30,157,31,221,31,134,31,42,31,182,31,145,31,145,30,145,29,145,28,239,31,19,31,182,31,182,30,15,31,166,31,119,31,243,31,203,31,203,30,57,31,57,30,57,29,31,31,157,31,157,30,192,31,200,31,44,31,26,31,26,30,246,31,215,31,164,31,6,31,6,30,140,31,140,30,219,31,130,31,243,31,4,31,73,31,64,31,5,31,5,30,52,31,52,30,132,31,249,31,249,30,121,31,21,31,98,31,146,31,24,31,4,31,133,31,133,30,161,31,161,30,119,31,119,30,54,31,170,31,170,30,85,31,189,31,183,31,234,31,164,31,29,31,29,30,133,31,133,30,133,29,203,31,203,30,119,31,119,30,16,31,241,31,69,31,113,31,101,31,77,31,77,30,77,29,3,31,139,31,187,31,88,31,88,30,31,31,68,31,123,31,123,30,87,31,82,31,188,31,188,30,188,29,252,31,4,31,4,30,144,31,144,30,125,31,200,31,162,31,251,31,83,31,248,31,234,31,73,31,73,30,132,31,161,31,231,31,155,31,21,31,34,31,34,30,122,31,127,31,30,31,96,31,102,31,223,31,183,31,152,31,218,31,250,31,50,31,50,30,195,31,195,30,234,31,128,31,50,31,200,31,126,31,4,31,153,31,160,31,160,30,170,31,144,31,240,31,18,31,60,31,65,31,1,31,3,31,3,30,3,29,15,31,15,30,15,29,162,31,22,31,22,30,173,31,104,31,104,30,218,31,219,31,62,31,177,31,221,31,221,30,241,31,204,31,174,31,174,30,114,31,121,31,251,31,117,31,58,31,148,31,148,30,148,29,87,31,87,30,235,31,10,31,223,31,13,31,63,31,96,31,231,31,48,31,235,31,26,31,140,31,70,31,59,31,127,31,121,31,121,30,108,31,167,31,167,30,110,31,110,30,137,31,230,31,163,31,28,31,120,31,158,31,96,31,87,31,87,30,54,31,70,31,95,31,163,31,200,31,183,31,183,30,51,31,39,31,15,31,130,31,188,31,188,30,188,29,164,31,61,31,61,30,61,29,94,31,55,31,2,31,69,31,69,30,74,31,161,31,190,31,190,30,76,31,155,31,155,30,155,29,7,31,209,31,26,31,75,31,194,31,77,31,233,31,251,31,229,31,145,31,156,31,133,31,23,31,7,31,61,31,17,31,139,31,127,31,140,31,140,30,92,31,94,31,42,31,119,31,185,31,105,31,24,31,249,31,132,31,132,30,61,31,228,31,219,31,121,31,121,30,191,31,28,31,228,31,228,30,228,29,249,31,66,31,131,31,222,31,193,31,193,30,226,31,102,31,117,31,117,30,182,31,99,31,167,31,167,30,162,31,105,31,129,31,237,31,41,31,130,31,29,31,131,31,131,30,105,31,76,31,94,31,94,30,244,31,131,31,88,31,98,31,14,31,14,30,47,31,68,31,141,31,232,31,144,31,10,31,42,31,77,31,130,31,217,31,40,31,100,31,1,31,205,31,205,30,209,31,209,30,209,31,83,31,83,30,32,31,84,31,160,31,155,31,145,31,167,31,247,31,209,31,154,31,244,31,140,31,232,31,99,31,4,31,105,31,214,31,205,31,254,31,254,30,176,31,176,30,241,31,102,31,85,31,161,31,244,31,121,31,44,31,203,31,203,30,151,31,116,31,18,31,76,31,186,31,188,31,188,30,39,31,39,30,202,31,204,31,204,30,204,29,204,28,204,27,41,31,128,31,244,31,176,31,114,31,229,31,60,31,254,31,187,31,10,31,45,31,172,31,172,31,175,31,204,31,173,31,164,31,61,31,61,30,61,29,250,31,89,31,89,30,240,31,67,31,75,31,63,31,63,30,51,31,123,31,82,31,137,31,17,31,159,31,159,30,82,31,246,31,5,31,5,30,22,31,49,31,49,30,139,31,201,31,193,31,147,31,16,31,156,31,129,31,129,30,224,31,160,31,111,31,47,31,58,31,255,31,8,31,123,31,37,31,37,30,37,29,29,31,29,30,24,31,40,31,201,31,214,31,80,31,244,31,244,30,237,31,237,30,237,29,234,31,106,31,106,30,106,29,106,28,76,31,29,31,37,31,6,31,163,31,128,31,128,30,128,29,128,28,32,31,15,31,71,31,184,31,184,30,104,31,104,30,4,31,160,31,93,31,81,31,174,31,58,31,223,31,223,30,147,31,17,31,178,31,235,31,235,30,235,29,19,31,19,30,147,31,170,31,121,31,83,31,42,31,237,31,237,30,86,31,75,31,169,31,58,31,58,30,103,31,201,31,73,31,159,31,41,31,58,31,58,30,88,31,46,31,16,31,16,30,16,29,86,31,235,31,50,31,127,31,127,30,42,31,246,31,246,30,220,31,183,31,189,31,189,30,129,31,189,31,98,31,226,31,226,30,117,31,57,31,57,30,97,31,244,31,202,31,162,31,121,31,30,31,220,31,176,31,138,31,104,31,147,31,147,30,201,31,42,31,42,30,42,29,101,31,101,30,159,31,23,31,248,31,216,31,129,31,136,31,204,31,36,31,156,31,170,31,61,31,129,31,174,31,49,31,124,31,66,31,124,31,36,31,211,31,137,31,44,31,220,31,91,31,86,31,105,31,58,31,58,30,215,31,179,31,179,30,179,29,22,31,22,30,181,31,5,31,208,31,208,30,11,31,214,31,68,31,68,30,35,31,35,30,17,31,227,31,186,31,186,30,186,29,186,28,239,31,94,31,160,31,13,31,201,31,111,31,111,30,12,31,207,31,161,31,219,31,219,30,239,31,213,31,40,31,40,30,192,31,144,31,98,31,98,30,122,31,66,31,98,31,20,31,5,31,96,31,24,31,119,31,119,30,184,31,237,31,253,31,160,31,71,31,116,31,7,31,114,31,133,31,165,31,165,30,68,31,241,31,201,31,149,31,94,31,123,31,245,31,53,31,53,30,25,31,25,30,9,31,244,31,244,30,114,31,114,30,172,31,141,31,141,30,129,31,240,31,166,31,139,31,169,31,140,31,175,31,175,30,175,29,120,31,120,30,14,31,14,30,94,31,164,31,164,30,116,31,96,31,152,31,46,31,46,30,42,31,246,31,103,31,179,31,10,31,217,31,14,31,14,30,98,31,98,30,95,31,80,31,87,31,68,31,68,30,68,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
