-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 664;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (151,0,186,0,0,0,0,0,107,0,0,0,255,0,0,0,0,0,60,0,0,0,0,0,21,0,188,0,150,0,0,0,76,0,123,0,0,0,248,0,109,0,226,0,0,0,11,0,164,0,220,0,70,0,0,0,239,0,184,0,242,0,34,0,79,0,78,0,105,0,106,0,0,0,219,0,119,0,173,0,199,0,88,0,104,0,35,0,240,0,55,0,48,0,0,0,216,0,95,0,75,0,222,0,210,0,248,0,30,0,184,0,10,0,207,0,176,0,0,0,235,0,32,0,30,0,180,0,138,0,75,0,10,0,0,0,132,0,230,0,107,0,205,0,133,0,145,0,0,0,253,0,93,0,138,0,214,0,30,0,0,0,0,0,34,0,86,0,0,0,0,0,0,0,77,0,157,0,62,0,51,0,117,0,45,0,175,0,26,0,80,0,0,0,194,0,0,0,2,0,211,0,149,0,106,0,187,0,223,0,12,0,7,0,168,0,250,0,131,0,10,0,130,0,161,0,255,0,221,0,60,0,95,0,7,0,141,0,0,0,127,0,227,0,152,0,198,0,211,0,110,0,162,0,177,0,118,0,169,0,26,0,12,0,0,0,131,0,32,0,0,0,0,0,0,0,213,0,6,0,123,0,25,0,12,0,84,0,211,0,143,0,185,0,4,0,56,0,182,0,180,0,193,0,102,0,10,0,83,0,108,0,0,0,0,0,71,0,132,0,98,0,187,0,51,0,192,0,90,0,41,0,194,0,0,0,47,0,4,0,207,0,219,0,42,0,122,0,0,0,19,0,0,0,230,0,0,0,219,0,82,0,138,0,237,0,47,0,202,0,86,0,77,0,160,0,0,0,63,0,136,0,0,0,86,0,182,0,78,0,220,0,222,0,203,0,122,0,234,0,11,0,237,0,179,0,198,0,172,0,113,0,195,0,35,0,15,0,170,0,68,0,156,0,85,0,129,0,63,0,154,0,246,0,10,0,0,0,109,0,0,0,253,0,53,0,247,0,132,0,196,0,186,0,206,0,0,0,186,0,176,0,81,0,43,0,194,0,0,0,0,0,0,0,0,0,2,0,220,0,124,0,130,0,0,0,97,0,199,0,190,0,141,0,112,0,46,0,194,0,202,0,133,0,108,0,55,0,12,0,29,0,126,0,118,0,0,0,138,0,82,0,0,0,77,0,0,0,74,0,231,0,15,0,53,0,156,0,158,0,179,0,56,0,0,0,56,0,194,0,54,0,28,0,87,0,7,0,0,0,127,0,55,0,0,0,50,0,14,0,35,0,63,0,169,0,215,0,250,0,134,0,199,0,210,0,26,0,146,0,95,0,161,0,221,0,145,0,5,0,0,0,0,0,191,0,111,0,0,0,251,0,133,0,84,0,71,0,189,0,0,0,8,0,0,0,0,0,43,0,7,0,16,0,145,0,57,0,0,0,30,0,157,0,208,0,212,0,137,0,0,0,0,0,0,0,82,0,138,0,77,0,76,0,136,0,107,0,227,0,4,0,204,0,205,0,10,0,230,0,248,0,0,0,156,0,36,0,55,0,93,0,0,0,196,0,0,0,63,0,0,0,38,0,0,0,120,0,68,0,227,0,62,0,0,0,59,0,5,0,171,0,33,0,71,0,0,0,30,0,244,0,241,0,183,0,173,0,122,0,0,0,208,0,129,0,121,0,0,0,0,0,67,0,131,0,207,0,0,0,0,0,248,0,187,0,89,0,112,0,233,0,149,0,133,0,0,0,34,0,233,0,0,0,151,0,29,0,191,0,0,0,45,0,0,0,203,0,126,0,153,0,250,0,189,0,208,0,168,0,233,0,194,0,241,0,41,0,248,0,246,0,49,0,224,0,106,0,142,0,0,0,199,0,100,0,34,0,115,0,201,0,235,0,0,0,112,0,161,0,18,0,0,0,210,0,228,0,165,0,0,0,78,0,181,0,206,0,218,0,0,0,10,0,27,0,100,0,234,0,26,0,35,0,47,0,174,0,111,0,41,0,83,0,79,0,0,0,159,0,12,0,17,0,69,0,92,0,115,0,0,0,0,0,65,0,0,0,121,0,119,0,28,0,0,0,210,0,0,0,215,0,219,0,48,0,29,0,10,0,47,0,128,0,234,0,144,0,0,0,33,0,0,0,115,0,56,0,0,0,108,0,63,0,0,0,137,0,0,0,227,0,205,0,0,0,116,0,55,0,181,0,82,0,51,0,58,0,138,0,228,0,210,0,247,0,14,0,183,0,14,0,0,0,103,0,86,0,1,0,207,0,147,0,115,0,245,0,201,0,135,0,220,0,129,0,64,0,230,0,167,0,51,0,197,0,4,0,247,0,0,0,54,0,251,0,0,0,245,0,67,0,248,0,93,0,186,0,0,0,0,0,0,0,112,0,0,0,0,0,0,0,157,0,239,0,73,0,0,0,16,0,30,0,131,0,178,0,204,0,223,0,166,0,49,0,49,0,0,0,250,0,90,0,165,0,0,0,199,0,0,0,107,0,88,0,172,0,247,0,27,0,23,0,85,0,190,0,0,0,147,0,97,0,202,0,116,0,4,0,154,0,0,0,120,0,254,0,0,0,19,0,0,0,0,0,135,0,202,0,6,0,179,0,135,0,108,0,154,0,81,0,187,0,237,0,74,0,0,0,125,0,230,0,172,0,0,0,191,0,63,0,120,0,253,0,112,0,188,0,113,0,204,0,48,0,81,0,107,0,207,0,73,0,51,0,114,0,229,0,80,0,97,0,222,0,158,0,56,0,240,0,103,0,43,0,151,0,228,0,192,0,99,0,200,0,63,0,170,0,100,0,208,0,127,0,0,0,96,0,5,0,162,0,157,0,22,0,30,0,36,0,199,0,248,0,0,0,0,0,176,0,0,0,127,0,0,0,70,0,250,0,216,0,45,0,117,0,230,0,0,0,15,0,226,0,26,0,68,0,22,0,51,0,0,0,131,0,218,0,124,0,0,0,184,0,251,0);
signal scenario_full  : scenario_type := (151,31,186,31,186,30,186,29,107,31,107,30,255,31,255,30,255,29,60,31,60,30,60,29,21,31,188,31,150,31,150,30,76,31,123,31,123,30,248,31,109,31,226,31,226,30,11,31,164,31,220,31,70,31,70,30,239,31,184,31,242,31,34,31,79,31,78,31,105,31,106,31,106,30,219,31,119,31,173,31,199,31,88,31,104,31,35,31,240,31,55,31,48,31,48,30,216,31,95,31,75,31,222,31,210,31,248,31,30,31,184,31,10,31,207,31,176,31,176,30,235,31,32,31,30,31,180,31,138,31,75,31,10,31,10,30,132,31,230,31,107,31,205,31,133,31,145,31,145,30,253,31,93,31,138,31,214,31,30,31,30,30,30,29,34,31,86,31,86,30,86,29,86,28,77,31,157,31,62,31,51,31,117,31,45,31,175,31,26,31,80,31,80,30,194,31,194,30,2,31,211,31,149,31,106,31,187,31,223,31,12,31,7,31,168,31,250,31,131,31,10,31,130,31,161,31,255,31,221,31,60,31,95,31,7,31,141,31,141,30,127,31,227,31,152,31,198,31,211,31,110,31,162,31,177,31,118,31,169,31,26,31,12,31,12,30,131,31,32,31,32,30,32,29,32,28,213,31,6,31,123,31,25,31,12,31,84,31,211,31,143,31,185,31,4,31,56,31,182,31,180,31,193,31,102,31,10,31,83,31,108,31,108,30,108,29,71,31,132,31,98,31,187,31,51,31,192,31,90,31,41,31,194,31,194,30,47,31,4,31,207,31,219,31,42,31,122,31,122,30,19,31,19,30,230,31,230,30,219,31,82,31,138,31,237,31,47,31,202,31,86,31,77,31,160,31,160,30,63,31,136,31,136,30,86,31,182,31,78,31,220,31,222,31,203,31,122,31,234,31,11,31,237,31,179,31,198,31,172,31,113,31,195,31,35,31,15,31,170,31,68,31,156,31,85,31,129,31,63,31,154,31,246,31,10,31,10,30,109,31,109,30,253,31,53,31,247,31,132,31,196,31,186,31,206,31,206,30,186,31,176,31,81,31,43,31,194,31,194,30,194,29,194,28,194,27,2,31,220,31,124,31,130,31,130,30,97,31,199,31,190,31,141,31,112,31,46,31,194,31,202,31,133,31,108,31,55,31,12,31,29,31,126,31,118,31,118,30,138,31,82,31,82,30,77,31,77,30,74,31,231,31,15,31,53,31,156,31,158,31,179,31,56,31,56,30,56,31,194,31,54,31,28,31,87,31,7,31,7,30,127,31,55,31,55,30,50,31,14,31,35,31,63,31,169,31,215,31,250,31,134,31,199,31,210,31,26,31,146,31,95,31,161,31,221,31,145,31,5,31,5,30,5,29,191,31,111,31,111,30,251,31,133,31,84,31,71,31,189,31,189,30,8,31,8,30,8,29,43,31,7,31,16,31,145,31,57,31,57,30,30,31,157,31,208,31,212,31,137,31,137,30,137,29,137,28,82,31,138,31,77,31,76,31,136,31,107,31,227,31,4,31,204,31,205,31,10,31,230,31,248,31,248,30,156,31,36,31,55,31,93,31,93,30,196,31,196,30,63,31,63,30,38,31,38,30,120,31,68,31,227,31,62,31,62,30,59,31,5,31,171,31,33,31,71,31,71,30,30,31,244,31,241,31,183,31,173,31,122,31,122,30,208,31,129,31,121,31,121,30,121,29,67,31,131,31,207,31,207,30,207,29,248,31,187,31,89,31,112,31,233,31,149,31,133,31,133,30,34,31,233,31,233,30,151,31,29,31,191,31,191,30,45,31,45,30,203,31,126,31,153,31,250,31,189,31,208,31,168,31,233,31,194,31,241,31,41,31,248,31,246,31,49,31,224,31,106,31,142,31,142,30,199,31,100,31,34,31,115,31,201,31,235,31,235,30,112,31,161,31,18,31,18,30,210,31,228,31,165,31,165,30,78,31,181,31,206,31,218,31,218,30,10,31,27,31,100,31,234,31,26,31,35,31,47,31,174,31,111,31,41,31,83,31,79,31,79,30,159,31,12,31,17,31,69,31,92,31,115,31,115,30,115,29,65,31,65,30,121,31,119,31,28,31,28,30,210,31,210,30,215,31,219,31,48,31,29,31,10,31,47,31,128,31,234,31,144,31,144,30,33,31,33,30,115,31,56,31,56,30,108,31,63,31,63,30,137,31,137,30,227,31,205,31,205,30,116,31,55,31,181,31,82,31,51,31,58,31,138,31,228,31,210,31,247,31,14,31,183,31,14,31,14,30,103,31,86,31,1,31,207,31,147,31,115,31,245,31,201,31,135,31,220,31,129,31,64,31,230,31,167,31,51,31,197,31,4,31,247,31,247,30,54,31,251,31,251,30,245,31,67,31,248,31,93,31,186,31,186,30,186,29,186,28,112,31,112,30,112,29,112,28,157,31,239,31,73,31,73,30,16,31,30,31,131,31,178,31,204,31,223,31,166,31,49,31,49,31,49,30,250,31,90,31,165,31,165,30,199,31,199,30,107,31,88,31,172,31,247,31,27,31,23,31,85,31,190,31,190,30,147,31,97,31,202,31,116,31,4,31,154,31,154,30,120,31,254,31,254,30,19,31,19,30,19,29,135,31,202,31,6,31,179,31,135,31,108,31,154,31,81,31,187,31,237,31,74,31,74,30,125,31,230,31,172,31,172,30,191,31,63,31,120,31,253,31,112,31,188,31,113,31,204,31,48,31,81,31,107,31,207,31,73,31,51,31,114,31,229,31,80,31,97,31,222,31,158,31,56,31,240,31,103,31,43,31,151,31,228,31,192,31,99,31,200,31,63,31,170,31,100,31,208,31,127,31,127,30,96,31,5,31,162,31,157,31,22,31,30,31,36,31,199,31,248,31,248,30,248,29,176,31,176,30,127,31,127,30,70,31,250,31,216,31,45,31,117,31,230,31,230,30,15,31,226,31,26,31,68,31,22,31,51,31,51,30,131,31,218,31,124,31,124,30,184,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
