-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 303;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (129,0,95,0,149,0,178,0,143,0,102,0,124,0,159,0,63,0,0,0,0,0,40,0,114,0,54,0,188,0,0,0,156,0,111,0,196,0,201,0,38,0,105,0,90,0,238,0,172,0,0,0,117,0,102,0,196,0,131,0,209,0,198,0,126,0,191,0,121,0,251,0,207,0,112,0,79,0,61,0,34,0,0,0,0,0,69,0,63,0,58,0,0,0,144,0,34,0,57,0,247,0,179,0,86,0,108,0,127,0,119,0,136,0,0,0,30,0,48,0,141,0,167,0,42,0,85,0,186,0,0,0,15,0,232,0,0,0,180,0,150,0,93,0,0,0,188,0,30,0,197,0,173,0,66,0,126,0,0,0,197,0,45,0,160,0,138,0,140,0,192,0,180,0,255,0,231,0,112,0,97,0,0,0,118,0,8,0,27,0,222,0,83,0,229,0,9,0,212,0,243,0,170,0,0,0,24,0,0,0,88,0,157,0,240,0,146,0,0,0,126,0,0,0,230,0,136,0,12,0,176,0,49,0,133,0,12,0,231,0,0,0,103,0,224,0,0,0,226,0,103,0,35,0,0,0,0,0,72,0,92,0,233,0,37,0,207,0,0,0,70,0,156,0,156,0,220,0,229,0,0,0,75,0,249,0,0,0,0,0,47,0,11,0,59,0,10,0,8,0,180,0,0,0,190,0,246,0,217,0,0,0,98,0,187,0,4,0,105,0,0,0,43,0,200,0,65,0,70,0,48,0,169,0,156,0,232,0,199,0,181,0,238,0,38,0,229,0,105,0,238,0,0,0,74,0,0,0,0,0,31,0,251,0,147,0,219,0,188,0,0,0,17,0,112,0,0,0,178,0,0,0,158,0,174,0,122,0,216,0,0,0,42,0,165,0,227,0,237,0,168,0,0,0,186,0,41,0,235,0,162,0,168,0,79,0,222,0,0,0,103,0,0,0,195,0,101,0,133,0,46,0,38,0,0,0,249,0,23,0,0,0,159,0,216,0,112,0,204,0,16,0,107,0,9,0,6,0,251,0,63,0,200,0,0,0,26,0,97,0,219,0,124,0,24,0,102,0,252,0,180,0,253,0,0,0,0,0,105,0,71,0,142,0,234,0,110,0,242,0,21,0,254,0,227,0,27,0,0,0,235,0,218,0,0,0,88,0,57,0,0,0,0,0,145,0,0,0,0,0,0,0,88,0,187,0,180,0,13,0,80,0,105,0,149,0,72,0,112,0,0,0,25,0,68,0,69,0,87,0,115,0,0,0,33,0,157,0,19,0,0,0,113,0,0,0,9,0,62,0,129,0,239,0,51,0,119,0,0,0,112,0,0,0,239,0,2,0,50,0,61,0,81,0,201,0);
signal scenario_full  : scenario_type := (129,31,95,31,149,31,178,31,143,31,102,31,124,31,159,31,63,31,63,30,63,29,40,31,114,31,54,31,188,31,188,30,156,31,111,31,196,31,201,31,38,31,105,31,90,31,238,31,172,31,172,30,117,31,102,31,196,31,131,31,209,31,198,31,126,31,191,31,121,31,251,31,207,31,112,31,79,31,61,31,34,31,34,30,34,29,69,31,63,31,58,31,58,30,144,31,34,31,57,31,247,31,179,31,86,31,108,31,127,31,119,31,136,31,136,30,30,31,48,31,141,31,167,31,42,31,85,31,186,31,186,30,15,31,232,31,232,30,180,31,150,31,93,31,93,30,188,31,30,31,197,31,173,31,66,31,126,31,126,30,197,31,45,31,160,31,138,31,140,31,192,31,180,31,255,31,231,31,112,31,97,31,97,30,118,31,8,31,27,31,222,31,83,31,229,31,9,31,212,31,243,31,170,31,170,30,24,31,24,30,88,31,157,31,240,31,146,31,146,30,126,31,126,30,230,31,136,31,12,31,176,31,49,31,133,31,12,31,231,31,231,30,103,31,224,31,224,30,226,31,103,31,35,31,35,30,35,29,72,31,92,31,233,31,37,31,207,31,207,30,70,31,156,31,156,31,220,31,229,31,229,30,75,31,249,31,249,30,249,29,47,31,11,31,59,31,10,31,8,31,180,31,180,30,190,31,246,31,217,31,217,30,98,31,187,31,4,31,105,31,105,30,43,31,200,31,65,31,70,31,48,31,169,31,156,31,232,31,199,31,181,31,238,31,38,31,229,31,105,31,238,31,238,30,74,31,74,30,74,29,31,31,251,31,147,31,219,31,188,31,188,30,17,31,112,31,112,30,178,31,178,30,158,31,174,31,122,31,216,31,216,30,42,31,165,31,227,31,237,31,168,31,168,30,186,31,41,31,235,31,162,31,168,31,79,31,222,31,222,30,103,31,103,30,195,31,101,31,133,31,46,31,38,31,38,30,249,31,23,31,23,30,159,31,216,31,112,31,204,31,16,31,107,31,9,31,6,31,251,31,63,31,200,31,200,30,26,31,97,31,219,31,124,31,24,31,102,31,252,31,180,31,253,31,253,30,253,29,105,31,71,31,142,31,234,31,110,31,242,31,21,31,254,31,227,31,27,31,27,30,235,31,218,31,218,30,88,31,57,31,57,30,57,29,145,31,145,30,145,29,145,28,88,31,187,31,180,31,13,31,80,31,105,31,149,31,72,31,112,31,112,30,25,31,68,31,69,31,87,31,115,31,115,30,33,31,157,31,19,31,19,30,113,31,113,30,9,31,62,31,129,31,239,31,51,31,119,31,119,30,112,31,112,30,239,31,2,31,50,31,61,31,81,31,201,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
