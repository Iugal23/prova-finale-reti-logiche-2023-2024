-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 330;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,0,0,13,0,0,0,0,0,56,0,46,0,0,0,119,0,97,0,198,0,132,0,251,0,152,0,36,0,26,0,100,0,0,0,79,0,157,0,103,0,0,0,151,0,47,0,101,0,251,0,50,0,230,0,208,0,189,0,14,0,139,0,0,0,0,0,175,0,4,0,0,0,208,0,215,0,96,0,245,0,7,0,174,0,169,0,93,0,232,0,151,0,16,0,20,0,211,0,157,0,181,0,0,0,111,0,0,0,0,0,225,0,101,0,7,0,90,0,23,0,183,0,214,0,93,0,77,0,163,0,219,0,207,0,196,0,198,0,15,0,146,0,0,0,154,0,72,0,0,0,27,0,0,0,171,0,183,0,141,0,121,0,151,0,241,0,231,0,0,0,222,0,171,0,223,0,43,0,0,0,196,0,38,0,192,0,79,0,86,0,157,0,0,0,49,0,112,0,192,0,0,0,0,0,54,0,159,0,185,0,0,0,231,0,91,0,0,0,253,0,233,0,249,0,117,0,158,0,130,0,0,0,89,0,25,0,159,0,68,0,139,0,35,0,156,0,0,0,179,0,108,0,216,0,91,0,55,0,113,0,189,0,0,0,182,0,18,0,127,0,178,0,207,0,115,0,120,0,244,0,92,0,0,0,26,0,0,0,166,0,240,0,0,0,0,0,22,0,193,0,11,0,187,0,116,0,53,0,24,0,53,0,57,0,201,0,206,0,0,0,21,0,0,0,87,0,0,0,126,0,0,0,91,0,0,0,137,0,0,0,0,0,255,0,203,0,0,0,252,0,50,0,49,0,197,0,0,0,16,0,196,0,221,0,56,0,240,0,229,0,56,0,187,0,0,0,110,0,82,0,212,0,138,0,163,0,0,0,0,0,8,0,22,0,0,0,165,0,29,0,67,0,238,0,198,0,237,0,116,0,23,0,209,0,42,0,34,0,49,0,64,0,0,0,125,0,237,0,50,0,164,0,0,0,209,0,41,0,0,0,172,0,150,0,136,0,62,0,0,0,140,0,118,0,0,0,137,0,3,0,20,0,68,0,170,0,247,0,130,0,16,0,57,0,174,0,178,0,200,0,78,0,0,0,254,0,0,0,211,0,148,0,17,0,245,0,103,0,0,0,175,0,132,0,0,0,206,0,0,0,11,0,47,0,154,0,165,0,218,0,113,0,191,0,22,0,222,0,160,0,12,0,0,0,203,0,14,0,0,0,0,0,136,0,242,0,151,0,60,0,90,0,92,0,82,0,139,0,0,0,73,0,135,0,35,0,77,0,177,0,117,0,200,0,227,0,163,0,143,0,0,0,3,0,29,0,0,0,19,0,0,0,37,0,1,0,59,0,0,0,0,0,41,0,0,0,226,0,0,0,137,0,22,0,237,0,0,0,50,0,165,0,28,0,0,0,161,0,9,0,91,0,0,0,0,0,228,0,0,0,173,0,0,0,21,0,219,0,0,0,146,0,0,0,77,0,93,0);
signal scenario_full  : scenario_type := (139,31,139,30,13,31,13,30,13,29,56,31,46,31,46,30,119,31,97,31,198,31,132,31,251,31,152,31,36,31,26,31,100,31,100,30,79,31,157,31,103,31,103,30,151,31,47,31,101,31,251,31,50,31,230,31,208,31,189,31,14,31,139,31,139,30,139,29,175,31,4,31,4,30,208,31,215,31,96,31,245,31,7,31,174,31,169,31,93,31,232,31,151,31,16,31,20,31,211,31,157,31,181,31,181,30,111,31,111,30,111,29,225,31,101,31,7,31,90,31,23,31,183,31,214,31,93,31,77,31,163,31,219,31,207,31,196,31,198,31,15,31,146,31,146,30,154,31,72,31,72,30,27,31,27,30,171,31,183,31,141,31,121,31,151,31,241,31,231,31,231,30,222,31,171,31,223,31,43,31,43,30,196,31,38,31,192,31,79,31,86,31,157,31,157,30,49,31,112,31,192,31,192,30,192,29,54,31,159,31,185,31,185,30,231,31,91,31,91,30,253,31,233,31,249,31,117,31,158,31,130,31,130,30,89,31,25,31,159,31,68,31,139,31,35,31,156,31,156,30,179,31,108,31,216,31,91,31,55,31,113,31,189,31,189,30,182,31,18,31,127,31,178,31,207,31,115,31,120,31,244,31,92,31,92,30,26,31,26,30,166,31,240,31,240,30,240,29,22,31,193,31,11,31,187,31,116,31,53,31,24,31,53,31,57,31,201,31,206,31,206,30,21,31,21,30,87,31,87,30,126,31,126,30,91,31,91,30,137,31,137,30,137,29,255,31,203,31,203,30,252,31,50,31,49,31,197,31,197,30,16,31,196,31,221,31,56,31,240,31,229,31,56,31,187,31,187,30,110,31,82,31,212,31,138,31,163,31,163,30,163,29,8,31,22,31,22,30,165,31,29,31,67,31,238,31,198,31,237,31,116,31,23,31,209,31,42,31,34,31,49,31,64,31,64,30,125,31,237,31,50,31,164,31,164,30,209,31,41,31,41,30,172,31,150,31,136,31,62,31,62,30,140,31,118,31,118,30,137,31,3,31,20,31,68,31,170,31,247,31,130,31,16,31,57,31,174,31,178,31,200,31,78,31,78,30,254,31,254,30,211,31,148,31,17,31,245,31,103,31,103,30,175,31,132,31,132,30,206,31,206,30,11,31,47,31,154,31,165,31,218,31,113,31,191,31,22,31,222,31,160,31,12,31,12,30,203,31,14,31,14,30,14,29,136,31,242,31,151,31,60,31,90,31,92,31,82,31,139,31,139,30,73,31,135,31,35,31,77,31,177,31,117,31,200,31,227,31,163,31,143,31,143,30,3,31,29,31,29,30,19,31,19,30,37,31,1,31,59,31,59,30,59,29,41,31,41,30,226,31,226,30,137,31,22,31,237,31,237,30,50,31,165,31,28,31,28,30,161,31,9,31,91,31,91,30,91,29,228,31,228,30,173,31,173,30,21,31,219,31,219,30,146,31,146,30,77,31,93,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
