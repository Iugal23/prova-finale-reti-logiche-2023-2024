-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_414 is
end project_tb_414;

architecture project_tb_arch_414 of project_tb_414 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 225;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,124,0,202,0,0,0,165,0,0,0,121,0,192,0,181,0,207,0,75,0,182,0,21,0,241,0,0,0,76,0,229,0,0,0,157,0,32,0,77,0,0,0,174,0,123,0,0,0,54,0,224,0,198,0,121,0,243,0,120,0,236,0,0,0,80,0,174,0,177,0,0,0,113,0,87,0,21,0,128,0,14,0,0,0,144,0,219,0,220,0,0,0,236,0,92,0,241,0,0,0,9,0,61,0,0,0,4,0,0,0,63,0,31,0,106,0,0,0,110,0,216,0,111,0,101,0,190,0,182,0,168,0,183,0,76,0,199,0,142,0,231,0,157,0,74,0,114,0,187,0,55,0,214,0,7,0,0,0,56,0,228,0,82,0,195,0,196,0,70,0,1,0,0,0,236,0,173,0,172,0,93,0,101,0,152,0,96,0,243,0,4,0,69,0,146,0,162,0,245,0,99,0,241,0,93,0,38,0,179,0,164,0,156,0,0,0,211,0,17,0,205,0,0,0,21,0,52,0,15,0,133,0,210,0,51,0,69,0,19,0,56,0,27,0,240,0,57,0,74,0,38,0,154,0,125,0,252,0,108,0,131,0,9,0,5,0,0,0,87,0,203,0,230,0,69,0,0,0,10,0,86,0,94,0,201,0,168,0,19,0,22,0,61,0,56,0,10,0,1,0,138,0,108,0,7,0,58,0,24,0,0,0,0,0,165,0,145,0,185,0,169,0,61,0,21,0,232,0,0,0,36,0,100,0,92,0,0,0,15,0,0,0,244,0,158,0,181,0,0,0,27,0,0,0,60,0,231,0,154,0,149,0,215,0,225,0,74,0,31,0,116,0,0,0,201,0,134,0,70,0,67,0,0,0,230,0,183,0,66,0,249,0,0,0,89,0,0,0,131,0,230,0,222,0,126,0,227,0,229,0,92,0,151,0,91,0,0,0,179,0,185,0,241,0,133,0,232,0,200,0,0,0,191,0,239,0,94,0,210,0,0,0,60,0,129,0,74,0);
signal scenario_full  : scenario_type := (0,0,124,31,202,31,202,30,165,31,165,30,121,31,192,31,181,31,207,31,75,31,182,31,21,31,241,31,241,30,76,31,229,31,229,30,157,31,32,31,77,31,77,30,174,31,123,31,123,30,54,31,224,31,198,31,121,31,243,31,120,31,236,31,236,30,80,31,174,31,177,31,177,30,113,31,87,31,21,31,128,31,14,31,14,30,144,31,219,31,220,31,220,30,236,31,92,31,241,31,241,30,9,31,61,31,61,30,4,31,4,30,63,31,31,31,106,31,106,30,110,31,216,31,111,31,101,31,190,31,182,31,168,31,183,31,76,31,199,31,142,31,231,31,157,31,74,31,114,31,187,31,55,31,214,31,7,31,7,30,56,31,228,31,82,31,195,31,196,31,70,31,1,31,1,30,236,31,173,31,172,31,93,31,101,31,152,31,96,31,243,31,4,31,69,31,146,31,162,31,245,31,99,31,241,31,93,31,38,31,179,31,164,31,156,31,156,30,211,31,17,31,205,31,205,30,21,31,52,31,15,31,133,31,210,31,51,31,69,31,19,31,56,31,27,31,240,31,57,31,74,31,38,31,154,31,125,31,252,31,108,31,131,31,9,31,5,31,5,30,87,31,203,31,230,31,69,31,69,30,10,31,86,31,94,31,201,31,168,31,19,31,22,31,61,31,56,31,10,31,1,31,138,31,108,31,7,31,58,31,24,31,24,30,24,29,165,31,145,31,185,31,169,31,61,31,21,31,232,31,232,30,36,31,100,31,92,31,92,30,15,31,15,30,244,31,158,31,181,31,181,30,27,31,27,30,60,31,231,31,154,31,149,31,215,31,225,31,74,31,31,31,116,31,116,30,201,31,134,31,70,31,67,31,67,30,230,31,183,31,66,31,249,31,249,30,89,31,89,30,131,31,230,31,222,31,126,31,227,31,229,31,92,31,151,31,91,31,91,30,179,31,185,31,241,31,133,31,232,31,200,31,200,30,191,31,239,31,94,31,210,31,210,30,60,31,129,31,74,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
