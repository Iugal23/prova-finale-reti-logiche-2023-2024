-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 520;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,193,0,136,0,48,0,253,0,200,0,217,0,2,0,94,0,0,0,26,0,77,0,178,0,38,0,93,0,232,0,137,0,51,0,226,0,0,0,106,0,114,0,190,0,165,0,91,0,0,0,189,0,165,0,52,0,253,0,169,0,243,0,0,0,99,0,164,0,89,0,220,0,98,0,26,0,0,0,187,0,0,0,0,0,95,0,21,0,80,0,0,0,134,0,236,0,0,0,238,0,231,0,126,0,48,0,12,0,87,0,0,0,180,0,121,0,148,0,229,0,247,0,0,0,35,0,12,0,37,0,45,0,157,0,0,0,1,0,117,0,147,0,12,0,252,0,138,0,0,0,63,0,218,0,119,0,123,0,40,0,25,0,136,0,90,0,49,0,182,0,61,0,190,0,128,0,183,0,179,0,101,0,88,0,235,0,216,0,87,0,0,0,116,0,0,0,16,0,236,0,96,0,69,0,0,0,136,0,177,0,110,0,67,0,93,0,181,0,0,0,172,0,199,0,0,0,134,0,0,0,251,0,20,0,111,0,33,0,123,0,0,0,107,0,225,0,152,0,2,0,43,0,7,0,205,0,0,0,107,0,179,0,81,0,54,0,134,0,217,0,84,0,224,0,167,0,56,0,35,0,0,0,145,0,0,0,7,0,70,0,0,0,0,0,26,0,0,0,219,0,205,0,141,0,65,0,59,0,65,0,34,0,71,0,108,0,222,0,63,0,196,0,237,0,34,0,0,0,170,0,16,0,0,0,238,0,161,0,144,0,225,0,168,0,50,0,237,0,123,0,208,0,136,0,0,0,144,0,93,0,131,0,230,0,0,0,44,0,25,0,121,0,102,0,201,0,0,0,0,0,0,0,246,0,88,0,144,0,53,0,230,0,0,0,101,0,0,0,186,0,112,0,248,0,137,0,74,0,201,0,3,0,0,0,111,0,73,0,49,0,57,0,202,0,139,0,39,0,135,0,0,0,39,0,174,0,84,0,250,0,45,0,253,0,86,0,157,0,88,0,254,0,0,0,203,0,229,0,110,0,72,0,208,0,0,0,93,0,141,0,0,0,0,0,160,0,130,0,0,0,0,0,125,0,0,0,103,0,121,0,82,0,219,0,16,0,233,0,184,0,0,0,0,0,236,0,204,0,140,0,169,0,0,0,15,0,0,0,0,0,41,0,42,0,77,0,185,0,246,0,15,0,121,0,174,0,209,0,32,0,188,0,253,0,229,0,147,0,238,0,194,0,98,0,176,0,0,0,219,0,12,0,57,0,0,0,37,0,19,0,133,0,172,0,52,0,0,0,37,0,68,0,249,0,209,0,30,0,214,0,0,0,87,0,87,0,0,0,60,0,119,0,189,0,189,0,43,0,29,0,0,0,159,0,12,0,10,0,8,0,185,0,85,0,157,0,231,0,134,0,123,0,202,0,0,0,72,0,97,0,13,0,159,0,7,0,222,0,0,0,0,0,249,0,35,0,109,0,0,0,109,0,9,0,48,0,0,0,0,0,104,0,76,0,168,0,205,0,84,0,0,0,0,0,211,0,0,0,73,0,138,0,16,0,13,0,182,0,0,0,5,0,32,0,70,0,223,0,219,0,191,0,197,0,0,0,183,0,153,0,100,0,234,0,169,0,85,0,236,0,194,0,239,0,60,0,32,0,114,0,91,0,229,0,0,0,108,0,0,0,188,0,177,0,251,0,72,0,222,0,137,0,31,0,0,0,0,0,39,0,0,0,89,0,126,0,204,0,247,0,181,0,139,0,132,0,153,0,155,0,82,0,220,0,141,0,172,0,157,0,55,0,193,0,35,0,222,0,202,0,0,0,250,0,216,0,0,0,7,0,118,0,190,0,32,0,207,0,0,0,0,0,155,0,0,0,189,0,18,0,0,0,0,0,28,0,53,0,0,0,181,0,123,0,0,0,254,0,53,0,0,0,253,0,24,0,0,0,213,0,221,0,42,0,72,0,192,0,0,0,242,0,130,0,43,0,165,0,116,0,54,0,20,0,158,0,148,0,43,0,0,0,0,0,39,0,15,0,197,0,201,0,18,0,143,0,233,0,107,0,9,0,133,0,221,0,4,0,0,0,171,0,51,0,0,0,0,0,192,0,111,0,36,0,214,0,39,0,0,0,46,0,231,0,55,0,59,0,151,0,32,0,25,0,171,0,172,0,118,0,4,0,121,0,26,0,50,0,143,0,132,0,60,0,0,0,16,0,200,0,79,0,0,0,216,0,0,0,156,0,184,0,73,0,219,0,39,0,0,0,48,0,119,0,0,0,177,0,239,0,135,0,0,0,0,0,0,0,220,0,99,0,0,0,0,0,72,0);
signal scenario_full  : scenario_type := (0,0,193,31,136,31,48,31,253,31,200,31,217,31,2,31,94,31,94,30,26,31,77,31,178,31,38,31,93,31,232,31,137,31,51,31,226,31,226,30,106,31,114,31,190,31,165,31,91,31,91,30,189,31,165,31,52,31,253,31,169,31,243,31,243,30,99,31,164,31,89,31,220,31,98,31,26,31,26,30,187,31,187,30,187,29,95,31,21,31,80,31,80,30,134,31,236,31,236,30,238,31,231,31,126,31,48,31,12,31,87,31,87,30,180,31,121,31,148,31,229,31,247,31,247,30,35,31,12,31,37,31,45,31,157,31,157,30,1,31,117,31,147,31,12,31,252,31,138,31,138,30,63,31,218,31,119,31,123,31,40,31,25,31,136,31,90,31,49,31,182,31,61,31,190,31,128,31,183,31,179,31,101,31,88,31,235,31,216,31,87,31,87,30,116,31,116,30,16,31,236,31,96,31,69,31,69,30,136,31,177,31,110,31,67,31,93,31,181,31,181,30,172,31,199,31,199,30,134,31,134,30,251,31,20,31,111,31,33,31,123,31,123,30,107,31,225,31,152,31,2,31,43,31,7,31,205,31,205,30,107,31,179,31,81,31,54,31,134,31,217,31,84,31,224,31,167,31,56,31,35,31,35,30,145,31,145,30,7,31,70,31,70,30,70,29,26,31,26,30,219,31,205,31,141,31,65,31,59,31,65,31,34,31,71,31,108,31,222,31,63,31,196,31,237,31,34,31,34,30,170,31,16,31,16,30,238,31,161,31,144,31,225,31,168,31,50,31,237,31,123,31,208,31,136,31,136,30,144,31,93,31,131,31,230,31,230,30,44,31,25,31,121,31,102,31,201,31,201,30,201,29,201,28,246,31,88,31,144,31,53,31,230,31,230,30,101,31,101,30,186,31,112,31,248,31,137,31,74,31,201,31,3,31,3,30,111,31,73,31,49,31,57,31,202,31,139,31,39,31,135,31,135,30,39,31,174,31,84,31,250,31,45,31,253,31,86,31,157,31,88,31,254,31,254,30,203,31,229,31,110,31,72,31,208,31,208,30,93,31,141,31,141,30,141,29,160,31,130,31,130,30,130,29,125,31,125,30,103,31,121,31,82,31,219,31,16,31,233,31,184,31,184,30,184,29,236,31,204,31,140,31,169,31,169,30,15,31,15,30,15,29,41,31,42,31,77,31,185,31,246,31,15,31,121,31,174,31,209,31,32,31,188,31,253,31,229,31,147,31,238,31,194,31,98,31,176,31,176,30,219,31,12,31,57,31,57,30,37,31,19,31,133,31,172,31,52,31,52,30,37,31,68,31,249,31,209,31,30,31,214,31,214,30,87,31,87,31,87,30,60,31,119,31,189,31,189,31,43,31,29,31,29,30,159,31,12,31,10,31,8,31,185,31,85,31,157,31,231,31,134,31,123,31,202,31,202,30,72,31,97,31,13,31,159,31,7,31,222,31,222,30,222,29,249,31,35,31,109,31,109,30,109,31,9,31,48,31,48,30,48,29,104,31,76,31,168,31,205,31,84,31,84,30,84,29,211,31,211,30,73,31,138,31,16,31,13,31,182,31,182,30,5,31,32,31,70,31,223,31,219,31,191,31,197,31,197,30,183,31,153,31,100,31,234,31,169,31,85,31,236,31,194,31,239,31,60,31,32,31,114,31,91,31,229,31,229,30,108,31,108,30,188,31,177,31,251,31,72,31,222,31,137,31,31,31,31,30,31,29,39,31,39,30,89,31,126,31,204,31,247,31,181,31,139,31,132,31,153,31,155,31,82,31,220,31,141,31,172,31,157,31,55,31,193,31,35,31,222,31,202,31,202,30,250,31,216,31,216,30,7,31,118,31,190,31,32,31,207,31,207,30,207,29,155,31,155,30,189,31,18,31,18,30,18,29,28,31,53,31,53,30,181,31,123,31,123,30,254,31,53,31,53,30,253,31,24,31,24,30,213,31,221,31,42,31,72,31,192,31,192,30,242,31,130,31,43,31,165,31,116,31,54,31,20,31,158,31,148,31,43,31,43,30,43,29,39,31,15,31,197,31,201,31,18,31,143,31,233,31,107,31,9,31,133,31,221,31,4,31,4,30,171,31,51,31,51,30,51,29,192,31,111,31,36,31,214,31,39,31,39,30,46,31,231,31,55,31,59,31,151,31,32,31,25,31,171,31,172,31,118,31,4,31,121,31,26,31,50,31,143,31,132,31,60,31,60,30,16,31,200,31,79,31,79,30,216,31,216,30,156,31,184,31,73,31,219,31,39,31,39,30,48,31,119,31,119,30,177,31,239,31,135,31,135,30,135,29,135,28,220,31,99,31,99,30,99,29,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
