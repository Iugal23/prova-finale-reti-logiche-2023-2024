-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 192;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (88,0,0,0,204,0,166,0,83,0,44,0,0,0,0,0,102,0,215,0,0,0,141,0,0,0,217,0,127,0,20,0,67,0,108,0,75,0,35,0,16,0,74,0,200,0,0,0,0,0,0,0,35,0,0,0,0,0,118,0,178,0,0,0,171,0,215,0,0,0,170,0,174,0,43,0,248,0,72,0,123,0,168,0,50,0,228,0,125,0,161,0,194,0,134,0,0,0,146,0,0,0,73,0,75,0,217,0,21,0,168,0,110,0,75,0,68,0,123,0,48,0,116,0,227,0,36,0,109,0,3,0,204,0,40,0,158,0,212,0,39,0,28,0,0,0,67,0,100,0,171,0,103,0,137,0,84,0,174,0,123,0,212,0,116,0,0,0,110,0,215,0,113,0,6,0,0,0,205,0,47,0,0,0,0,0,176,0,147,0,96,0,39,0,0,0,216,0,0,0,78,0,53,0,0,0,216,0,251,0,28,0,90,0,0,0,0,0,13,0,0,0,0,0,0,0,71,0,159,0,78,0,231,0,0,0,13,0,165,0,156,0,0,0,5,0,63,0,116,0,36,0,0,0,139,0,103,0,62,0,147,0,136,0,109,0,70,0,136,0,0,0,232,0,192,0,122,0,23,0,11,0,0,0,165,0,5,0,17,0,176,0,137,0,219,0,145,0,53,0,155,0,143,0,0,0,165,0,197,0,85,0,193,0,233,0,18,0,0,0,0,0,233,0,79,0,57,0,0,0,0,0,223,0,31,0,121,0,229,0,25,0,138,0,227,0,132,0,162,0,230,0,2,0,0,0,0,0,173,0,0,0,30,0,0,0,0,0,112,0,221,0,0,0,33,0,0,0,0,0,4,0,108,0);
signal scenario_full  : scenario_type := (88,31,88,30,204,31,166,31,83,31,44,31,44,30,44,29,102,31,215,31,215,30,141,31,141,30,217,31,127,31,20,31,67,31,108,31,75,31,35,31,16,31,74,31,200,31,200,30,200,29,200,28,35,31,35,30,35,29,118,31,178,31,178,30,171,31,215,31,215,30,170,31,174,31,43,31,248,31,72,31,123,31,168,31,50,31,228,31,125,31,161,31,194,31,134,31,134,30,146,31,146,30,73,31,75,31,217,31,21,31,168,31,110,31,75,31,68,31,123,31,48,31,116,31,227,31,36,31,109,31,3,31,204,31,40,31,158,31,212,31,39,31,28,31,28,30,67,31,100,31,171,31,103,31,137,31,84,31,174,31,123,31,212,31,116,31,116,30,110,31,215,31,113,31,6,31,6,30,205,31,47,31,47,30,47,29,176,31,147,31,96,31,39,31,39,30,216,31,216,30,78,31,53,31,53,30,216,31,251,31,28,31,90,31,90,30,90,29,13,31,13,30,13,29,13,28,71,31,159,31,78,31,231,31,231,30,13,31,165,31,156,31,156,30,5,31,63,31,116,31,36,31,36,30,139,31,103,31,62,31,147,31,136,31,109,31,70,31,136,31,136,30,232,31,192,31,122,31,23,31,11,31,11,30,165,31,5,31,17,31,176,31,137,31,219,31,145,31,53,31,155,31,143,31,143,30,165,31,197,31,85,31,193,31,233,31,18,31,18,30,18,29,233,31,79,31,57,31,57,30,57,29,223,31,31,31,121,31,229,31,25,31,138,31,227,31,132,31,162,31,230,31,2,31,2,30,2,29,173,31,173,30,30,31,30,30,30,29,112,31,221,31,221,30,33,31,33,30,33,29,4,31,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
