-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 491;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (78,0,232,0,90,0,254,0,1,0,39,0,244,0,249,0,0,0,204,0,216,0,64,0,4,0,0,0,0,0,67,0,155,0,186,0,140,0,200,0,240,0,0,0,166,0,13,0,134,0,68,0,56,0,28,0,26,0,35,0,116,0,0,0,33,0,43,0,212,0,32,0,183,0,108,0,0,0,104,0,241,0,82,0,33,0,157,0,166,0,33,0,230,0,26,0,0,0,166,0,85,0,237,0,207,0,252,0,193,0,45,0,75,0,86,0,141,0,109,0,244,0,119,0,126,0,123,0,112,0,110,0,235,0,139,0,154,0,0,0,78,0,94,0,0,0,169,0,80,0,0,0,106,0,179,0,91,0,0,0,76,0,29,0,0,0,241,0,26,0,0,0,138,0,255,0,187,0,24,0,0,0,0,0,150,0,41,0,169,0,157,0,116,0,138,0,120,0,97,0,225,0,87,0,46,0,0,0,40,0,123,0,0,0,33,0,0,0,94,0,0,0,120,0,156,0,182,0,207,0,226,0,0,0,91,0,65,0,29,0,217,0,0,0,234,0,13,0,230,0,168,0,191,0,28,0,0,0,169,0,135,0,77,0,176,0,231,0,132,0,0,0,92,0,241,0,57,0,201,0,162,0,0,0,139,0,215,0,98,0,157,0,0,0,76,0,151,0,119,0,64,0,143,0,0,0,0,0,8,0,48,0,37,0,89,0,0,0,97,0,17,0,87,0,69,0,90,0,92,0,196,0,0,0,11,0,233,0,29,0,0,0,195,0,192,0,0,0,223,0,0,0,99,0,71,0,47,0,126,0,91,0,138,0,0,0,70,0,176,0,60,0,68,0,12,0,0,0,48,0,0,0,79,0,6,0,69,0,186,0,172,0,169,0,0,0,89,0,63,0,80,0,92,0,192,0,79,0,135,0,150,0,23,0,97,0,0,0,20,0,6,0,162,0,242,0,0,0,0,0,20,0,18,0,30,0,33,0,103,0,0,0,69,0,78,0,0,0,0,0,238,0,138,0,35,0,117,0,0,0,0,0,0,0,0,0,103,0,0,0,74,0,65,0,0,0,83,0,0,0,0,0,153,0,219,0,21,0,0,0,247,0,0,0,164,0,43,0,10,0,147,0,30,0,179,0,47,0,67,0,31,0,0,0,0,0,153,0,119,0,200,0,0,0,94,0,7,0,0,0,0,0,113,0,154,0,0,0,206,0,89,0,204,0,239,0,234,0,110,0,218,0,0,0,111,0,0,0,218,0,0,0,205,0,251,0,0,0,120,0,37,0,0,0,175,0,0,0,179,0,225,0,0,0,203,0,145,0,95,0,50,0,76,0,232,0,114,0,0,0,3,0,130,0,4,0,8,0,181,0,233,0,0,0,45,0,57,0,113,0,3,0,0,0,232,0,216,0,112,0,73,0,0,0,155,0,143,0,134,0,117,0,253,0,0,0,197,0,118,0,131,0,0,0,110,0,131,0,175,0,234,0,66,0,0,0,244,0,0,0,195,0,40,0,67,0,12,0,80,0,17,0,0,0,0,0,85,0,155,0,101,0,180,0,194,0,0,0,131,0,231,0,106,0,93,0,0,0,145,0,236,0,189,0,0,0,183,0,0,0,49,0,184,0,62,0,176,0,178,0,103,0,206,0,220,0,112,0,193,0,107,0,233,0,231,0,178,0,139,0,47,0,210,0,82,0,243,0,170,0,199,0,0,0,241,0,0,0,201,0,122,0,19,0,16,0,219,0,184,0,133,0,196,0,50,0,0,0,146,0,255,0,116,0,82,0,194,0,117,0,14,0,0,0,214,0,55,0,0,0,65,0,243,0,177,0,84,0,0,0,208,0,228,0,0,0,0,0,144,0,231,0,0,0,88,0,25,0,93,0,31,0,222,0,0,0,0,0,40,0,98,0,181,0,120,0,164,0,90,0,0,0,0,0,233,0,83,0,18,0,123,0,236,0,13,0,0,0,43,0,44,0,179,0,24,0,93,0,42,0,237,0,30,0,121,0,249,0,15,0,253,0,235,0,0,0,169,0,175,0,108,0,67,0,247,0,0,0,0,0,232,0,22,0,142,0,137,0,142,0,0,0,155,0,198,0,53,0,165,0,204,0,0,0,0,0,0,0,0,0,181,0,0,0,34,0,103,0,32,0,228,0,121,0,35,0,0,0,211,0,10,0,153,0,0,0,50,0,139,0,21,0);
signal scenario_full  : scenario_type := (78,31,232,31,90,31,254,31,1,31,39,31,244,31,249,31,249,30,204,31,216,31,64,31,4,31,4,30,4,29,67,31,155,31,186,31,140,31,200,31,240,31,240,30,166,31,13,31,134,31,68,31,56,31,28,31,26,31,35,31,116,31,116,30,33,31,43,31,212,31,32,31,183,31,108,31,108,30,104,31,241,31,82,31,33,31,157,31,166,31,33,31,230,31,26,31,26,30,166,31,85,31,237,31,207,31,252,31,193,31,45,31,75,31,86,31,141,31,109,31,244,31,119,31,126,31,123,31,112,31,110,31,235,31,139,31,154,31,154,30,78,31,94,31,94,30,169,31,80,31,80,30,106,31,179,31,91,31,91,30,76,31,29,31,29,30,241,31,26,31,26,30,138,31,255,31,187,31,24,31,24,30,24,29,150,31,41,31,169,31,157,31,116,31,138,31,120,31,97,31,225,31,87,31,46,31,46,30,40,31,123,31,123,30,33,31,33,30,94,31,94,30,120,31,156,31,182,31,207,31,226,31,226,30,91,31,65,31,29,31,217,31,217,30,234,31,13,31,230,31,168,31,191,31,28,31,28,30,169,31,135,31,77,31,176,31,231,31,132,31,132,30,92,31,241,31,57,31,201,31,162,31,162,30,139,31,215,31,98,31,157,31,157,30,76,31,151,31,119,31,64,31,143,31,143,30,143,29,8,31,48,31,37,31,89,31,89,30,97,31,17,31,87,31,69,31,90,31,92,31,196,31,196,30,11,31,233,31,29,31,29,30,195,31,192,31,192,30,223,31,223,30,99,31,71,31,47,31,126,31,91,31,138,31,138,30,70,31,176,31,60,31,68,31,12,31,12,30,48,31,48,30,79,31,6,31,69,31,186,31,172,31,169,31,169,30,89,31,63,31,80,31,92,31,192,31,79,31,135,31,150,31,23,31,97,31,97,30,20,31,6,31,162,31,242,31,242,30,242,29,20,31,18,31,30,31,33,31,103,31,103,30,69,31,78,31,78,30,78,29,238,31,138,31,35,31,117,31,117,30,117,29,117,28,117,27,103,31,103,30,74,31,65,31,65,30,83,31,83,30,83,29,153,31,219,31,21,31,21,30,247,31,247,30,164,31,43,31,10,31,147,31,30,31,179,31,47,31,67,31,31,31,31,30,31,29,153,31,119,31,200,31,200,30,94,31,7,31,7,30,7,29,113,31,154,31,154,30,206,31,89,31,204,31,239,31,234,31,110,31,218,31,218,30,111,31,111,30,218,31,218,30,205,31,251,31,251,30,120,31,37,31,37,30,175,31,175,30,179,31,225,31,225,30,203,31,145,31,95,31,50,31,76,31,232,31,114,31,114,30,3,31,130,31,4,31,8,31,181,31,233,31,233,30,45,31,57,31,113,31,3,31,3,30,232,31,216,31,112,31,73,31,73,30,155,31,143,31,134,31,117,31,253,31,253,30,197,31,118,31,131,31,131,30,110,31,131,31,175,31,234,31,66,31,66,30,244,31,244,30,195,31,40,31,67,31,12,31,80,31,17,31,17,30,17,29,85,31,155,31,101,31,180,31,194,31,194,30,131,31,231,31,106,31,93,31,93,30,145,31,236,31,189,31,189,30,183,31,183,30,49,31,184,31,62,31,176,31,178,31,103,31,206,31,220,31,112,31,193,31,107,31,233,31,231,31,178,31,139,31,47,31,210,31,82,31,243,31,170,31,199,31,199,30,241,31,241,30,201,31,122,31,19,31,16,31,219,31,184,31,133,31,196,31,50,31,50,30,146,31,255,31,116,31,82,31,194,31,117,31,14,31,14,30,214,31,55,31,55,30,65,31,243,31,177,31,84,31,84,30,208,31,228,31,228,30,228,29,144,31,231,31,231,30,88,31,25,31,93,31,31,31,222,31,222,30,222,29,40,31,98,31,181,31,120,31,164,31,90,31,90,30,90,29,233,31,83,31,18,31,123,31,236,31,13,31,13,30,43,31,44,31,179,31,24,31,93,31,42,31,237,31,30,31,121,31,249,31,15,31,253,31,235,31,235,30,169,31,175,31,108,31,67,31,247,31,247,30,247,29,232,31,22,31,142,31,137,31,142,31,142,30,155,31,198,31,53,31,165,31,204,31,204,30,204,29,204,28,204,27,181,31,181,30,34,31,103,31,32,31,228,31,121,31,35,31,35,30,211,31,10,31,153,31,153,30,50,31,139,31,21,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
