-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_290 is
end project_tb_290;

architecture project_tb_arch_290 of project_tb_290 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 862;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (176,0,145,0,162,0,39,0,116,0,0,0,0,0,167,0,146,0,242,0,66,0,136,0,241,0,0,0,0,0,66,0,17,0,18,0,159,0,226,0,254,0,0,0,238,0,7,0,104,0,122,0,64,0,91,0,68,0,0,0,241,0,100,0,190,0,79,0,0,0,0,0,249,0,99,0,0,0,54,0,135,0,254,0,149,0,0,0,45,0,89,0,240,0,12,0,196,0,115,0,231,0,43,0,122,0,49,0,155,0,0,0,0,0,221,0,21,0,0,0,93,0,225,0,111,0,0,0,0,0,36,0,209,0,0,0,111,0,75,0,61,0,225,0,51,0,0,0,74,0,236,0,0,0,21,0,33,0,91,0,233,0,34,0,64,0,0,0,0,0,0,0,109,0,0,0,238,0,0,0,254,0,221,0,109,0,51,0,50,0,151,0,0,0,0,0,183,0,70,0,80,0,123,0,149,0,53,0,53,0,243,0,87,0,90,0,119,0,235,0,122,0,154,0,0,0,45,0,72,0,0,0,195,0,89,0,226,0,125,0,217,0,199,0,0,0,204,0,246,0,38,0,11,0,177,0,5,0,171,0,0,0,95,0,234,0,86,0,92,0,49,0,80,0,0,0,241,0,76,0,13,0,255,0,46,0,0,0,80,0,144,0,189,0,74,0,225,0,0,0,16,0,222,0,0,0,98,0,0,0,112,0,0,0,243,0,11,0,151,0,0,0,126,0,56,0,172,0,0,0,0,0,54,0,0,0,172,0,82,0,209,0,43,0,0,0,32,0,84,0,0,0,72,0,48,0,162,0,130,0,237,0,230,0,83,0,147,0,79,0,24,0,87,0,45,0,183,0,244,0,143,0,128,0,145,0,174,0,8,0,22,0,168,0,94,0,0,0,69,0,139,0,14,0,0,0,76,0,52,0,132,0,3,0,225,0,232,0,157,0,232,0,182,0,146,0,0,0,0,0,11,0,127,0,49,0,0,0,0,0,252,0,206,0,125,0,62,0,25,0,0,0,255,0,32,0,25,0,130,0,0,0,0,0,0,0,7,0,99,0,0,0,14,0,149,0,237,0,87,0,0,0,142,0,0,0,136,0,164,0,14,0,0,0,19,0,0,0,158,0,0,0,206,0,7,0,87,0,0,0,249,0,123,0,97,0,204,0,86,0,208,0,59,0,143,0,251,0,58,0,96,0,114,0,195,0,0,0,209,0,93,0,208,0,255,0,169,0,183,0,52,0,192,0,107,0,84,0,209,0,191,0,47,0,113,0,216,0,0,0,30,0,83,0,37,0,83,0,100,0,164,0,0,0,0,0,0,0,112,0,13,0,16,0,191,0,0,0,213,0,0,0,50,0,71,0,245,0,0,0,1,0,7,0,139,0,171,0,0,0,102,0,48,0,141,0,223,0,201,0,129,0,102,0,130,0,94,0,0,0,0,0,88,0,0,0,194,0,185,0,145,0,130,0,72,0,48,0,83,0,169,0,30,0,0,0,0,0,174,0,0,0,193,0,0,0,238,0,251,0,141,0,142,0,99,0,204,0,176,0,8,0,11,0,84,0,63,0,91,0,170,0,0,0,0,0,135,0,70,0,194,0,0,0,0,0,242,0,120,0,61,0,9,0,187,0,114,0,0,0,170,0,137,0,113,0,82,0,62,0,0,0,232,0,0,0,173,0,112,0,141,0,193,0,0,0,143,0,112,0,77,0,23,0,200,0,16,0,0,0,246,0,115,0,144,0,230,0,0,0,188,0,180,0,0,0,190,0,91,0,196,0,59,0,97,0,0,0,74,0,161,0,95,0,55,0,0,0,89,0,0,0,124,0,240,0,221,0,20,0,138,0,121,0,93,0,30,0,125,0,0,0,133,0,110,0,231,0,0,0,68,0,35,0,165,0,0,0,225,0,65,0,0,0,229,0,165,0,96,0,85,0,137,0,183,0,216,0,0,0,171,0,99,0,194,0,225,0,11,0,0,0,0,0,21,0,69,0,22,0,77,0,251,0,21,0,61,0,125,0,127,0,161,0,122,0,159,0,56,0,139,0,0,0,185,0,216,0,20,0,241,0,128,0,184,0,195,0,228,0,0,0,115,0,219,0,193,0,0,0,36,0,72,0,205,0,41,0,174,0,97,0,73,0,215,0,204,0,13,0,0,0,31,0,19,0,6,0,61,0,129,0,252,0,220,0,0,0,34,0,33,0,0,0,0,0,79,0,113,0,32,0,233,0,14,0,164,0,0,0,168,0,2,0,219,0,0,0,24,0,0,0,254,0,195,0,33,0,112,0,150,0,33,0,77,0,189,0,251,0,0,0,189,0,0,0,212,0,47,0,172,0,223,0,145,0,230,0,0,0,117,0,0,0,18,0,3,0,25,0,83,0,51,0,108,0,166,0,0,0,31,0,0,0,0,0,141,0,156,0,235,0,67,0,4,0,185,0,60,0,134,0,169,0,126,0,0,0,55,0,224,0,178,0,169,0,0,0,0,0,128,0,170,0,254,0,41,0,0,0,0,0,0,0,211,0,44,0,179,0,185,0,172,0,7,0,199,0,241,0,190,0,0,0,10,0,9,0,211,0,0,0,63,0,239,0,243,0,163,0,62,0,0,0,176,0,88,0,18,0,0,0,0,0,233,0,24,0,43,0,253,0,153,0,15,0,70,0,84,0,0,0,0,0,166,0,164,0,175,0,0,0,0,0,94,0,25,0,0,0,229,0,134,0,212,0,13,0,0,0,177,0,31,0,181,0,3,0,144,0,97,0,85,0,0,0,191,0,0,0,207,0,147,0,68,0,0,0,231,0,0,0,0,0,131,0,0,0,161,0,48,0,143,0,0,0,251,0,162,0,0,0,0,0,7,0,135,0,191,0,217,0,246,0,252,0,0,0,148,0,2,0,197,0,80,0,0,0,0,0,30,0,0,0,236,0,172,0,46,0,0,0,0,0,173,0,0,0,152,0,55,0,45,0,101,0,0,0,0,0,40,0,244,0,122,0,0,0,69,0,173,0,229,0,217,0,215,0,157,0,251,0,40,0,0,0,0,0,0,0,0,0,164,0,31,0,136,0,31,0,15,0,114,0,153,0,0,0,201,0,14,0,172,0,41,0,65,0,157,0,0,0,225,0,89,0,223,0,0,0,0,0,0,0,0,0,0,0,118,0,59,0,165,0,0,0,36,0,22,0,233,0,94,0,238,0,0,0,0,0,176,0,34,0,63,0,53,0,190,0,233,0,210,0,52,0,111,0,97,0,119,0,157,0,134,0,208,0,0,0,101,0,0,0,128,0,0,0,66,0,0,0,91,0,85,0,102,0,43,0,95,0,32,0,99,0,208,0,247,0,245,0,140,0,95,0,139,0,172,0,0,0,169,0,54,0,0,0,180,0,0,0,0,0,41,0,96,0,198,0,54,0,64,0,190,0,29,0,0,0,188,0,0,0,88,0,180,0,203,0,154,0,60,0,215,0,0,0,26,0,154,0,85,0,69,0,66,0,249,0,58,0,222,0,40,0,111,0,144,0,56,0,94,0,164,0,0,0,0,0,0,0,0,0,200,0,248,0,40,0,254,0,133,0,187,0,81,0,186,0,52,0,142,0,109,0,107,0,0,0,219,0,114,0,86,0,166,0,0,0,2,0,208,0,231,0,144,0,135,0,205,0,0,0,184,0,179,0,191,0,245,0,49,0,0,0,222,0,162,0,195,0,114,0,149,0,0,0,46,0,153,0,137,0,254,0,15,0,181,0,230,0,254,0,26,0,36,0,82,0,7,0,151,0,0,0,192,0,9,0,215,0,0,0,81,0,188,0,27,0,150,0,68,0,246,0,24,0,73,0,52,0,3,0,209,0,242,0,72,0,0,0,122,0);
signal scenario_full  : scenario_type := (176,31,145,31,162,31,39,31,116,31,116,30,116,29,167,31,146,31,242,31,66,31,136,31,241,31,241,30,241,29,66,31,17,31,18,31,159,31,226,31,254,31,254,30,238,31,7,31,104,31,122,31,64,31,91,31,68,31,68,30,241,31,100,31,190,31,79,31,79,30,79,29,249,31,99,31,99,30,54,31,135,31,254,31,149,31,149,30,45,31,89,31,240,31,12,31,196,31,115,31,231,31,43,31,122,31,49,31,155,31,155,30,155,29,221,31,21,31,21,30,93,31,225,31,111,31,111,30,111,29,36,31,209,31,209,30,111,31,75,31,61,31,225,31,51,31,51,30,74,31,236,31,236,30,21,31,33,31,91,31,233,31,34,31,64,31,64,30,64,29,64,28,109,31,109,30,238,31,238,30,254,31,221,31,109,31,51,31,50,31,151,31,151,30,151,29,183,31,70,31,80,31,123,31,149,31,53,31,53,31,243,31,87,31,90,31,119,31,235,31,122,31,154,31,154,30,45,31,72,31,72,30,195,31,89,31,226,31,125,31,217,31,199,31,199,30,204,31,246,31,38,31,11,31,177,31,5,31,171,31,171,30,95,31,234,31,86,31,92,31,49,31,80,31,80,30,241,31,76,31,13,31,255,31,46,31,46,30,80,31,144,31,189,31,74,31,225,31,225,30,16,31,222,31,222,30,98,31,98,30,112,31,112,30,243,31,11,31,151,31,151,30,126,31,56,31,172,31,172,30,172,29,54,31,54,30,172,31,82,31,209,31,43,31,43,30,32,31,84,31,84,30,72,31,48,31,162,31,130,31,237,31,230,31,83,31,147,31,79,31,24,31,87,31,45,31,183,31,244,31,143,31,128,31,145,31,174,31,8,31,22,31,168,31,94,31,94,30,69,31,139,31,14,31,14,30,76,31,52,31,132,31,3,31,225,31,232,31,157,31,232,31,182,31,146,31,146,30,146,29,11,31,127,31,49,31,49,30,49,29,252,31,206,31,125,31,62,31,25,31,25,30,255,31,32,31,25,31,130,31,130,30,130,29,130,28,7,31,99,31,99,30,14,31,149,31,237,31,87,31,87,30,142,31,142,30,136,31,164,31,14,31,14,30,19,31,19,30,158,31,158,30,206,31,7,31,87,31,87,30,249,31,123,31,97,31,204,31,86,31,208,31,59,31,143,31,251,31,58,31,96,31,114,31,195,31,195,30,209,31,93,31,208,31,255,31,169,31,183,31,52,31,192,31,107,31,84,31,209,31,191,31,47,31,113,31,216,31,216,30,30,31,83,31,37,31,83,31,100,31,164,31,164,30,164,29,164,28,112,31,13,31,16,31,191,31,191,30,213,31,213,30,50,31,71,31,245,31,245,30,1,31,7,31,139,31,171,31,171,30,102,31,48,31,141,31,223,31,201,31,129,31,102,31,130,31,94,31,94,30,94,29,88,31,88,30,194,31,185,31,145,31,130,31,72,31,48,31,83,31,169,31,30,31,30,30,30,29,174,31,174,30,193,31,193,30,238,31,251,31,141,31,142,31,99,31,204,31,176,31,8,31,11,31,84,31,63,31,91,31,170,31,170,30,170,29,135,31,70,31,194,31,194,30,194,29,242,31,120,31,61,31,9,31,187,31,114,31,114,30,170,31,137,31,113,31,82,31,62,31,62,30,232,31,232,30,173,31,112,31,141,31,193,31,193,30,143,31,112,31,77,31,23,31,200,31,16,31,16,30,246,31,115,31,144,31,230,31,230,30,188,31,180,31,180,30,190,31,91,31,196,31,59,31,97,31,97,30,74,31,161,31,95,31,55,31,55,30,89,31,89,30,124,31,240,31,221,31,20,31,138,31,121,31,93,31,30,31,125,31,125,30,133,31,110,31,231,31,231,30,68,31,35,31,165,31,165,30,225,31,65,31,65,30,229,31,165,31,96,31,85,31,137,31,183,31,216,31,216,30,171,31,99,31,194,31,225,31,11,31,11,30,11,29,21,31,69,31,22,31,77,31,251,31,21,31,61,31,125,31,127,31,161,31,122,31,159,31,56,31,139,31,139,30,185,31,216,31,20,31,241,31,128,31,184,31,195,31,228,31,228,30,115,31,219,31,193,31,193,30,36,31,72,31,205,31,41,31,174,31,97,31,73,31,215,31,204,31,13,31,13,30,31,31,19,31,6,31,61,31,129,31,252,31,220,31,220,30,34,31,33,31,33,30,33,29,79,31,113,31,32,31,233,31,14,31,164,31,164,30,168,31,2,31,219,31,219,30,24,31,24,30,254,31,195,31,33,31,112,31,150,31,33,31,77,31,189,31,251,31,251,30,189,31,189,30,212,31,47,31,172,31,223,31,145,31,230,31,230,30,117,31,117,30,18,31,3,31,25,31,83,31,51,31,108,31,166,31,166,30,31,31,31,30,31,29,141,31,156,31,235,31,67,31,4,31,185,31,60,31,134,31,169,31,126,31,126,30,55,31,224,31,178,31,169,31,169,30,169,29,128,31,170,31,254,31,41,31,41,30,41,29,41,28,211,31,44,31,179,31,185,31,172,31,7,31,199,31,241,31,190,31,190,30,10,31,9,31,211,31,211,30,63,31,239,31,243,31,163,31,62,31,62,30,176,31,88,31,18,31,18,30,18,29,233,31,24,31,43,31,253,31,153,31,15,31,70,31,84,31,84,30,84,29,166,31,164,31,175,31,175,30,175,29,94,31,25,31,25,30,229,31,134,31,212,31,13,31,13,30,177,31,31,31,181,31,3,31,144,31,97,31,85,31,85,30,191,31,191,30,207,31,147,31,68,31,68,30,231,31,231,30,231,29,131,31,131,30,161,31,48,31,143,31,143,30,251,31,162,31,162,30,162,29,7,31,135,31,191,31,217,31,246,31,252,31,252,30,148,31,2,31,197,31,80,31,80,30,80,29,30,31,30,30,236,31,172,31,46,31,46,30,46,29,173,31,173,30,152,31,55,31,45,31,101,31,101,30,101,29,40,31,244,31,122,31,122,30,69,31,173,31,229,31,217,31,215,31,157,31,251,31,40,31,40,30,40,29,40,28,40,27,164,31,31,31,136,31,31,31,15,31,114,31,153,31,153,30,201,31,14,31,172,31,41,31,65,31,157,31,157,30,225,31,89,31,223,31,223,30,223,29,223,28,223,27,223,26,118,31,59,31,165,31,165,30,36,31,22,31,233,31,94,31,238,31,238,30,238,29,176,31,34,31,63,31,53,31,190,31,233,31,210,31,52,31,111,31,97,31,119,31,157,31,134,31,208,31,208,30,101,31,101,30,128,31,128,30,66,31,66,30,91,31,85,31,102,31,43,31,95,31,32,31,99,31,208,31,247,31,245,31,140,31,95,31,139,31,172,31,172,30,169,31,54,31,54,30,180,31,180,30,180,29,41,31,96,31,198,31,54,31,64,31,190,31,29,31,29,30,188,31,188,30,88,31,180,31,203,31,154,31,60,31,215,31,215,30,26,31,154,31,85,31,69,31,66,31,249,31,58,31,222,31,40,31,111,31,144,31,56,31,94,31,164,31,164,30,164,29,164,28,164,27,200,31,248,31,40,31,254,31,133,31,187,31,81,31,186,31,52,31,142,31,109,31,107,31,107,30,219,31,114,31,86,31,166,31,166,30,2,31,208,31,231,31,144,31,135,31,205,31,205,30,184,31,179,31,191,31,245,31,49,31,49,30,222,31,162,31,195,31,114,31,149,31,149,30,46,31,153,31,137,31,254,31,15,31,181,31,230,31,254,31,26,31,36,31,82,31,7,31,151,31,151,30,192,31,9,31,215,31,215,30,81,31,188,31,27,31,150,31,68,31,246,31,24,31,73,31,52,31,3,31,209,31,242,31,72,31,72,30,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
