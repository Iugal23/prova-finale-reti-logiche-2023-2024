-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 369;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (11,0,104,0,108,0,0,0,152,0,146,0,242,0,179,0,157,0,156,0,58,0,219,0,0,0,2,0,254,0,19,0,0,0,216,0,142,0,45,0,0,0,0,0,120,0,162,0,118,0,16,0,33,0,77,0,0,0,178,0,215,0,110,0,168,0,0,0,166,0,87,0,93,0,178,0,149,0,0,0,18,0,32,0,0,0,30,0,235,0,37,0,44,0,252,0,16,0,251,0,0,0,125,0,73,0,7,0,63,0,219,0,0,0,142,0,204,0,209,0,7,0,0,0,15,0,0,0,0,0,11,0,28,0,224,0,158,0,0,0,75,0,0,0,152,0,177,0,101,0,231,0,121,0,190,0,214,0,13,0,127,0,216,0,245,0,210,0,78,0,237,0,109,0,0,0,106,0,229,0,128,0,106,0,36,0,0,0,0,0,0,0,0,0,245,0,1,0,36,0,182,0,173,0,241,0,249,0,77,0,59,0,23,0,238,0,0,0,0,0,17,0,80,0,242,0,0,0,151,0,121,0,164,0,47,0,165,0,185,0,27,0,32,0,247,0,26,0,188,0,76,0,214,0,179,0,12,0,0,0,137,0,205,0,231,0,31,0,237,0,69,0,63,0,0,0,40,0,0,0,0,0,20,0,52,0,65,0,0,0,8,0,17,0,0,0,212,0,100,0,0,0,0,0,66,0,147,0,54,0,59,0,0,0,81,0,157,0,55,0,33,0,0,0,18,0,47,0,92,0,142,0,78,0,23,0,186,0,182,0,169,0,28,0,141,0,210,0,158,0,71,0,69,0,0,0,188,0,252,0,0,0,53,0,0,0,46,0,73,0,149,0,44,0,0,0,155,0,0,0,168,0,200,0,237,0,132,0,201,0,222,0,0,0,85,0,209,0,0,0,153,0,56,0,42,0,0,0,97,0,83,0,0,0,12,0,221,0,164,0,139,0,0,0,0,0,82,0,115,0,124,0,72,0,252,0,147,0,119,0,196,0,104,0,105,0,207,0,0,0,73,0,68,0,152,0,0,0,79,0,132,0,62,0,218,0,81,0,47,0,0,0,144,0,207,0,239,0,253,0,176,0,179,0,116,0,0,0,0,0,249,0,17,0,225,0,197,0,23,0,147,0,118,0,162,0,96,0,144,0,0,0,52,0,253,0,2,0,0,0,4,0,75,0,21,0,0,0,132,0,194,0,100,0,139,0,141,0,138,0,6,0,189,0,60,0,0,0,71,0,0,0,0,0,2,0,0,0,118,0,140,0,166,0,81,0,222,0,58,0,186,0,194,0,223,0,159,0,31,0,0,0,125,0,47,0,0,0,2,0,0,0,200,0,102,0,148,0,91,0,0,0,101,0,114,0,92,0,33,0,0,0,242,0,141,0,178,0,106,0,125,0,87,0,95,0,5,0,0,0,45,0,0,0,26,0,163,0,120,0,101,0,185,0,0,0,124,0,115,0,188,0,0,0,255,0,178,0,46,0,71,0,83,0,9,0,0,0,227,0,118,0,0,0,61,0,184,0,52,0,65,0,131,0,247,0,120,0,171,0,75,0,88,0,188,0,72,0,139,0,140,0,231,0,227,0,0,0,192,0,244,0,195,0,61,0,0,0,162,0,77,0,49,0,216,0,89,0,51,0,0,0,0,0,143,0,246,0);
signal scenario_full  : scenario_type := (11,31,104,31,108,31,108,30,152,31,146,31,242,31,179,31,157,31,156,31,58,31,219,31,219,30,2,31,254,31,19,31,19,30,216,31,142,31,45,31,45,30,45,29,120,31,162,31,118,31,16,31,33,31,77,31,77,30,178,31,215,31,110,31,168,31,168,30,166,31,87,31,93,31,178,31,149,31,149,30,18,31,32,31,32,30,30,31,235,31,37,31,44,31,252,31,16,31,251,31,251,30,125,31,73,31,7,31,63,31,219,31,219,30,142,31,204,31,209,31,7,31,7,30,15,31,15,30,15,29,11,31,28,31,224,31,158,31,158,30,75,31,75,30,152,31,177,31,101,31,231,31,121,31,190,31,214,31,13,31,127,31,216,31,245,31,210,31,78,31,237,31,109,31,109,30,106,31,229,31,128,31,106,31,36,31,36,30,36,29,36,28,36,27,245,31,1,31,36,31,182,31,173,31,241,31,249,31,77,31,59,31,23,31,238,31,238,30,238,29,17,31,80,31,242,31,242,30,151,31,121,31,164,31,47,31,165,31,185,31,27,31,32,31,247,31,26,31,188,31,76,31,214,31,179,31,12,31,12,30,137,31,205,31,231,31,31,31,237,31,69,31,63,31,63,30,40,31,40,30,40,29,20,31,52,31,65,31,65,30,8,31,17,31,17,30,212,31,100,31,100,30,100,29,66,31,147,31,54,31,59,31,59,30,81,31,157,31,55,31,33,31,33,30,18,31,47,31,92,31,142,31,78,31,23,31,186,31,182,31,169,31,28,31,141,31,210,31,158,31,71,31,69,31,69,30,188,31,252,31,252,30,53,31,53,30,46,31,73,31,149,31,44,31,44,30,155,31,155,30,168,31,200,31,237,31,132,31,201,31,222,31,222,30,85,31,209,31,209,30,153,31,56,31,42,31,42,30,97,31,83,31,83,30,12,31,221,31,164,31,139,31,139,30,139,29,82,31,115,31,124,31,72,31,252,31,147,31,119,31,196,31,104,31,105,31,207,31,207,30,73,31,68,31,152,31,152,30,79,31,132,31,62,31,218,31,81,31,47,31,47,30,144,31,207,31,239,31,253,31,176,31,179,31,116,31,116,30,116,29,249,31,17,31,225,31,197,31,23,31,147,31,118,31,162,31,96,31,144,31,144,30,52,31,253,31,2,31,2,30,4,31,75,31,21,31,21,30,132,31,194,31,100,31,139,31,141,31,138,31,6,31,189,31,60,31,60,30,71,31,71,30,71,29,2,31,2,30,118,31,140,31,166,31,81,31,222,31,58,31,186,31,194,31,223,31,159,31,31,31,31,30,125,31,47,31,47,30,2,31,2,30,200,31,102,31,148,31,91,31,91,30,101,31,114,31,92,31,33,31,33,30,242,31,141,31,178,31,106,31,125,31,87,31,95,31,5,31,5,30,45,31,45,30,26,31,163,31,120,31,101,31,185,31,185,30,124,31,115,31,188,31,188,30,255,31,178,31,46,31,71,31,83,31,9,31,9,30,227,31,118,31,118,30,61,31,184,31,52,31,65,31,131,31,247,31,120,31,171,31,75,31,88,31,188,31,72,31,139,31,140,31,231,31,227,31,227,30,192,31,244,31,195,31,61,31,61,30,162,31,77,31,49,31,216,31,89,31,51,31,51,30,51,29,143,31,246,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
