-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 336;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,0,0,75,0,251,0,81,0,231,0,90,0,66,0,168,0,0,0,113,0,180,0,17,0,126,0,0,0,255,0,198,0,221,0,249,0,167,0,21,0,0,0,0,0,0,0,0,0,0,0,2,0,45,0,235,0,89,0,101,0,10,0,24,0,84,0,162,0,223,0,28,0,212,0,183,0,0,0,0,0,77,0,244,0,0,0,245,0,54,0,7,0,20,0,177,0,159,0,0,0,0,0,0,0,82,0,232,0,5,0,120,0,94,0,0,0,243,0,66,0,137,0,129,0,165,0,62,0,74,0,0,0,0,0,201,0,0,0,99,0,0,0,113,0,232,0,40,0,0,0,0,0,19,0,224,0,229,0,90,0,39,0,83,0,0,0,61,0,19,0,0,0,0,0,194,0,42,0,86,0,22,0,29,0,0,0,0,0,0,0,72,0,216,0,142,0,0,0,0,0,13,0,190,0,61,0,163,0,0,0,222,0,167,0,210,0,0,0,59,0,21,0,0,0,137,0,16,0,162,0,0,0,110,0,76,0,51,0,88,0,0,0,0,0,150,0,55,0,251,0,87,0,15,0,0,0,5,0,75,0,10,0,157,0,157,0,0,0,155,0,57,0,185,0,117,0,215,0,174,0,0,0,0,0,212,0,152,0,30,0,0,0,222,0,239,0,34,0,62,0,164,0,0,0,60,0,154,0,0,0,0,0,248,0,0,0,192,0,0,0,209,0,0,0,0,0,220,0,215,0,49,0,26,0,20,0,25,0,246,0,147,0,74,0,91,0,0,0,0,0,164,0,0,0,0,0,170,0,34,0,0,0,96,0,231,0,45,0,184,0,0,0,168,0,0,0,14,0,128,0,148,0,123,0,191,0,214,0,180,0,216,0,246,0,235,0,105,0,0,0,0,0,77,0,69,0,223,0,0,0,138,0,197,0,17,0,246,0,225,0,46,0,59,0,97,0,0,0,53,0,230,0,0,0,0,0,31,0,247,0,5,0,135,0,92,0,218,0,83,0,66,0,8,0,0,0,101,0,131,0,255,0,0,0,0,0,0,0,175,0,252,0,94,0,0,0,216,0,49,0,0,0,243,0,133,0,226,0,215,0,0,0,0,0,76,0,7,0,63,0,73,0,62,0,215,0,175,0,3,0,151,0,164,0,136,0,0,0,0,0,0,0,157,0,28,0,84,0,88,0,144,0,0,0,45,0,74,0,178,0,73,0,128,0,183,0,70,0,81,0,191,0,114,0,156,0,86,0,0,0,245,0,0,0,231,0,0,0,191,0,54,0,180,0,44,0,194,0,0,0,0,0,0,0,226,0,69,0,1,0,56,0,180,0,229,0,246,0,150,0,0,0,234,0,69,0,0,0,219,0,100,0,74,0,0,0,0,0,247,0,244,0,66,0,255,0,67,0,0,0,150,0,250,0,0,0,159,0,236,0,33,0,28,0,195,0,62,0,226,0,199,0,72,0,89,0,108,0,203,0,0,0,239,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,0,0,75,31,251,31,81,31,231,31,90,31,66,31,168,31,168,30,113,31,180,31,17,31,126,31,126,30,255,31,198,31,221,31,249,31,167,31,21,31,21,30,21,29,21,28,21,27,21,26,2,31,45,31,235,31,89,31,101,31,10,31,24,31,84,31,162,31,223,31,28,31,212,31,183,31,183,30,183,29,77,31,244,31,244,30,245,31,54,31,7,31,20,31,177,31,159,31,159,30,159,29,159,28,82,31,232,31,5,31,120,31,94,31,94,30,243,31,66,31,137,31,129,31,165,31,62,31,74,31,74,30,74,29,201,31,201,30,99,31,99,30,113,31,232,31,40,31,40,30,40,29,19,31,224,31,229,31,90,31,39,31,83,31,83,30,61,31,19,31,19,30,19,29,194,31,42,31,86,31,22,31,29,31,29,30,29,29,29,28,72,31,216,31,142,31,142,30,142,29,13,31,190,31,61,31,163,31,163,30,222,31,167,31,210,31,210,30,59,31,21,31,21,30,137,31,16,31,162,31,162,30,110,31,76,31,51,31,88,31,88,30,88,29,150,31,55,31,251,31,87,31,15,31,15,30,5,31,75,31,10,31,157,31,157,31,157,30,155,31,57,31,185,31,117,31,215,31,174,31,174,30,174,29,212,31,152,31,30,31,30,30,222,31,239,31,34,31,62,31,164,31,164,30,60,31,154,31,154,30,154,29,248,31,248,30,192,31,192,30,209,31,209,30,209,29,220,31,215,31,49,31,26,31,20,31,25,31,246,31,147,31,74,31,91,31,91,30,91,29,164,31,164,30,164,29,170,31,34,31,34,30,96,31,231,31,45,31,184,31,184,30,168,31,168,30,14,31,128,31,148,31,123,31,191,31,214,31,180,31,216,31,246,31,235,31,105,31,105,30,105,29,77,31,69,31,223,31,223,30,138,31,197,31,17,31,246,31,225,31,46,31,59,31,97,31,97,30,53,31,230,31,230,30,230,29,31,31,247,31,5,31,135,31,92,31,218,31,83,31,66,31,8,31,8,30,101,31,131,31,255,31,255,30,255,29,255,28,175,31,252,31,94,31,94,30,216,31,49,31,49,30,243,31,133,31,226,31,215,31,215,30,215,29,76,31,7,31,63,31,73,31,62,31,215,31,175,31,3,31,151,31,164,31,136,31,136,30,136,29,136,28,157,31,28,31,84,31,88,31,144,31,144,30,45,31,74,31,178,31,73,31,128,31,183,31,70,31,81,31,191,31,114,31,156,31,86,31,86,30,245,31,245,30,231,31,231,30,191,31,54,31,180,31,44,31,194,31,194,30,194,29,194,28,226,31,69,31,1,31,56,31,180,31,229,31,246,31,150,31,150,30,234,31,69,31,69,30,219,31,100,31,74,31,74,30,74,29,247,31,244,31,66,31,255,31,67,31,67,30,150,31,250,31,250,30,159,31,236,31,33,31,28,31,195,31,62,31,226,31,199,31,72,31,89,31,108,31,203,31,203,30,239,31,239,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
