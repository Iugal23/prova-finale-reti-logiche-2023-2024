-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 227;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (127,0,154,0,230,0,175,0,194,0,222,0,192,0,79,0,0,0,0,0,221,0,146,0,136,0,112,0,178,0,206,0,115,0,160,0,189,0,132,0,134,0,18,0,0,0,253,0,0,0,173,0,102,0,98,0,198,0,34,0,120,0,50,0,0,0,161,0,66,0,0,0,188,0,0,0,81,0,106,0,18,0,79,0,137,0,246,0,254,0,193,0,249,0,6,0,21,0,36,0,170,0,58,0,5,0,119,0,130,0,86,0,93,0,0,0,2,0,193,0,102,0,0,0,120,0,170,0,4,0,0,0,25,0,171,0,4,0,0,0,0,0,0,0,161,0,35,0,202,0,0,0,8,0,63,0,89,0,0,0,55,0,41,0,170,0,217,0,72,0,114,0,0,0,169,0,26,0,182,0,0,0,232,0,198,0,146,0,162,0,148,0,0,0,203,0,149,0,254,0,20,0,50,0,0,0,0,0,0,0,36,0,125,0,128,0,0,0,152,0,13,0,135,0,120,0,151,0,158,0,0,0,154,0,0,0,91,0,79,0,0,0,14,0,75,0,178,0,39,0,31,0,0,0,37,0,134,0,189,0,0,0,65,0,178,0,0,0,13,0,61,0,0,0,0,0,0,0,16,0,0,0,203,0,54,0,3,0,54,0,0,0,0,0,11,0,31,0,79,0,74,0,169,0,82,0,16,0,185,0,0,0,48,0,166,0,103,0,35,0,130,0,195,0,192,0,147,0,0,0,150,0,110,0,62,0,171,0,162,0,93,0,174,0,143,0,135,0,51,0,75,0,250,0,38,0,45,0,123,0,65,0,49,0,190,0,232,0,76,0,233,0,153,0,189,0,0,0,239,0,51,0,0,0,161,0,233,0,254,0,126,0,4,0,135,0,46,0,0,0,208,0,194,0,26,0,76,0,168,0,0,0,20,0,0,0,200,0,57,0,13,0,24,0,185,0,106,0,251,0,213,0,77,0,0,0,10,0,12,0,126,0,65,0,164,0,234,0,0,0,179,0,136,0);
signal scenario_full  : scenario_type := (127,31,154,31,230,31,175,31,194,31,222,31,192,31,79,31,79,30,79,29,221,31,146,31,136,31,112,31,178,31,206,31,115,31,160,31,189,31,132,31,134,31,18,31,18,30,253,31,253,30,173,31,102,31,98,31,198,31,34,31,120,31,50,31,50,30,161,31,66,31,66,30,188,31,188,30,81,31,106,31,18,31,79,31,137,31,246,31,254,31,193,31,249,31,6,31,21,31,36,31,170,31,58,31,5,31,119,31,130,31,86,31,93,31,93,30,2,31,193,31,102,31,102,30,120,31,170,31,4,31,4,30,25,31,171,31,4,31,4,30,4,29,4,28,161,31,35,31,202,31,202,30,8,31,63,31,89,31,89,30,55,31,41,31,170,31,217,31,72,31,114,31,114,30,169,31,26,31,182,31,182,30,232,31,198,31,146,31,162,31,148,31,148,30,203,31,149,31,254,31,20,31,50,31,50,30,50,29,50,28,36,31,125,31,128,31,128,30,152,31,13,31,135,31,120,31,151,31,158,31,158,30,154,31,154,30,91,31,79,31,79,30,14,31,75,31,178,31,39,31,31,31,31,30,37,31,134,31,189,31,189,30,65,31,178,31,178,30,13,31,61,31,61,30,61,29,61,28,16,31,16,30,203,31,54,31,3,31,54,31,54,30,54,29,11,31,31,31,79,31,74,31,169,31,82,31,16,31,185,31,185,30,48,31,166,31,103,31,35,31,130,31,195,31,192,31,147,31,147,30,150,31,110,31,62,31,171,31,162,31,93,31,174,31,143,31,135,31,51,31,75,31,250,31,38,31,45,31,123,31,65,31,49,31,190,31,232,31,76,31,233,31,153,31,189,31,189,30,239,31,51,31,51,30,161,31,233,31,254,31,126,31,4,31,135,31,46,31,46,30,208,31,194,31,26,31,76,31,168,31,168,30,20,31,20,30,200,31,57,31,13,31,24,31,185,31,106,31,251,31,213,31,77,31,77,30,10,31,12,31,126,31,65,31,164,31,234,31,234,30,179,31,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
