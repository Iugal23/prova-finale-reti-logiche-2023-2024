-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 947;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,252,0,101,0,200,0,90,0,56,0,8,0,71,0,87,0,0,0,31,0,157,0,0,0,35,0,133,0,53,0,0,0,232,0,206,0,59,0,104,0,155,0,201,0,95,0,0,0,45,0,246,0,98,0,219,0,222,0,0,0,106,0,0,0,86,0,182,0,18,0,247,0,169,0,0,0,103,0,107,0,55,0,143,0,74,0,239,0,208,0,23,0,182,0,184,0,138,0,201,0,105,0,102,0,18,0,11,0,0,0,119,0,3,0,33,0,130,0,246,0,228,0,168,0,117,0,9,0,112,0,145,0,177,0,120,0,0,0,137,0,223,0,4,0,243,0,248,0,87,0,33,0,59,0,18,0,246,0,138,0,189,0,116,0,195,0,215,0,95,0,220,0,197,0,108,0,232,0,0,0,72,0,76,0,220,0,192,0,56,0,0,0,0,0,143,0,234,0,97,0,198,0,213,0,195,0,7,0,0,0,129,0,42,0,166,0,135,0,111,0,77,0,0,0,193,0,0,0,69,0,217,0,0,0,0,0,140,0,0,0,222,0,182,0,143,0,0,0,70,0,0,0,0,0,254,0,193,0,221,0,233,0,234,0,97,0,87,0,234,0,0,0,80,0,0,0,18,0,86,0,65,0,26,0,175,0,155,0,48,0,175,0,0,0,16,0,191,0,17,0,69,0,153,0,43,0,57,0,47,0,41,0,74,0,123,0,0,0,220,0,0,0,175,0,139,0,32,0,168,0,114,0,245,0,0,0,161,0,192,0,185,0,20,0,168,0,193,0,121,0,252,0,209,0,69,0,208,0,172,0,0,0,77,0,195,0,250,0,75,0,108,0,2,0,65,0,0,0,70,0,111,0,0,0,60,0,152,0,139,0,62,0,208,0,103,0,60,0,79,0,231,0,0,0,0,0,180,0,60,0,73,0,203,0,7,0,81,0,111,0,0,0,154,0,201,0,233,0,185,0,0,0,125,0,103,0,181,0,148,0,243,0,0,0,136,0,205,0,2,0,185,0,8,0,193,0,166,0,0,0,75,0,0,0,213,0,246,0,0,0,193,0,86,0,0,0,38,0,0,0,209,0,80,0,65,0,129,0,189,0,83,0,150,0,0,0,0,0,0,0,8,0,8,0,6,0,60,0,178,0,0,0,12,0,0,0,0,0,95,0,0,0,28,0,0,0,17,0,87,0,0,0,103,0,119,0,13,0,164,0,126,0,0,0,78,0,0,0,237,0,252,0,242,0,240,0,213,0,154,0,30,0,243,0,151,0,128,0,185,0,157,0,143,0,247,0,0,0,0,0,247,0,49,0,74,0,192,0,102,0,252,0,245,0,197,0,8,0,186,0,38,0,62,0,254,0,240,0,49,0,161,0,112,0,26,0,101,0,146,0,0,0,226,0,0,0,36,0,242,0,112,0,123,0,145,0,23,0,29,0,0,0,0,0,0,0,0,0,32,0,255,0,170,0,144,0,0,0,120,0,22,0,0,0,216,0,54,0,0,0,28,0,205,0,201,0,140,0,0,0,100,0,227,0,22,0,178,0,158,0,0,0,83,0,0,0,26,0,128,0,0,0,0,0,156,0,104,0,189,0,160,0,67,0,0,0,116,0,34,0,187,0,164,0,25,0,129,0,0,0,7,0,0,0,0,0,74,0,207,0,102,0,0,0,199,0,0,0,162,0,158,0,103,0,3,0,155,0,120,0,166,0,136,0,62,0,81,0,43,0,64,0,149,0,246,0,104,0,46,0,222,0,96,0,0,0,76,0,79,0,12,0,215,0,19,0,186,0,87,0,0,0,64,0,74,0,134,0,0,0,138,0,213,0,239,0,89,0,0,0,158,0,242,0,148,0,35,0,0,0,10,0,233,0,252,0,0,0,230,0,58,0,114,0,93,0,119,0,157,0,183,0,0,0,0,0,0,0,25,0,65,0,194,0,52,0,255,0,167,0,29,0,123,0,0,0,146,0,205,0,141,0,202,0,116,0,6,0,255,0,0,0,179,0,0,0,210,0,0,0,253,0,144,0,0,0,56,0,65,0,142,0,4,0,104,0,238,0,220,0,52,0,17,0,0,0,30,0,184,0,166,0,50,0,230,0,34,0,69,0,29,0,245,0,115,0,197,0,0,0,63,0,12,0,0,0,169,0,245,0,248,0,204,0,0,0,0,0,192,0,216,0,145,0,121,0,110,0,56,0,253,0,0,0,241,0,154,0,30,0,68,0,100,0,156,0,239,0,0,0,0,0,0,0,119,0,35,0,50,0,240,0,80,0,0,0,0,0,0,0,0,0,37,0,131,0,0,0,50,0,175,0,219,0,130,0,169,0,0,0,0,0,120,0,60,0,0,0,99,0,174,0,143,0,69,0,52,0,17,0,196,0,0,0,0,0,70,0,0,0,96,0,217,0,15,0,6,0,90,0,0,0,162,0,121,0,237,0,65,0,154,0,45,0,90,0,156,0,242,0,0,0,176,0,188,0,205,0,133,0,108,0,183,0,67,0,45,0,0,0,171,0,121,0,26,0,0,0,158,0,216,0,139,0,129,0,42,0,118,0,0,0,207,0,130,0,0,0,212,0,247,0,202,0,160,0,221,0,250,0,0,0,47,0,15,0,0,0,101,0,15,0,219,0,255,0,130,0,42,0,62,0,93,0,0,0,0,0,14,0,29,0,24,0,111,0,18,0,145,0,39,0,0,0,71,0,0,0,120,0,121,0,189,0,132,0,87,0,129,0,155,0,21,0,133,0,100,0,250,0,194,0,8,0,139,0,0,0,166,0,47,0,213,0,0,0,76,0,48,0,236,0,54,0,218,0,19,0,4,0,44,0,172,0,87,0,207,0,77,0,176,0,152,0,142,0,0,0,66,0,117,0,186,0,0,0,88,0,0,0,116,0,0,0,130,0,94,0,18,0,231,0,0,0,0,0,189,0,201,0,241,0,0,0,0,0,97,0,73,0,0,0,0,0,0,0,249,0,0,0,71,0,170,0,213,0,211,0,176,0,156,0,0,0,55,0,46,0,248,0,212,0,43,0,209,0,0,0,0,0,215,0,10,0,0,0,0,0,254,0,9,0,67,0,157,0,0,0,0,0,0,0,31,0,174,0,163,0,184,0,48,0,0,0,133,0,219,0,0,0,229,0,0,0,57,0,211,0,188,0,0,0,235,0,147,0,0,0,48,0,64,0,228,0,199,0,116,0,0,0,133,0,0,0,44,0,168,0,255,0,244,0,19,0,162,0,158,0,175,0,19,0,66,0,174,0,231,0,99,0,149,0,226,0,0,0,0,0,121,0,218,0,109,0,160,0,0,0,115,0,0,0,0,0,64,0,182,0,220,0,108,0,108,0,46,0,0,0,0,0,0,0,0,0,0,0,25,0,244,0,141,0,0,0,195,0,243,0,0,0,104,0,85,0,192,0,165,0,214,0,181,0,45,0,70,0,13,0,11,0,227,0,203,0,0,0,254,0,233,0,40,0,95,0,207,0,54,0,85,0,237,0,0,0,86,0,149,0,21,0,188,0,106,0,10,0,48,0,27,0,82,0,167,0,180,0,0,0,0,0,0,0,138,0,138,0,105,0,0,0,0,0,0,0,122,0,104,0,125,0,144,0,173,0,0,0,195,0,0,0,151,0,19,0,16,0,0,0,0,0,97,0,0,0,175,0,75,0,144,0,55,0,216,0,0,0,221,0,247,0,29,0,136,0,158,0,0,0,156,0,231,0,83,0,202,0,136,0,122,0,104,0,30,0,95,0,128,0,223,0,100,0,0,0,49,0,0,0,83,0,9,0,0,0,33,0,98,0,173,0,120,0,177,0,53,0,115,0,0,0,242,0,156,0,149,0,30,0,220,0,0,0,107,0,239,0,6,0,0,0,222,0,188,0,0,0,0,0,137,0,71,0,111,0,140,0,251,0,67,0,0,0,63,0,187,0,146,0,0,0,10,0,0,0,0,0,173,0,194,0,18,0,167,0,0,0,169,0,149,0,102,0,182,0,90,0,0,0,184,0,121,0,105,0,184,0,93,0,170,0,0,0,104,0,151,0,200,0,103,0,52,0,0,0,11,0,34,0,50,0,51,0,140,0,18,0,235,0,189,0,63,0,12,0,182,0,118,0,56,0,37,0,91,0,40,0,39,0,0,0,200,0,12,0,102,0,108,0,121,0,212,0,46,0,32,0,245,0,0,0,0,0,10,0,199,0,0,0,225,0,27,0,72,0,7,0,108,0,149,0,73,0);
signal scenario_full  : scenario_type := (95,31,252,31,101,31,200,31,90,31,56,31,8,31,71,31,87,31,87,30,31,31,157,31,157,30,35,31,133,31,53,31,53,30,232,31,206,31,59,31,104,31,155,31,201,31,95,31,95,30,45,31,246,31,98,31,219,31,222,31,222,30,106,31,106,30,86,31,182,31,18,31,247,31,169,31,169,30,103,31,107,31,55,31,143,31,74,31,239,31,208,31,23,31,182,31,184,31,138,31,201,31,105,31,102,31,18,31,11,31,11,30,119,31,3,31,33,31,130,31,246,31,228,31,168,31,117,31,9,31,112,31,145,31,177,31,120,31,120,30,137,31,223,31,4,31,243,31,248,31,87,31,33,31,59,31,18,31,246,31,138,31,189,31,116,31,195,31,215,31,95,31,220,31,197,31,108,31,232,31,232,30,72,31,76,31,220,31,192,31,56,31,56,30,56,29,143,31,234,31,97,31,198,31,213,31,195,31,7,31,7,30,129,31,42,31,166,31,135,31,111,31,77,31,77,30,193,31,193,30,69,31,217,31,217,30,217,29,140,31,140,30,222,31,182,31,143,31,143,30,70,31,70,30,70,29,254,31,193,31,221,31,233,31,234,31,97,31,87,31,234,31,234,30,80,31,80,30,18,31,86,31,65,31,26,31,175,31,155,31,48,31,175,31,175,30,16,31,191,31,17,31,69,31,153,31,43,31,57,31,47,31,41,31,74,31,123,31,123,30,220,31,220,30,175,31,139,31,32,31,168,31,114,31,245,31,245,30,161,31,192,31,185,31,20,31,168,31,193,31,121,31,252,31,209,31,69,31,208,31,172,31,172,30,77,31,195,31,250,31,75,31,108,31,2,31,65,31,65,30,70,31,111,31,111,30,60,31,152,31,139,31,62,31,208,31,103,31,60,31,79,31,231,31,231,30,231,29,180,31,60,31,73,31,203,31,7,31,81,31,111,31,111,30,154,31,201,31,233,31,185,31,185,30,125,31,103,31,181,31,148,31,243,31,243,30,136,31,205,31,2,31,185,31,8,31,193,31,166,31,166,30,75,31,75,30,213,31,246,31,246,30,193,31,86,31,86,30,38,31,38,30,209,31,80,31,65,31,129,31,189,31,83,31,150,31,150,30,150,29,150,28,8,31,8,31,6,31,60,31,178,31,178,30,12,31,12,30,12,29,95,31,95,30,28,31,28,30,17,31,87,31,87,30,103,31,119,31,13,31,164,31,126,31,126,30,78,31,78,30,237,31,252,31,242,31,240,31,213,31,154,31,30,31,243,31,151,31,128,31,185,31,157,31,143,31,247,31,247,30,247,29,247,31,49,31,74,31,192,31,102,31,252,31,245,31,197,31,8,31,186,31,38,31,62,31,254,31,240,31,49,31,161,31,112,31,26,31,101,31,146,31,146,30,226,31,226,30,36,31,242,31,112,31,123,31,145,31,23,31,29,31,29,30,29,29,29,28,29,27,32,31,255,31,170,31,144,31,144,30,120,31,22,31,22,30,216,31,54,31,54,30,28,31,205,31,201,31,140,31,140,30,100,31,227,31,22,31,178,31,158,31,158,30,83,31,83,30,26,31,128,31,128,30,128,29,156,31,104,31,189,31,160,31,67,31,67,30,116,31,34,31,187,31,164,31,25,31,129,31,129,30,7,31,7,30,7,29,74,31,207,31,102,31,102,30,199,31,199,30,162,31,158,31,103,31,3,31,155,31,120,31,166,31,136,31,62,31,81,31,43,31,64,31,149,31,246,31,104,31,46,31,222,31,96,31,96,30,76,31,79,31,12,31,215,31,19,31,186,31,87,31,87,30,64,31,74,31,134,31,134,30,138,31,213,31,239,31,89,31,89,30,158,31,242,31,148,31,35,31,35,30,10,31,233,31,252,31,252,30,230,31,58,31,114,31,93,31,119,31,157,31,183,31,183,30,183,29,183,28,25,31,65,31,194,31,52,31,255,31,167,31,29,31,123,31,123,30,146,31,205,31,141,31,202,31,116,31,6,31,255,31,255,30,179,31,179,30,210,31,210,30,253,31,144,31,144,30,56,31,65,31,142,31,4,31,104,31,238,31,220,31,52,31,17,31,17,30,30,31,184,31,166,31,50,31,230,31,34,31,69,31,29,31,245,31,115,31,197,31,197,30,63,31,12,31,12,30,169,31,245,31,248,31,204,31,204,30,204,29,192,31,216,31,145,31,121,31,110,31,56,31,253,31,253,30,241,31,154,31,30,31,68,31,100,31,156,31,239,31,239,30,239,29,239,28,119,31,35,31,50,31,240,31,80,31,80,30,80,29,80,28,80,27,37,31,131,31,131,30,50,31,175,31,219,31,130,31,169,31,169,30,169,29,120,31,60,31,60,30,99,31,174,31,143,31,69,31,52,31,17,31,196,31,196,30,196,29,70,31,70,30,96,31,217,31,15,31,6,31,90,31,90,30,162,31,121,31,237,31,65,31,154,31,45,31,90,31,156,31,242,31,242,30,176,31,188,31,205,31,133,31,108,31,183,31,67,31,45,31,45,30,171,31,121,31,26,31,26,30,158,31,216,31,139,31,129,31,42,31,118,31,118,30,207,31,130,31,130,30,212,31,247,31,202,31,160,31,221,31,250,31,250,30,47,31,15,31,15,30,101,31,15,31,219,31,255,31,130,31,42,31,62,31,93,31,93,30,93,29,14,31,29,31,24,31,111,31,18,31,145,31,39,31,39,30,71,31,71,30,120,31,121,31,189,31,132,31,87,31,129,31,155,31,21,31,133,31,100,31,250,31,194,31,8,31,139,31,139,30,166,31,47,31,213,31,213,30,76,31,48,31,236,31,54,31,218,31,19,31,4,31,44,31,172,31,87,31,207,31,77,31,176,31,152,31,142,31,142,30,66,31,117,31,186,31,186,30,88,31,88,30,116,31,116,30,130,31,94,31,18,31,231,31,231,30,231,29,189,31,201,31,241,31,241,30,241,29,97,31,73,31,73,30,73,29,73,28,249,31,249,30,71,31,170,31,213,31,211,31,176,31,156,31,156,30,55,31,46,31,248,31,212,31,43,31,209,31,209,30,209,29,215,31,10,31,10,30,10,29,254,31,9,31,67,31,157,31,157,30,157,29,157,28,31,31,174,31,163,31,184,31,48,31,48,30,133,31,219,31,219,30,229,31,229,30,57,31,211,31,188,31,188,30,235,31,147,31,147,30,48,31,64,31,228,31,199,31,116,31,116,30,133,31,133,30,44,31,168,31,255,31,244,31,19,31,162,31,158,31,175,31,19,31,66,31,174,31,231,31,99,31,149,31,226,31,226,30,226,29,121,31,218,31,109,31,160,31,160,30,115,31,115,30,115,29,64,31,182,31,220,31,108,31,108,31,46,31,46,30,46,29,46,28,46,27,46,26,25,31,244,31,141,31,141,30,195,31,243,31,243,30,104,31,85,31,192,31,165,31,214,31,181,31,45,31,70,31,13,31,11,31,227,31,203,31,203,30,254,31,233,31,40,31,95,31,207,31,54,31,85,31,237,31,237,30,86,31,149,31,21,31,188,31,106,31,10,31,48,31,27,31,82,31,167,31,180,31,180,30,180,29,180,28,138,31,138,31,105,31,105,30,105,29,105,28,122,31,104,31,125,31,144,31,173,31,173,30,195,31,195,30,151,31,19,31,16,31,16,30,16,29,97,31,97,30,175,31,75,31,144,31,55,31,216,31,216,30,221,31,247,31,29,31,136,31,158,31,158,30,156,31,231,31,83,31,202,31,136,31,122,31,104,31,30,31,95,31,128,31,223,31,100,31,100,30,49,31,49,30,83,31,9,31,9,30,33,31,98,31,173,31,120,31,177,31,53,31,115,31,115,30,242,31,156,31,149,31,30,31,220,31,220,30,107,31,239,31,6,31,6,30,222,31,188,31,188,30,188,29,137,31,71,31,111,31,140,31,251,31,67,31,67,30,63,31,187,31,146,31,146,30,10,31,10,30,10,29,173,31,194,31,18,31,167,31,167,30,169,31,149,31,102,31,182,31,90,31,90,30,184,31,121,31,105,31,184,31,93,31,170,31,170,30,104,31,151,31,200,31,103,31,52,31,52,30,11,31,34,31,50,31,51,31,140,31,18,31,235,31,189,31,63,31,12,31,182,31,118,31,56,31,37,31,91,31,40,31,39,31,39,30,200,31,12,31,102,31,108,31,121,31,212,31,46,31,32,31,245,31,245,30,245,29,10,31,199,31,199,30,225,31,27,31,72,31,7,31,108,31,149,31,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
