-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 471;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,148,0,113,0,100,0,224,0,0,0,205,0,0,0,49,0,36,0,70,0,23,0,110,0,39,0,66,0,0,0,252,0,112,0,71,0,232,0,37,0,0,0,54,0,202,0,119,0,209,0,0,0,209,0,25,0,112,0,0,0,204,0,12,0,0,0,27,0,151,0,66,0,149,0,0,0,6,0,14,0,0,0,0,0,116,0,0,0,235,0,63,0,0,0,87,0,129,0,246,0,32,0,122,0,12,0,52,0,195,0,114,0,243,0,113,0,107,0,0,0,0,0,196,0,174,0,207,0,8,0,0,0,17,0,223,0,47,0,202,0,0,0,233,0,0,0,185,0,126,0,87,0,42,0,40,0,58,0,21,0,121,0,164,0,24,0,82,0,9,0,65,0,138,0,0,0,19,0,14,0,48,0,82,0,243,0,0,0,74,0,101,0,151,0,17,0,247,0,0,0,251,0,48,0,192,0,27,0,172,0,107,0,0,0,26,0,212,0,14,0,206,0,102,0,19,0,106,0,156,0,118,0,28,0,67,0,187,0,192,0,216,0,34,0,203,0,187,0,0,0,247,0,101,0,167,0,73,0,152,0,0,0,0,0,234,0,215,0,238,0,4,0,231,0,35,0,98,0,251,0,133,0,145,0,10,0,234,0,25,0,59,0,0,0,107,0,160,0,50,0,152,0,160,0,0,0,0,0,209,0,200,0,228,0,106,0,36,0,0,0,118,0,64,0,52,0,9,0,0,0,45,0,0,0,199,0,26,0,173,0,0,0,124,0,0,0,12,0,130,0,87,0,58,0,27,0,49,0,242,0,165,0,221,0,29,0,17,0,206,0,72,0,153,0,9,0,73,0,157,0,75,0,0,0,174,0,255,0,75,0,30,0,195,0,83,0,168,0,96,0,171,0,201,0,0,0,0,0,0,0,11,0,0,0,193,0,57,0,160,0,0,0,44,0,89,0,91,0,32,0,111,0,97,0,81,0,235,0,0,0,14,0,176,0,131,0,36,0,0,0,208,0,240,0,145,0,22,0,253,0,106,0,131,0,119,0,39,0,31,0,247,0,67,0,122,0,205,0,0,0,0,0,54,0,80,0,172,0,134,0,0,0,222,0,140,0,211,0,244,0,53,0,136,0,208,0,65,0,143,0,119,0,0,0,143,0,0,0,73,0,0,0,25,0,64,0,66,0,0,0,93,0,175,0,18,0,229,0,206,0,0,0,83,0,138,0,238,0,194,0,216,0,244,0,32,0,119,0,0,0,91,0,74,0,12,0,5,0,125,0,96,0,125,0,248,0,0,0,74,0,190,0,143,0,80,0,103,0,6,0,149,0,143,0,211,0,86,0,142,0,176,0,243,0,60,0,0,0,250,0,0,0,81,0,0,0,0,0,166,0,228,0,17,0,82,0,172,0,0,0,0,0,229,0,88,0,126,0,10,0,154,0,67,0,208,0,0,0,44,0,134,0,211,0,248,0,138,0,148,0,108,0,0,0,31,0,3,0,165,0,222,0,11,0,0,0,50,0,117,0,56,0,0,0,0,0,196,0,182,0,39,0,0,0,7,0,195,0,0,0,145,0,113,0,25,0,76,0,208,0,22,0,0,0,58,0,245,0,0,0,0,0,0,0,0,0,17,0,0,0,0,0,189,0,120,0,252,0,75,0,0,0,102,0,76,0,22,0,36,0,112,0,245,0,99,0,41,0,0,0,39,0,221,0,120,0,246,0,252,0,0,0,0,0,0,0,245,0,72,0,0,0,21,0,76,0,0,0,0,0,11,0,81,0,156,0,187,0,13,0,181,0,216,0,107,0,225,0,50,0,12,0,119,0,0,0,130,0,48,0,95,0,172,0,26,0,42,0,0,0,164,0,251,0,43,0,245,0,0,0,250,0,0,0,0,0,247,0,116,0,248,0,254,0,191,0,92,0,38,0,140,0,147,0,166,0,215,0,155,0,188,0,21,0,123,0,107,0,216,0,0,0,152,0,205,0,199,0,163,0,0,0,95,0,170,0,91,0,0,0,0,0,159,0,242,0,126,0,46,0,129,0,164,0,212,0,127,0,189,0,2,0,216,0,231,0,17,0,116,0,116,0,128,0,130,0,0,0,0,0);
signal scenario_full  : scenario_type := (149,31,148,31,113,31,100,31,224,31,224,30,205,31,205,30,49,31,36,31,70,31,23,31,110,31,39,31,66,31,66,30,252,31,112,31,71,31,232,31,37,31,37,30,54,31,202,31,119,31,209,31,209,30,209,31,25,31,112,31,112,30,204,31,12,31,12,30,27,31,151,31,66,31,149,31,149,30,6,31,14,31,14,30,14,29,116,31,116,30,235,31,63,31,63,30,87,31,129,31,246,31,32,31,122,31,12,31,52,31,195,31,114,31,243,31,113,31,107,31,107,30,107,29,196,31,174,31,207,31,8,31,8,30,17,31,223,31,47,31,202,31,202,30,233,31,233,30,185,31,126,31,87,31,42,31,40,31,58,31,21,31,121,31,164,31,24,31,82,31,9,31,65,31,138,31,138,30,19,31,14,31,48,31,82,31,243,31,243,30,74,31,101,31,151,31,17,31,247,31,247,30,251,31,48,31,192,31,27,31,172,31,107,31,107,30,26,31,212,31,14,31,206,31,102,31,19,31,106,31,156,31,118,31,28,31,67,31,187,31,192,31,216,31,34,31,203,31,187,31,187,30,247,31,101,31,167,31,73,31,152,31,152,30,152,29,234,31,215,31,238,31,4,31,231,31,35,31,98,31,251,31,133,31,145,31,10,31,234,31,25,31,59,31,59,30,107,31,160,31,50,31,152,31,160,31,160,30,160,29,209,31,200,31,228,31,106,31,36,31,36,30,118,31,64,31,52,31,9,31,9,30,45,31,45,30,199,31,26,31,173,31,173,30,124,31,124,30,12,31,130,31,87,31,58,31,27,31,49,31,242,31,165,31,221,31,29,31,17,31,206,31,72,31,153,31,9,31,73,31,157,31,75,31,75,30,174,31,255,31,75,31,30,31,195,31,83,31,168,31,96,31,171,31,201,31,201,30,201,29,201,28,11,31,11,30,193,31,57,31,160,31,160,30,44,31,89,31,91,31,32,31,111,31,97,31,81,31,235,31,235,30,14,31,176,31,131,31,36,31,36,30,208,31,240,31,145,31,22,31,253,31,106,31,131,31,119,31,39,31,31,31,247,31,67,31,122,31,205,31,205,30,205,29,54,31,80,31,172,31,134,31,134,30,222,31,140,31,211,31,244,31,53,31,136,31,208,31,65,31,143,31,119,31,119,30,143,31,143,30,73,31,73,30,25,31,64,31,66,31,66,30,93,31,175,31,18,31,229,31,206,31,206,30,83,31,138,31,238,31,194,31,216,31,244,31,32,31,119,31,119,30,91,31,74,31,12,31,5,31,125,31,96,31,125,31,248,31,248,30,74,31,190,31,143,31,80,31,103,31,6,31,149,31,143,31,211,31,86,31,142,31,176,31,243,31,60,31,60,30,250,31,250,30,81,31,81,30,81,29,166,31,228,31,17,31,82,31,172,31,172,30,172,29,229,31,88,31,126,31,10,31,154,31,67,31,208,31,208,30,44,31,134,31,211,31,248,31,138,31,148,31,108,31,108,30,31,31,3,31,165,31,222,31,11,31,11,30,50,31,117,31,56,31,56,30,56,29,196,31,182,31,39,31,39,30,7,31,195,31,195,30,145,31,113,31,25,31,76,31,208,31,22,31,22,30,58,31,245,31,245,30,245,29,245,28,245,27,17,31,17,30,17,29,189,31,120,31,252,31,75,31,75,30,102,31,76,31,22,31,36,31,112,31,245,31,99,31,41,31,41,30,39,31,221,31,120,31,246,31,252,31,252,30,252,29,252,28,245,31,72,31,72,30,21,31,76,31,76,30,76,29,11,31,81,31,156,31,187,31,13,31,181,31,216,31,107,31,225,31,50,31,12,31,119,31,119,30,130,31,48,31,95,31,172,31,26,31,42,31,42,30,164,31,251,31,43,31,245,31,245,30,250,31,250,30,250,29,247,31,116,31,248,31,254,31,191,31,92,31,38,31,140,31,147,31,166,31,215,31,155,31,188,31,21,31,123,31,107,31,216,31,216,30,152,31,205,31,199,31,163,31,163,30,95,31,170,31,91,31,91,30,91,29,159,31,242,31,126,31,46,31,129,31,164,31,212,31,127,31,189,31,2,31,216,31,231,31,17,31,116,31,116,31,128,31,130,31,130,30,130,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
