-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 874;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (55,0,38,0,57,0,243,0,0,0,0,0,96,0,23,0,0,0,101,0,68,0,42,0,18,0,38,0,158,0,164,0,250,0,24,0,27,0,109,0,55,0,0,0,0,0,219,0,21,0,171,0,131,0,207,0,39,0,139,0,0,0,143,0,70,0,0,0,156,0,195,0,240,0,3,0,186,0,237,0,80,0,241,0,8,0,187,0,0,0,140,0,190,0,215,0,121,0,223,0,0,0,181,0,121,0,149,0,210,0,200,0,50,0,245,0,0,0,162,0,138,0,0,0,181,0,223,0,30,0,187,0,121,0,66,0,140,0,178,0,165,0,102,0,1,0,216,0,44,0,221,0,0,0,38,0,0,0,150,0,17,0,175,0,59,0,193,0,249,0,249,0,71,0,0,0,115,0,0,0,51,0,124,0,191,0,167,0,172,0,28,0,97,0,0,0,0,0,0,0,62,0,0,0,62,0,235,0,126,0,0,0,223,0,222,0,204,0,223,0,14,0,67,0,191,0,0,0,64,0,134,0,203,0,128,0,82,0,118,0,30,0,198,0,210,0,208,0,105,0,213,0,180,0,17,0,205,0,31,0,222,0,67,0,8,0,47,0,119,0,167,0,124,0,107,0,243,0,0,0,4,0,232,0,164,0,43,0,61,0,177,0,137,0,0,0,33,0,1,0,0,0,24,0,206,0,193,0,204,0,66,0,144,0,0,0,28,0,72,0,163,0,3,0,193,0,12,0,120,0,181,0,137,0,144,0,63,0,167,0,232,0,159,0,214,0,170,0,14,0,122,0,87,0,140,0,155,0,53,0,138,0,79,0,9,0,104,0,87,0,141,0,40,0,100,0,126,0,142,0,147,0,94,0,64,0,0,0,198,0,174,0,81,0,194,0,102,0,25,0,172,0,190,0,0,0,0,0,0,0,0,0,170,0,0,0,172,0,0,0,67,0,180,0,240,0,108,0,95,0,0,0,254,0,213,0,0,0,247,0,92,0,176,0,129,0,0,0,231,0,89,0,0,0,128,0,251,0,160,0,0,0,130,0,218,0,154,0,245,0,0,0,155,0,238,0,0,0,32,0,180,0,58,0,132,0,115,0,176,0,138,0,0,0,0,0,221,0,100,0,207,0,101,0,69,0,78,0,0,0,251,0,113,0,244,0,78,0,178,0,16,0,141,0,105,0,160,0,47,0,38,0,238,0,34,0,4,0,208,0,0,0,180,0,194,0,169,0,217,0,40,0,0,0,38,0,231,0,215,0,196,0,0,0,20,0,132,0,0,0,0,0,13,0,162,0,117,0,157,0,39,0,90,0,186,0,141,0,231,0,37,0,216,0,240,0,64,0,147,0,0,0,150,0,0,0,205,0,10,0,45,0,162,0,115,0,115,0,246,0,241,0,202,0,97,0,254,0,85,0,170,0,0,0,42,0,146,0,234,0,70,0,62,0,96,0,187,0,199,0,208,0,122,0,0,0,40,0,203,0,247,0,26,0,0,0,94,0,157,0,209,0,28,0,0,0,47,0,5,0,136,0,214,0,186,0,0,0,140,0,130,0,159,0,203,0,70,0,185,0,119,0,242,0,4,0,0,0,229,0,232,0,206,0,207,0,0,0,174,0,39,0,13,0,128,0,16,0,211,0,147,0,134,0,18,0,233,0,116,0,0,0,14,0,160,0,0,0,0,0,193,0,88,0,81,0,174,0,0,0,0,0,45,0,0,0,165,0,149,0,232,0,117,0,20,0,69,0,35,0,167,0,168,0,58,0,212,0,79,0,0,0,15,0,0,0,116,0,214,0,186,0,36,0,115,0,213,0,50,0,10,0,233,0,0,0,0,0,2,0,246,0,92,0,168,0,118,0,58,0,33,0,228,0,204,0,134,0,62,0,71,0,0,0,63,0,197,0,149,0,129,0,51,0,210,0,203,0,0,0,0,0,45,0,254,0,207,0,0,0,7,0,114,0,0,0,145,0,0,0,120,0,3,0,206,0,108,0,124,0,0,0,0,0,0,0,140,0,0,0,197,0,0,0,181,0,154,0,201,0,0,0,185,0,153,0,103,0,0,0,36,0,241,0,193,0,225,0,144,0,194,0,0,0,41,0,232,0,154,0,33,0,11,0,70,0,110,0,99,0,67,0,220,0,112,0,108,0,0,0,169,0,178,0,0,0,53,0,44,0,237,0,137,0,87,0,98,0,251,0,0,0,232,0,195,0,0,0,174,0,27,0,0,0,100,0,43,0,33,0,152,0,122,0,6,0,153,0,6,0,65,0,92,0,132,0,91,0,155,0,58,0,136,0,43,0,85,0,73,0,0,0,176,0,14,0,19,0,83,0,236,0,0,0,62,0,160,0,22,0,92,0,226,0,0,0,15,0,141,0,0,0,55,0,170,0,0,0,233,0,180,0,215,0,0,0,231,0,130,0,32,0,80,0,188,0,0,0,31,0,192,0,0,0,254,0,17,0,0,0,89,0,50,0,129,0,154,0,118,0,0,0,149,0,155,0,33,0,27,0,33,0,210,0,179,0,109,0,202,0,47,0,117,0,0,0,0,0,0,0,219,0,204,0,0,0,11,0,122,0,0,0,0,0,109,0,188,0,138,0,175,0,135,0,67,0,195,0,8,0,0,0,147,0,254,0,217,0,130,0,153,0,68,0,250,0,184,0,115,0,242,0,203,0,221,0,213,0,245,0,101,0,212,0,41,0,111,0,0,0,0,0,36,0,75,0,162,0,163,0,203,0,86,0,92,0,0,0,9,0,0,0,0,0,57,0,213,0,0,0,73,0,0,0,41,0,235,0,239,0,14,0,15,0,241,0,135,0,0,0,247,0,252,0,168,0,54,0,153,0,0,0,240,0,2,0,0,0,0,0,218,0,7,0,0,0,76,0,5,0,0,0,65,0,177,0,0,0,53,0,223,0,0,0,0,0,127,0,0,0,49,0,19,0,209,0,237,0,232,0,0,0,200,0,0,0,0,0,161,0,0,0,182,0,0,0,62,0,111,0,221,0,17,0,35,0,212,0,0,0,0,0,241,0,70,0,250,0,126,0,60,0,138,0,52,0,220,0,0,0,118,0,0,0,83,0,115,0,149,0,138,0,220,0,197,0,5,0,84,0,189,0,0,0,103,0,218,0,232,0,223,0,34,0,149,0,182,0,133,0,30,0,199,0,185,0,0,0,30,0,131,0,90,0,82,0,247,0,76,0,42,0,0,0,150,0,174,0,211,0,115,0,202,0,125,0,200,0,0,0,0,0,143,0,64,0,109,0,233,0,0,0,136,0,208,0,251,0,1,0,158,0,56,0,236,0,121,0,0,0,94,0,140,0,78,0,100,0,198,0,26,0,239,0,222,0,152,0,170,0,155,0,210,0,228,0,249,0,187,0,145,0,26,0,178,0,255,0,30,0,180,0,0,0,130,0,173,0,222,0,50,0,203,0,112,0,63,0,0,0,236,0,0,0,131,0,100,0,0,0,208,0,0,0,0,0,236,0,75,0,0,0,219,0,74,0,173,0,0,0,246,0,4,0,39,0,161,0,20,0,0,0,234,0,122,0,193,0,0,0,0,0,176,0,78,0,180,0,92,0,51,0,0,0,0,0,36,0,122,0,90,0,77,0,20,0,169,0,0,0,44,0,0,0,0,0,0,0,167,0,188,0,0,0,246,0,0,0,205,0,64,0,179,0,0,0,198,0,222,0,199,0,251,0,123,0,171,0,194,0,61,0,36,0,244,0,239,0,209,0,244,0,60,0,225,0,167,0,229,0,0,0,246,0,123,0,42,0,63,0,139,0,95,0,42,0,97,0,78,0,219,0,0,0,248,0,18,0,177,0,6,0,0,0,0,0,0,0,0,0,194,0,134,0,233,0,173,0,124,0,0,0,0,0,190,0,13,0,117,0,10,0,237,0,95,0,2,0);
signal scenario_full  : scenario_type := (55,31,38,31,57,31,243,31,243,30,243,29,96,31,23,31,23,30,101,31,68,31,42,31,18,31,38,31,158,31,164,31,250,31,24,31,27,31,109,31,55,31,55,30,55,29,219,31,21,31,171,31,131,31,207,31,39,31,139,31,139,30,143,31,70,31,70,30,156,31,195,31,240,31,3,31,186,31,237,31,80,31,241,31,8,31,187,31,187,30,140,31,190,31,215,31,121,31,223,31,223,30,181,31,121,31,149,31,210,31,200,31,50,31,245,31,245,30,162,31,138,31,138,30,181,31,223,31,30,31,187,31,121,31,66,31,140,31,178,31,165,31,102,31,1,31,216,31,44,31,221,31,221,30,38,31,38,30,150,31,17,31,175,31,59,31,193,31,249,31,249,31,71,31,71,30,115,31,115,30,51,31,124,31,191,31,167,31,172,31,28,31,97,31,97,30,97,29,97,28,62,31,62,30,62,31,235,31,126,31,126,30,223,31,222,31,204,31,223,31,14,31,67,31,191,31,191,30,64,31,134,31,203,31,128,31,82,31,118,31,30,31,198,31,210,31,208,31,105,31,213,31,180,31,17,31,205,31,31,31,222,31,67,31,8,31,47,31,119,31,167,31,124,31,107,31,243,31,243,30,4,31,232,31,164,31,43,31,61,31,177,31,137,31,137,30,33,31,1,31,1,30,24,31,206,31,193,31,204,31,66,31,144,31,144,30,28,31,72,31,163,31,3,31,193,31,12,31,120,31,181,31,137,31,144,31,63,31,167,31,232,31,159,31,214,31,170,31,14,31,122,31,87,31,140,31,155,31,53,31,138,31,79,31,9,31,104,31,87,31,141,31,40,31,100,31,126,31,142,31,147,31,94,31,64,31,64,30,198,31,174,31,81,31,194,31,102,31,25,31,172,31,190,31,190,30,190,29,190,28,190,27,170,31,170,30,172,31,172,30,67,31,180,31,240,31,108,31,95,31,95,30,254,31,213,31,213,30,247,31,92,31,176,31,129,31,129,30,231,31,89,31,89,30,128,31,251,31,160,31,160,30,130,31,218,31,154,31,245,31,245,30,155,31,238,31,238,30,32,31,180,31,58,31,132,31,115,31,176,31,138,31,138,30,138,29,221,31,100,31,207,31,101,31,69,31,78,31,78,30,251,31,113,31,244,31,78,31,178,31,16,31,141,31,105,31,160,31,47,31,38,31,238,31,34,31,4,31,208,31,208,30,180,31,194,31,169,31,217,31,40,31,40,30,38,31,231,31,215,31,196,31,196,30,20,31,132,31,132,30,132,29,13,31,162,31,117,31,157,31,39,31,90,31,186,31,141,31,231,31,37,31,216,31,240,31,64,31,147,31,147,30,150,31,150,30,205,31,10,31,45,31,162,31,115,31,115,31,246,31,241,31,202,31,97,31,254,31,85,31,170,31,170,30,42,31,146,31,234,31,70,31,62,31,96,31,187,31,199,31,208,31,122,31,122,30,40,31,203,31,247,31,26,31,26,30,94,31,157,31,209,31,28,31,28,30,47,31,5,31,136,31,214,31,186,31,186,30,140,31,130,31,159,31,203,31,70,31,185,31,119,31,242,31,4,31,4,30,229,31,232,31,206,31,207,31,207,30,174,31,39,31,13,31,128,31,16,31,211,31,147,31,134,31,18,31,233,31,116,31,116,30,14,31,160,31,160,30,160,29,193,31,88,31,81,31,174,31,174,30,174,29,45,31,45,30,165,31,149,31,232,31,117,31,20,31,69,31,35,31,167,31,168,31,58,31,212,31,79,31,79,30,15,31,15,30,116,31,214,31,186,31,36,31,115,31,213,31,50,31,10,31,233,31,233,30,233,29,2,31,246,31,92,31,168,31,118,31,58,31,33,31,228,31,204,31,134,31,62,31,71,31,71,30,63,31,197,31,149,31,129,31,51,31,210,31,203,31,203,30,203,29,45,31,254,31,207,31,207,30,7,31,114,31,114,30,145,31,145,30,120,31,3,31,206,31,108,31,124,31,124,30,124,29,124,28,140,31,140,30,197,31,197,30,181,31,154,31,201,31,201,30,185,31,153,31,103,31,103,30,36,31,241,31,193,31,225,31,144,31,194,31,194,30,41,31,232,31,154,31,33,31,11,31,70,31,110,31,99,31,67,31,220,31,112,31,108,31,108,30,169,31,178,31,178,30,53,31,44,31,237,31,137,31,87,31,98,31,251,31,251,30,232,31,195,31,195,30,174,31,27,31,27,30,100,31,43,31,33,31,152,31,122,31,6,31,153,31,6,31,65,31,92,31,132,31,91,31,155,31,58,31,136,31,43,31,85,31,73,31,73,30,176,31,14,31,19,31,83,31,236,31,236,30,62,31,160,31,22,31,92,31,226,31,226,30,15,31,141,31,141,30,55,31,170,31,170,30,233,31,180,31,215,31,215,30,231,31,130,31,32,31,80,31,188,31,188,30,31,31,192,31,192,30,254,31,17,31,17,30,89,31,50,31,129,31,154,31,118,31,118,30,149,31,155,31,33,31,27,31,33,31,210,31,179,31,109,31,202,31,47,31,117,31,117,30,117,29,117,28,219,31,204,31,204,30,11,31,122,31,122,30,122,29,109,31,188,31,138,31,175,31,135,31,67,31,195,31,8,31,8,30,147,31,254,31,217,31,130,31,153,31,68,31,250,31,184,31,115,31,242,31,203,31,221,31,213,31,245,31,101,31,212,31,41,31,111,31,111,30,111,29,36,31,75,31,162,31,163,31,203,31,86,31,92,31,92,30,9,31,9,30,9,29,57,31,213,31,213,30,73,31,73,30,41,31,235,31,239,31,14,31,15,31,241,31,135,31,135,30,247,31,252,31,168,31,54,31,153,31,153,30,240,31,2,31,2,30,2,29,218,31,7,31,7,30,76,31,5,31,5,30,65,31,177,31,177,30,53,31,223,31,223,30,223,29,127,31,127,30,49,31,19,31,209,31,237,31,232,31,232,30,200,31,200,30,200,29,161,31,161,30,182,31,182,30,62,31,111,31,221,31,17,31,35,31,212,31,212,30,212,29,241,31,70,31,250,31,126,31,60,31,138,31,52,31,220,31,220,30,118,31,118,30,83,31,115,31,149,31,138,31,220,31,197,31,5,31,84,31,189,31,189,30,103,31,218,31,232,31,223,31,34,31,149,31,182,31,133,31,30,31,199,31,185,31,185,30,30,31,131,31,90,31,82,31,247,31,76,31,42,31,42,30,150,31,174,31,211,31,115,31,202,31,125,31,200,31,200,30,200,29,143,31,64,31,109,31,233,31,233,30,136,31,208,31,251,31,1,31,158,31,56,31,236,31,121,31,121,30,94,31,140,31,78,31,100,31,198,31,26,31,239,31,222,31,152,31,170,31,155,31,210,31,228,31,249,31,187,31,145,31,26,31,178,31,255,31,30,31,180,31,180,30,130,31,173,31,222,31,50,31,203,31,112,31,63,31,63,30,236,31,236,30,131,31,100,31,100,30,208,31,208,30,208,29,236,31,75,31,75,30,219,31,74,31,173,31,173,30,246,31,4,31,39,31,161,31,20,31,20,30,234,31,122,31,193,31,193,30,193,29,176,31,78,31,180,31,92,31,51,31,51,30,51,29,36,31,122,31,90,31,77,31,20,31,169,31,169,30,44,31,44,30,44,29,44,28,167,31,188,31,188,30,246,31,246,30,205,31,64,31,179,31,179,30,198,31,222,31,199,31,251,31,123,31,171,31,194,31,61,31,36,31,244,31,239,31,209,31,244,31,60,31,225,31,167,31,229,31,229,30,246,31,123,31,42,31,63,31,139,31,95,31,42,31,97,31,78,31,219,31,219,30,248,31,18,31,177,31,6,31,6,30,6,29,6,28,6,27,194,31,134,31,233,31,173,31,124,31,124,30,124,29,190,31,13,31,117,31,10,31,237,31,95,31,2,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
