-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_398 is
end project_tb_398;

architecture project_tb_arch_398 of project_tb_398 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 685;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,64,0,247,0,182,0,183,0,199,0,205,0,39,0,46,0,201,0,171,0,0,0,17,0,49,0,85,0,156,0,96,0,131,0,191,0,241,0,126,0,0,0,142,0,0,0,0,0,248,0,254,0,212,0,189,0,130,0,189,0,180,0,104,0,45,0,0,0,226,0,246,0,8,0,168,0,196,0,208,0,133,0,0,0,44,0,98,0,39,0,0,0,196,0,0,0,147,0,191,0,48,0,64,0,246,0,62,0,0,0,0,0,214,0,82,0,221,0,75,0,0,0,242,0,158,0,118,0,171,0,192,0,159,0,201,0,35,0,0,0,0,0,105,0,99,0,253,0,160,0,72,0,41,0,219,0,126,0,11,0,121,0,118,0,0,0,168,0,174,0,43,0,0,0,66,0,36,0,0,0,34,0,112,0,159,0,22,0,0,0,31,0,81,0,88,0,176,0,123,0,188,0,185,0,227,0,103,0,100,0,238,0,94,0,131,0,0,0,73,0,23,0,83,0,115,0,163,0,212,0,0,0,213,0,0,0,113,0,81,0,0,0,0,0,13,0,233,0,180,0,152,0,0,0,159,0,61,0,250,0,0,0,88,0,165,0,62,0,227,0,162,0,0,0,177,0,13,0,175,0,165,0,21,0,0,0,243,0,0,0,216,0,191,0,22,0,164,0,171,0,15,0,0,0,0,0,134,0,223,0,0,0,0,0,80,0,0,0,76,0,0,0,122,0,137,0,209,0,103,0,171,0,113,0,155,0,0,0,76,0,184,0,29,0,216,0,0,0,0,0,34,0,87,0,223,0,0,0,0,0,147,0,236,0,124,0,18,0,31,0,170,0,222,0,0,0,37,0,151,0,31,0,43,0,233,0,120,0,0,0,159,0,172,0,0,0,151,0,78,0,29,0,178,0,135,0,145,0,229,0,219,0,233,0,180,0,0,0,236,0,0,0,16,0,21,0,133,0,49,0,0,0,87,0,58,0,230,0,99,0,0,0,52,0,80,0,248,0,98,0,133,0,74,0,0,0,0,0,232,0,58,0,251,0,0,0,241,0,119,0,0,0,47,0,0,0,19,0,43,0,81,0,39,0,21,0,231,0,120,0,81,0,190,0,47,0,213,0,59,0,128,0,195,0,254,0,169,0,57,0,238,0,36,0,0,0,193,0,246,0,27,0,0,0,227,0,171,0,18,0,111,0,142,0,138,0,251,0,103,0,0,0,113,0,0,0,73,0,96,0,55,0,0,0,97,0,41,0,228,0,0,0,0,0,17,0,255,0,106,0,48,0,228,0,99,0,0,0,213,0,169,0,108,0,254,0,183,0,95,0,80,0,25,0,0,0,77,0,135,0,236,0,0,0,0,0,0,0,75,0,0,0,113,0,122,0,0,0,79,0,0,0,0,0,174,0,45,0,169,0,104,0,142,0,167,0,11,0,63,0,253,0,75,0,89,0,45,0,153,0,97,0,14,0,145,0,248,0,115,0,52,0,10,0,151,0,116,0,112,0,251,0,152,0,159,0,0,0,17,0,0,0,211,0,141,0,148,0,0,0,191,0,119,0,9,0,253,0,21,0,1,0,62,0,131,0,248,0,172,0,6,0,0,0,0,0,217,0,0,0,131,0,76,0,104,0,61,0,148,0,0,0,0,0,64,0,0,0,0,0,202,0,118,0,37,0,94,0,55,0,204,0,201,0,0,0,47,0,254,0,205,0,130,0,109,0,0,0,118,0,121,0,124,0,127,0,0,0,249,0,0,0,0,0,37,0,200,0,0,0,9,0,0,0,227,0,197,0,125,0,180,0,0,0,93,0,145,0,56,0,0,0,102,0,0,0,88,0,8,0,142,0,128,0,143,0,239,0,39,0,55,0,0,0,140,0,119,0,165,0,0,0,160,0,246,0,95,0,0,0,134,0,0,0,91,0,41,0,201,0,129,0,227,0,0,0,254,0,82,0,82,0,98,0,0,0,0,0,103,0,46,0,22,0,176,0,145,0,152,0,0,0,159,0,64,0,6,0,195,0,112,0,0,0,157,0,0,0,0,0,29,0,228,0,85,0,83,0,17,0,0,0,108,0,96,0,56,0,199,0,0,0,255,0,176,0,188,0,83,0,153,0,0,0,0,0,244,0,105,0,192,0,123,0,11,0,132,0,238,0,53,0,181,0,162,0,250,0,37,0,136,0,141,0,176,0,213,0,188,0,33,0,0,0,216,0,0,0,111,0,125,0,34,0,0,0,137,0,209,0,74,0,176,0,252,0,52,0,177,0,30,0,103,0,189,0,180,0,5,0,0,0,179,0,174,0,63,0,232,0,216,0,50,0,111,0,0,0,70,0,0,0,245,0,108,0,0,0,0,0,165,0,0,0,0,0,0,0,229,0,216,0,27,0,0,0,162,0,217,0,212,0,173,0,91,0,239,0,178,0,230,0,121,0,182,0,0,0,173,0,47,0,46,0,0,0,181,0,243,0,220,0,204,0,243,0,106,0,156,0,114,0,156,0,133,0,0,0,189,0,0,0,171,0,216,0,72,0,0,0,0,0,74,0,72,0,104,0,16,0,149,0,242,0,96,0,43,0,60,0,228,0,251,0,201,0,0,0,0,0,34,0,0,0,0,0,151,0,0,0,0,0,69,0,0,0,221,0,255,0,206,0,222,0,209,0,75,0,163,0,200,0,167,0,171,0,182,0,80,0,8,0,0,0,0,0,30,0,0,0,168,0,180,0,253,0,90,0,0,0,10,0,246,0,0,0,6,0,231,0,62,0,166,0,223,0,37,0,213,0,58,0,0,0,31,0,12,0,0,0,252,0,112,0,0,0,60,0,0,0,64,0,142,0,102,0,38,0,0,0,15,0,71,0,0,0,193,0,0,0,80,0,0,0,120,0,52,0,45,0,88,0,0,0,95,0,31,0,10,0,0,0,197,0,47,0,0,0,170,0,168,0,0,0,25,0,114,0,0,0,6,0,138,0,200,0,190,0,225,0,168,0,0,0,84,0,185,0,0,0,59,0,199,0,190,0,83,0,36,0,38,0,87,0,116,0,16,0,175,0,0,0,28,0,20,0,164,0);
signal scenario_full  : scenario_type := (34,31,64,31,247,31,182,31,183,31,199,31,205,31,39,31,46,31,201,31,171,31,171,30,17,31,49,31,85,31,156,31,96,31,131,31,191,31,241,31,126,31,126,30,142,31,142,30,142,29,248,31,254,31,212,31,189,31,130,31,189,31,180,31,104,31,45,31,45,30,226,31,246,31,8,31,168,31,196,31,208,31,133,31,133,30,44,31,98,31,39,31,39,30,196,31,196,30,147,31,191,31,48,31,64,31,246,31,62,31,62,30,62,29,214,31,82,31,221,31,75,31,75,30,242,31,158,31,118,31,171,31,192,31,159,31,201,31,35,31,35,30,35,29,105,31,99,31,253,31,160,31,72,31,41,31,219,31,126,31,11,31,121,31,118,31,118,30,168,31,174,31,43,31,43,30,66,31,36,31,36,30,34,31,112,31,159,31,22,31,22,30,31,31,81,31,88,31,176,31,123,31,188,31,185,31,227,31,103,31,100,31,238,31,94,31,131,31,131,30,73,31,23,31,83,31,115,31,163,31,212,31,212,30,213,31,213,30,113,31,81,31,81,30,81,29,13,31,233,31,180,31,152,31,152,30,159,31,61,31,250,31,250,30,88,31,165,31,62,31,227,31,162,31,162,30,177,31,13,31,175,31,165,31,21,31,21,30,243,31,243,30,216,31,191,31,22,31,164,31,171,31,15,31,15,30,15,29,134,31,223,31,223,30,223,29,80,31,80,30,76,31,76,30,122,31,137,31,209,31,103,31,171,31,113,31,155,31,155,30,76,31,184,31,29,31,216,31,216,30,216,29,34,31,87,31,223,31,223,30,223,29,147,31,236,31,124,31,18,31,31,31,170,31,222,31,222,30,37,31,151,31,31,31,43,31,233,31,120,31,120,30,159,31,172,31,172,30,151,31,78,31,29,31,178,31,135,31,145,31,229,31,219,31,233,31,180,31,180,30,236,31,236,30,16,31,21,31,133,31,49,31,49,30,87,31,58,31,230,31,99,31,99,30,52,31,80,31,248,31,98,31,133,31,74,31,74,30,74,29,232,31,58,31,251,31,251,30,241,31,119,31,119,30,47,31,47,30,19,31,43,31,81,31,39,31,21,31,231,31,120,31,81,31,190,31,47,31,213,31,59,31,128,31,195,31,254,31,169,31,57,31,238,31,36,31,36,30,193,31,246,31,27,31,27,30,227,31,171,31,18,31,111,31,142,31,138,31,251,31,103,31,103,30,113,31,113,30,73,31,96,31,55,31,55,30,97,31,41,31,228,31,228,30,228,29,17,31,255,31,106,31,48,31,228,31,99,31,99,30,213,31,169,31,108,31,254,31,183,31,95,31,80,31,25,31,25,30,77,31,135,31,236,31,236,30,236,29,236,28,75,31,75,30,113,31,122,31,122,30,79,31,79,30,79,29,174,31,45,31,169,31,104,31,142,31,167,31,11,31,63,31,253,31,75,31,89,31,45,31,153,31,97,31,14,31,145,31,248,31,115,31,52,31,10,31,151,31,116,31,112,31,251,31,152,31,159,31,159,30,17,31,17,30,211,31,141,31,148,31,148,30,191,31,119,31,9,31,253,31,21,31,1,31,62,31,131,31,248,31,172,31,6,31,6,30,6,29,217,31,217,30,131,31,76,31,104,31,61,31,148,31,148,30,148,29,64,31,64,30,64,29,202,31,118,31,37,31,94,31,55,31,204,31,201,31,201,30,47,31,254,31,205,31,130,31,109,31,109,30,118,31,121,31,124,31,127,31,127,30,249,31,249,30,249,29,37,31,200,31,200,30,9,31,9,30,227,31,197,31,125,31,180,31,180,30,93,31,145,31,56,31,56,30,102,31,102,30,88,31,8,31,142,31,128,31,143,31,239,31,39,31,55,31,55,30,140,31,119,31,165,31,165,30,160,31,246,31,95,31,95,30,134,31,134,30,91,31,41,31,201,31,129,31,227,31,227,30,254,31,82,31,82,31,98,31,98,30,98,29,103,31,46,31,22,31,176,31,145,31,152,31,152,30,159,31,64,31,6,31,195,31,112,31,112,30,157,31,157,30,157,29,29,31,228,31,85,31,83,31,17,31,17,30,108,31,96,31,56,31,199,31,199,30,255,31,176,31,188,31,83,31,153,31,153,30,153,29,244,31,105,31,192,31,123,31,11,31,132,31,238,31,53,31,181,31,162,31,250,31,37,31,136,31,141,31,176,31,213,31,188,31,33,31,33,30,216,31,216,30,111,31,125,31,34,31,34,30,137,31,209,31,74,31,176,31,252,31,52,31,177,31,30,31,103,31,189,31,180,31,5,31,5,30,179,31,174,31,63,31,232,31,216,31,50,31,111,31,111,30,70,31,70,30,245,31,108,31,108,30,108,29,165,31,165,30,165,29,165,28,229,31,216,31,27,31,27,30,162,31,217,31,212,31,173,31,91,31,239,31,178,31,230,31,121,31,182,31,182,30,173,31,47,31,46,31,46,30,181,31,243,31,220,31,204,31,243,31,106,31,156,31,114,31,156,31,133,31,133,30,189,31,189,30,171,31,216,31,72,31,72,30,72,29,74,31,72,31,104,31,16,31,149,31,242,31,96,31,43,31,60,31,228,31,251,31,201,31,201,30,201,29,34,31,34,30,34,29,151,31,151,30,151,29,69,31,69,30,221,31,255,31,206,31,222,31,209,31,75,31,163,31,200,31,167,31,171,31,182,31,80,31,8,31,8,30,8,29,30,31,30,30,168,31,180,31,253,31,90,31,90,30,10,31,246,31,246,30,6,31,231,31,62,31,166,31,223,31,37,31,213,31,58,31,58,30,31,31,12,31,12,30,252,31,112,31,112,30,60,31,60,30,64,31,142,31,102,31,38,31,38,30,15,31,71,31,71,30,193,31,193,30,80,31,80,30,120,31,52,31,45,31,88,31,88,30,95,31,31,31,10,31,10,30,197,31,47,31,47,30,170,31,168,31,168,30,25,31,114,31,114,30,6,31,138,31,200,31,190,31,225,31,168,31,168,30,84,31,185,31,185,30,59,31,199,31,190,31,83,31,36,31,38,31,87,31,116,31,16,31,175,31,175,30,28,31,20,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
