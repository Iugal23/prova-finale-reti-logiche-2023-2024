-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 599;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (178,0,189,0,0,0,45,0,224,0,0,0,2,0,42,0,181,0,224,0,156,0,22,0,42,0,161,0,0,0,87,0,207,0,85,0,255,0,17,0,109,0,129,0,79,0,0,0,34,0,51,0,0,0,0,0,0,0,0,0,83,0,13,0,68,0,36,0,193,0,0,0,0,0,0,0,78,0,178,0,77,0,26,0,136,0,0,0,108,0,37,0,0,0,59,0,181,0,0,0,72,0,148,0,0,0,125,0,36,0,129,0,85,0,101,0,24,0,21,0,197,0,188,0,174,0,248,0,0,0,84,0,0,0,47,0,73,0,190,0,185,0,219,0,114,0,60,0,152,0,0,0,0,0,162,0,224,0,67,0,107,0,2,0,39,0,62,0,49,0,0,0,183,0,65,0,159,0,138,0,71,0,0,0,0,0,103,0,166,0,47,0,19,0,97,0,223,0,65,0,56,0,83,0,25,0,94,0,117,0,218,0,30,0,21,0,0,0,0,0,0,0,75,0,74,0,60,0,0,0,120,0,0,0,0,0,159,0,0,0,200,0,108,0,190,0,219,0,198,0,122,0,30,0,69,0,28,0,63,0,55,0,179,0,0,0,4,0,155,0,36,0,249,0,127,0,123,0,96,0,123,0,254,0,176,0,237,0,168,0,83,0,0,0,192,0,42,0,67,0,222,0,0,0,123,0,127,0,30,0,153,0,35,0,237,0,0,0,43,0,119,0,84,0,122,0,182,0,0,0,0,0,0,0,138,0,172,0,106,0,78,0,166,0,45,0,0,0,0,0,160,0,119,0,0,0,103,0,249,0,37,0,78,0,33,0,49,0,0,0,40,0,165,0,0,0,3,0,0,0,8,0,80,0,166,0,12,0,28,0,0,0,64,0,223,0,124,0,242,0,133,0,249,0,248,0,180,0,0,0,20,0,0,0,199,0,86,0,253,0,126,0,112,0,163,0,126,0,17,0,145,0,222,0,55,0,13,0,223,0,182,0,115,0,0,0,0,0,133,0,249,0,197,0,194,0,117,0,62,0,0,0,195,0,114,0,5,0,0,0,0,0,5,0,0,0,71,0,169,0,0,0,237,0,0,0,187,0,157,0,10,0,180,0,123,0,247,0,161,0,65,0,0,0,2,0,41,0,68,0,16,0,92,0,86,0,0,0,243,0,74,0,159,0,62,0,238,0,79,0,0,0,50,0,0,0,140,0,0,0,245,0,193,0,237,0,139,0,154,0,0,0,0,0,206,0,239,0,252,0,33,0,0,0,216,0,58,0,31,0,95,0,114,0,73,0,0,0,0,0,188,0,77,0,27,0,156,0,86,0,175,0,204,0,77,0,0,0,72,0,0,0,168,0,230,0,155,0,2,0,216,0,234,0,130,0,10,0,1,0,174,0,0,0,0,0,78,0,25,0,195,0,74,0,70,0,243,0,11,0,231,0,35,0,2,0,195,0,226,0,0,0,0,0,202,0,0,0,0,0,188,0,4,0,72,0,129,0,136,0,61,0,80,0,42,0,71,0,125,0,232,0,162,0,205,0,180,0,233,0,250,0,0,0,219,0,171,0,167,0,30,0,146,0,18,0,0,0,0,0,0,0,112,0,142,0,61,0,0,0,195,0,195,0,96,0,0,0,230,0,185,0,26,0,81,0,243,0,156,0,215,0,188,0,62,0,255,0,223,0,36,0,205,0,206,0,84,0,87,0,0,0,207,0,207,0,7,0,62,0,0,0,180,0,109,0,136,0,0,0,67,0,115,0,11,0,206,0,0,0,125,0,8,0,145,0,107,0,42,0,247,0,23,0,225,0,178,0,91,0,76,0,56,0,196,0,189,0,134,0,154,0,0,0,234,0,0,0,14,0,62,0,54,0,0,0,84,0,55,0,106,0,197,0,116,0,56,0,28,0,130,0,0,0,118,0,0,0,226,0,73,0,239,0,235,0,0,0,233,0,199,0,0,0,20,0,169,0,47,0,0,0,49,0,0,0,33,0,30,0,41,0,179,0,46,0,54,0,1,0,24,0,0,0,211,0,244,0,139,0,215,0,26,0,168,0,20,0,130,0,0,0,155,0,0,0,145,0,149,0,240,0,0,0,79,0,0,0,226,0,0,0,240,0,0,0,105,0,191,0,111,0,0,0,0,0,82,0,116,0,8,0,27,0,123,0,192,0,84,0,216,0,190,0,235,0,0,0,0,0,0,0,30,0,94,0,157,0,13,0,204,0,246,0,234,0,0,0,153,0,149,0,145,0,0,0,51,0,137,0,56,0,195,0,132,0,228,0,90,0,253,0,101,0,36,0,217,0,67,0,224,0,8,0,0,0,0,0,233,0,211,0,0,0,0,0,149,0,160,0,83,0,193,0,207,0,63,0,139,0,3,0,244,0,47,0,53,0,0,0,241,0,201,0,0,0,200,0,162,0,203,0,156,0,156,0,151,0,218,0,222,0,18,0,138,0,113,0,17,0,0,0,0,0,80,0,147,0,63,0,194,0,0,0,205,0,193,0,249,0,175,0,12,0,48,0,195,0,83,0,42,0,89,0,90,0,0,0,186,0,161,0,58,0,183,0,87,0,218,0,19,0,89,0,27,0,153,0,130,0,236,0,31,0,0,0,22,0,0,0,0,0,27,0,251,0,254,0,0,0,231,0,118,0,103,0,0,0,0,0,0,0,45,0,70,0,0,0);
signal scenario_full  : scenario_type := (178,31,189,31,189,30,45,31,224,31,224,30,2,31,42,31,181,31,224,31,156,31,22,31,42,31,161,31,161,30,87,31,207,31,85,31,255,31,17,31,109,31,129,31,79,31,79,30,34,31,51,31,51,30,51,29,51,28,51,27,83,31,13,31,68,31,36,31,193,31,193,30,193,29,193,28,78,31,178,31,77,31,26,31,136,31,136,30,108,31,37,31,37,30,59,31,181,31,181,30,72,31,148,31,148,30,125,31,36,31,129,31,85,31,101,31,24,31,21,31,197,31,188,31,174,31,248,31,248,30,84,31,84,30,47,31,73,31,190,31,185,31,219,31,114,31,60,31,152,31,152,30,152,29,162,31,224,31,67,31,107,31,2,31,39,31,62,31,49,31,49,30,183,31,65,31,159,31,138,31,71,31,71,30,71,29,103,31,166,31,47,31,19,31,97,31,223,31,65,31,56,31,83,31,25,31,94,31,117,31,218,31,30,31,21,31,21,30,21,29,21,28,75,31,74,31,60,31,60,30,120,31,120,30,120,29,159,31,159,30,200,31,108,31,190,31,219,31,198,31,122,31,30,31,69,31,28,31,63,31,55,31,179,31,179,30,4,31,155,31,36,31,249,31,127,31,123,31,96,31,123,31,254,31,176,31,237,31,168,31,83,31,83,30,192,31,42,31,67,31,222,31,222,30,123,31,127,31,30,31,153,31,35,31,237,31,237,30,43,31,119,31,84,31,122,31,182,31,182,30,182,29,182,28,138,31,172,31,106,31,78,31,166,31,45,31,45,30,45,29,160,31,119,31,119,30,103,31,249,31,37,31,78,31,33,31,49,31,49,30,40,31,165,31,165,30,3,31,3,30,8,31,80,31,166,31,12,31,28,31,28,30,64,31,223,31,124,31,242,31,133,31,249,31,248,31,180,31,180,30,20,31,20,30,199,31,86,31,253,31,126,31,112,31,163,31,126,31,17,31,145,31,222,31,55,31,13,31,223,31,182,31,115,31,115,30,115,29,133,31,249,31,197,31,194,31,117,31,62,31,62,30,195,31,114,31,5,31,5,30,5,29,5,31,5,30,71,31,169,31,169,30,237,31,237,30,187,31,157,31,10,31,180,31,123,31,247,31,161,31,65,31,65,30,2,31,41,31,68,31,16,31,92,31,86,31,86,30,243,31,74,31,159,31,62,31,238,31,79,31,79,30,50,31,50,30,140,31,140,30,245,31,193,31,237,31,139,31,154,31,154,30,154,29,206,31,239,31,252,31,33,31,33,30,216,31,58,31,31,31,95,31,114,31,73,31,73,30,73,29,188,31,77,31,27,31,156,31,86,31,175,31,204,31,77,31,77,30,72,31,72,30,168,31,230,31,155,31,2,31,216,31,234,31,130,31,10,31,1,31,174,31,174,30,174,29,78,31,25,31,195,31,74,31,70,31,243,31,11,31,231,31,35,31,2,31,195,31,226,31,226,30,226,29,202,31,202,30,202,29,188,31,4,31,72,31,129,31,136,31,61,31,80,31,42,31,71,31,125,31,232,31,162,31,205,31,180,31,233,31,250,31,250,30,219,31,171,31,167,31,30,31,146,31,18,31,18,30,18,29,18,28,112,31,142,31,61,31,61,30,195,31,195,31,96,31,96,30,230,31,185,31,26,31,81,31,243,31,156,31,215,31,188,31,62,31,255,31,223,31,36,31,205,31,206,31,84,31,87,31,87,30,207,31,207,31,7,31,62,31,62,30,180,31,109,31,136,31,136,30,67,31,115,31,11,31,206,31,206,30,125,31,8,31,145,31,107,31,42,31,247,31,23,31,225,31,178,31,91,31,76,31,56,31,196,31,189,31,134,31,154,31,154,30,234,31,234,30,14,31,62,31,54,31,54,30,84,31,55,31,106,31,197,31,116,31,56,31,28,31,130,31,130,30,118,31,118,30,226,31,73,31,239,31,235,31,235,30,233,31,199,31,199,30,20,31,169,31,47,31,47,30,49,31,49,30,33,31,30,31,41,31,179,31,46,31,54,31,1,31,24,31,24,30,211,31,244,31,139,31,215,31,26,31,168,31,20,31,130,31,130,30,155,31,155,30,145,31,149,31,240,31,240,30,79,31,79,30,226,31,226,30,240,31,240,30,105,31,191,31,111,31,111,30,111,29,82,31,116,31,8,31,27,31,123,31,192,31,84,31,216,31,190,31,235,31,235,30,235,29,235,28,30,31,94,31,157,31,13,31,204,31,246,31,234,31,234,30,153,31,149,31,145,31,145,30,51,31,137,31,56,31,195,31,132,31,228,31,90,31,253,31,101,31,36,31,217,31,67,31,224,31,8,31,8,30,8,29,233,31,211,31,211,30,211,29,149,31,160,31,83,31,193,31,207,31,63,31,139,31,3,31,244,31,47,31,53,31,53,30,241,31,201,31,201,30,200,31,162,31,203,31,156,31,156,31,151,31,218,31,222,31,18,31,138,31,113,31,17,31,17,30,17,29,80,31,147,31,63,31,194,31,194,30,205,31,193,31,249,31,175,31,12,31,48,31,195,31,83,31,42,31,89,31,90,31,90,30,186,31,161,31,58,31,183,31,87,31,218,31,19,31,89,31,27,31,153,31,130,31,236,31,31,31,31,30,22,31,22,30,22,29,27,31,251,31,254,31,254,30,231,31,118,31,103,31,103,30,103,29,103,28,45,31,70,31,70,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
