-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_528 is
end project_tb_528;

architecture project_tb_arch_528 of project_tb_528 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 828;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (167,0,172,0,127,0,158,0,0,0,201,0,0,0,176,0,32,0,146,0,130,0,189,0,177,0,118,0,39,0,28,0,71,0,111,0,70,0,122,0,162,0,46,0,0,0,17,0,52,0,162,0,77,0,120,0,139,0,48,0,151,0,42,0,184,0,165,0,95,0,149,0,14,0,56,0,105,0,139,0,0,0,27,0,0,0,0,0,186,0,224,0,20,0,23,0,61,0,0,0,120,0,197,0,0,0,247,0,224,0,84,0,0,0,212,0,0,0,210,0,0,0,137,0,0,0,55,0,102,0,197,0,0,0,117,0,251,0,71,0,182,0,20,0,250,0,64,0,76,0,0,0,219,0,159,0,0,0,4,0,16,0,134,0,237,0,0,0,197,0,120,0,82,0,130,0,162,0,215,0,70,0,19,0,194,0,40,0,110,0,104,0,0,0,155,0,250,0,65,0,151,0,0,0,214,0,43,0,180,0,153,0,0,0,212,0,211,0,220,0,152,0,1,0,63,0,255,0,147,0,0,0,147,0,115,0,221,0,87,0,0,0,0,0,120,0,93,0,179,0,110,0,18,0,140,0,151,0,212,0,0,0,49,0,0,0,211,0,190,0,45,0,88,0,69,0,13,0,130,0,150,0,47,0,0,0,37,0,178,0,92,0,186,0,0,0,47,0,254,0,143,0,121,0,206,0,217,0,206,0,230,0,27,0,28,0,82,0,178,0,31,0,0,0,243,0,0,0,248,0,139,0,0,0,208,0,0,0,0,0,32,0,32,0,108,0,56,0,164,0,89,0,72,0,52,0,129,0,195,0,248,0,0,0,0,0,25,0,199,0,151,0,151,0,83,0,61,0,147,0,229,0,141,0,22,0,0,0,182,0,184,0,14,0,124,0,57,0,87,0,227,0,92,0,87,0,180,0,146,0,0,0,30,0,0,0,0,0,36,0,143,0,20,0,228,0,20,0,0,0,56,0,164,0,186,0,198,0,181,0,0,0,0,0,130,0,94,0,0,0,217,0,0,0,0,0,102,0,91,0,244,0,90,0,0,0,0,0,23,0,112,0,83,0,14,0,0,0,234,0,121,0,186,0,185,0,145,0,230,0,142,0,235,0,7,0,0,0,106,0,192,0,0,0,245,0,97,0,58,0,171,0,182,0,0,0,0,0,236,0,138,0,81,0,61,0,118,0,213,0,0,0,219,0,0,0,33,0,29,0,125,0,221,0,251,0,74,0,10,0,111,0,28,0,0,0,123,0,1,0,121,0,232,0,38,0,246,0,0,0,90,0,0,0,0,0,124,0,202,0,33,0,166,0,46,0,76,0,169,0,235,0,105,0,255,0,123,0,1,0,74,0,140,0,102,0,0,0,185,0,0,0,247,0,69,0,0,0,12,0,0,0,212,0,10,0,0,0,251,0,27,0,0,0,196,0,33,0,0,0,0,0,2,0,15,0,86,0,71,0,133,0,152,0,131,0,167,0,222,0,182,0,123,0,249,0,57,0,0,0,161,0,0,0,97,0,143,0,21,0,170,0,250,0,126,0,105,0,19,0,213,0,68,0,0,0,140,0,32,0,28,0,148,0,229,0,118,0,175,0,0,0,145,0,249,0,0,0,83,0,64,0,205,0,110,0,169,0,162,0,0,0,201,0,49,0,94,0,57,0,218,0,249,0,250,0,169,0,67,0,0,0,1,0,73,0,99,0,137,0,67,0,240,0,95,0,32,0,34,0,134,0,48,0,19,0,0,0,49,0,0,0,123,0,217,0,153,0,31,0,120,0,227,0,116,0,108,0,152,0,253,0,0,0,190,0,14,0,8,0,35,0,88,0,62,0,167,0,142,0,129,0,142,0,181,0,76,0,252,0,120,0,0,0,63,0,0,0,53,0,100,0,230,0,0,0,112,0,246,0,0,0,15,0,177,0,163,0,143,0,0,0,157,0,0,0,0,0,0,0,64,0,251,0,220,0,255,0,3,0,180,0,158,0,116,0,230,0,18,0,84,0,2,0,64,0,0,0,0,0,0,0,17,0,217,0,2,0,192,0,3,0,218,0,250,0,52,0,0,0,73,0,19,0,109,0,0,0,207,0,0,0,74,0,105,0,207,0,94,0,33,0,51,0,137,0,159,0,105,0,187,0,0,0,156,0,209,0,223,0,0,0,62,0,0,0,184,0,217,0,19,0,0,0,148,0,106,0,52,0,5,0,173,0,27,0,30,0,0,0,202,0,29,0,119,0,19,0,15,0,36,0,57,0,146,0,153,0,46,0,163,0,55,0,32,0,233,0,78,0,170,0,94,0,177,0,20,0,188,0,245,0,184,0,0,0,0,0,23,0,143,0,142,0,54,0,158,0,8,0,136,0,152,0,0,0,51,0,199,0,0,0,249,0,116,0,219,0,69,0,0,0,102,0,27,0,58,0,14,0,142,0,182,0,240,0,215,0,0,0,0,0,168,0,0,0,229,0,0,0,214,0,121,0,233,0,6,0,169,0,142,0,85,0,172,0,74,0,90,0,0,0,111,0,0,0,154,0,83,0,13,0,252,0,248,0,227,0,127,0,188,0,0,0,94,0,246,0,92,0,58,0,106,0,0,0,219,0,61,0,202,0,9,0,181,0,235,0,136,0,248,0,115,0,133,0,21,0,62,0,69,0,51,0,0,0,172,0,23,0,103,0,56,0,67,0,13,0,0,0,0,0,141,0,212,0,225,0,70,0,168,0,73,0,86,0,126,0,105,0,0,0,103,0,117,0,123,0,203,0,4,0,216,0,132,0,227,0,195,0,0,0,0,0,141,0,14,0,55,0,167,0,0,0,206,0,161,0,112,0,22,0,177,0,170,0,255,0,14,0,236,0,4,0,182,0,232,0,98,0,0,0,0,0,187,0,0,0,0,0,122,0,134,0,165,0,244,0,54,0,0,0,91,0,209,0,0,0,29,0,201,0,0,0,111,0,234,0,106,0,51,0,84,0,51,0,59,0,0,0,215,0,231,0,0,0,122,0,48,0,214,0,111,0,20,0,122,0,75,0,96,0,237,0,145,0,80,0,210,0,150,0,69,0,8,0,162,0,144,0,212,0,247,0,0,0,0,0,0,0,0,0,234,0,49,0,232,0,83,0,54,0,124,0,16,0,0,0,184,0,196,0,191,0,218,0,0,0,0,0,228,0,193,0,59,0,45,0,0,0,152,0,38,0,34,0,31,0,125,0,0,0,0,0,88,0,45,0,164,0,251,0,0,0,123,0,26,0,50,0,27,0,92,0,144,0,93,0,89,0,242,0,231,0,69,0,0,0,0,0,241,0,223,0,89,0,213,0,103,0,0,0,163,0,132,0,11,0,0,0,247,0,237,0,5,0,0,0,135,0,63,0,22,0,4,0,116,0,189,0,234,0,0,0,227,0,100,0,0,0,21,0,0,0,0,0,0,0,140,0,8,0,216,0,101,0,40,0,18,0,0,0,181,0,27,0,64,0,19,0,158,0,14,0,183,0,0,0,209,0,66,0,242,0,188,0,130,0,118,0,58,0,0,0,0,0,163,0,195,0,146,0,11,0,57,0,77,0,0,0,219,0,0,0,157,0,220,0,41,0,0,0,105,0,0,0,123,0,67,0,241,0,180,0,76,0,156,0,161,0,129,0,91,0,0,0,9,0,185,0,111,0,0,0,0,0,39,0,223,0,110,0,0,0,34,0,208,0,128,0,188,0,0,0,211,0);
signal scenario_full  : scenario_type := (167,31,172,31,127,31,158,31,158,30,201,31,201,30,176,31,32,31,146,31,130,31,189,31,177,31,118,31,39,31,28,31,71,31,111,31,70,31,122,31,162,31,46,31,46,30,17,31,52,31,162,31,77,31,120,31,139,31,48,31,151,31,42,31,184,31,165,31,95,31,149,31,14,31,56,31,105,31,139,31,139,30,27,31,27,30,27,29,186,31,224,31,20,31,23,31,61,31,61,30,120,31,197,31,197,30,247,31,224,31,84,31,84,30,212,31,212,30,210,31,210,30,137,31,137,30,55,31,102,31,197,31,197,30,117,31,251,31,71,31,182,31,20,31,250,31,64,31,76,31,76,30,219,31,159,31,159,30,4,31,16,31,134,31,237,31,237,30,197,31,120,31,82,31,130,31,162,31,215,31,70,31,19,31,194,31,40,31,110,31,104,31,104,30,155,31,250,31,65,31,151,31,151,30,214,31,43,31,180,31,153,31,153,30,212,31,211,31,220,31,152,31,1,31,63,31,255,31,147,31,147,30,147,31,115,31,221,31,87,31,87,30,87,29,120,31,93,31,179,31,110,31,18,31,140,31,151,31,212,31,212,30,49,31,49,30,211,31,190,31,45,31,88,31,69,31,13,31,130,31,150,31,47,31,47,30,37,31,178,31,92,31,186,31,186,30,47,31,254,31,143,31,121,31,206,31,217,31,206,31,230,31,27,31,28,31,82,31,178,31,31,31,31,30,243,31,243,30,248,31,139,31,139,30,208,31,208,30,208,29,32,31,32,31,108,31,56,31,164,31,89,31,72,31,52,31,129,31,195,31,248,31,248,30,248,29,25,31,199,31,151,31,151,31,83,31,61,31,147,31,229,31,141,31,22,31,22,30,182,31,184,31,14,31,124,31,57,31,87,31,227,31,92,31,87,31,180,31,146,31,146,30,30,31,30,30,30,29,36,31,143,31,20,31,228,31,20,31,20,30,56,31,164,31,186,31,198,31,181,31,181,30,181,29,130,31,94,31,94,30,217,31,217,30,217,29,102,31,91,31,244,31,90,31,90,30,90,29,23,31,112,31,83,31,14,31,14,30,234,31,121,31,186,31,185,31,145,31,230,31,142,31,235,31,7,31,7,30,106,31,192,31,192,30,245,31,97,31,58,31,171,31,182,31,182,30,182,29,236,31,138,31,81,31,61,31,118,31,213,31,213,30,219,31,219,30,33,31,29,31,125,31,221,31,251,31,74,31,10,31,111,31,28,31,28,30,123,31,1,31,121,31,232,31,38,31,246,31,246,30,90,31,90,30,90,29,124,31,202,31,33,31,166,31,46,31,76,31,169,31,235,31,105,31,255,31,123,31,1,31,74,31,140,31,102,31,102,30,185,31,185,30,247,31,69,31,69,30,12,31,12,30,212,31,10,31,10,30,251,31,27,31,27,30,196,31,33,31,33,30,33,29,2,31,15,31,86,31,71,31,133,31,152,31,131,31,167,31,222,31,182,31,123,31,249,31,57,31,57,30,161,31,161,30,97,31,143,31,21,31,170,31,250,31,126,31,105,31,19,31,213,31,68,31,68,30,140,31,32,31,28,31,148,31,229,31,118,31,175,31,175,30,145,31,249,31,249,30,83,31,64,31,205,31,110,31,169,31,162,31,162,30,201,31,49,31,94,31,57,31,218,31,249,31,250,31,169,31,67,31,67,30,1,31,73,31,99,31,137,31,67,31,240,31,95,31,32,31,34,31,134,31,48,31,19,31,19,30,49,31,49,30,123,31,217,31,153,31,31,31,120,31,227,31,116,31,108,31,152,31,253,31,253,30,190,31,14,31,8,31,35,31,88,31,62,31,167,31,142,31,129,31,142,31,181,31,76,31,252,31,120,31,120,30,63,31,63,30,53,31,100,31,230,31,230,30,112,31,246,31,246,30,15,31,177,31,163,31,143,31,143,30,157,31,157,30,157,29,157,28,64,31,251,31,220,31,255,31,3,31,180,31,158,31,116,31,230,31,18,31,84,31,2,31,64,31,64,30,64,29,64,28,17,31,217,31,2,31,192,31,3,31,218,31,250,31,52,31,52,30,73,31,19,31,109,31,109,30,207,31,207,30,74,31,105,31,207,31,94,31,33,31,51,31,137,31,159,31,105,31,187,31,187,30,156,31,209,31,223,31,223,30,62,31,62,30,184,31,217,31,19,31,19,30,148,31,106,31,52,31,5,31,173,31,27,31,30,31,30,30,202,31,29,31,119,31,19,31,15,31,36,31,57,31,146,31,153,31,46,31,163,31,55,31,32,31,233,31,78,31,170,31,94,31,177,31,20,31,188,31,245,31,184,31,184,30,184,29,23,31,143,31,142,31,54,31,158,31,8,31,136,31,152,31,152,30,51,31,199,31,199,30,249,31,116,31,219,31,69,31,69,30,102,31,27,31,58,31,14,31,142,31,182,31,240,31,215,31,215,30,215,29,168,31,168,30,229,31,229,30,214,31,121,31,233,31,6,31,169,31,142,31,85,31,172,31,74,31,90,31,90,30,111,31,111,30,154,31,83,31,13,31,252,31,248,31,227,31,127,31,188,31,188,30,94,31,246,31,92,31,58,31,106,31,106,30,219,31,61,31,202,31,9,31,181,31,235,31,136,31,248,31,115,31,133,31,21,31,62,31,69,31,51,31,51,30,172,31,23,31,103,31,56,31,67,31,13,31,13,30,13,29,141,31,212,31,225,31,70,31,168,31,73,31,86,31,126,31,105,31,105,30,103,31,117,31,123,31,203,31,4,31,216,31,132,31,227,31,195,31,195,30,195,29,141,31,14,31,55,31,167,31,167,30,206,31,161,31,112,31,22,31,177,31,170,31,255,31,14,31,236,31,4,31,182,31,232,31,98,31,98,30,98,29,187,31,187,30,187,29,122,31,134,31,165,31,244,31,54,31,54,30,91,31,209,31,209,30,29,31,201,31,201,30,111,31,234,31,106,31,51,31,84,31,51,31,59,31,59,30,215,31,231,31,231,30,122,31,48,31,214,31,111,31,20,31,122,31,75,31,96,31,237,31,145,31,80,31,210,31,150,31,69,31,8,31,162,31,144,31,212,31,247,31,247,30,247,29,247,28,247,27,234,31,49,31,232,31,83,31,54,31,124,31,16,31,16,30,184,31,196,31,191,31,218,31,218,30,218,29,228,31,193,31,59,31,45,31,45,30,152,31,38,31,34,31,31,31,125,31,125,30,125,29,88,31,45,31,164,31,251,31,251,30,123,31,26,31,50,31,27,31,92,31,144,31,93,31,89,31,242,31,231,31,69,31,69,30,69,29,241,31,223,31,89,31,213,31,103,31,103,30,163,31,132,31,11,31,11,30,247,31,237,31,5,31,5,30,135,31,63,31,22,31,4,31,116,31,189,31,234,31,234,30,227,31,100,31,100,30,21,31,21,30,21,29,21,28,140,31,8,31,216,31,101,31,40,31,18,31,18,30,181,31,27,31,64,31,19,31,158,31,14,31,183,31,183,30,209,31,66,31,242,31,188,31,130,31,118,31,58,31,58,30,58,29,163,31,195,31,146,31,11,31,57,31,77,31,77,30,219,31,219,30,157,31,220,31,41,31,41,30,105,31,105,30,123,31,67,31,241,31,180,31,76,31,156,31,161,31,129,31,91,31,91,30,9,31,185,31,111,31,111,30,111,29,39,31,223,31,110,31,110,30,34,31,208,31,128,31,188,31,188,30,211,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
