-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 336;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (62,0,0,0,124,0,169,0,0,0,228,0,50,0,0,0,251,0,79,0,58,0,0,0,0,0,22,0,96,0,201,0,131,0,0,0,0,0,0,0,111,0,0,0,173,0,0,0,66,0,0,0,0,0,117,0,149,0,138,0,187,0,86,0,111,0,0,0,96,0,0,0,0,0,220,0,200,0,169,0,0,0,58,0,120,0,246,0,0,0,94,0,134,0,48,0,151,0,89,0,0,0,252,0,107,0,228,0,210,0,19,0,31,0,17,0,116,0,45,0,27,0,61,0,0,0,0,0,0,0,21,0,238,0,96,0,147,0,47,0,0,0,0,0,0,0,0,0,8,0,143,0,168,0,85,0,60,0,204,0,20,0,113,0,124,0,43,0,74,0,0,0,199,0,0,0,47,0,0,0,178,0,234,0,0,0,135,0,26,0,0,0,133,0,245,0,0,0,235,0,140,0,52,0,233,0,0,0,192,0,3,0,151,0,0,0,0,0,224,0,0,0,40,0,197,0,143,0,127,0,108,0,165,0,113,0,0,0,164,0,3,0,92,0,212,0,110,0,168,0,125,0,239,0,237,0,0,0,169,0,168,0,0,0,58,0,126,0,223,0,197,0,65,0,82,0,177,0,21,0,78,0,111,0,206,0,0,0,64,0,24,0,4,0,250,0,148,0,13,0,88,0,96,0,124,0,0,0,68,0,97,0,0,0,187,0,91,0,33,0,0,0,132,0,201,0,49,0,48,0,95,0,177,0,63,0,252,0,191,0,116,0,252,0,129,0,2,0,5,0,222,0,62,0,216,0,0,0,0,0,78,0,15,0,242,0,73,0,149,0,146,0,25,0,140,0,99,0,64,0,127,0,0,0,165,0,141,0,0,0,167,0,57,0,84,0,0,0,223,0,117,0,73,0,125,0,142,0,41,0,211,0,17,0,124,0,0,0,164,0,179,0,145,0,200,0,0,0,0,0,47,0,51,0,80,0,20,0,115,0,47,0,110,0,175,0,229,0,63,0,163,0,131,0,65,0,141,0,0,0,87,0,105,0,216,0,220,0,248,0,207,0,0,0,147,0,101,0,202,0,115,0,0,0,51,0,0,0,70,0,216,0,125,0,0,0,61,0,225,0,158,0,167,0,86,0,115,0,102,0,250,0,1,0,0,0,220,0,49,0,61,0,0,0,0,0,255,0,232,0,195,0,246,0,185,0,174,0,243,0,161,0,177,0,59,0,0,0,212,0,0,0,237,0,0,0,116,0,250,0,63,0,213,0,223,0,65,0,198,0,38,0,139,0,52,0,246,0,0,0,215,0,41,0,189,0,0,0,0,0,36,0,87,0,125,0,239,0,47,0,187,0,0,0,187,0,0,0,25,0,26,0,253,0,78,0,123,0,0,0,255,0,45,0,139,0,3,0,96,0,79,0,190,0,222,0,235,0,28,0,115,0,45,0,161,0,167,0,10,0,99,0,239,0,0,0,119,0,106,0,186,0,23,0,235,0,13,0,58,0,180,0);
signal scenario_full  : scenario_type := (62,31,62,30,124,31,169,31,169,30,228,31,50,31,50,30,251,31,79,31,58,31,58,30,58,29,22,31,96,31,201,31,131,31,131,30,131,29,131,28,111,31,111,30,173,31,173,30,66,31,66,30,66,29,117,31,149,31,138,31,187,31,86,31,111,31,111,30,96,31,96,30,96,29,220,31,200,31,169,31,169,30,58,31,120,31,246,31,246,30,94,31,134,31,48,31,151,31,89,31,89,30,252,31,107,31,228,31,210,31,19,31,31,31,17,31,116,31,45,31,27,31,61,31,61,30,61,29,61,28,21,31,238,31,96,31,147,31,47,31,47,30,47,29,47,28,47,27,8,31,143,31,168,31,85,31,60,31,204,31,20,31,113,31,124,31,43,31,74,31,74,30,199,31,199,30,47,31,47,30,178,31,234,31,234,30,135,31,26,31,26,30,133,31,245,31,245,30,235,31,140,31,52,31,233,31,233,30,192,31,3,31,151,31,151,30,151,29,224,31,224,30,40,31,197,31,143,31,127,31,108,31,165,31,113,31,113,30,164,31,3,31,92,31,212,31,110,31,168,31,125,31,239,31,237,31,237,30,169,31,168,31,168,30,58,31,126,31,223,31,197,31,65,31,82,31,177,31,21,31,78,31,111,31,206,31,206,30,64,31,24,31,4,31,250,31,148,31,13,31,88,31,96,31,124,31,124,30,68,31,97,31,97,30,187,31,91,31,33,31,33,30,132,31,201,31,49,31,48,31,95,31,177,31,63,31,252,31,191,31,116,31,252,31,129,31,2,31,5,31,222,31,62,31,216,31,216,30,216,29,78,31,15,31,242,31,73,31,149,31,146,31,25,31,140,31,99,31,64,31,127,31,127,30,165,31,141,31,141,30,167,31,57,31,84,31,84,30,223,31,117,31,73,31,125,31,142,31,41,31,211,31,17,31,124,31,124,30,164,31,179,31,145,31,200,31,200,30,200,29,47,31,51,31,80,31,20,31,115,31,47,31,110,31,175,31,229,31,63,31,163,31,131,31,65,31,141,31,141,30,87,31,105,31,216,31,220,31,248,31,207,31,207,30,147,31,101,31,202,31,115,31,115,30,51,31,51,30,70,31,216,31,125,31,125,30,61,31,225,31,158,31,167,31,86,31,115,31,102,31,250,31,1,31,1,30,220,31,49,31,61,31,61,30,61,29,255,31,232,31,195,31,246,31,185,31,174,31,243,31,161,31,177,31,59,31,59,30,212,31,212,30,237,31,237,30,116,31,250,31,63,31,213,31,223,31,65,31,198,31,38,31,139,31,52,31,246,31,246,30,215,31,41,31,189,31,189,30,189,29,36,31,87,31,125,31,239,31,47,31,187,31,187,30,187,31,187,30,25,31,26,31,253,31,78,31,123,31,123,30,255,31,45,31,139,31,3,31,96,31,79,31,190,31,222,31,235,31,28,31,115,31,45,31,161,31,167,31,10,31,99,31,239,31,239,30,119,31,106,31,186,31,23,31,235,31,13,31,58,31,180,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
