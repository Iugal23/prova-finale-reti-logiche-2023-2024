-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_521 is
end project_tb_521;

architecture project_tb_arch_521 of project_tb_521 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 934;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (77,0,0,0,142,0,198,0,74,0,135,0,0,0,97,0,161,0,0,0,0,0,90,0,119,0,4,0,164,0,171,0,0,0,108,0,0,0,182,0,241,0,0,0,69,0,182,0,109,0,92,0,138,0,187,0,249,0,0,0,133,0,61,0,233,0,20,0,61,0,101,0,0,0,139,0,182,0,57,0,225,0,131,0,0,0,217,0,196,0,211,0,144,0,0,0,247,0,198,0,49,0,44,0,168,0,202,0,80,0,105,0,49,0,14,0,250,0,115,0,0,0,223,0,15,0,0,0,7,0,120,0,58,0,177,0,0,0,0,0,255,0,0,0,0,0,255,0,254,0,3,0,244,0,214,0,0,0,86,0,129,0,194,0,96,0,0,0,7,0,120,0,0,0,73,0,123,0,23,0,195,0,207,0,137,0,253,0,0,0,2,0,173,0,140,0,124,0,42,0,243,0,174,0,199,0,178,0,62,0,191,0,0,0,220,0,243,0,0,0,0,0,76,0,202,0,0,0,139,0,32,0,105,0,0,0,82,0,20,0,46,0,6,0,30,0,68,0,223,0,0,0,0,0,86,0,150,0,35,0,172,0,0,0,232,0,97,0,231,0,227,0,180,0,249,0,200,0,179,0,34,0,18,0,61,0,150,0,94,0,8,0,154,0,107,0,122,0,33,0,0,0,224,0,32,0,0,0,104,0,161,0,205,0,74,0,211,0,192,0,0,0,147,0,78,0,0,0,109,0,255,0,177,0,28,0,132,0,150,0,0,0,159,0,145,0,210,0,0,0,29,0,241,0,238,0,141,0,160,0,63,0,182,0,151,0,190,0,0,0,31,0,87,0,111,0,176,0,111,0,34,0,187,0,0,0,191,0,154,0,0,0,40,0,21,0,66,0,95,0,12,0,50,0,144,0,126,0,0,0,0,0,64,0,117,0,0,0,10,0,71,0,86,0,167,0,1,0,187,0,23,0,0,0,165,0,57,0,100,0,0,0,116,0,251,0,71,0,0,0,235,0,0,0,103,0,211,0,242,0,9,0,213,0,134,0,106,0,141,0,0,0,161,0,46,0,126,0,0,0,15,0,221,0,211,0,109,0,122,0,250,0,240,0,33,0,186,0,0,0,216,0,0,0,185,0,188,0,31,0,0,0,0,0,19,0,94,0,0,0,25,0,0,0,0,0,0,0,217,0,125,0,144,0,29,0,77,0,99,0,154,0,89,0,68,0,168,0,9,0,230,0,0,0,78,0,55,0,187,0,0,0,198,0,205,0,101,0,0,0,185,0,205,0,79,0,0,0,0,0,214,0,0,0,0,0,13,0,35,0,0,0,0,0,194,0,7,0,0,0,238,0,0,0,235,0,28,0,0,0,184,0,0,0,47,0,0,0,77,0,130,0,70,0,176,0,142,0,0,0,49,0,232,0,0,0,78,0,241,0,108,0,119,0,6,0,184,0,23,0,0,0,0,0,0,0,53,0,180,0,184,0,33,0,243,0,70,0,121,0,0,0,33,0,41,0,0,0,154,0,254,0,93,0,91,0,164,0,113,0,162,0,0,0,140,0,0,0,116,0,169,0,45,0,189,0,229,0,164,0,148,0,145,0,0,0,44,0,0,0,11,0,202,0,245,0,109,0,50,0,241,0,106,0,198,0,0,0,228,0,0,0,212,0,0,0,59,0,40,0,113,0,142,0,103,0,4,0,204,0,185,0,153,0,135,0,215,0,53,0,116,0,195,0,201,0,92,0,2,0,224,0,222,0,0,0,0,0,48,0,193,0,250,0,171,0,21,0,119,0,0,0,148,0,197,0,87,0,13,0,0,0,0,0,183,0,17,0,40,0,105,0,244,0,0,0,59,0,0,0,116,0,50,0,154,0,0,0,102,0,0,0,218,0,232,0,34,0,234,0,164,0,180,0,228,0,212,0,28,0,142,0,0,0,63,0,149,0,0,0,0,0,241,0,130,0,175,0,16,0,18,0,0,0,59,0,77,0,0,0,66,0,134,0,11,0,195,0,145,0,216,0,0,0,0,0,9,0,107,0,0,0,91,0,118,0,0,0,135,0,30,0,0,0,79,0,28,0,0,0,39,0,59,0,61,0,205,0,0,0,159,0,250,0,150,0,67,0,0,0,111,0,126,0,30,0,0,0,238,0,194,0,0,0,24,0,21,0,152,0,0,0,134,0,139,0,196,0,96,0,58,0,171,0,158,0,213,0,0,0,0,0,244,0,105,0,213,0,209,0,198,0,248,0,145,0,0,0,183,0,91,0,234,0,26,0,229,0,243,0,239,0,40,0,0,0,28,0,1,0,81,0,61,0,132,0,0,0,254,0,85,0,0,0,37,0,96,0,237,0,0,0,118,0,42,0,0,0,255,0,228,0,160,0,178,0,86,0,0,0,131,0,0,0,162,0,0,0,0,0,0,0,172,0,30,0,253,0,67,0,109,0,159,0,99,0,47,0,0,0,86,0,103,0,240,0,47,0,53,0,108,0,207,0,102,0,156,0,47,0,69,0,0,0,94,0,251,0,0,0,199,0,0,0,37,0,48,0,122,0,18,0,87,0,161,0,0,0,74,0,124,0,32,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,185,0,164,0,26,0,203,0,121,0,0,0,0,0,0,0,0,0,0,0,60,0,44,0,103,0,204,0,114,0,182,0,216,0,254,0,212,0,127,0,88,0,46,0,136,0,115,0,71,0,195,0,98,0,11,0,42,0,85,0,69,0,5,0,231,0,29,0,232,0,0,0,3,0,236,0,11,0,164,0,182,0,168,0,64,0,255,0,66,0,133,0,184,0,239,0,158,0,0,0,175,0,187,0,0,0,71,0,250,0,254,0,120,0,51,0,0,0,0,0,164,0,255,0,0,0,63,0,70,0,123,0,0,0,0,0,243,0,0,0,226,0,68,0,206,0,140,0,254,0,0,0,141,0,204,0,65,0,89,0,93,0,162,0,8,0,91,0,162,0,0,0,0,0,39,0,193,0,126,0,156,0,89,0,0,0,39,0,58,0,67,0,12,0,52,0,6,0,39,0,60,0,163,0,254,0,0,0,119,0,113,0,0,0,142,0,175,0,59,0,14,0,0,0,141,0,226,0,133,0,141,0,183,0,136,0,226,0,137,0,46,0,254,0,0,0,237,0,196,0,0,0,165,0,61,0,0,0,144,0,141,0,59,0,58,0,17,0,234,0,0,0,46,0,27,0,0,0,96,0,124,0,0,0,0,0,104,0,215,0,92,0,22,0,0,0,25,0,170,0,24,0,11,0,9,0,88,0,92,0,0,0,247,0,111,0,83,0,0,0,5,0,139,0,124,0,189,0,6,0,7,0,46,0,39,0,101,0,238,0,0,0,56,0,183,0,142,0,158,0,117,0,0,0,27,0,0,0,111,0,50,0,163,0,122,0,224,0,147,0,219,0,0,0,0,0,176,0,58,0,63,0,134,0,33,0,124,0,0,0,85,0,226,0,0,0,201,0,16,0,226,0,228,0,8,0,248,0,29,0,0,0,125,0,0,0,203,0,111,0,192,0,7,0,0,0,0,0,189,0,27,0,0,0,196,0,86,0,245,0,0,0,132,0,79,0,207,0,59,0,0,0,7,0,0,0,138,0,0,0,214,0,4,0,238,0,167,0,8,0,154,0,255,0,164,0,163,0,84,0,99,0,0,0,223,0,82,0,16,0,222,0,89,0,0,0,0,0,225,0,54,0,127,0,101,0,0,0,125,0,52,0,211,0,197,0,192,0,131,0,12,0,0,0,133,0,215,0,178,0,62,0,60,0,82,0,222,0,72,0,182,0,204,0,179,0,0,0,0,0,124,0,178,0,220,0,185,0,132,0,255,0,80,0,159,0,56,0,220,0,158,0,121,0,0,0,72,0,103,0,150,0,51,0,0,0,0,0,0,0,0,0,0,0,110,0,50,0,126,0,0,0,229,0,0,0,212,0,243,0,64,0,97,0,161,0,251,0,0,0,252,0,139,0,255,0,211,0,191,0,184,0,122,0,146,0,50,0,130,0,213,0,0,0,255,0,0,0,237,0,254,0,209,0,237,0,122,0,151,0,0,0,117,0,180,0,145,0,117,0,40,0,144,0,84,0,137,0,190,0,0,0,20,0,0,0,44,0,0,0,124,0,0,0,4,0,137,0);
signal scenario_full  : scenario_type := (77,31,77,30,142,31,198,31,74,31,135,31,135,30,97,31,161,31,161,30,161,29,90,31,119,31,4,31,164,31,171,31,171,30,108,31,108,30,182,31,241,31,241,30,69,31,182,31,109,31,92,31,138,31,187,31,249,31,249,30,133,31,61,31,233,31,20,31,61,31,101,31,101,30,139,31,182,31,57,31,225,31,131,31,131,30,217,31,196,31,211,31,144,31,144,30,247,31,198,31,49,31,44,31,168,31,202,31,80,31,105,31,49,31,14,31,250,31,115,31,115,30,223,31,15,31,15,30,7,31,120,31,58,31,177,31,177,30,177,29,255,31,255,30,255,29,255,31,254,31,3,31,244,31,214,31,214,30,86,31,129,31,194,31,96,31,96,30,7,31,120,31,120,30,73,31,123,31,23,31,195,31,207,31,137,31,253,31,253,30,2,31,173,31,140,31,124,31,42,31,243,31,174,31,199,31,178,31,62,31,191,31,191,30,220,31,243,31,243,30,243,29,76,31,202,31,202,30,139,31,32,31,105,31,105,30,82,31,20,31,46,31,6,31,30,31,68,31,223,31,223,30,223,29,86,31,150,31,35,31,172,31,172,30,232,31,97,31,231,31,227,31,180,31,249,31,200,31,179,31,34,31,18,31,61,31,150,31,94,31,8,31,154,31,107,31,122,31,33,31,33,30,224,31,32,31,32,30,104,31,161,31,205,31,74,31,211,31,192,31,192,30,147,31,78,31,78,30,109,31,255,31,177,31,28,31,132,31,150,31,150,30,159,31,145,31,210,31,210,30,29,31,241,31,238,31,141,31,160,31,63,31,182,31,151,31,190,31,190,30,31,31,87,31,111,31,176,31,111,31,34,31,187,31,187,30,191,31,154,31,154,30,40,31,21,31,66,31,95,31,12,31,50,31,144,31,126,31,126,30,126,29,64,31,117,31,117,30,10,31,71,31,86,31,167,31,1,31,187,31,23,31,23,30,165,31,57,31,100,31,100,30,116,31,251,31,71,31,71,30,235,31,235,30,103,31,211,31,242,31,9,31,213,31,134,31,106,31,141,31,141,30,161,31,46,31,126,31,126,30,15,31,221,31,211,31,109,31,122,31,250,31,240,31,33,31,186,31,186,30,216,31,216,30,185,31,188,31,31,31,31,30,31,29,19,31,94,31,94,30,25,31,25,30,25,29,25,28,217,31,125,31,144,31,29,31,77,31,99,31,154,31,89,31,68,31,168,31,9,31,230,31,230,30,78,31,55,31,187,31,187,30,198,31,205,31,101,31,101,30,185,31,205,31,79,31,79,30,79,29,214,31,214,30,214,29,13,31,35,31,35,30,35,29,194,31,7,31,7,30,238,31,238,30,235,31,28,31,28,30,184,31,184,30,47,31,47,30,77,31,130,31,70,31,176,31,142,31,142,30,49,31,232,31,232,30,78,31,241,31,108,31,119,31,6,31,184,31,23,31,23,30,23,29,23,28,53,31,180,31,184,31,33,31,243,31,70,31,121,31,121,30,33,31,41,31,41,30,154,31,254,31,93,31,91,31,164,31,113,31,162,31,162,30,140,31,140,30,116,31,169,31,45,31,189,31,229,31,164,31,148,31,145,31,145,30,44,31,44,30,11,31,202,31,245,31,109,31,50,31,241,31,106,31,198,31,198,30,228,31,228,30,212,31,212,30,59,31,40,31,113,31,142,31,103,31,4,31,204,31,185,31,153,31,135,31,215,31,53,31,116,31,195,31,201,31,92,31,2,31,224,31,222,31,222,30,222,29,48,31,193,31,250,31,171,31,21,31,119,31,119,30,148,31,197,31,87,31,13,31,13,30,13,29,183,31,17,31,40,31,105,31,244,31,244,30,59,31,59,30,116,31,50,31,154,31,154,30,102,31,102,30,218,31,232,31,34,31,234,31,164,31,180,31,228,31,212,31,28,31,142,31,142,30,63,31,149,31,149,30,149,29,241,31,130,31,175,31,16,31,18,31,18,30,59,31,77,31,77,30,66,31,134,31,11,31,195,31,145,31,216,31,216,30,216,29,9,31,107,31,107,30,91,31,118,31,118,30,135,31,30,31,30,30,79,31,28,31,28,30,39,31,59,31,61,31,205,31,205,30,159,31,250,31,150,31,67,31,67,30,111,31,126,31,30,31,30,30,238,31,194,31,194,30,24,31,21,31,152,31,152,30,134,31,139,31,196,31,96,31,58,31,171,31,158,31,213,31,213,30,213,29,244,31,105,31,213,31,209,31,198,31,248,31,145,31,145,30,183,31,91,31,234,31,26,31,229,31,243,31,239,31,40,31,40,30,28,31,1,31,81,31,61,31,132,31,132,30,254,31,85,31,85,30,37,31,96,31,237,31,237,30,118,31,42,31,42,30,255,31,228,31,160,31,178,31,86,31,86,30,131,31,131,30,162,31,162,30,162,29,162,28,172,31,30,31,253,31,67,31,109,31,159,31,99,31,47,31,47,30,86,31,103,31,240,31,47,31,53,31,108,31,207,31,102,31,156,31,47,31,69,31,69,30,94,31,251,31,251,30,199,31,199,30,37,31,48,31,122,31,18,31,87,31,161,31,161,30,74,31,124,31,32,31,32,30,32,29,32,28,32,27,32,26,32,25,32,24,32,23,185,31,164,31,26,31,203,31,121,31,121,30,121,29,121,28,121,27,121,26,60,31,44,31,103,31,204,31,114,31,182,31,216,31,254,31,212,31,127,31,88,31,46,31,136,31,115,31,71,31,195,31,98,31,11,31,42,31,85,31,69,31,5,31,231,31,29,31,232,31,232,30,3,31,236,31,11,31,164,31,182,31,168,31,64,31,255,31,66,31,133,31,184,31,239,31,158,31,158,30,175,31,187,31,187,30,71,31,250,31,254,31,120,31,51,31,51,30,51,29,164,31,255,31,255,30,63,31,70,31,123,31,123,30,123,29,243,31,243,30,226,31,68,31,206,31,140,31,254,31,254,30,141,31,204,31,65,31,89,31,93,31,162,31,8,31,91,31,162,31,162,30,162,29,39,31,193,31,126,31,156,31,89,31,89,30,39,31,58,31,67,31,12,31,52,31,6,31,39,31,60,31,163,31,254,31,254,30,119,31,113,31,113,30,142,31,175,31,59,31,14,31,14,30,141,31,226,31,133,31,141,31,183,31,136,31,226,31,137,31,46,31,254,31,254,30,237,31,196,31,196,30,165,31,61,31,61,30,144,31,141,31,59,31,58,31,17,31,234,31,234,30,46,31,27,31,27,30,96,31,124,31,124,30,124,29,104,31,215,31,92,31,22,31,22,30,25,31,170,31,24,31,11,31,9,31,88,31,92,31,92,30,247,31,111,31,83,31,83,30,5,31,139,31,124,31,189,31,6,31,7,31,46,31,39,31,101,31,238,31,238,30,56,31,183,31,142,31,158,31,117,31,117,30,27,31,27,30,111,31,50,31,163,31,122,31,224,31,147,31,219,31,219,30,219,29,176,31,58,31,63,31,134,31,33,31,124,31,124,30,85,31,226,31,226,30,201,31,16,31,226,31,228,31,8,31,248,31,29,31,29,30,125,31,125,30,203,31,111,31,192,31,7,31,7,30,7,29,189,31,27,31,27,30,196,31,86,31,245,31,245,30,132,31,79,31,207,31,59,31,59,30,7,31,7,30,138,31,138,30,214,31,4,31,238,31,167,31,8,31,154,31,255,31,164,31,163,31,84,31,99,31,99,30,223,31,82,31,16,31,222,31,89,31,89,30,89,29,225,31,54,31,127,31,101,31,101,30,125,31,52,31,211,31,197,31,192,31,131,31,12,31,12,30,133,31,215,31,178,31,62,31,60,31,82,31,222,31,72,31,182,31,204,31,179,31,179,30,179,29,124,31,178,31,220,31,185,31,132,31,255,31,80,31,159,31,56,31,220,31,158,31,121,31,121,30,72,31,103,31,150,31,51,31,51,30,51,29,51,28,51,27,51,26,110,31,50,31,126,31,126,30,229,31,229,30,212,31,243,31,64,31,97,31,161,31,251,31,251,30,252,31,139,31,255,31,211,31,191,31,184,31,122,31,146,31,50,31,130,31,213,31,213,30,255,31,255,30,237,31,254,31,209,31,237,31,122,31,151,31,151,30,117,31,180,31,145,31,117,31,40,31,144,31,84,31,137,31,190,31,190,30,20,31,20,30,44,31,44,30,124,31,124,30,4,31,137,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
