-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 746;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,138,0,0,0,48,0,9,0,134,0,29,0,147,0,103,0,199,0,3,0,12,0,0,0,0,0,175,0,118,0,0,0,0,0,0,0,255,0,88,0,0,0,0,0,97,0,50,0,115,0,36,0,134,0,0,0,33,0,40,0,238,0,55,0,168,0,2,0,44,0,181,0,79,0,244,0,59,0,0,0,0,0,219,0,208,0,142,0,168,0,0,0,57,0,159,0,137,0,91,0,14,0,125,0,55,0,139,0,83,0,0,0,225,0,213,0,208,0,92,0,0,0,138,0,99,0,166,0,34,0,56,0,97,0,24,0,0,0,234,0,21,0,0,0,0,0,48,0,0,0,230,0,255,0,105,0,21,0,0,0,236,0,109,0,65,0,108,0,193,0,206,0,67,0,76,0,172,0,0,0,254,0,0,0,89,0,0,0,30,0,33,0,135,0,239,0,174,0,215,0,252,0,9,0,223,0,164,0,109,0,4,0,0,0,203,0,238,0,0,0,32,0,134,0,59,0,130,0,105,0,130,0,0,0,101,0,83,0,85,0,109,0,0,0,0,0,29,0,210,0,192,0,0,0,0,0,29,0,18,0,203,0,0,0,0,0,164,0,202,0,74,0,65,0,0,0,29,0,0,0,81,0,155,0,96,0,88,0,114,0,10,0,228,0,47,0,150,0,220,0,219,0,254,0,120,0,241,0,135,0,104,0,249,0,186,0,186,0,186,0,63,0,212,0,0,0,229,0,179,0,11,0,0,0,147,0,51,0,174,0,0,0,111,0,125,0,16,0,0,0,83,0,178,0,21,0,153,0,0,0,134,0,47,0,26,0,42,0,121,0,0,0,0,0,141,0,230,0,141,0,242,0,0,0,13,0,234,0,76,0,0,0,162,0,156,0,52,0,198,0,0,0,39,0,0,0,199,0,210,0,126,0,81,0,222,0,0,0,202,0,0,0,140,0,165,0,44,0,150,0,132,0,39,0,254,0,244,0,216,0,121,0,199,0,240,0,240,0,0,0,102,0,79,0,0,0,0,0,106,0,0,0,136,0,186,0,70,0,97,0,11,0,125,0,178,0,73,0,250,0,113,0,0,0,189,0,123,0,76,0,188,0,133,0,157,0,156,0,152,0,223,0,235,0,157,0,105,0,247,0,171,0,44,0,40,0,65,0,188,0,96,0,102,0,213,0,117,0,204,0,0,0,254,0,134,0,0,0,25,0,171,0,0,0,229,0,128,0,126,0,90,0,97,0,234,0,230,0,0,0,185,0,53,0,214,0,198,0,34,0,120,0,246,0,243,0,218,0,0,0,0,0,38,0,116,0,186,0,79,0,204,0,0,0,192,0,75,0,93,0,0,0,208,0,246,0,63,0,128,0,0,0,2,0,224,0,26,0,193,0,146,0,0,0,32,0,16,0,86,0,146,0,157,0,188,0,53,0,5,0,153,0,6,0,252,0,94,0,0,0,127,0,151,0,245,0,124,0,30,0,0,0,240,0,252,0,241,0,0,0,100,0,106,0,0,0,185,0,128,0,67,0,251,0,187,0,247,0,49,0,231,0,163,0,60,0,201,0,0,0,236,0,194,0,235,0,248,0,111,0,168,0,251,0,204,0,0,0,239,0,0,0,86,0,0,0,0,0,30,0,121,0,124,0,0,0,49,0,108,0,103,0,121,0,107,0,26,0,203,0,138,0,175,0,170,0,0,0,105,0,0,0,71,0,0,0,0,0,125,0,84,0,220,0,0,0,27,0,40,0,0,0,43,0,220,0,73,0,234,0,0,0,0,0,99,0,159,0,130,0,27,0,71,0,0,0,115,0,138,0,82,0,211,0,0,0,0,0,221,0,86,0,0,0,254,0,3,0,86,0,0,0,1,0,0,0,163,0,98,0,51,0,0,0,194,0,151,0,122,0,86,0,50,0,0,0,159,0,143,0,0,0,152,0,223,0,151,0,61,0,0,0,189,0,61,0,0,0,218,0,0,0,120,0,127,0,0,0,0,0,220,0,190,0,129,0,174,0,51,0,30,0,187,0,74,0,0,0,167,0,144,0,35,0,147,0,186,0,0,0,253,0,208,0,0,0,87,0,107,0,102,0,0,0,0,0,223,0,95,0,139,0,232,0,201,0,60,0,226,0,87,0,75,0,96,0,158,0,191,0,161,0,0,0,97,0,55,0,21,0,29,0,194,0,124,0,42,0,72,0,217,0,161,0,123,0,0,0,137,0,21,0,250,0,154,0,30,0,186,0,48,0,11,0,0,0,0,0,46,0,0,0,187,0,121,0,110,0,0,0,241,0,144,0,93,0,159,0,231,0,215,0,199,0,33,0,3,0,156,0,68,0,64,0,52,0,130,0,165,0,28,0,0,0,207,0,99,0,88,0,253,0,0,0,236,0,70,0,161,0,21,0,254,0,33,0,10,0,217,0,230,0,97,0,31,0,0,0,210,0,199,0,0,0,59,0,231,0,0,0,4,0,152,0,174,0,228,0,140,0,47,0,177,0,68,0,36,0,83,0,0,0,210,0,0,0,193,0,136,0,139,0,166,0,196,0,129,0,251,0,201,0,132,0,169,0,27,0,247,0,105,0,219,0,0,0,158,0,252,0,76,0,206,0,142,0,216,0,168,0,28,0,105,0,83,0,209,0,23,0,0,0,42,0,147,0,0,0,6,0,184,0,120,0,245,0,4,0,20,0,155,0,133,0,121,0,7,0,157,0,51,0,68,0,214,0,62,0,0,0,11,0,218,0,234,0,185,0,64,0,153,0,134,0,79,0,0,0,216,0,179,0,0,0,153,0,208,0,113,0,34,0,63,0,137,0,0,0,168,0,231,0,239,0,139,0,163,0,93,0,0,0,23,0,181,0,118,0,0,0,179,0,76,0,117,0,73,0,0,0,0,0,138,0,0,0,48,0,25,0,90,0,60,0,0,0,207,0,146,0,223,0,192,0,0,0,58,0,100,0,185,0,84,0,12,0,122,0,51,0,237,0,0,0,0,0,0,0,0,0,252,0,4,0,203,0,0,0,96,0,49,0,46,0,64,0,53,0,69,0,217,0,246,0,0,0,0,0,128,0,82,0,4,0,73,0,171,0,0,0,238,0,183,0,188,0,242,0,242,0,225,0,166,0,91,0,190,0,210,0,79,0,9,0,0,0,187,0,62,0,0,0,86,0,119,0,199,0,0,0,128,0,36,0,24,0,109,0,207,0,69,0,147,0,193,0,112,0,119,0,210,0,0,0,168,0,106,0,109,0,99,0,0,0,4,0,220,0,45,0,15,0,0,0,22,0,150,0,44,0,81,0,205,0,81,0,239,0,225,0,116,0,0,0,66,0,87,0,0,0);
signal scenario_full  : scenario_type := (0,0,138,31,138,30,48,31,9,31,134,31,29,31,147,31,103,31,199,31,3,31,12,31,12,30,12,29,175,31,118,31,118,30,118,29,118,28,255,31,88,31,88,30,88,29,97,31,50,31,115,31,36,31,134,31,134,30,33,31,40,31,238,31,55,31,168,31,2,31,44,31,181,31,79,31,244,31,59,31,59,30,59,29,219,31,208,31,142,31,168,31,168,30,57,31,159,31,137,31,91,31,14,31,125,31,55,31,139,31,83,31,83,30,225,31,213,31,208,31,92,31,92,30,138,31,99,31,166,31,34,31,56,31,97,31,24,31,24,30,234,31,21,31,21,30,21,29,48,31,48,30,230,31,255,31,105,31,21,31,21,30,236,31,109,31,65,31,108,31,193,31,206,31,67,31,76,31,172,31,172,30,254,31,254,30,89,31,89,30,30,31,33,31,135,31,239,31,174,31,215,31,252,31,9,31,223,31,164,31,109,31,4,31,4,30,203,31,238,31,238,30,32,31,134,31,59,31,130,31,105,31,130,31,130,30,101,31,83,31,85,31,109,31,109,30,109,29,29,31,210,31,192,31,192,30,192,29,29,31,18,31,203,31,203,30,203,29,164,31,202,31,74,31,65,31,65,30,29,31,29,30,81,31,155,31,96,31,88,31,114,31,10,31,228,31,47,31,150,31,220,31,219,31,254,31,120,31,241,31,135,31,104,31,249,31,186,31,186,31,186,31,63,31,212,31,212,30,229,31,179,31,11,31,11,30,147,31,51,31,174,31,174,30,111,31,125,31,16,31,16,30,83,31,178,31,21,31,153,31,153,30,134,31,47,31,26,31,42,31,121,31,121,30,121,29,141,31,230,31,141,31,242,31,242,30,13,31,234,31,76,31,76,30,162,31,156,31,52,31,198,31,198,30,39,31,39,30,199,31,210,31,126,31,81,31,222,31,222,30,202,31,202,30,140,31,165,31,44,31,150,31,132,31,39,31,254,31,244,31,216,31,121,31,199,31,240,31,240,31,240,30,102,31,79,31,79,30,79,29,106,31,106,30,136,31,186,31,70,31,97,31,11,31,125,31,178,31,73,31,250,31,113,31,113,30,189,31,123,31,76,31,188,31,133,31,157,31,156,31,152,31,223,31,235,31,157,31,105,31,247,31,171,31,44,31,40,31,65,31,188,31,96,31,102,31,213,31,117,31,204,31,204,30,254,31,134,31,134,30,25,31,171,31,171,30,229,31,128,31,126,31,90,31,97,31,234,31,230,31,230,30,185,31,53,31,214,31,198,31,34,31,120,31,246,31,243,31,218,31,218,30,218,29,38,31,116,31,186,31,79,31,204,31,204,30,192,31,75,31,93,31,93,30,208,31,246,31,63,31,128,31,128,30,2,31,224,31,26,31,193,31,146,31,146,30,32,31,16,31,86,31,146,31,157,31,188,31,53,31,5,31,153,31,6,31,252,31,94,31,94,30,127,31,151,31,245,31,124,31,30,31,30,30,240,31,252,31,241,31,241,30,100,31,106,31,106,30,185,31,128,31,67,31,251,31,187,31,247,31,49,31,231,31,163,31,60,31,201,31,201,30,236,31,194,31,235,31,248,31,111,31,168,31,251,31,204,31,204,30,239,31,239,30,86,31,86,30,86,29,30,31,121,31,124,31,124,30,49,31,108,31,103,31,121,31,107,31,26,31,203,31,138,31,175,31,170,31,170,30,105,31,105,30,71,31,71,30,71,29,125,31,84,31,220,31,220,30,27,31,40,31,40,30,43,31,220,31,73,31,234,31,234,30,234,29,99,31,159,31,130,31,27,31,71,31,71,30,115,31,138,31,82,31,211,31,211,30,211,29,221,31,86,31,86,30,254,31,3,31,86,31,86,30,1,31,1,30,163,31,98,31,51,31,51,30,194,31,151,31,122,31,86,31,50,31,50,30,159,31,143,31,143,30,152,31,223,31,151,31,61,31,61,30,189,31,61,31,61,30,218,31,218,30,120,31,127,31,127,30,127,29,220,31,190,31,129,31,174,31,51,31,30,31,187,31,74,31,74,30,167,31,144,31,35,31,147,31,186,31,186,30,253,31,208,31,208,30,87,31,107,31,102,31,102,30,102,29,223,31,95,31,139,31,232,31,201,31,60,31,226,31,87,31,75,31,96,31,158,31,191,31,161,31,161,30,97,31,55,31,21,31,29,31,194,31,124,31,42,31,72,31,217,31,161,31,123,31,123,30,137,31,21,31,250,31,154,31,30,31,186,31,48,31,11,31,11,30,11,29,46,31,46,30,187,31,121,31,110,31,110,30,241,31,144,31,93,31,159,31,231,31,215,31,199,31,33,31,3,31,156,31,68,31,64,31,52,31,130,31,165,31,28,31,28,30,207,31,99,31,88,31,253,31,253,30,236,31,70,31,161,31,21,31,254,31,33,31,10,31,217,31,230,31,97,31,31,31,31,30,210,31,199,31,199,30,59,31,231,31,231,30,4,31,152,31,174,31,228,31,140,31,47,31,177,31,68,31,36,31,83,31,83,30,210,31,210,30,193,31,136,31,139,31,166,31,196,31,129,31,251,31,201,31,132,31,169,31,27,31,247,31,105,31,219,31,219,30,158,31,252,31,76,31,206,31,142,31,216,31,168,31,28,31,105,31,83,31,209,31,23,31,23,30,42,31,147,31,147,30,6,31,184,31,120,31,245,31,4,31,20,31,155,31,133,31,121,31,7,31,157,31,51,31,68,31,214,31,62,31,62,30,11,31,218,31,234,31,185,31,64,31,153,31,134,31,79,31,79,30,216,31,179,31,179,30,153,31,208,31,113,31,34,31,63,31,137,31,137,30,168,31,231,31,239,31,139,31,163,31,93,31,93,30,23,31,181,31,118,31,118,30,179,31,76,31,117,31,73,31,73,30,73,29,138,31,138,30,48,31,25,31,90,31,60,31,60,30,207,31,146,31,223,31,192,31,192,30,58,31,100,31,185,31,84,31,12,31,122,31,51,31,237,31,237,30,237,29,237,28,237,27,252,31,4,31,203,31,203,30,96,31,49,31,46,31,64,31,53,31,69,31,217,31,246,31,246,30,246,29,128,31,82,31,4,31,73,31,171,31,171,30,238,31,183,31,188,31,242,31,242,31,225,31,166,31,91,31,190,31,210,31,79,31,9,31,9,30,187,31,62,31,62,30,86,31,119,31,199,31,199,30,128,31,36,31,24,31,109,31,207,31,69,31,147,31,193,31,112,31,119,31,210,31,210,30,168,31,106,31,109,31,99,31,99,30,4,31,220,31,45,31,15,31,15,30,22,31,150,31,44,31,81,31,205,31,81,31,239,31,225,31,116,31,116,30,66,31,87,31,87,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
