-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_10 is
end project_tb_10;

architecture project_tb_arch_10 of project_tb_10 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 688;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (101,0,157,0,249,0,0,0,248,0,166,0,39,0,44,0,0,0,14,0,175,0,141,0,37,0,185,0,68,0,87,0,184,0,144,0,216,0,179,0,48,0,66,0,17,0,186,0,147,0,149,0,161,0,123,0,7,0,168,0,71,0,127,0,0,0,61,0,89,0,187,0,0,0,96,0,98,0,146,0,138,0,194,0,131,0,86,0,252,0,211,0,175,0,190,0,69,0,230,0,5,0,125,0,0,0,26,0,211,0,33,0,235,0,168,0,120,0,240,0,9,0,143,0,0,0,209,0,104,0,236,0,42,0,162,0,67,0,181,0,209,0,45,0,225,0,0,0,0,0,237,0,39,0,52,0,58,0,48,0,24,0,9,0,167,0,117,0,0,0,106,0,115,0,0,0,0,0,112,0,108,0,98,0,0,0,0,0,166,0,82,0,98,0,100,0,0,0,0,0,0,0,0,0,0,0,40,0,220,0,24,0,162,0,58,0,26,0,119,0,220,0,177,0,197,0,199,0,20,0,0,0,149,0,0,0,0,0,110,0,217,0,0,0,148,0,0,0,119,0,186,0,126,0,105,0,115,0,23,0,105,0,11,0,164,0,14,0,86,0,8,0,0,0,101,0,20,0,0,0,31,0,228,0,118,0,236,0,179,0,244,0,164,0,113,0,0,0,196,0,100,0,196,0,74,0,95,0,159,0,38,0,20,0,193,0,157,0,109,0,173,0,103,0,109,0,0,0,9,0,174,0,115,0,158,0,0,0,0,0,238,0,206,0,66,0,87,0,254,0,237,0,192,0,0,0,105,0,0,0,222,0,238,0,116,0,0,0,207,0,39,0,0,0,181,0,67,0,178,0,2,0,0,0,23,0,188,0,100,0,224,0,113,0,105,0,109,0,49,0,40,0,152,0,151,0,0,0,184,0,3,0,0,0,191,0,83,0,177,0,234,0,0,0,152,0,36,0,127,0,94,0,177,0,207,0,0,0,107,0,154,0,124,0,168,0,0,0,147,0,50,0,0,0,157,0,247,0,60,0,0,0,21,0,181,0,185,0,185,0,131,0,199,0,99,0,92,0,0,0,240,0,0,0,0,0,0,0,244,0,177,0,16,0,0,0,134,0,163,0,102,0,33,0,135,0,232,0,0,0,39,0,0,0,172,0,166,0,220,0,31,0,86,0,92,0,254,0,122,0,190,0,61,0,0,0,0,0,0,0,34,0,86,0,214,0,0,0,210,0,12,0,54,0,0,0,28,0,183,0,181,0,59,0,172,0,24,0,67,0,0,0,197,0,0,0,17,0,101,0,48,0,0,0,0,0,121,0,136,0,47,0,229,0,65,0,191,0,138,0,0,0,1,0,28,0,177,0,77,0,0,0,50,0,150,0,180,0,0,0,162,0,0,0,11,0,0,0,0,0,19,0,17,0,78,0,0,0,126,0,98,0,207,0,0,0,0,0,124,0,142,0,217,0,0,0,9,0,198,0,0,0,215,0,0,0,119,0,151,0,80,0,117,0,165,0,43,0,68,0,0,0,32,0,128,0,31,0,87,0,209,0,0,0,191,0,0,0,65,0,229,0,26,0,44,0,0,0,0,0,198,0,75,0,206,0,33,0,0,0,74,0,95,0,46,0,255,0,142,0,65,0,0,0,0,0,63,0,5,0,216,0,156,0,135,0,79,0,107,0,156,0,50,0,169,0,110,0,98,0,40,0,156,0,82,0,212,0,102,0,191,0,216,0,42,0,222,0,85,0,79,0,23,0,205,0,0,0,48,0,194,0,0,0,84,0,181,0,10,0,105,0,0,0,212,0,173,0,0,0,0,0,0,0,14,0,0,0,178,0,81,0,26,0,157,0,101,0,0,0,0,0,130,0,245,0,115,0,44,0,208,0,139,0,0,0,122,0,74,0,13,0,116,0,213,0,249,0,0,0,224,0,0,0,0,0,0,0,104,0,111,0,206,0,28,0,231,0,148,0,118,0,161,0,10,0,0,0,0,0,129,0,122,0,175,0,53,0,13,0,32,0,35,0,0,0,197,0,0,0,74,0,71,0,0,0,195,0,9,0,0,0,192,0,126,0,0,0,150,0,87,0,130,0,253,0,145,0,148,0,158,0,16,0,231,0,0,0,198,0,249,0,0,0,50,0,109,0,248,0,235,0,246,0,91,0,153,0,116,0,40,0,141,0,151,0,7,0,204,0,121,0,219,0,184,0,27,0,159,0,165,0,0,0,152,0,113,0,193,0,76,0,47,0,176,0,131,0,0,0,74,0,6,0,60,0,0,0,138,0,188,0,71,0,41,0,5,0,61,0,55,0,0,0,244,0,0,0,0,0,195,0,212,0,0,0,162,0,55,0,92,0,236,0,21,0,163,0,185,0,24,0,0,0,167,0,0,0,202,0,141,0,0,0,0,0,101,0,0,0,0,0,0,0,42,0,104,0,35,0,255,0,172,0,88,0,36,0,0,0,0,0,94,0,45,0,41,0,143,0,248,0,0,0,0,0,1,0,247,0,224,0,84,0,199,0,208,0,111,0,241,0,181,0,92,0,155,0,144,0,0,0,83,0,100,0,6,0,177,0,0,0,218,0,144,0,233,0,111,0,0,0,73,0,16,0,110,0,235,0,0,0,62,0,218,0,0,0,174,0,0,0,101,0,112,0,36,0,51,0,253,0,14,0,118,0,0,0,49,0,45,0,19,0,230,0,71,0,115,0,240,0,40,0,51,0,0,0,102,0,127,0,143,0,16,0,1,0,0,0,0,0,211,0,65,0,32,0,246,0,132,0,0,0,74,0,254,0,0,0,94,0,0,0,198,0,133,0,165,0,163,0,0,0,156,0,103,0,0,0,210,0,82,0,41,0,254,0,0,0,98,0,137,0,181,0,0,0,168,0,55,0,5,0,48,0,139,0,0,0,243,0,0,0,100,0,0,0,220,0,138,0,225,0,177,0,0,0,147,0,146,0,252,0,0,0,190,0,212,0,0,0,0,0,22,0,95,0,88,0,134,0,86,0,138,0,39,0,0,0,79,0,0,0,125,0,2,0,0,0,30,0,120,0,176,0,146,0,63,0,0,0,121,0,0,0);
signal scenario_full  : scenario_type := (101,31,157,31,249,31,249,30,248,31,166,31,39,31,44,31,44,30,14,31,175,31,141,31,37,31,185,31,68,31,87,31,184,31,144,31,216,31,179,31,48,31,66,31,17,31,186,31,147,31,149,31,161,31,123,31,7,31,168,31,71,31,127,31,127,30,61,31,89,31,187,31,187,30,96,31,98,31,146,31,138,31,194,31,131,31,86,31,252,31,211,31,175,31,190,31,69,31,230,31,5,31,125,31,125,30,26,31,211,31,33,31,235,31,168,31,120,31,240,31,9,31,143,31,143,30,209,31,104,31,236,31,42,31,162,31,67,31,181,31,209,31,45,31,225,31,225,30,225,29,237,31,39,31,52,31,58,31,48,31,24,31,9,31,167,31,117,31,117,30,106,31,115,31,115,30,115,29,112,31,108,31,98,31,98,30,98,29,166,31,82,31,98,31,100,31,100,30,100,29,100,28,100,27,100,26,40,31,220,31,24,31,162,31,58,31,26,31,119,31,220,31,177,31,197,31,199,31,20,31,20,30,149,31,149,30,149,29,110,31,217,31,217,30,148,31,148,30,119,31,186,31,126,31,105,31,115,31,23,31,105,31,11,31,164,31,14,31,86,31,8,31,8,30,101,31,20,31,20,30,31,31,228,31,118,31,236,31,179,31,244,31,164,31,113,31,113,30,196,31,100,31,196,31,74,31,95,31,159,31,38,31,20,31,193,31,157,31,109,31,173,31,103,31,109,31,109,30,9,31,174,31,115,31,158,31,158,30,158,29,238,31,206,31,66,31,87,31,254,31,237,31,192,31,192,30,105,31,105,30,222,31,238,31,116,31,116,30,207,31,39,31,39,30,181,31,67,31,178,31,2,31,2,30,23,31,188,31,100,31,224,31,113,31,105,31,109,31,49,31,40,31,152,31,151,31,151,30,184,31,3,31,3,30,191,31,83,31,177,31,234,31,234,30,152,31,36,31,127,31,94,31,177,31,207,31,207,30,107,31,154,31,124,31,168,31,168,30,147,31,50,31,50,30,157,31,247,31,60,31,60,30,21,31,181,31,185,31,185,31,131,31,199,31,99,31,92,31,92,30,240,31,240,30,240,29,240,28,244,31,177,31,16,31,16,30,134,31,163,31,102,31,33,31,135,31,232,31,232,30,39,31,39,30,172,31,166,31,220,31,31,31,86,31,92,31,254,31,122,31,190,31,61,31,61,30,61,29,61,28,34,31,86,31,214,31,214,30,210,31,12,31,54,31,54,30,28,31,183,31,181,31,59,31,172,31,24,31,67,31,67,30,197,31,197,30,17,31,101,31,48,31,48,30,48,29,121,31,136,31,47,31,229,31,65,31,191,31,138,31,138,30,1,31,28,31,177,31,77,31,77,30,50,31,150,31,180,31,180,30,162,31,162,30,11,31,11,30,11,29,19,31,17,31,78,31,78,30,126,31,98,31,207,31,207,30,207,29,124,31,142,31,217,31,217,30,9,31,198,31,198,30,215,31,215,30,119,31,151,31,80,31,117,31,165,31,43,31,68,31,68,30,32,31,128,31,31,31,87,31,209,31,209,30,191,31,191,30,65,31,229,31,26,31,44,31,44,30,44,29,198,31,75,31,206,31,33,31,33,30,74,31,95,31,46,31,255,31,142,31,65,31,65,30,65,29,63,31,5,31,216,31,156,31,135,31,79,31,107,31,156,31,50,31,169,31,110,31,98,31,40,31,156,31,82,31,212,31,102,31,191,31,216,31,42,31,222,31,85,31,79,31,23,31,205,31,205,30,48,31,194,31,194,30,84,31,181,31,10,31,105,31,105,30,212,31,173,31,173,30,173,29,173,28,14,31,14,30,178,31,81,31,26,31,157,31,101,31,101,30,101,29,130,31,245,31,115,31,44,31,208,31,139,31,139,30,122,31,74,31,13,31,116,31,213,31,249,31,249,30,224,31,224,30,224,29,224,28,104,31,111,31,206,31,28,31,231,31,148,31,118,31,161,31,10,31,10,30,10,29,129,31,122,31,175,31,53,31,13,31,32,31,35,31,35,30,197,31,197,30,74,31,71,31,71,30,195,31,9,31,9,30,192,31,126,31,126,30,150,31,87,31,130,31,253,31,145,31,148,31,158,31,16,31,231,31,231,30,198,31,249,31,249,30,50,31,109,31,248,31,235,31,246,31,91,31,153,31,116,31,40,31,141,31,151,31,7,31,204,31,121,31,219,31,184,31,27,31,159,31,165,31,165,30,152,31,113,31,193,31,76,31,47,31,176,31,131,31,131,30,74,31,6,31,60,31,60,30,138,31,188,31,71,31,41,31,5,31,61,31,55,31,55,30,244,31,244,30,244,29,195,31,212,31,212,30,162,31,55,31,92,31,236,31,21,31,163,31,185,31,24,31,24,30,167,31,167,30,202,31,141,31,141,30,141,29,101,31,101,30,101,29,101,28,42,31,104,31,35,31,255,31,172,31,88,31,36,31,36,30,36,29,94,31,45,31,41,31,143,31,248,31,248,30,248,29,1,31,247,31,224,31,84,31,199,31,208,31,111,31,241,31,181,31,92,31,155,31,144,31,144,30,83,31,100,31,6,31,177,31,177,30,218,31,144,31,233,31,111,31,111,30,73,31,16,31,110,31,235,31,235,30,62,31,218,31,218,30,174,31,174,30,101,31,112,31,36,31,51,31,253,31,14,31,118,31,118,30,49,31,45,31,19,31,230,31,71,31,115,31,240,31,40,31,51,31,51,30,102,31,127,31,143,31,16,31,1,31,1,30,1,29,211,31,65,31,32,31,246,31,132,31,132,30,74,31,254,31,254,30,94,31,94,30,198,31,133,31,165,31,163,31,163,30,156,31,103,31,103,30,210,31,82,31,41,31,254,31,254,30,98,31,137,31,181,31,181,30,168,31,55,31,5,31,48,31,139,31,139,30,243,31,243,30,100,31,100,30,220,31,138,31,225,31,177,31,177,30,147,31,146,31,252,31,252,30,190,31,212,31,212,30,212,29,22,31,95,31,88,31,134,31,86,31,138,31,39,31,39,30,79,31,79,30,125,31,2,31,2,30,30,31,120,31,176,31,146,31,63,31,63,30,121,31,121,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
