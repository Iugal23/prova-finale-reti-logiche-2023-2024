-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_257 is
end project_tb_257;

architecture project_tb_arch_257 of project_tb_257 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 926;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (26,0,15,0,100,0,225,0,94,0,0,0,63,0,49,0,0,0,59,0,229,0,70,0,0,0,0,0,246,0,0,0,127,0,251,0,104,0,174,0,158,0,178,0,233,0,140,0,45,0,157,0,202,0,148,0,253,0,167,0,54,0,204,0,142,0,74,0,129,0,0,0,223,0,157,0,193,0,0,0,70,0,216,0,72,0,49,0,0,0,0,0,164,0,188,0,96,0,34,0,84,0,0,0,39,0,60,0,180,0,213,0,0,0,0,0,236,0,15,0,41,0,39,0,221,0,66,0,220,0,0,0,115,0,200,0,2,0,16,0,49,0,130,0,0,0,0,0,0,0,20,0,0,0,147,0,0,0,161,0,59,0,151,0,65,0,0,0,229,0,0,0,250,0,101,0,0,0,73,0,46,0,40,0,26,0,226,0,56,0,100,0,0,0,58,0,166,0,11,0,218,0,85,0,213,0,0,0,133,0,15,0,178,0,96,0,135,0,35,0,233,0,3,0,93,0,209,0,52,0,0,0,131,0,239,0,0,0,0,0,148,0,248,0,78,0,96,0,120,0,218,0,244,0,0,0,92,0,38,0,0,0,250,0,0,0,36,0,175,0,0,0,184,0,49,0,11,0,242,0,148,0,233,0,246,0,197,0,96,0,161,0,227,0,196,0,155,0,162,0,162,0,224,0,219,0,120,0,0,0,0,0,104,0,127,0,0,0,0,0,0,0,224,0,158,0,22,0,224,0,28,0,0,0,94,0,164,0,170,0,117,0,228,0,0,0,181,0,14,0,142,0,16,0,0,0,170,0,203,0,224,0,0,0,145,0,175,0,7,0,121,0,96,0,140,0,0,0,54,0,83,0,195,0,0,0,192,0,40,0,189,0,50,0,70,0,0,0,248,0,156,0,141,0,182,0,204,0,235,0,250,0,0,0,117,0,255,0,0,0,180,0,64,0,0,0,100,0,10,0,156,0,67,0,197,0,79,0,0,0,129,0,149,0,34,0,155,0,127,0,0,0,126,0,209,0,242,0,0,0,144,0,226,0,23,0,87,0,68,0,213,0,10,0,97,0,247,0,14,0,60,0,0,0,204,0,67,0,137,0,135,0,148,0,204,0,0,0,0,0,0,0,3,0,90,0,0,0,209,0,131,0,244,0,181,0,159,0,224,0,89,0,0,0,169,0,83,0,0,0,210,0,255,0,0,0,139,0,243,0,108,0,228,0,164,0,215,0,5,0,0,0,233,0,0,0,84,0,0,0,176,0,0,0,48,0,165,0,249,0,111,0,98,0,0,0,60,0,203,0,0,0,63,0,59,0,144,0,0,0,84,0,148,0,0,0,114,0,201,0,70,0,177,0,95,0,128,0,3,0,209,0,79,0,0,0,2,0,241,0,131,0,230,0,97,0,119,0,158,0,108,0,240,0,0,0,221,0,49,0,0,0,122,0,171,0,165,0,121,0,0,0,0,0,0,0,0,0,0,0,75,0,105,0,0,0,0,0,180,0,117,0,0,0,131,0,161,0,166,0,201,0,235,0,125,0,207,0,226,0,203,0,0,0,0,0,142,0,0,0,30,0,44,0,46,0,0,0,142,0,234,0,23,0,0,0,134,0,127,0,165,0,194,0,55,0,114,0,158,0,68,0,26,0,210,0,81,0,107,0,89,0,154,0,12,0,131,0,212,0,158,0,0,0,65,0,13,0,83,0,85,0,189,0,187,0,82,0,125,0,178,0,191,0,106,0,7,0,140,0,0,0,184,0,135,0,184,0,42,0,40,0,241,0,0,0,248,0,233,0,63,0,0,0,198,0,246,0,164,0,84,0,84,0,23,0,41,0,124,0,0,0,154,0,34,0,0,0,219,0,138,0,166,0,95,0,0,0,246,0,143,0,234,0,58,0,32,0,0,0,150,0,114,0,189,0,6,0,35,0,0,0,176,0,0,0,154,0,157,0,133,0,151,0,0,0,0,0,100,0,15,0,38,0,147,0,206,0,66,0,143,0,128,0,3,0,214,0,85,0,0,0,30,0,222,0,13,0,66,0,163,0,96,0,224,0,0,0,126,0,134,0,235,0,151,0,35,0,165,0,135,0,191,0,120,0,0,0,131,0,151,0,99,0,26,0,179,0,107,0,0,0,85,0,204,0,0,0,103,0,10,0,237,0,95,0,68,0,2,0,14,0,23,0,137,0,0,0,28,0,249,0,171,0,1,0,23,0,0,0,154,0,205,0,184,0,0,0,115,0,76,0,67,0,207,0,166,0,0,0,0,0,238,0,105,0,45,0,46,0,146,0,233,0,207,0,125,0,226,0,199,0,0,0,95,0,81,0,65,0,22,0,222,0,142,0,0,0,0,0,177,0,77,0,172,0,64,0,252,0,0,0,57,0,112,0,16,0,235,0,166,0,241,0,237,0,185,0,218,0,25,0,241,0,22,0,229,0,0,0,125,0,231,0,100,0,1,0,0,0,116,0,76,0,0,0,216,0,0,0,131,0,201,0,0,0,2,0,174,0,0,0,240,0,188,0,81,0,0,0,31,0,152,0,147,0,146,0,140,0,82,0,245,0,0,0,0,0,188,0,0,0,0,0,35,0,0,0,228,0,154,0,158,0,77,0,226,0,0,0,183,0,243,0,125,0,26,0,124,0,53,0,48,0,206,0,55,0,65,0,21,0,166,0,186,0,159,0,0,0,0,0,119,0,59,0,61,0,198,0,38,0,51,0,62,0,93,0,24,0,248,0,113,0,0,0,219,0,170,0,0,0,123,0,0,0,232,0,32,0,22,0,30,0,52,0,0,0,205,0,13,0,103,0,255,0,192,0,32,0,190,0,105,0,9,0,30,0,68,0,143,0,19,0,0,0,247,0,160,0,81,0,0,0,236,0,146,0,222,0,75,0,106,0,152,0,144,0,0,0,60,0,64,0,44,0,228,0,0,0,95,0,244,0,143,0,50,0,120,0,107,0,4,0,0,0,107,0,4,0,29,0,61,0,253,0,123,0,132,0,60,0,9,0,94,0,0,0,121,0,183,0,0,0,155,0,87,0,147,0,207,0,62,0,248,0,144,0,0,0,0,0,115,0,248,0,7,0,15,0,160,0,39,0,8,0,165,0,82,0,142,0,147,0,118,0,12,0,0,0,48,0,0,0,128,0,182,0,97,0,0,0,237,0,7,0,19,0,15,0,0,0,0,0,109,0,121,0,136,0,130,0,158,0,0,0,67,0,86,0,156,0,150,0,177,0,0,0,57,0,115,0,0,0,179,0,90,0,58,0,239,0,0,0,126,0,232,0,0,0,17,0,21,0,74,0,37,0,36,0,0,0,22,0,20,0,232,0,181,0,31,0,230,0,140,0,3,0,189,0,96,0,18,0,92,0,106,0,200,0,1,0,0,0,103,0,127,0,0,0,0,0,174,0,241,0,137,0,246,0,171,0,144,0,36,0,53,0,153,0,50,0,142,0,0,0,143,0,0,0,48,0,63,0,95,0,16,0,0,0,167,0,89,0,30,0,37,0,22,0,0,0,222,0,243,0,11,0,66,0,0,0,0,0,127,0,97,0,89,0,36,0,109,0,0,0,0,0,0,0,0,0,130,0,168,0,0,0,119,0,138,0,34,0,247,0,174,0,113,0,184,0,106,0,187,0,199,0,0,0,251,0,174,0,120,0,0,0,35,0,205,0,173,0,77,0,140,0,207,0,37,0,0,0,70,0,114,0,167,0,0,0,169,0,66,0,55,0,153,0,18,0,75,0,86,0,165,0,183,0,0,0,223,0,245,0,187,0,51,0,70,0,0,0,140,0,222,0,0,0,165,0,32,0,164,0,0,0,0,0,0,0,196,0,0,0,235,0,207,0,0,0,99,0,122,0,110,0,0,0,236,0,63,0,151,0,95,0,231,0,6,0,220,0,34,0,159,0,0,0,189,0,48,0,114,0,111,0,88,0,111,0,0,0,0,0,31,0,205,0,0,0,238,0,71,0,0,0,194,0,149,0,235,0,0,0,119,0,144,0,124,0,40,0,193,0,143,0,0,0,40,0,255,0,218,0,62,0,195,0,43,0,168,0,187,0,184,0,254,0,50,0,0,0,238,0,186,0,245,0,0,0,22,0,0,0,1,0,197,0,92,0,33,0,0,0,0,0,125,0,0,0);
signal scenario_full  : scenario_type := (26,31,15,31,100,31,225,31,94,31,94,30,63,31,49,31,49,30,59,31,229,31,70,31,70,30,70,29,246,31,246,30,127,31,251,31,104,31,174,31,158,31,178,31,233,31,140,31,45,31,157,31,202,31,148,31,253,31,167,31,54,31,204,31,142,31,74,31,129,31,129,30,223,31,157,31,193,31,193,30,70,31,216,31,72,31,49,31,49,30,49,29,164,31,188,31,96,31,34,31,84,31,84,30,39,31,60,31,180,31,213,31,213,30,213,29,236,31,15,31,41,31,39,31,221,31,66,31,220,31,220,30,115,31,200,31,2,31,16,31,49,31,130,31,130,30,130,29,130,28,20,31,20,30,147,31,147,30,161,31,59,31,151,31,65,31,65,30,229,31,229,30,250,31,101,31,101,30,73,31,46,31,40,31,26,31,226,31,56,31,100,31,100,30,58,31,166,31,11,31,218,31,85,31,213,31,213,30,133,31,15,31,178,31,96,31,135,31,35,31,233,31,3,31,93,31,209,31,52,31,52,30,131,31,239,31,239,30,239,29,148,31,248,31,78,31,96,31,120,31,218,31,244,31,244,30,92,31,38,31,38,30,250,31,250,30,36,31,175,31,175,30,184,31,49,31,11,31,242,31,148,31,233,31,246,31,197,31,96,31,161,31,227,31,196,31,155,31,162,31,162,31,224,31,219,31,120,31,120,30,120,29,104,31,127,31,127,30,127,29,127,28,224,31,158,31,22,31,224,31,28,31,28,30,94,31,164,31,170,31,117,31,228,31,228,30,181,31,14,31,142,31,16,31,16,30,170,31,203,31,224,31,224,30,145,31,175,31,7,31,121,31,96,31,140,31,140,30,54,31,83,31,195,31,195,30,192,31,40,31,189,31,50,31,70,31,70,30,248,31,156,31,141,31,182,31,204,31,235,31,250,31,250,30,117,31,255,31,255,30,180,31,64,31,64,30,100,31,10,31,156,31,67,31,197,31,79,31,79,30,129,31,149,31,34,31,155,31,127,31,127,30,126,31,209,31,242,31,242,30,144,31,226,31,23,31,87,31,68,31,213,31,10,31,97,31,247,31,14,31,60,31,60,30,204,31,67,31,137,31,135,31,148,31,204,31,204,30,204,29,204,28,3,31,90,31,90,30,209,31,131,31,244,31,181,31,159,31,224,31,89,31,89,30,169,31,83,31,83,30,210,31,255,31,255,30,139,31,243,31,108,31,228,31,164,31,215,31,5,31,5,30,233,31,233,30,84,31,84,30,176,31,176,30,48,31,165,31,249,31,111,31,98,31,98,30,60,31,203,31,203,30,63,31,59,31,144,31,144,30,84,31,148,31,148,30,114,31,201,31,70,31,177,31,95,31,128,31,3,31,209,31,79,31,79,30,2,31,241,31,131,31,230,31,97,31,119,31,158,31,108,31,240,31,240,30,221,31,49,31,49,30,122,31,171,31,165,31,121,31,121,30,121,29,121,28,121,27,121,26,75,31,105,31,105,30,105,29,180,31,117,31,117,30,131,31,161,31,166,31,201,31,235,31,125,31,207,31,226,31,203,31,203,30,203,29,142,31,142,30,30,31,44,31,46,31,46,30,142,31,234,31,23,31,23,30,134,31,127,31,165,31,194,31,55,31,114,31,158,31,68,31,26,31,210,31,81,31,107,31,89,31,154,31,12,31,131,31,212,31,158,31,158,30,65,31,13,31,83,31,85,31,189,31,187,31,82,31,125,31,178,31,191,31,106,31,7,31,140,31,140,30,184,31,135,31,184,31,42,31,40,31,241,31,241,30,248,31,233,31,63,31,63,30,198,31,246,31,164,31,84,31,84,31,23,31,41,31,124,31,124,30,154,31,34,31,34,30,219,31,138,31,166,31,95,31,95,30,246,31,143,31,234,31,58,31,32,31,32,30,150,31,114,31,189,31,6,31,35,31,35,30,176,31,176,30,154,31,157,31,133,31,151,31,151,30,151,29,100,31,15,31,38,31,147,31,206,31,66,31,143,31,128,31,3,31,214,31,85,31,85,30,30,31,222,31,13,31,66,31,163,31,96,31,224,31,224,30,126,31,134,31,235,31,151,31,35,31,165,31,135,31,191,31,120,31,120,30,131,31,151,31,99,31,26,31,179,31,107,31,107,30,85,31,204,31,204,30,103,31,10,31,237,31,95,31,68,31,2,31,14,31,23,31,137,31,137,30,28,31,249,31,171,31,1,31,23,31,23,30,154,31,205,31,184,31,184,30,115,31,76,31,67,31,207,31,166,31,166,30,166,29,238,31,105,31,45,31,46,31,146,31,233,31,207,31,125,31,226,31,199,31,199,30,95,31,81,31,65,31,22,31,222,31,142,31,142,30,142,29,177,31,77,31,172,31,64,31,252,31,252,30,57,31,112,31,16,31,235,31,166,31,241,31,237,31,185,31,218,31,25,31,241,31,22,31,229,31,229,30,125,31,231,31,100,31,1,31,1,30,116,31,76,31,76,30,216,31,216,30,131,31,201,31,201,30,2,31,174,31,174,30,240,31,188,31,81,31,81,30,31,31,152,31,147,31,146,31,140,31,82,31,245,31,245,30,245,29,188,31,188,30,188,29,35,31,35,30,228,31,154,31,158,31,77,31,226,31,226,30,183,31,243,31,125,31,26,31,124,31,53,31,48,31,206,31,55,31,65,31,21,31,166,31,186,31,159,31,159,30,159,29,119,31,59,31,61,31,198,31,38,31,51,31,62,31,93,31,24,31,248,31,113,31,113,30,219,31,170,31,170,30,123,31,123,30,232,31,32,31,22,31,30,31,52,31,52,30,205,31,13,31,103,31,255,31,192,31,32,31,190,31,105,31,9,31,30,31,68,31,143,31,19,31,19,30,247,31,160,31,81,31,81,30,236,31,146,31,222,31,75,31,106,31,152,31,144,31,144,30,60,31,64,31,44,31,228,31,228,30,95,31,244,31,143,31,50,31,120,31,107,31,4,31,4,30,107,31,4,31,29,31,61,31,253,31,123,31,132,31,60,31,9,31,94,31,94,30,121,31,183,31,183,30,155,31,87,31,147,31,207,31,62,31,248,31,144,31,144,30,144,29,115,31,248,31,7,31,15,31,160,31,39,31,8,31,165,31,82,31,142,31,147,31,118,31,12,31,12,30,48,31,48,30,128,31,182,31,97,31,97,30,237,31,7,31,19,31,15,31,15,30,15,29,109,31,121,31,136,31,130,31,158,31,158,30,67,31,86,31,156,31,150,31,177,31,177,30,57,31,115,31,115,30,179,31,90,31,58,31,239,31,239,30,126,31,232,31,232,30,17,31,21,31,74,31,37,31,36,31,36,30,22,31,20,31,232,31,181,31,31,31,230,31,140,31,3,31,189,31,96,31,18,31,92,31,106,31,200,31,1,31,1,30,103,31,127,31,127,30,127,29,174,31,241,31,137,31,246,31,171,31,144,31,36,31,53,31,153,31,50,31,142,31,142,30,143,31,143,30,48,31,63,31,95,31,16,31,16,30,167,31,89,31,30,31,37,31,22,31,22,30,222,31,243,31,11,31,66,31,66,30,66,29,127,31,97,31,89,31,36,31,109,31,109,30,109,29,109,28,109,27,130,31,168,31,168,30,119,31,138,31,34,31,247,31,174,31,113,31,184,31,106,31,187,31,199,31,199,30,251,31,174,31,120,31,120,30,35,31,205,31,173,31,77,31,140,31,207,31,37,31,37,30,70,31,114,31,167,31,167,30,169,31,66,31,55,31,153,31,18,31,75,31,86,31,165,31,183,31,183,30,223,31,245,31,187,31,51,31,70,31,70,30,140,31,222,31,222,30,165,31,32,31,164,31,164,30,164,29,164,28,196,31,196,30,235,31,207,31,207,30,99,31,122,31,110,31,110,30,236,31,63,31,151,31,95,31,231,31,6,31,220,31,34,31,159,31,159,30,189,31,48,31,114,31,111,31,88,31,111,31,111,30,111,29,31,31,205,31,205,30,238,31,71,31,71,30,194,31,149,31,235,31,235,30,119,31,144,31,124,31,40,31,193,31,143,31,143,30,40,31,255,31,218,31,62,31,195,31,43,31,168,31,187,31,184,31,254,31,50,31,50,30,238,31,186,31,245,31,245,30,22,31,22,30,1,31,197,31,92,31,33,31,33,30,33,29,125,31,125,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
