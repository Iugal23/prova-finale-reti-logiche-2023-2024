-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 276;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,155,0,62,0,0,0,195,0,180,0,134,0,127,0,75,0,7,0,231,0,87,0,137,0,255,0,60,0,169,0,52,0,191,0,85,0,65,0,199,0,0,0,42,0,121,0,41,0,216,0,55,0,35,0,223,0,36,0,0,0,0,0,88,0,242,0,237,0,212,0,42,0,11,0,198,0,208,0,236,0,31,0,134,0,52,0,180,0,188,0,0,0,242,0,217,0,0,0,203,0,220,0,0,0,105,0,0,0,206,0,213,0,0,0,187,0,0,0,194,0,0,0,0,0,65,0,0,0,156,0,135,0,36,0,0,0,54,0,223,0,191,0,207,0,155,0,0,0,0,0,0,0,219,0,227,0,79,0,92,0,18,0,0,0,235,0,166,0,150,0,110,0,248,0,62,0,213,0,14,0,19,0,134,0,0,0,252,0,133,0,0,0,60,0,77,0,19,0,61,0,111,0,238,0,0,0,199,0,252,0,111,0,202,0,204,0,88,0,0,0,155,0,164,0,219,0,16,0,80,0,243,0,132,0,0,0,158,0,100,0,44,0,42,0,204,0,191,0,215,0,209,0,137,0,30,0,112,0,133,0,156,0,0,0,21,0,87,0,98,0,17,0,187,0,76,0,0,0,241,0,0,0,140,0,51,0,136,0,57,0,223,0,0,0,91,0,214,0,14,0,118,0,189,0,0,0,240,0,37,0,130,0,20,0,25,0,34,0,175,0,110,0,0,0,0,0,203,0,0,0,246,0,0,0,0,0,8,0,144,0,147,0,166,0,0,0,122,0,44,0,168,0,29,0,0,0,0,0,243,0,113,0,83,0,0,0,248,0,231,0,0,0,0,0,158,0,0,0,0,0,32,0,86,0,80,0,39,0,254,0,0,0,251,0,77,0,0,0,57,0,1,0,0,0,84,0,71,0,0,0,217,0,59,0,24,0,176,0,151,0,108,0,0,0,142,0,0,0,0,0,247,0,147,0,242,0,98,0,26,0,55,0,208,0,237,0,0,0,177,0,185,0,74,0,69,0,187,0,71,0,96,0,171,0,202,0,110,0,56,0,241,0,40,0,1,0,33,0,62,0,0,0,33,0,30,0,188,0,102,0,33,0,80,0,119,0,43,0,139,0,149,0,0,0,119,0,44,0,0,0,67,0,238,0,198,0,0,0,189,0,81,0,172,0,75,0,0,0,51,0,177,0,230,0,146,0,22,0,12,0,16,0,223,0,252,0,72,0,194,0);
signal scenario_full  : scenario_type := (0,0,155,31,62,31,62,30,195,31,180,31,134,31,127,31,75,31,7,31,231,31,87,31,137,31,255,31,60,31,169,31,52,31,191,31,85,31,65,31,199,31,199,30,42,31,121,31,41,31,216,31,55,31,35,31,223,31,36,31,36,30,36,29,88,31,242,31,237,31,212,31,42,31,11,31,198,31,208,31,236,31,31,31,134,31,52,31,180,31,188,31,188,30,242,31,217,31,217,30,203,31,220,31,220,30,105,31,105,30,206,31,213,31,213,30,187,31,187,30,194,31,194,30,194,29,65,31,65,30,156,31,135,31,36,31,36,30,54,31,223,31,191,31,207,31,155,31,155,30,155,29,155,28,219,31,227,31,79,31,92,31,18,31,18,30,235,31,166,31,150,31,110,31,248,31,62,31,213,31,14,31,19,31,134,31,134,30,252,31,133,31,133,30,60,31,77,31,19,31,61,31,111,31,238,31,238,30,199,31,252,31,111,31,202,31,204,31,88,31,88,30,155,31,164,31,219,31,16,31,80,31,243,31,132,31,132,30,158,31,100,31,44,31,42,31,204,31,191,31,215,31,209,31,137,31,30,31,112,31,133,31,156,31,156,30,21,31,87,31,98,31,17,31,187,31,76,31,76,30,241,31,241,30,140,31,51,31,136,31,57,31,223,31,223,30,91,31,214,31,14,31,118,31,189,31,189,30,240,31,37,31,130,31,20,31,25,31,34,31,175,31,110,31,110,30,110,29,203,31,203,30,246,31,246,30,246,29,8,31,144,31,147,31,166,31,166,30,122,31,44,31,168,31,29,31,29,30,29,29,243,31,113,31,83,31,83,30,248,31,231,31,231,30,231,29,158,31,158,30,158,29,32,31,86,31,80,31,39,31,254,31,254,30,251,31,77,31,77,30,57,31,1,31,1,30,84,31,71,31,71,30,217,31,59,31,24,31,176,31,151,31,108,31,108,30,142,31,142,30,142,29,247,31,147,31,242,31,98,31,26,31,55,31,208,31,237,31,237,30,177,31,185,31,74,31,69,31,187,31,71,31,96,31,171,31,202,31,110,31,56,31,241,31,40,31,1,31,33,31,62,31,62,30,33,31,30,31,188,31,102,31,33,31,80,31,119,31,43,31,139,31,149,31,149,30,119,31,44,31,44,30,67,31,238,31,198,31,198,30,189,31,81,31,172,31,75,31,75,30,51,31,177,31,230,31,146,31,22,31,12,31,16,31,223,31,252,31,72,31,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
