-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_622 is
end project_tb_622;

architecture project_tb_arch_622 of project_tb_622 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 814;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,199,0,26,0,239,0,0,0,0,0,57,0,241,0,34,0,73,0,84,0,188,0,0,0,76,0,131,0,193,0,120,0,0,0,103,0,26,0,255,0,13,0,105,0,149,0,69,0,118,0,8,0,172,0,101,0,179,0,62,0,181,0,0,0,98,0,91,0,0,0,0,0,123,0,0,0,0,0,0,0,0,0,0,0,199,0,59,0,96,0,92,0,225,0,200,0,203,0,102,0,16,0,148,0,158,0,143,0,182,0,218,0,73,0,97,0,0,0,0,0,194,0,58,0,8,0,223,0,0,0,119,0,0,0,121,0,37,0,0,0,0,0,225,0,159,0,128,0,0,0,233,0,117,0,0,0,41,0,104,0,132,0,0,0,245,0,32,0,116,0,102,0,97,0,163,0,102,0,179,0,215,0,0,0,165,0,184,0,0,0,38,0,149,0,72,0,198,0,0,0,144,0,0,0,9,0,124,0,2,0,86,0,61,0,57,0,7,0,144,0,247,0,175,0,0,0,168,0,45,0,0,0,0,0,148,0,185,0,247,0,91,0,0,0,142,0,158,0,202,0,235,0,0,0,165,0,84,0,63,0,41,0,20,0,192,0,0,0,197,0,8,0,44,0,5,0,26,0,0,0,87,0,0,0,97,0,97,0,0,0,190,0,245,0,0,0,21,0,82,0,236,0,29,0,147,0,238,0,77,0,23,0,32,0,0,0,193,0,66,0,0,0,144,0,195,0,149,0,201,0,242,0,55,0,0,0,0,0,185,0,46,0,253,0,73,0,0,0,155,0,100,0,215,0,98,0,152,0,177,0,175,0,178,0,11,0,233,0,218,0,58,0,20,0,77,0,245,0,210,0,231,0,59,0,54,0,203,0,103,0,148,0,154,0,0,0,183,0,250,0,130,0,159,0,0,0,169,0,0,0,99,0,61,0,9,0,0,0,23,0,128,0,0,0,215,0,74,0,14,0,0,0,0,0,0,0,6,0,71,0,117,0,152,0,0,0,62,0,197,0,125,0,66,0,0,0,0,0,39,0,157,0,83,0,33,0,0,0,240,0,0,0,138,0,42,0,177,0,163,0,233,0,86,0,88,0,213,0,145,0,0,0,187,0,42,0,200,0,68,0,45,0,110,0,144,0,59,0,0,0,187,0,45,0,50,0,50,0,49,0,0,0,198,0,127,0,122,0,184,0,182,0,246,0,189,0,229,0,25,0,41,0,0,0,126,0,35,0,212,0,0,0,73,0,180,0,162,0,120,0,96,0,248,0,220,0,0,0,0,0,193,0,167,0,147,0,247,0,25,0,5,0,84,0,0,0,45,0,84,0,122,0,109,0,61,0,95,0,9,0,23,0,79,0,14,0,157,0,236,0,0,0,156,0,0,0,0,0,82,0,102,0,0,0,84,0,176,0,228,0,18,0,61,0,233,0,128,0,220,0,54,0,0,0,0,0,46,0,43,0,75,0,0,0,168,0,247,0,0,0,54,0,89,0,21,0,255,0,0,0,166,0,213,0,0,0,39,0,171,0,149,0,16,0,0,0,218,0,107,0,90,0,164,0,178,0,0,0,35,0,133,0,11,0,58,0,0,0,241,0,211,0,116,0,203,0,23,0,0,0,144,0,83,0,44,0,118,0,2,0,82,0,218,0,0,0,157,0,123,0,103,0,59,0,44,0,195,0,54,0,227,0,51,0,141,0,0,0,61,0,30,0,60,0,212,0,113,0,109,0,2,0,87,0,194,0,133,0,0,0,132,0,198,0,0,0,83,0,145,0,142,0,166,0,6,0,0,0,42,0,105,0,193,0,171,0,0,0,218,0,182,0,78,0,56,0,186,0,0,0,0,0,184,0,98,0,244,0,165,0,28,0,208,0,0,0,181,0,0,0,88,0,192,0,67,0,80,0,93,0,0,0,0,0,218,0,240,0,88,0,234,0,74,0,0,0,73,0,153,0,160,0,22,0,255,0,138,0,116,0,0,0,98,0,252,0,166,0,225,0,255,0,242,0,124,0,85,0,202,0,20,0,174,0,58,0,55,0,228,0,0,0,207,0,173,0,122,0,113,0,0,0,191,0,89,0,47,0,85,0,141,0,0,0,155,0,0,0,0,0,182,0,143,0,178,0,85,0,119,0,140,0,196,0,141,0,18,0,139,0,222,0,235,0,168,0,132,0,204,0,244,0,64,0,128,0,101,0,47,0,75,0,225,0,204,0,0,0,190,0,0,0,125,0,145,0,0,0,159,0,224,0,0,0,152,0,0,0,159,0,0,0,0,0,31,0,61,0,0,0,141,0,219,0,0,0,30,0,0,0,108,0,169,0,27,0,179,0,86,0,0,0,0,0,0,0,0,0,81,0,0,0,238,0,174,0,52,0,0,0,229,0,19,0,190,0,0,0,187,0,149,0,187,0,145,0,209,0,23,0,0,0,164,0,34,0,247,0,0,0,0,0,125,0,11,0,82,0,133,0,209,0,0,0,92,0,228,0,8,0,35,0,0,0,205,0,147,0,138,0,0,0,0,0,130,0,91,0,83,0,146,0,249,0,190,0,80,0,68,0,67,0,61,0,238,0,19,0,0,0,98,0,25,0,58,0,114,0,0,0,135,0,17,0,0,0,109,0,231,0,54,0,122,0,114,0,0,0,50,0,201,0,95,0,167,0,208,0,0,0,137,0,238,0,228,0,0,0,230,0,90,0,73,0,42,0,157,0,102,0,235,0,166,0,0,0,0,0,91,0,245,0,96,0,44,0,228,0,238,0,0,0,112,0,205,0,247,0,98,0,0,0,6,0,0,0,0,0,202,0,110,0,178,0,243,0,221,0,115,0,182,0,215,0,217,0,72,0,197,0,144,0,66,0,37,0,111,0,161,0,113,0,166,0,246,0,203,0,0,0,0,0,57,0,183,0,71,0,146,0,0,0,163,0,0,0,45,0,254,0,34,0,126,0,226,0,0,0,166,0,86,0,73,0,6,0,103,0,120,0,169,0,0,0,205,0,167,0,124,0,0,0,158,0,0,0,0,0,167,0,51,0,0,0,0,0,219,0,0,0,89,0,37,0,15,0,50,0,0,0,155,0,132,0,0,0,21,0,124,0,183,0,104,0,74,0,3,0,0,0,106,0,250,0,109,0,91,0,0,0,0,0,0,0,203,0,182,0,113,0,191,0,0,0,5,0,212,0,35,0,0,0,205,0,0,0,121,0,0,0,133,0,58,0,214,0,212,0,0,0,0,0,174,0,33,0,11,0,172,0,47,0,31,0,13,0,123,0,2,0,0,0,0,0,0,0,124,0,0,0,244,0,31,0,69,0,197,0,112,0,0,0,199,0,27,0,83,0,136,0,52,0,28,0,0,0,160,0,0,0,232,0,218,0,0,0,39,0,102,0,88,0,206,0,88,0,206,0,0,0,165,0,225,0,125,0,83,0,62,0,228,0,77,0,20,0,148,0,233,0,153,0,67,0,16,0,27,0,37,0,27,0,0,0,179,0,161,0,87,0,168,0,238,0,105,0,76,0,183,0,148,0,45,0,133,0,29,0,20,0,227,0,208,0,0,0,0,0,0,0,59,0,6,0,124,0,170,0,120,0,0,0,96,0,80,0,143,0,212,0,98,0,0,0,243,0,207,0,243,0,118,0,0,0,154,0);
signal scenario_full  : scenario_type := (169,31,199,31,26,31,239,31,239,30,239,29,57,31,241,31,34,31,73,31,84,31,188,31,188,30,76,31,131,31,193,31,120,31,120,30,103,31,26,31,255,31,13,31,105,31,149,31,69,31,118,31,8,31,172,31,101,31,179,31,62,31,181,31,181,30,98,31,91,31,91,30,91,29,123,31,123,30,123,29,123,28,123,27,123,26,199,31,59,31,96,31,92,31,225,31,200,31,203,31,102,31,16,31,148,31,158,31,143,31,182,31,218,31,73,31,97,31,97,30,97,29,194,31,58,31,8,31,223,31,223,30,119,31,119,30,121,31,37,31,37,30,37,29,225,31,159,31,128,31,128,30,233,31,117,31,117,30,41,31,104,31,132,31,132,30,245,31,32,31,116,31,102,31,97,31,163,31,102,31,179,31,215,31,215,30,165,31,184,31,184,30,38,31,149,31,72,31,198,31,198,30,144,31,144,30,9,31,124,31,2,31,86,31,61,31,57,31,7,31,144,31,247,31,175,31,175,30,168,31,45,31,45,30,45,29,148,31,185,31,247,31,91,31,91,30,142,31,158,31,202,31,235,31,235,30,165,31,84,31,63,31,41,31,20,31,192,31,192,30,197,31,8,31,44,31,5,31,26,31,26,30,87,31,87,30,97,31,97,31,97,30,190,31,245,31,245,30,21,31,82,31,236,31,29,31,147,31,238,31,77,31,23,31,32,31,32,30,193,31,66,31,66,30,144,31,195,31,149,31,201,31,242,31,55,31,55,30,55,29,185,31,46,31,253,31,73,31,73,30,155,31,100,31,215,31,98,31,152,31,177,31,175,31,178,31,11,31,233,31,218,31,58,31,20,31,77,31,245,31,210,31,231,31,59,31,54,31,203,31,103,31,148,31,154,31,154,30,183,31,250,31,130,31,159,31,159,30,169,31,169,30,99,31,61,31,9,31,9,30,23,31,128,31,128,30,215,31,74,31,14,31,14,30,14,29,14,28,6,31,71,31,117,31,152,31,152,30,62,31,197,31,125,31,66,31,66,30,66,29,39,31,157,31,83,31,33,31,33,30,240,31,240,30,138,31,42,31,177,31,163,31,233,31,86,31,88,31,213,31,145,31,145,30,187,31,42,31,200,31,68,31,45,31,110,31,144,31,59,31,59,30,187,31,45,31,50,31,50,31,49,31,49,30,198,31,127,31,122,31,184,31,182,31,246,31,189,31,229,31,25,31,41,31,41,30,126,31,35,31,212,31,212,30,73,31,180,31,162,31,120,31,96,31,248,31,220,31,220,30,220,29,193,31,167,31,147,31,247,31,25,31,5,31,84,31,84,30,45,31,84,31,122,31,109,31,61,31,95,31,9,31,23,31,79,31,14,31,157,31,236,31,236,30,156,31,156,30,156,29,82,31,102,31,102,30,84,31,176,31,228,31,18,31,61,31,233,31,128,31,220,31,54,31,54,30,54,29,46,31,43,31,75,31,75,30,168,31,247,31,247,30,54,31,89,31,21,31,255,31,255,30,166,31,213,31,213,30,39,31,171,31,149,31,16,31,16,30,218,31,107,31,90,31,164,31,178,31,178,30,35,31,133,31,11,31,58,31,58,30,241,31,211,31,116,31,203,31,23,31,23,30,144,31,83,31,44,31,118,31,2,31,82,31,218,31,218,30,157,31,123,31,103,31,59,31,44,31,195,31,54,31,227,31,51,31,141,31,141,30,61,31,30,31,60,31,212,31,113,31,109,31,2,31,87,31,194,31,133,31,133,30,132,31,198,31,198,30,83,31,145,31,142,31,166,31,6,31,6,30,42,31,105,31,193,31,171,31,171,30,218,31,182,31,78,31,56,31,186,31,186,30,186,29,184,31,98,31,244,31,165,31,28,31,208,31,208,30,181,31,181,30,88,31,192,31,67,31,80,31,93,31,93,30,93,29,218,31,240,31,88,31,234,31,74,31,74,30,73,31,153,31,160,31,22,31,255,31,138,31,116,31,116,30,98,31,252,31,166,31,225,31,255,31,242,31,124,31,85,31,202,31,20,31,174,31,58,31,55,31,228,31,228,30,207,31,173,31,122,31,113,31,113,30,191,31,89,31,47,31,85,31,141,31,141,30,155,31,155,30,155,29,182,31,143,31,178,31,85,31,119,31,140,31,196,31,141,31,18,31,139,31,222,31,235,31,168,31,132,31,204,31,244,31,64,31,128,31,101,31,47,31,75,31,225,31,204,31,204,30,190,31,190,30,125,31,145,31,145,30,159,31,224,31,224,30,152,31,152,30,159,31,159,30,159,29,31,31,61,31,61,30,141,31,219,31,219,30,30,31,30,30,108,31,169,31,27,31,179,31,86,31,86,30,86,29,86,28,86,27,81,31,81,30,238,31,174,31,52,31,52,30,229,31,19,31,190,31,190,30,187,31,149,31,187,31,145,31,209,31,23,31,23,30,164,31,34,31,247,31,247,30,247,29,125,31,11,31,82,31,133,31,209,31,209,30,92,31,228,31,8,31,35,31,35,30,205,31,147,31,138,31,138,30,138,29,130,31,91,31,83,31,146,31,249,31,190,31,80,31,68,31,67,31,61,31,238,31,19,31,19,30,98,31,25,31,58,31,114,31,114,30,135,31,17,31,17,30,109,31,231,31,54,31,122,31,114,31,114,30,50,31,201,31,95,31,167,31,208,31,208,30,137,31,238,31,228,31,228,30,230,31,90,31,73,31,42,31,157,31,102,31,235,31,166,31,166,30,166,29,91,31,245,31,96,31,44,31,228,31,238,31,238,30,112,31,205,31,247,31,98,31,98,30,6,31,6,30,6,29,202,31,110,31,178,31,243,31,221,31,115,31,182,31,215,31,217,31,72,31,197,31,144,31,66,31,37,31,111,31,161,31,113,31,166,31,246,31,203,31,203,30,203,29,57,31,183,31,71,31,146,31,146,30,163,31,163,30,45,31,254,31,34,31,126,31,226,31,226,30,166,31,86,31,73,31,6,31,103,31,120,31,169,31,169,30,205,31,167,31,124,31,124,30,158,31,158,30,158,29,167,31,51,31,51,30,51,29,219,31,219,30,89,31,37,31,15,31,50,31,50,30,155,31,132,31,132,30,21,31,124,31,183,31,104,31,74,31,3,31,3,30,106,31,250,31,109,31,91,31,91,30,91,29,91,28,203,31,182,31,113,31,191,31,191,30,5,31,212,31,35,31,35,30,205,31,205,30,121,31,121,30,133,31,58,31,214,31,212,31,212,30,212,29,174,31,33,31,11,31,172,31,47,31,31,31,13,31,123,31,2,31,2,30,2,29,2,28,124,31,124,30,244,31,31,31,69,31,197,31,112,31,112,30,199,31,27,31,83,31,136,31,52,31,28,31,28,30,160,31,160,30,232,31,218,31,218,30,39,31,102,31,88,31,206,31,88,31,206,31,206,30,165,31,225,31,125,31,83,31,62,31,228,31,77,31,20,31,148,31,233,31,153,31,67,31,16,31,27,31,37,31,27,31,27,30,179,31,161,31,87,31,168,31,238,31,105,31,76,31,183,31,148,31,45,31,133,31,29,31,20,31,227,31,208,31,208,30,208,29,208,28,59,31,6,31,124,31,170,31,120,31,120,30,96,31,80,31,143,31,212,31,98,31,98,30,243,31,207,31,243,31,118,31,118,30,154,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
