-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_459 is
end project_tb_459;

architecture project_tb_arch_459 of project_tb_459 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 190;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (150,0,0,0,120,0,31,0,252,0,166,0,71,0,245,0,219,0,0,0,0,0,118,0,0,0,249,0,136,0,0,0,61,0,148,0,201,0,225,0,17,0,13,0,235,0,0,0,0,0,51,0,198,0,141,0,196,0,0,0,0,0,229,0,219,0,173,0,0,0,167,0,247,0,0,0,0,0,113,0,140,0,0,0,76,0,0,0,77,0,187,0,219,0,0,0,107,0,200,0,116,0,0,0,12,0,54,0,252,0,0,0,176,0,169,0,212,0,14,0,94,0,47,0,84,0,102,0,242,0,0,0,0,0,221,0,24,0,240,0,0,0,4,0,3,0,0,0,137,0,45,0,0,0,0,0,125,0,217,0,3,0,77,0,0,0,64,0,106,0,80,0,224,0,238,0,88,0,115,0,102,0,165,0,200,0,164,0,0,0,234,0,155,0,62,0,122,0,155,0,58,0,210,0,0,0,114,0,220,0,196,0,0,0,137,0,29,0,102,0,119,0,0,0,230,0,74,0,255,0,221,0,0,0,26,0,117,0,59,0,220,0,83,0,191,0,237,0,211,0,233,0,177,0,225,0,249,0,0,0,137,0,14,0,145,0,204,0,186,0,0,0,151,0,162,0,127,0,243,0,0,0,93,0,0,0,158,0,71,0,6,0,196,0,106,0,150,0,254,0,31,0,13,0,1,0,159,0,46,0,98,0,110,0,180,0,208,0,0,0,241,0,143,0,127,0,191,0,0,0,0,0,110,0,0,0,104,0,16,0,230,0,54,0,204,0,0,0,0,0,173,0,151,0,115,0,0,0,0,0,0,0,38,0,144,0,110,0,6,0,218,0,190,0,253,0,109,0,0,0);
signal scenario_full  : scenario_type := (150,31,150,30,120,31,31,31,252,31,166,31,71,31,245,31,219,31,219,30,219,29,118,31,118,30,249,31,136,31,136,30,61,31,148,31,201,31,225,31,17,31,13,31,235,31,235,30,235,29,51,31,198,31,141,31,196,31,196,30,196,29,229,31,219,31,173,31,173,30,167,31,247,31,247,30,247,29,113,31,140,31,140,30,76,31,76,30,77,31,187,31,219,31,219,30,107,31,200,31,116,31,116,30,12,31,54,31,252,31,252,30,176,31,169,31,212,31,14,31,94,31,47,31,84,31,102,31,242,31,242,30,242,29,221,31,24,31,240,31,240,30,4,31,3,31,3,30,137,31,45,31,45,30,45,29,125,31,217,31,3,31,77,31,77,30,64,31,106,31,80,31,224,31,238,31,88,31,115,31,102,31,165,31,200,31,164,31,164,30,234,31,155,31,62,31,122,31,155,31,58,31,210,31,210,30,114,31,220,31,196,31,196,30,137,31,29,31,102,31,119,31,119,30,230,31,74,31,255,31,221,31,221,30,26,31,117,31,59,31,220,31,83,31,191,31,237,31,211,31,233,31,177,31,225,31,249,31,249,30,137,31,14,31,145,31,204,31,186,31,186,30,151,31,162,31,127,31,243,31,243,30,93,31,93,30,158,31,71,31,6,31,196,31,106,31,150,31,254,31,31,31,13,31,1,31,159,31,46,31,98,31,110,31,180,31,208,31,208,30,241,31,143,31,127,31,191,31,191,30,191,29,110,31,110,30,104,31,16,31,230,31,54,31,204,31,204,30,204,29,173,31,151,31,115,31,115,30,115,29,115,28,38,31,144,31,110,31,6,31,218,31,190,31,253,31,109,31,109,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
