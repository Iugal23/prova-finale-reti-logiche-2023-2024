-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 824;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (234,0,191,0,38,0,88,0,107,0,181,0,166,0,130,0,29,0,0,0,0,0,65,0,246,0,0,0,126,0,123,0,31,0,223,0,150,0,121,0,49,0,0,0,96,0,0,0,233,0,134,0,63,0,0,0,14,0,170,0,142,0,96,0,91,0,138,0,93,0,121,0,0,0,112,0,0,0,224,0,254,0,0,0,153,0,58,0,74,0,221,0,28,0,0,0,138,0,191,0,135,0,0,0,138,0,195,0,94,0,75,0,0,0,0,0,95,0,173,0,54,0,10,0,5,0,87,0,0,0,112,0,100,0,230,0,139,0,180,0,180,0,237,0,0,0,0,0,33,0,168,0,255,0,0,0,26,0,0,0,216,0,244,0,105,0,210,0,119,0,0,0,23,0,124,0,0,0,54,0,108,0,5,0,94,0,176,0,104,0,62,0,106,0,28,0,251,0,30,0,0,0,78,0,111,0,12,0,121,0,76,0,131,0,117,0,101,0,16,0,25,0,237,0,0,0,231,0,251,0,205,0,17,0,238,0,182,0,183,0,209,0,206,0,144,0,15,0,0,0,33,0,0,0,144,0,0,0,166,0,22,0,31,0,255,0,243,0,42,0,253,0,0,0,16,0,212,0,190,0,29,0,204,0,23,0,0,0,239,0,226,0,48,0,230,0,160,0,99,0,193,0,149,0,44,0,6,0,135,0,0,0,129,0,0,0,203,0,106,0,111,0,127,0,223,0,0,0,188,0,0,0,31,0,30,0,16,0,35,0,0,0,248,0,0,0,40,0,82,0,0,0,49,0,0,0,91,0,175,0,251,0,0,0,34,0,0,0,123,0,43,0,180,0,130,0,47,0,0,0,97,0,160,0,143,0,230,0,0,0,72,0,201,0,126,0,137,0,15,0,241,0,31,0,39,0,91,0,89,0,82,0,142,0,240,0,0,0,149,0,74,0,105,0,0,0,0,0,241,0,254,0,121,0,0,0,223,0,207,0,42,0,17,0,0,0,34,0,78,0,101,0,194,0,105,0,0,0,36,0,78,0,45,0,200,0,61,0,162,0,110,0,143,0,232,0,176,0,0,0,11,0,100,0,79,0,0,0,32,0,177,0,131,0,255,0,162,0,88,0,90,0,186,0,94,0,36,0,179,0,0,0,179,0,96,0,1,0,0,0,0,0,16,0,0,0,106,0,0,0,47,0,153,0,181,0,94,0,0,0,244,0,176,0,0,0,153,0,75,0,249,0,249,0,0,0,172,0,223,0,64,0,128,0,117,0,0,0,105,0,45,0,171,0,0,0,14,0,22,0,0,0,201,0,198,0,20,0,69,0,43,0,230,0,55,0,83,0,237,0,224,0,88,0,86,0,206,0,213,0,163,0,123,0,100,0,124,0,158,0,168,0,101,0,170,0,188,0,212,0,188,0,0,0,0,0,0,0,21,0,0,0,9,0,0,0,0,0,104,0,86,0,0,0,170,0,43,0,156,0,54,0,151,0,0,0,69,0,17,0,0,0,194,0,50,0,163,0,0,0,79,0,188,0,20,0,114,0,210,0,209,0,203,0,14,0,104,0,150,0,52,0,72,0,16,0,26,0,0,0,152,0,0,0,3,0,239,0,178,0,128,0,1,0,0,0,0,0,177,0,128,0,8,0,58,0,0,0,66,0,224,0,46,0,173,0,94,0,86,0,48,0,179,0,79,0,206,0,75,0,0,0,112,0,9,0,200,0,85,0,0,0,0,0,0,0,128,0,0,0,77,0,157,0,0,0,0,0,16,0,68,0,15,0,0,0,187,0,225,0,94,0,103,0,124,0,209,0,0,0,179,0,58,0,129,0,0,0,108,0,21,0,15,0,243,0,0,0,216,0,99,0,210,0,159,0,36,0,204,0,42,0,135,0,96,0,142,0,10,0,0,0,0,0,140,0,58,0,155,0,115,0,226,0,204,0,140,0,244,0,162,0,214,0,8,0,222,0,212,0,106,0,102,0,18,0,65,0,204,0,98,0,215,0,0,0,36,0,154,0,0,0,230,0,49,0,0,0,10,0,0,0,108,0,215,0,212,0,95,0,182,0,154,0,5,0,251,0,0,0,165,0,41,0,232,0,0,0,241,0,49,0,173,0,112,0,51,0,0,0,72,0,60,0,0,0,191,0,85,0,0,0,3,0,8,0,161,0,30,0,153,0,19,0,151,0,140,0,0,0,155,0,215,0,199,0,0,0,167,0,55,0,43,0,115,0,140,0,0,0,78,0,0,0,0,0,165,0,98,0,207,0,103,0,83,0,153,0,23,0,46,0,214,0,186,0,185,0,160,0,17,0,112,0,145,0,41,0,156,0,0,0,0,0,97,0,0,0,118,0,131,0,0,0,101,0,192,0,42,0,0,0,37,0,0,0,194,0,58,0,76,0,194,0,247,0,71,0,219,0,75,0,205,0,66,0,149,0,201,0,80,0,100,0,157,0,6,0,175,0,237,0,171,0,51,0,41,0,177,0,192,0,168,0,137,0,97,0,0,0,187,0,247,0,218,0,137,0,0,0,38,0,0,0,208,0,34,0,44,0,147,0,195,0,0,0,94,0,223,0,111,0,239,0,45,0,1,0,24,0,0,0,234,0,0,0,114,0,175,0,79,0,120,0,18,0,191,0,0,0,0,0,115,0,244,0,75,0,134,0,108,0,202,0,19,0,22,0,0,0,165,0,108,0,213,0,0,0,39,0,56,0,136,0,32,0,175,0,0,0,98,0,240,0,0,0,58,0,0,0,0,0,160,0,21,0,115,0,81,0,59,0,59,0,21,0,208,0,0,0,167,0,119,0,0,0,243,0,0,0,211,0,0,0,75,0,38,0,17,0,241,0,0,0,140,0,156,0,152,0,78,0,70,0,0,0,235,0,27,0,102,0,162,0,157,0,0,0,224,0,0,0,0,0,14,0,32,0,209,0,101,0,170,0,117,0,246,0,80,0,205,0,190,0,0,0,87,0,118,0,32,0,165,0,0,0,0,0,91,0,238,0,3,0,232,0,243,0,0,0,10,0,44,0,46,0,177,0,20,0,0,0,173,0,0,0,0,0,161,0,148,0,0,0,172,0,0,0,2,0,237,0,38,0,200,0,0,0,205,0,143,0,167,0,132,0,74,0,133,0,243,0,248,0,2,0,119,0,170,0,0,0,0,0,212,0,26,0,129,0,149,0,194,0,137,0,0,0,156,0,231,0,246,0,191,0,37,0,209,0,192,0,0,0,0,0,139,0,149,0,32,0,182,0,0,0,242,0,0,0,156,0,73,0,197,0,0,0,127,0,242,0,31,0,158,0,130,0,0,0,75,0,77,0,35,0,0,0,0,0,7,0,207,0,0,0,244,0,140,0,232,0,53,0,220,0,0,0,27,0,147,0,241,0,180,0,49,0,0,0,88,0,222,0,0,0,29,0,43,0,231,0,0,0,158,0,198,0,254,0,1,0,0,0,44,0,1,0,161,0,157,0,126,0,137,0,0,0,12,0,113,0,34,0,0,0,7,0,133,0,188,0,154,0,0,0,81,0,150,0,164,0,0,0,0,0,64,0,64,0,192,0,138,0,1,0,31,0,249,0,142,0,61,0,80,0,242,0,0,0,237,0,83,0,171,0,0,0,148,0,68,0,213,0,45,0,20,0,188,0,108,0,71,0,165,0,247,0,92,0,245,0,0,0,0,0,15,0);
signal scenario_full  : scenario_type := (234,31,191,31,38,31,88,31,107,31,181,31,166,31,130,31,29,31,29,30,29,29,65,31,246,31,246,30,126,31,123,31,31,31,223,31,150,31,121,31,49,31,49,30,96,31,96,30,233,31,134,31,63,31,63,30,14,31,170,31,142,31,96,31,91,31,138,31,93,31,121,31,121,30,112,31,112,30,224,31,254,31,254,30,153,31,58,31,74,31,221,31,28,31,28,30,138,31,191,31,135,31,135,30,138,31,195,31,94,31,75,31,75,30,75,29,95,31,173,31,54,31,10,31,5,31,87,31,87,30,112,31,100,31,230,31,139,31,180,31,180,31,237,31,237,30,237,29,33,31,168,31,255,31,255,30,26,31,26,30,216,31,244,31,105,31,210,31,119,31,119,30,23,31,124,31,124,30,54,31,108,31,5,31,94,31,176,31,104,31,62,31,106,31,28,31,251,31,30,31,30,30,78,31,111,31,12,31,121,31,76,31,131,31,117,31,101,31,16,31,25,31,237,31,237,30,231,31,251,31,205,31,17,31,238,31,182,31,183,31,209,31,206,31,144,31,15,31,15,30,33,31,33,30,144,31,144,30,166,31,22,31,31,31,255,31,243,31,42,31,253,31,253,30,16,31,212,31,190,31,29,31,204,31,23,31,23,30,239,31,226,31,48,31,230,31,160,31,99,31,193,31,149,31,44,31,6,31,135,31,135,30,129,31,129,30,203,31,106,31,111,31,127,31,223,31,223,30,188,31,188,30,31,31,30,31,16,31,35,31,35,30,248,31,248,30,40,31,82,31,82,30,49,31,49,30,91,31,175,31,251,31,251,30,34,31,34,30,123,31,43,31,180,31,130,31,47,31,47,30,97,31,160,31,143,31,230,31,230,30,72,31,201,31,126,31,137,31,15,31,241,31,31,31,39,31,91,31,89,31,82,31,142,31,240,31,240,30,149,31,74,31,105,31,105,30,105,29,241,31,254,31,121,31,121,30,223,31,207,31,42,31,17,31,17,30,34,31,78,31,101,31,194,31,105,31,105,30,36,31,78,31,45,31,200,31,61,31,162,31,110,31,143,31,232,31,176,31,176,30,11,31,100,31,79,31,79,30,32,31,177,31,131,31,255,31,162,31,88,31,90,31,186,31,94,31,36,31,179,31,179,30,179,31,96,31,1,31,1,30,1,29,16,31,16,30,106,31,106,30,47,31,153,31,181,31,94,31,94,30,244,31,176,31,176,30,153,31,75,31,249,31,249,31,249,30,172,31,223,31,64,31,128,31,117,31,117,30,105,31,45,31,171,31,171,30,14,31,22,31,22,30,201,31,198,31,20,31,69,31,43,31,230,31,55,31,83,31,237,31,224,31,88,31,86,31,206,31,213,31,163,31,123,31,100,31,124,31,158,31,168,31,101,31,170,31,188,31,212,31,188,31,188,30,188,29,188,28,21,31,21,30,9,31,9,30,9,29,104,31,86,31,86,30,170,31,43,31,156,31,54,31,151,31,151,30,69,31,17,31,17,30,194,31,50,31,163,31,163,30,79,31,188,31,20,31,114,31,210,31,209,31,203,31,14,31,104,31,150,31,52,31,72,31,16,31,26,31,26,30,152,31,152,30,3,31,239,31,178,31,128,31,1,31,1,30,1,29,177,31,128,31,8,31,58,31,58,30,66,31,224,31,46,31,173,31,94,31,86,31,48,31,179,31,79,31,206,31,75,31,75,30,112,31,9,31,200,31,85,31,85,30,85,29,85,28,128,31,128,30,77,31,157,31,157,30,157,29,16,31,68,31,15,31,15,30,187,31,225,31,94,31,103,31,124,31,209,31,209,30,179,31,58,31,129,31,129,30,108,31,21,31,15,31,243,31,243,30,216,31,99,31,210,31,159,31,36,31,204,31,42,31,135,31,96,31,142,31,10,31,10,30,10,29,140,31,58,31,155,31,115,31,226,31,204,31,140,31,244,31,162,31,214,31,8,31,222,31,212,31,106,31,102,31,18,31,65,31,204,31,98,31,215,31,215,30,36,31,154,31,154,30,230,31,49,31,49,30,10,31,10,30,108,31,215,31,212,31,95,31,182,31,154,31,5,31,251,31,251,30,165,31,41,31,232,31,232,30,241,31,49,31,173,31,112,31,51,31,51,30,72,31,60,31,60,30,191,31,85,31,85,30,3,31,8,31,161,31,30,31,153,31,19,31,151,31,140,31,140,30,155,31,215,31,199,31,199,30,167,31,55,31,43,31,115,31,140,31,140,30,78,31,78,30,78,29,165,31,98,31,207,31,103,31,83,31,153,31,23,31,46,31,214,31,186,31,185,31,160,31,17,31,112,31,145,31,41,31,156,31,156,30,156,29,97,31,97,30,118,31,131,31,131,30,101,31,192,31,42,31,42,30,37,31,37,30,194,31,58,31,76,31,194,31,247,31,71,31,219,31,75,31,205,31,66,31,149,31,201,31,80,31,100,31,157,31,6,31,175,31,237,31,171,31,51,31,41,31,177,31,192,31,168,31,137,31,97,31,97,30,187,31,247,31,218,31,137,31,137,30,38,31,38,30,208,31,34,31,44,31,147,31,195,31,195,30,94,31,223,31,111,31,239,31,45,31,1,31,24,31,24,30,234,31,234,30,114,31,175,31,79,31,120,31,18,31,191,31,191,30,191,29,115,31,244,31,75,31,134,31,108,31,202,31,19,31,22,31,22,30,165,31,108,31,213,31,213,30,39,31,56,31,136,31,32,31,175,31,175,30,98,31,240,31,240,30,58,31,58,30,58,29,160,31,21,31,115,31,81,31,59,31,59,31,21,31,208,31,208,30,167,31,119,31,119,30,243,31,243,30,211,31,211,30,75,31,38,31,17,31,241,31,241,30,140,31,156,31,152,31,78,31,70,31,70,30,235,31,27,31,102,31,162,31,157,31,157,30,224,31,224,30,224,29,14,31,32,31,209,31,101,31,170,31,117,31,246,31,80,31,205,31,190,31,190,30,87,31,118,31,32,31,165,31,165,30,165,29,91,31,238,31,3,31,232,31,243,31,243,30,10,31,44,31,46,31,177,31,20,31,20,30,173,31,173,30,173,29,161,31,148,31,148,30,172,31,172,30,2,31,237,31,38,31,200,31,200,30,205,31,143,31,167,31,132,31,74,31,133,31,243,31,248,31,2,31,119,31,170,31,170,30,170,29,212,31,26,31,129,31,149,31,194,31,137,31,137,30,156,31,231,31,246,31,191,31,37,31,209,31,192,31,192,30,192,29,139,31,149,31,32,31,182,31,182,30,242,31,242,30,156,31,73,31,197,31,197,30,127,31,242,31,31,31,158,31,130,31,130,30,75,31,77,31,35,31,35,30,35,29,7,31,207,31,207,30,244,31,140,31,232,31,53,31,220,31,220,30,27,31,147,31,241,31,180,31,49,31,49,30,88,31,222,31,222,30,29,31,43,31,231,31,231,30,158,31,198,31,254,31,1,31,1,30,44,31,1,31,161,31,157,31,126,31,137,31,137,30,12,31,113,31,34,31,34,30,7,31,133,31,188,31,154,31,154,30,81,31,150,31,164,31,164,30,164,29,64,31,64,31,192,31,138,31,1,31,31,31,249,31,142,31,61,31,80,31,242,31,242,30,237,31,83,31,171,31,171,30,148,31,68,31,213,31,45,31,20,31,188,31,108,31,71,31,165,31,247,31,92,31,245,31,245,30,245,29,15,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
