-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 720;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (211,0,100,0,163,0,188,0,77,0,57,0,0,0,90,0,28,0,140,0,253,0,29,0,114,0,132,0,139,0,111,0,167,0,100,0,211,0,117,0,0,0,223,0,0,0,0,0,29,0,106,0,49,0,0,0,153,0,250,0,182,0,184,0,158,0,0,0,182,0,110,0,161,0,164,0,0,0,76,0,32,0,254,0,84,0,81,0,55,0,159,0,215,0,213,0,77,0,104,0,132,0,0,0,202,0,253,0,208,0,45,0,248,0,10,0,181,0,172,0,0,0,114,0,0,0,171,0,5,0,41,0,123,0,0,0,102,0,0,0,241,0,0,0,170,0,230,0,33,0,180,0,73,0,0,0,88,0,5,0,183,0,71,0,37,0,0,0,0,0,109,0,86,0,108,0,0,0,105,0,239,0,177,0,0,0,60,0,0,0,208,0,0,0,212,0,179,0,255,0,137,0,53,0,81,0,0,0,0,0,53,0,11,0,234,0,0,0,98,0,221,0,216,0,151,0,55,0,145,0,61,0,11,0,217,0,147,0,198,0,239,0,39,0,177,0,102,0,0,0,0,0,161,0,179,0,6,0,172,0,1,0,133,0,229,0,6,0,0,0,22,0,158,0,16,0,208,0,255,0,0,0,35,0,61,0,126,0,0,0,91,0,244,0,57,0,0,0,0,0,235,0,71,0,201,0,77,0,48,0,79,0,223,0,135,0,154,0,225,0,36,0,85,0,91,0,167,0,79,0,211,0,177,0,0,0,49,0,114,0,0,0,218,0,247,0,52,0,3,0,208,0,116,0,210,0,0,0,169,0,18,0,183,0,250,0,0,0,84,0,234,0,0,0,104,0,222,0,0,0,116,0,192,0,234,0,52,0,232,0,33,0,185,0,168,0,7,0,0,0,84,0,117,0,57,0,0,0,221,0,245,0,63,0,159,0,0,0,131,0,227,0,0,0,115,0,96,0,189,0,63,0,191,0,33,0,132,0,0,0,185,0,79,0,152,0,0,0,0,0,163,0,0,0,89,0,190,0,74,0,81,0,134,0,187,0,238,0,74,0,53,0,24,0,41,0,179,0,223,0,41,0,90,0,132,0,46,0,30,0,10,0,169,0,190,0,0,0,125,0,0,0,0,0,133,0,179,0,237,0,5,0,171,0,199,0,206,0,119,0,45,0,121,0,0,0,58,0,241,0,158,0,235,0,0,0,242,0,20,0,251,0,254,0,40,0,168,0,41,0,0,0,242,0,73,0,224,0,216,0,199,0,212,0,60,0,37,0,121,0,36,0,43,0,0,0,0,0,19,0,1,0,205,0,196,0,42,0,219,0,180,0,87,0,231,0,9,0,0,0,79,0,0,0,0,0,86,0,0,0,183,0,230,0,42,0,198,0,0,0,229,0,213,0,0,0,39,0,70,0,190,0,135,0,162,0,21,0,0,0,49,0,170,0,48,0,121,0,230,0,52,0,0,0,54,0,36,0,108,0,0,0,0,0,74,0,25,0,138,0,92,0,251,0,52,0,162,0,0,0,0,0,231,0,0,0,62,0,39,0,0,0,0,0,0,0,0,0,0,0,180,0,0,0,0,0,172,0,0,0,247,0,195,0,0,0,188,0,227,0,39,0,4,0,0,0,0,0,65,0,225,0,26,0,0,0,0,0,106,0,108,0,215,0,58,0,0,0,178,0,141,0,214,0,200,0,121,0,0,0,0,0,216,0,194,0,0,0,0,0,169,0,105,0,0,0,121,0,132,0,0,0,189,0,1,0,157,0,172,0,12,0,0,0,234,0,219,0,191,0,201,0,252,0,97,0,126,0,0,0,0,0,246,0,50,0,0,0,5,0,0,0,0,0,186,0,70,0,182,0,225,0,0,0,223,0,198,0,0,0,149,0,241,0,187,0,0,0,19,0,0,0,220,0,0,0,223,0,145,0,234,0,57,0,195,0,246,0,106,0,194,0,52,0,194,0,203,0,113,0,1,0,161,0,24,0,0,0,200,0,57,0,100,0,0,0,82,0,178,0,0,0,0,0,0,0,152,0,0,0,58,0,177,0,55,0,27,0,47,0,221,0,0,0,0,0,119,0,9,0,11,0,57,0,168,0,99,0,14,0,182,0,244,0,118,0,227,0,215,0,232,0,179,0,54,0,202,0,242,0,135,0,68,0,104,0,207,0,44,0,0,0,69,0,34,0,0,0,177,0,203,0,232,0,192,0,197,0,217,0,113,0,253,0,20,0,46,0,0,0,159,0,0,0,0,0,41,0,136,0,141,0,240,0,20,0,192,0,0,0,0,0,27,0,0,0,212,0,172,0,139,0,64,0,143,0,11,0,63,0,159,0,166,0,32,0,0,0,111,0,155,0,134,0,0,0,198,0,0,0,108,0,162,0,113,0,181,0,110,0,15,0,80,0,64,0,27,0,249,0,127,0,244,0,0,0,0,0,129,0,168,0,0,0,26,0,0,0,29,0,140,0,236,0,0,0,234,0,199,0,193,0,73,0,140,0,199,0,141,0,14,0,0,0,114,0,0,0,55,0,48,0,168,0,60,0,8,0,69,0,147,0,158,0,139,0,185,0,136,0,14,0,64,0,193,0,134,0,37,0,185,0,113,0,66,0,151,0,187,0,53,0,196,0,169,0,28,0,247,0,149,0,0,0,0,0,211,0,120,0,85,0,0,0,0,0,174,0,50,0,225,0,77,0,30,0,119,0,222,0,0,0,59,0,235,0,51,0,95,0,154,0,0,0,61,0,28,0,144,0,111,0,94,0,134,0,0,0,69,0,98,0,111,0,211,0,0,0,164,0,254,0,115,0,14,0,5,0,22,0,81,0,172,0,215,0,17,0,139,0,74,0,0,0,97,0,0,0,46,0,0,0,0,0,198,0,237,0,42,0,0,0,0,0,104,0,0,0,208,0,3,0,0,0,118,0,0,0,240,0,250,0,185,0,28,0,0,0,85,0,217,0,103,0,84,0,0,0,19,0,238,0,194,0,202,0,227,0,194,0,41,0,110,0,0,0,187,0,221,0,167,0,199,0,0,0,161,0,250,0,93,0,122,0,185,0,178,0,74,0,47,0,0,0,189,0,248,0,253,0,193,0,190,0,232,0,0,0,244,0,0,0,124,0,208,0,184,0,0,0,55,0,168,0,213,0,0,0,155,0,4,0,192,0,138,0,88,0,0,0,24,0,5,0,116,0,253,0,113,0,235,0,243,0,0,0,85,0,184,0);
signal scenario_full  : scenario_type := (211,31,100,31,163,31,188,31,77,31,57,31,57,30,90,31,28,31,140,31,253,31,29,31,114,31,132,31,139,31,111,31,167,31,100,31,211,31,117,31,117,30,223,31,223,30,223,29,29,31,106,31,49,31,49,30,153,31,250,31,182,31,184,31,158,31,158,30,182,31,110,31,161,31,164,31,164,30,76,31,32,31,254,31,84,31,81,31,55,31,159,31,215,31,213,31,77,31,104,31,132,31,132,30,202,31,253,31,208,31,45,31,248,31,10,31,181,31,172,31,172,30,114,31,114,30,171,31,5,31,41,31,123,31,123,30,102,31,102,30,241,31,241,30,170,31,230,31,33,31,180,31,73,31,73,30,88,31,5,31,183,31,71,31,37,31,37,30,37,29,109,31,86,31,108,31,108,30,105,31,239,31,177,31,177,30,60,31,60,30,208,31,208,30,212,31,179,31,255,31,137,31,53,31,81,31,81,30,81,29,53,31,11,31,234,31,234,30,98,31,221,31,216,31,151,31,55,31,145,31,61,31,11,31,217,31,147,31,198,31,239,31,39,31,177,31,102,31,102,30,102,29,161,31,179,31,6,31,172,31,1,31,133,31,229,31,6,31,6,30,22,31,158,31,16,31,208,31,255,31,255,30,35,31,61,31,126,31,126,30,91,31,244,31,57,31,57,30,57,29,235,31,71,31,201,31,77,31,48,31,79,31,223,31,135,31,154,31,225,31,36,31,85,31,91,31,167,31,79,31,211,31,177,31,177,30,49,31,114,31,114,30,218,31,247,31,52,31,3,31,208,31,116,31,210,31,210,30,169,31,18,31,183,31,250,31,250,30,84,31,234,31,234,30,104,31,222,31,222,30,116,31,192,31,234,31,52,31,232,31,33,31,185,31,168,31,7,31,7,30,84,31,117,31,57,31,57,30,221,31,245,31,63,31,159,31,159,30,131,31,227,31,227,30,115,31,96,31,189,31,63,31,191,31,33,31,132,31,132,30,185,31,79,31,152,31,152,30,152,29,163,31,163,30,89,31,190,31,74,31,81,31,134,31,187,31,238,31,74,31,53,31,24,31,41,31,179,31,223,31,41,31,90,31,132,31,46,31,30,31,10,31,169,31,190,31,190,30,125,31,125,30,125,29,133,31,179,31,237,31,5,31,171,31,199,31,206,31,119,31,45,31,121,31,121,30,58,31,241,31,158,31,235,31,235,30,242,31,20,31,251,31,254,31,40,31,168,31,41,31,41,30,242,31,73,31,224,31,216,31,199,31,212,31,60,31,37,31,121,31,36,31,43,31,43,30,43,29,19,31,1,31,205,31,196,31,42,31,219,31,180,31,87,31,231,31,9,31,9,30,79,31,79,30,79,29,86,31,86,30,183,31,230,31,42,31,198,31,198,30,229,31,213,31,213,30,39,31,70,31,190,31,135,31,162,31,21,31,21,30,49,31,170,31,48,31,121,31,230,31,52,31,52,30,54,31,36,31,108,31,108,30,108,29,74,31,25,31,138,31,92,31,251,31,52,31,162,31,162,30,162,29,231,31,231,30,62,31,39,31,39,30,39,29,39,28,39,27,39,26,180,31,180,30,180,29,172,31,172,30,247,31,195,31,195,30,188,31,227,31,39,31,4,31,4,30,4,29,65,31,225,31,26,31,26,30,26,29,106,31,108,31,215,31,58,31,58,30,178,31,141,31,214,31,200,31,121,31,121,30,121,29,216,31,194,31,194,30,194,29,169,31,105,31,105,30,121,31,132,31,132,30,189,31,1,31,157,31,172,31,12,31,12,30,234,31,219,31,191,31,201,31,252,31,97,31,126,31,126,30,126,29,246,31,50,31,50,30,5,31,5,30,5,29,186,31,70,31,182,31,225,31,225,30,223,31,198,31,198,30,149,31,241,31,187,31,187,30,19,31,19,30,220,31,220,30,223,31,145,31,234,31,57,31,195,31,246,31,106,31,194,31,52,31,194,31,203,31,113,31,1,31,161,31,24,31,24,30,200,31,57,31,100,31,100,30,82,31,178,31,178,30,178,29,178,28,152,31,152,30,58,31,177,31,55,31,27,31,47,31,221,31,221,30,221,29,119,31,9,31,11,31,57,31,168,31,99,31,14,31,182,31,244,31,118,31,227,31,215,31,232,31,179,31,54,31,202,31,242,31,135,31,68,31,104,31,207,31,44,31,44,30,69,31,34,31,34,30,177,31,203,31,232,31,192,31,197,31,217,31,113,31,253,31,20,31,46,31,46,30,159,31,159,30,159,29,41,31,136,31,141,31,240,31,20,31,192,31,192,30,192,29,27,31,27,30,212,31,172,31,139,31,64,31,143,31,11,31,63,31,159,31,166,31,32,31,32,30,111,31,155,31,134,31,134,30,198,31,198,30,108,31,162,31,113,31,181,31,110,31,15,31,80,31,64,31,27,31,249,31,127,31,244,31,244,30,244,29,129,31,168,31,168,30,26,31,26,30,29,31,140,31,236,31,236,30,234,31,199,31,193,31,73,31,140,31,199,31,141,31,14,31,14,30,114,31,114,30,55,31,48,31,168,31,60,31,8,31,69,31,147,31,158,31,139,31,185,31,136,31,14,31,64,31,193,31,134,31,37,31,185,31,113,31,66,31,151,31,187,31,53,31,196,31,169,31,28,31,247,31,149,31,149,30,149,29,211,31,120,31,85,31,85,30,85,29,174,31,50,31,225,31,77,31,30,31,119,31,222,31,222,30,59,31,235,31,51,31,95,31,154,31,154,30,61,31,28,31,144,31,111,31,94,31,134,31,134,30,69,31,98,31,111,31,211,31,211,30,164,31,254,31,115,31,14,31,5,31,22,31,81,31,172,31,215,31,17,31,139,31,74,31,74,30,97,31,97,30,46,31,46,30,46,29,198,31,237,31,42,31,42,30,42,29,104,31,104,30,208,31,3,31,3,30,118,31,118,30,240,31,250,31,185,31,28,31,28,30,85,31,217,31,103,31,84,31,84,30,19,31,238,31,194,31,202,31,227,31,194,31,41,31,110,31,110,30,187,31,221,31,167,31,199,31,199,30,161,31,250,31,93,31,122,31,185,31,178,31,74,31,47,31,47,30,189,31,248,31,253,31,193,31,190,31,232,31,232,30,244,31,244,30,124,31,208,31,184,31,184,30,55,31,168,31,213,31,213,30,155,31,4,31,192,31,138,31,88,31,88,30,24,31,5,31,116,31,253,31,113,31,235,31,243,31,243,30,85,31,184,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
