-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_881 is
end project_tb_881;

architecture project_tb_arch_881 of project_tb_881 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 264;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,110,0,44,0,0,0,252,0,110,0,0,0,0,0,63,0,210,0,86,0,0,0,84,0,166,0,248,0,227,0,233,0,9,0,83,0,95,0,23,0,0,0,187,0,201,0,81,0,84,0,183,0,75,0,4,0,149,0,0,0,81,0,0,0,234,0,159,0,0,0,104,0,0,0,154,0,0,0,69,0,127,0,137,0,139,0,20,0,77,0,102,0,176,0,227,0,0,0,50,0,101,0,105,0,124,0,255,0,112,0,67,0,79,0,87,0,0,0,89,0,45,0,45,0,56,0,255,0,108,0,61,0,50,0,87,0,0,0,0,0,49,0,244,0,194,0,89,0,82,0,52,0,0,0,0,0,67,0,0,0,0,0,154,0,72,0,208,0,190,0,197,0,234,0,199,0,102,0,85,0,144,0,46,0,130,0,194,0,143,0,195,0,0,0,0,0,184,0,149,0,86,0,0,0,114,0,58,0,145,0,106,0,107,0,57,0,141,0,0,0,0,0,0,0,0,0,32,0,126,0,0,0,0,0,143,0,68,0,52,0,198,0,132,0,209,0,233,0,209,0,9,0,54,0,0,0,131,0,0,0,0,0,190,0,200,0,208,0,170,0,177,0,145,0,194,0,104,0,206,0,25,0,0,0,119,0,213,0,0,0,26,0,0,0,243,0,9,0,216,0,139,0,151,0,129,0,0,0,55,0,0,0,0,0,236,0,111,0,245,0,187,0,232,0,170,0,203,0,230,0,87,0,49,0,168,0,236,0,175,0,180,0,237,0,0,0,174,0,45,0,0,0,0,0,105,0,212,0,0,0,140,0,224,0,3,0,162,0,40,0,47,0,147,0,238,0,0,0,132,0,0,0,0,0,0,0,132,0,183,0,249,0,172,0,159,0,230,0,0,0,48,0,168,0,90,0,150,0,0,0,214,0,222,0,149,0,112,0,129,0,102,0,0,0,108,0,86,0,145,0,0,0,90,0,217,0,0,0,250,0,0,0,225,0,20,0,239,0,162,0,188,0,85,0,101,0,16,0,244,0,0,0,57,0,118,0,145,0,66,0,29,0,0,0,220,0,0,0,94,0,113,0,199,0,144,0,129,0,8,0,215,0,0,0,253,0,205,0,130,0,95,0,133,0,109,0,0,0,14,0,60,0,207,0,107,0,230,0,130,0,106,0,0,0,123,0);
signal scenario_full  : scenario_type := (105,31,110,31,44,31,44,30,252,31,110,31,110,30,110,29,63,31,210,31,86,31,86,30,84,31,166,31,248,31,227,31,233,31,9,31,83,31,95,31,23,31,23,30,187,31,201,31,81,31,84,31,183,31,75,31,4,31,149,31,149,30,81,31,81,30,234,31,159,31,159,30,104,31,104,30,154,31,154,30,69,31,127,31,137,31,139,31,20,31,77,31,102,31,176,31,227,31,227,30,50,31,101,31,105,31,124,31,255,31,112,31,67,31,79,31,87,31,87,30,89,31,45,31,45,31,56,31,255,31,108,31,61,31,50,31,87,31,87,30,87,29,49,31,244,31,194,31,89,31,82,31,52,31,52,30,52,29,67,31,67,30,67,29,154,31,72,31,208,31,190,31,197,31,234,31,199,31,102,31,85,31,144,31,46,31,130,31,194,31,143,31,195,31,195,30,195,29,184,31,149,31,86,31,86,30,114,31,58,31,145,31,106,31,107,31,57,31,141,31,141,30,141,29,141,28,141,27,32,31,126,31,126,30,126,29,143,31,68,31,52,31,198,31,132,31,209,31,233,31,209,31,9,31,54,31,54,30,131,31,131,30,131,29,190,31,200,31,208,31,170,31,177,31,145,31,194,31,104,31,206,31,25,31,25,30,119,31,213,31,213,30,26,31,26,30,243,31,9,31,216,31,139,31,151,31,129,31,129,30,55,31,55,30,55,29,236,31,111,31,245,31,187,31,232,31,170,31,203,31,230,31,87,31,49,31,168,31,236,31,175,31,180,31,237,31,237,30,174,31,45,31,45,30,45,29,105,31,212,31,212,30,140,31,224,31,3,31,162,31,40,31,47,31,147,31,238,31,238,30,132,31,132,30,132,29,132,28,132,31,183,31,249,31,172,31,159,31,230,31,230,30,48,31,168,31,90,31,150,31,150,30,214,31,222,31,149,31,112,31,129,31,102,31,102,30,108,31,86,31,145,31,145,30,90,31,217,31,217,30,250,31,250,30,225,31,20,31,239,31,162,31,188,31,85,31,101,31,16,31,244,31,244,30,57,31,118,31,145,31,66,31,29,31,29,30,220,31,220,30,94,31,113,31,199,31,144,31,129,31,8,31,215,31,215,30,253,31,205,31,130,31,95,31,133,31,109,31,109,30,14,31,60,31,207,31,107,31,230,31,130,31,106,31,106,30,123,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
