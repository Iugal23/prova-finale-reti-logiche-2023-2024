-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 685;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,103,0,92,0,197,0,243,0,0,0,215,0,249,0,0,0,0,0,0,0,55,0,187,0,0,0,217,0,0,0,2,0,0,0,57,0,88,0,0,0,243,0,4,0,199,0,195,0,0,0,190,0,143,0,247,0,153,0,252,0,221,0,177,0,69,0,10,0,246,0,0,0,27,0,25,0,25,0,179,0,165,0,27,0,0,0,239,0,67,0,206,0,5,0,192,0,225,0,0,0,0,0,171,0,178,0,127,0,0,0,238,0,78,0,33,0,195,0,3,0,150,0,45,0,186,0,144,0,35,0,18,0,240,0,196,0,194,0,19,0,248,0,142,0,237,0,240,0,172,0,56,0,36,0,0,0,40,0,0,0,0,0,122,0,124,0,165,0,244,0,159,0,216,0,160,0,4,0,220,0,0,0,30,0,217,0,245,0,126,0,109,0,102,0,121,0,96,0,0,0,1,0,191,0,61,0,0,0,180,0,57,0,179,0,0,0,33,0,78,0,118,0,0,0,213,0,90,0,23,0,0,0,59,0,32,0,130,0,232,0,234,0,14,0,162,0,159,0,143,0,109,0,147,0,130,0,0,0,208,0,0,0,45,0,159,0,254,0,79,0,121,0,238,0,108,0,59,0,124,0,37,0,242,0,0,0,0,0,35,0,97,0,14,0,40,0,90,0,16,0,42,0,156,0,0,0,41,0,230,0,138,0,0,0,102,0,10,0,116,0,0,0,231,0,129,0,0,0,58,0,246,0,144,0,0,0,55,0,23,0,59,0,70,0,113,0,12,0,172,0,95,0,229,0,36,0,67,0,121,0,95,0,22,0,15,0,207,0,177,0,0,0,25,0,51,0,71,0,227,0,147,0,158,0,143,0,50,0,0,0,95,0,211,0,217,0,223,0,156,0,68,0,0,0,35,0,35,0,30,0,0,0,46,0,84,0,45,0,0,0,32,0,208,0,202,0,223,0,251,0,114,0,146,0,97,0,159,0,195,0,19,0,106,0,32,0,63,0,206,0,159,0,0,0,127,0,98,0,185,0,241,0,225,0,160,0,0,0,0,0,106,0,202,0,124,0,41,0,46,0,0,0,90,0,217,0,194,0,4,0,243,0,0,0,171,0,206,0,78,0,187,0,117,0,65,0,0,0,0,0,31,0,154,0,163,0,0,0,124,0,67,0,177,0,0,0,0,0,0,0,6,0,152,0,168,0,0,0,153,0,176,0,37,0,119,0,0,0,120,0,195,0,199,0,25,0,199,0,0,0,126,0,254,0,82,0,133,0,226,0,197,0,233,0,36,0,0,0,0,0,219,0,39,0,0,0,222,0,23,0,190,0,19,0,0,0,0,0,0,0,245,0,0,0,173,0,234,0,0,0,65,0,105,0,56,0,119,0,0,0,244,0,172,0,59,0,0,0,193,0,98,0,116,0,96,0,178,0,66,0,17,0,72,0,144,0,124,0,119,0,51,0,0,0,92,0,0,0,110,0,84,0,0,0,238,0,131,0,115,0,0,0,117,0,163,0,61,0,45,0,34,0,0,0,106,0,127,0,7,0,0,0,79,0,51,0,175,0,62,0,0,0,252,0,126,0,248,0,202,0,0,0,54,0,69,0,63,0,193,0,75,0,0,0,201,0,125,0,100,0,130,0,210,0,65,0,92,0,22,0,0,0,221,0,104,0,133,0,214,0,136,0,202,0,226,0,0,0,222,0,162,0,115,0,7,0,249,0,192,0,0,0,0,0,17,0,0,0,62,0,10,0,116,0,211,0,113,0,138,0,233,0,45,0,144,0,192,0,127,0,0,0,62,0,0,0,0,0,114,0,0,0,115,0,31,0,225,0,0,0,209,0,42,0,44,0,173,0,159,0,164,0,0,0,61,0,112,0,101,0,0,0,83,0,132,0,253,0,120,0,253,0,236,0,0,0,136,0,1,0,71,0,0,0,172,0,135,0,24,0,83,0,0,0,85,0,41,0,229,0,231,0,0,0,158,0,44,0,33,0,234,0,203,0,185,0,225,0,242,0,0,0,208,0,57,0,117,0,0,0,206,0,0,0,207,0,158,0,5,0,0,0,163,0,231,0,0,0,74,0,0,0,0,0,0,0,0,0,202,0,0,0,0,0,0,0,96,0,0,0,254,0,193,0,57,0,16,0,39,0,199,0,193,0,43,0,0,0,229,0,177,0,188,0,52,0,0,0,60,0,246,0,123,0,226,0,0,0,162,0,207,0,35,0,229,0,162,0,94,0,25,0,0,0,105,0,8,0,48,0,191,0,0,0,242,0,0,0,250,0,208,0,76,0,125,0,22,0,67,0,0,0,18,0,81,0,7,0,0,0,160,0,0,0,183,0,88,0,139,0,46,0,213,0,159,0,215,0,0,0,61,0,101,0,0,0,72,0,43,0,229,0,138,0,0,0,151,0,113,0,148,0,86,0,42,0,0,0,0,0,139,0,156,0,170,0,0,0,0,0,0,0,142,0,134,0,120,0,136,0,115,0,127,0,219,0,9,0,127,0,0,0,213,0,0,0,5,0,116,0,85,0,247,0,185,0,112,0,65,0,0,0,150,0,170,0,187,0,146,0,0,0,239,0,181,0,211,0,225,0,0,0,230,0,207,0,10,0,0,0,7,0,0,0,68,0,14,0,129,0,0,0,93,0,0,0,120,0,0,0,35,0,91,0,0,0,254,0,235,0,57,0,145,0,130,0,51,0,67,0,0,0,0,0,163,0,141,0,202,0,232,0,179,0,141,0,138,0,16,0,140,0,60,0,79,0,132,0,118,0,12,0,61,0,153,0,42,0,227,0,34,0,136,0,95,0,237,0,0,0,69,0,178,0,6,0,90,0,110,0,182,0,0,0,208,0,167,0,221,0,106,0,190,0,41,0,0,0,77,0,72,0,0,0,44,0,43,0,6,0,163,0,0,0,206,0,0,0,131,0,0,0,137,0,141,0,0,0,171,0,64,0,80,0,0,0,64,0,148,0,221,0,70,0,0,0,179,0,160,0,243,0,155,0,55,0,0,0,0,0,0,0,100,0,82,0,20,0,0,0,236,0,49,0,56,0,80,0);
signal scenario_full  : scenario_type := (0,0,103,31,92,31,197,31,243,31,243,30,215,31,249,31,249,30,249,29,249,28,55,31,187,31,187,30,217,31,217,30,2,31,2,30,57,31,88,31,88,30,243,31,4,31,199,31,195,31,195,30,190,31,143,31,247,31,153,31,252,31,221,31,177,31,69,31,10,31,246,31,246,30,27,31,25,31,25,31,179,31,165,31,27,31,27,30,239,31,67,31,206,31,5,31,192,31,225,31,225,30,225,29,171,31,178,31,127,31,127,30,238,31,78,31,33,31,195,31,3,31,150,31,45,31,186,31,144,31,35,31,18,31,240,31,196,31,194,31,19,31,248,31,142,31,237,31,240,31,172,31,56,31,36,31,36,30,40,31,40,30,40,29,122,31,124,31,165,31,244,31,159,31,216,31,160,31,4,31,220,31,220,30,30,31,217,31,245,31,126,31,109,31,102,31,121,31,96,31,96,30,1,31,191,31,61,31,61,30,180,31,57,31,179,31,179,30,33,31,78,31,118,31,118,30,213,31,90,31,23,31,23,30,59,31,32,31,130,31,232,31,234,31,14,31,162,31,159,31,143,31,109,31,147,31,130,31,130,30,208,31,208,30,45,31,159,31,254,31,79,31,121,31,238,31,108,31,59,31,124,31,37,31,242,31,242,30,242,29,35,31,97,31,14,31,40,31,90,31,16,31,42,31,156,31,156,30,41,31,230,31,138,31,138,30,102,31,10,31,116,31,116,30,231,31,129,31,129,30,58,31,246,31,144,31,144,30,55,31,23,31,59,31,70,31,113,31,12,31,172,31,95,31,229,31,36,31,67,31,121,31,95,31,22,31,15,31,207,31,177,31,177,30,25,31,51,31,71,31,227,31,147,31,158,31,143,31,50,31,50,30,95,31,211,31,217,31,223,31,156,31,68,31,68,30,35,31,35,31,30,31,30,30,46,31,84,31,45,31,45,30,32,31,208,31,202,31,223,31,251,31,114,31,146,31,97,31,159,31,195,31,19,31,106,31,32,31,63,31,206,31,159,31,159,30,127,31,98,31,185,31,241,31,225,31,160,31,160,30,160,29,106,31,202,31,124,31,41,31,46,31,46,30,90,31,217,31,194,31,4,31,243,31,243,30,171,31,206,31,78,31,187,31,117,31,65,31,65,30,65,29,31,31,154,31,163,31,163,30,124,31,67,31,177,31,177,30,177,29,177,28,6,31,152,31,168,31,168,30,153,31,176,31,37,31,119,31,119,30,120,31,195,31,199,31,25,31,199,31,199,30,126,31,254,31,82,31,133,31,226,31,197,31,233,31,36,31,36,30,36,29,219,31,39,31,39,30,222,31,23,31,190,31,19,31,19,30,19,29,19,28,245,31,245,30,173,31,234,31,234,30,65,31,105,31,56,31,119,31,119,30,244,31,172,31,59,31,59,30,193,31,98,31,116,31,96,31,178,31,66,31,17,31,72,31,144,31,124,31,119,31,51,31,51,30,92,31,92,30,110,31,84,31,84,30,238,31,131,31,115,31,115,30,117,31,163,31,61,31,45,31,34,31,34,30,106,31,127,31,7,31,7,30,79,31,51,31,175,31,62,31,62,30,252,31,126,31,248,31,202,31,202,30,54,31,69,31,63,31,193,31,75,31,75,30,201,31,125,31,100,31,130,31,210,31,65,31,92,31,22,31,22,30,221,31,104,31,133,31,214,31,136,31,202,31,226,31,226,30,222,31,162,31,115,31,7,31,249,31,192,31,192,30,192,29,17,31,17,30,62,31,10,31,116,31,211,31,113,31,138,31,233,31,45,31,144,31,192,31,127,31,127,30,62,31,62,30,62,29,114,31,114,30,115,31,31,31,225,31,225,30,209,31,42,31,44,31,173,31,159,31,164,31,164,30,61,31,112,31,101,31,101,30,83,31,132,31,253,31,120,31,253,31,236,31,236,30,136,31,1,31,71,31,71,30,172,31,135,31,24,31,83,31,83,30,85,31,41,31,229,31,231,31,231,30,158,31,44,31,33,31,234,31,203,31,185,31,225,31,242,31,242,30,208,31,57,31,117,31,117,30,206,31,206,30,207,31,158,31,5,31,5,30,163,31,231,31,231,30,74,31,74,30,74,29,74,28,74,27,202,31,202,30,202,29,202,28,96,31,96,30,254,31,193,31,57,31,16,31,39,31,199,31,193,31,43,31,43,30,229,31,177,31,188,31,52,31,52,30,60,31,246,31,123,31,226,31,226,30,162,31,207,31,35,31,229,31,162,31,94,31,25,31,25,30,105,31,8,31,48,31,191,31,191,30,242,31,242,30,250,31,208,31,76,31,125,31,22,31,67,31,67,30,18,31,81,31,7,31,7,30,160,31,160,30,183,31,88,31,139,31,46,31,213,31,159,31,215,31,215,30,61,31,101,31,101,30,72,31,43,31,229,31,138,31,138,30,151,31,113,31,148,31,86,31,42,31,42,30,42,29,139,31,156,31,170,31,170,30,170,29,170,28,142,31,134,31,120,31,136,31,115,31,127,31,219,31,9,31,127,31,127,30,213,31,213,30,5,31,116,31,85,31,247,31,185,31,112,31,65,31,65,30,150,31,170,31,187,31,146,31,146,30,239,31,181,31,211,31,225,31,225,30,230,31,207,31,10,31,10,30,7,31,7,30,68,31,14,31,129,31,129,30,93,31,93,30,120,31,120,30,35,31,91,31,91,30,254,31,235,31,57,31,145,31,130,31,51,31,67,31,67,30,67,29,163,31,141,31,202,31,232,31,179,31,141,31,138,31,16,31,140,31,60,31,79,31,132,31,118,31,12,31,61,31,153,31,42,31,227,31,34,31,136,31,95,31,237,31,237,30,69,31,178,31,6,31,90,31,110,31,182,31,182,30,208,31,167,31,221,31,106,31,190,31,41,31,41,30,77,31,72,31,72,30,44,31,43,31,6,31,163,31,163,30,206,31,206,30,131,31,131,30,137,31,141,31,141,30,171,31,64,31,80,31,80,30,64,31,148,31,221,31,70,31,70,30,179,31,160,31,243,31,155,31,55,31,55,30,55,29,55,28,100,31,82,31,20,31,20,30,236,31,49,31,56,31,80,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
