-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_69 is
end project_tb_69;

architecture project_tb_arch_69 of project_tb_69 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 329;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,14,0,0,0,22,0,182,0,170,0,208,0,0,0,224,0,62,0,233,0,58,0,0,0,0,0,0,0,205,0,237,0,11,0,64,0,104,0,0,0,0,0,202,0,168,0,230,0,243,0,140,0,150,0,146,0,71,0,38,0,54,0,92,0,0,0,22,0,0,0,98,0,0,0,149,0,68,0,0,0,203,0,20,0,188,0,232,0,236,0,52,0,187,0,205,0,91,0,193,0,22,0,98,0,236,0,218,0,155,0,188,0,19,0,243,0,78,0,155,0,226,0,0,0,147,0,103,0,218,0,119,0,53,0,116,0,130,0,151,0,112,0,210,0,103,0,183,0,76,0,129,0,146,0,72,0,0,0,49,0,73,0,110,0,248,0,70,0,109,0,229,0,152,0,79,0,0,0,0,0,7,0,217,0,68,0,111,0,32,0,191,0,161,0,39,0,40,0,252,0,0,0,0,0,170,0,53,0,120,0,39,0,138,0,7,0,0,0,0,0,202,0,36,0,163,0,19,0,49,0,214,0,0,0,25,0,85,0,148,0,0,0,102,0,13,0,0,0,214,0,243,0,0,0,112,0,125,0,31,0,199,0,166,0,6,0,72,0,87,0,97,0,174,0,95,0,172,0,5,0,46,0,95,0,185,0,0,0,182,0,158,0,0,0,48,0,0,0,93,0,208,0,0,0,250,0,250,0,117,0,94,0,47,0,169,0,176,0,3,0,104,0,210,0,41,0,0,0,138,0,247,0,110,0,0,0,111,0,0,0,179,0,91,0,155,0,102,0,0,0,226,0,105,0,31,0,77,0,54,0,119,0,157,0,172,0,190,0,95,0,54,0,101,0,0,0,169,0,73,0,0,0,220,0,97,0,236,0,140,0,193,0,126,0,27,0,0,0,108,0,141,0,152,0,0,0,187,0,215,0,38,0,162,0,33,0,152,0,0,0,124,0,26,0,245,0,0,0,54,0,111,0,32,0,83,0,221,0,0,0,87,0,138,0,222,0,184,0,0,0,230,0,32,0,73,0,0,0,145,0,30,0,0,0,196,0,0,0,231,0,160,0,223,0,46,0,120,0,203,0,0,0,84,0,0,0,103,0,0,0,96,0,144,0,128,0,124,0,0,0,0,0,62,0,212,0,0,0,160,0,140,0,0,0,253,0,144,0,87,0,135,0,189,0,64,0,0,0,132,0,254,0,119,0,55,0,251,0,146,0,210,0,198,0,85,0,254,0,41,0,98,0,0,0,0,0,55,0,192,0,242,0,137,0,59,0,210,0,102,0,85,0,217,0,123,0,98,0,224,0,41,0,225,0,194,0,243,0,134,0,143,0,50,0,0,0,0,0,237,0,0,0,228,0,134,0,0,0,203,0,249,0,207,0,133,0,0,0,88,0,204,0,16,0,14,0,23,0,185,0,0,0,0,0,128,0,209,0,61,0,104,0,98,0,251,0,2,0,0,0,246,0,0,0,111,0);
signal scenario_full  : scenario_type := (201,31,14,31,14,30,22,31,182,31,170,31,208,31,208,30,224,31,62,31,233,31,58,31,58,30,58,29,58,28,205,31,237,31,11,31,64,31,104,31,104,30,104,29,202,31,168,31,230,31,243,31,140,31,150,31,146,31,71,31,38,31,54,31,92,31,92,30,22,31,22,30,98,31,98,30,149,31,68,31,68,30,203,31,20,31,188,31,232,31,236,31,52,31,187,31,205,31,91,31,193,31,22,31,98,31,236,31,218,31,155,31,188,31,19,31,243,31,78,31,155,31,226,31,226,30,147,31,103,31,218,31,119,31,53,31,116,31,130,31,151,31,112,31,210,31,103,31,183,31,76,31,129,31,146,31,72,31,72,30,49,31,73,31,110,31,248,31,70,31,109,31,229,31,152,31,79,31,79,30,79,29,7,31,217,31,68,31,111,31,32,31,191,31,161,31,39,31,40,31,252,31,252,30,252,29,170,31,53,31,120,31,39,31,138,31,7,31,7,30,7,29,202,31,36,31,163,31,19,31,49,31,214,31,214,30,25,31,85,31,148,31,148,30,102,31,13,31,13,30,214,31,243,31,243,30,112,31,125,31,31,31,199,31,166,31,6,31,72,31,87,31,97,31,174,31,95,31,172,31,5,31,46,31,95,31,185,31,185,30,182,31,158,31,158,30,48,31,48,30,93,31,208,31,208,30,250,31,250,31,117,31,94,31,47,31,169,31,176,31,3,31,104,31,210,31,41,31,41,30,138,31,247,31,110,31,110,30,111,31,111,30,179,31,91,31,155,31,102,31,102,30,226,31,105,31,31,31,77,31,54,31,119,31,157,31,172,31,190,31,95,31,54,31,101,31,101,30,169,31,73,31,73,30,220,31,97,31,236,31,140,31,193,31,126,31,27,31,27,30,108,31,141,31,152,31,152,30,187,31,215,31,38,31,162,31,33,31,152,31,152,30,124,31,26,31,245,31,245,30,54,31,111,31,32,31,83,31,221,31,221,30,87,31,138,31,222,31,184,31,184,30,230,31,32,31,73,31,73,30,145,31,30,31,30,30,196,31,196,30,231,31,160,31,223,31,46,31,120,31,203,31,203,30,84,31,84,30,103,31,103,30,96,31,144,31,128,31,124,31,124,30,124,29,62,31,212,31,212,30,160,31,140,31,140,30,253,31,144,31,87,31,135,31,189,31,64,31,64,30,132,31,254,31,119,31,55,31,251,31,146,31,210,31,198,31,85,31,254,31,41,31,98,31,98,30,98,29,55,31,192,31,242,31,137,31,59,31,210,31,102,31,85,31,217,31,123,31,98,31,224,31,41,31,225,31,194,31,243,31,134,31,143,31,50,31,50,30,50,29,237,31,237,30,228,31,134,31,134,30,203,31,249,31,207,31,133,31,133,30,88,31,204,31,16,31,14,31,23,31,185,31,185,30,185,29,128,31,209,31,61,31,104,31,98,31,251,31,2,31,2,30,246,31,246,30,111,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
