-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 165;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (66,0,149,0,242,0,166,0,204,0,196,0,11,0,47,0,61,0,155,0,199,0,0,0,80,0,3,0,0,0,0,0,0,0,45,0,0,0,13,0,38,0,154,0,0,0,18,0,0,0,198,0,0,0,251,0,240,0,14,0,29,0,128,0,0,0,117,0,244,0,179,0,79,0,237,0,62,0,237,0,135,0,6,0,95,0,251,0,0,0,37,0,222,0,204,0,236,0,30,0,75,0,71,0,31,0,147,0,29,0,0,0,140,0,90,0,176,0,253,0,54,0,155,0,74,0,68,0,83,0,68,0,8,0,0,0,164,0,0,0,81,0,206,0,0,0,243,0,17,0,36,0,28,0,0,0,0,0,0,0,237,0,104,0,250,0,6,0,5,0,195,0,0,0,0,0,76,0,0,0,234,0,232,0,117,0,173,0,0,0,200,0,40,0,0,0,110,0,129,0,83,0,0,0,121,0,0,0,0,0,113,0,114,0,119,0,154,0,92,0,246,0,195,0,134,0,201,0,4,0,147,0,193,0,147,0,0,0,13,0,228,0,160,0,88,0,0,0,113,0,239,0,112,0,22,0,200,0,0,0,0,0,0,0,0,0,69,0,228,0,222,0,246,0,9,0,98,0,66,0,0,0,95,0,73,0,0,0,21,0,203,0,30,0,0,0,177,0,48,0,189,0,0,0,62,0,15,0,37,0,12,0,215,0,0,0,0,0,110,0,175,0,0,0,122,0,235,0,67,0);
signal scenario_full  : scenario_type := (66,31,149,31,242,31,166,31,204,31,196,31,11,31,47,31,61,31,155,31,199,31,199,30,80,31,3,31,3,30,3,29,3,28,45,31,45,30,13,31,38,31,154,31,154,30,18,31,18,30,198,31,198,30,251,31,240,31,14,31,29,31,128,31,128,30,117,31,244,31,179,31,79,31,237,31,62,31,237,31,135,31,6,31,95,31,251,31,251,30,37,31,222,31,204,31,236,31,30,31,75,31,71,31,31,31,147,31,29,31,29,30,140,31,90,31,176,31,253,31,54,31,155,31,74,31,68,31,83,31,68,31,8,31,8,30,164,31,164,30,81,31,206,31,206,30,243,31,17,31,36,31,28,31,28,30,28,29,28,28,237,31,104,31,250,31,6,31,5,31,195,31,195,30,195,29,76,31,76,30,234,31,232,31,117,31,173,31,173,30,200,31,40,31,40,30,110,31,129,31,83,31,83,30,121,31,121,30,121,29,113,31,114,31,119,31,154,31,92,31,246,31,195,31,134,31,201,31,4,31,147,31,193,31,147,31,147,30,13,31,228,31,160,31,88,31,88,30,113,31,239,31,112,31,22,31,200,31,200,30,200,29,200,28,200,27,69,31,228,31,222,31,246,31,9,31,98,31,66,31,66,30,95,31,73,31,73,30,21,31,203,31,30,31,30,30,177,31,48,31,189,31,189,30,62,31,15,31,37,31,12,31,215,31,215,30,215,29,110,31,175,31,175,30,122,31,235,31,67,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
