-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 496;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,222,0,10,0,188,0,118,0,25,0,171,0,0,0,164,0,0,0,129,0,19,0,137,0,19,0,19,0,0,0,154,0,154,0,0,0,9,0,0,0,202,0,253,0,0,0,38,0,88,0,4,0,0,0,0,0,233,0,0,0,0,0,200,0,167,0,78,0,5,0,0,0,195,0,0,0,94,0,117,0,0,0,0,0,105,0,139,0,11,0,125,0,132,0,195,0,0,0,150,0,87,0,55,0,174,0,17,0,253,0,91,0,0,0,113,0,0,0,87,0,31,0,0,0,229,0,67,0,157,0,195,0,0,0,180,0,246,0,137,0,0,0,189,0,56,0,0,0,79,0,214,0,88,0,81,0,113,0,0,0,169,0,169,0,54,0,158,0,0,0,73,0,252,0,83,0,44,0,115,0,91,0,135,0,0,0,168,0,76,0,254,0,98,0,174,0,122,0,0,0,66,0,197,0,170,0,140,0,126,0,149,0,250,0,0,0,93,0,26,0,149,0,247,0,0,0,0,0,70,0,73,0,97,0,209,0,129,0,177,0,26,0,246,0,196,0,35,0,190,0,234,0,214,0,73,0,155,0,82,0,44,0,159,0,228,0,174,0,3,0,0,0,205,0,223,0,134,0,253,0,74,0,60,0,10,0,6,0,197,0,213,0,0,0,155,0,53,0,193,0,88,0,14,0,235,0,153,0,135,0,81,0,123,0,167,0,217,0,145,0,246,0,140,0,107,0,0,0,230,0,249,0,237,0,59,0,60,0,3,0,23,0,199,0,0,0,254,0,39,0,215,0,0,0,146,0,246,0,69,0,102,0,102,0,112,0,197,0,21,0,90,0,0,0,213,0,180,0,182,0,25,0,137,0,120,0,223,0,116,0,159,0,195,0,23,0,0,0,192,0,151,0,136,0,101,0,198,0,194,0,0,0,28,0,121,0,128,0,164,0,36,0,157,0,112,0,0,0,73,0,0,0,217,0,253,0,246,0,161,0,0,0,106,0,0,0,185,0,75,0,34,0,153,0,70,0,223,0,221,0,238,0,116,0,0,0,248,0,47,0,72,0,43,0,18,0,134,0,114,0,0,0,224,0,131,0,83,0,0,0,174,0,82,0,119,0,0,0,248,0,253,0,0,0,0,0,0,0,94,0,67,0,0,0,22,0,191,0,224,0,235,0,141,0,48,0,0,0,0,0,97,0,237,0,188,0,48,0,0,0,15,0,156,0,9,0,210,0,249,0,0,0,119,0,0,0,54,0,0,0,0,0,179,0,203,0,24,0,251,0,107,0,231,0,0,0,129,0,106,0,0,0,224,0,77,0,0,0,201,0,130,0,28,0,16,0,79,0,0,0,0,0,188,0,141,0,221,0,0,0,214,0,80,0,0,0,135,0,232,0,221,0,0,0,58,0,244,0,128,0,0,0,26,0,193,0,112,0,75,0,23,0,67,0,0,0,119,0,119,0,152,0,128,0,4,0,215,0,83,0,0,0,179,0,41,0,0,0,110,0,156,0,159,0,138,0,2,0,241,0,0,0,181,0,172,0,128,0,112,0,230,0,210,0,94,0,0,0,165,0,164,0,51,0,0,0,186,0,205,0,0,0,0,0,0,0,100,0,40,0,143,0,230,0,165,0,251,0,108,0,137,0,0,0,217,0,129,0,189,0,20,0,14,0,0,0,255,0,186,0,36,0,113,0,145,0,124,0,80,0,106,0,235,0,151,0,121,0,155,0,202,0,162,0,59,0,26,0,0,0,182,0,27,0,0,0,158,0,179,0,236,0,122,0,0,0,155,0,114,0,6,0,132,0,131,0,0,0,0,0,0,0,247,0,71,0,0,0,0,0,3,0,70,0,31,0,0,0,59,0,155,0,1,0,167,0,76,0,198,0,145,0,0,0,95,0,230,0,96,0,67,0,101,0,211,0,80,0,223,0,69,0,162,0,162,0,152,0,15,0,0,0,248,0,0,0,220,0,167,0,93,0,83,0,194,0,75,0,224,0,23,0,157,0,91,0,29,0,57,0,87,0,224,0,238,0,167,0,212,0,0,0,11,0,198,0,185,0,0,0,6,0,0,0,145,0,108,0,255,0,18,0,40,0,70,0,111,0,124,0,73,0,77,0,44,0,73,0,245,0,51,0,0,0,49,0,210,0,1,0,155,0,0,0,194,0,229,0,0,0,0,0,172,0,118,0,49,0,39,0,143,0,116,0,250,0,246,0,233,0);
signal scenario_full  : scenario_type := (24,31,222,31,10,31,188,31,118,31,25,31,171,31,171,30,164,31,164,30,129,31,19,31,137,31,19,31,19,31,19,30,154,31,154,31,154,30,9,31,9,30,202,31,253,31,253,30,38,31,88,31,4,31,4,30,4,29,233,31,233,30,233,29,200,31,167,31,78,31,5,31,5,30,195,31,195,30,94,31,117,31,117,30,117,29,105,31,139,31,11,31,125,31,132,31,195,31,195,30,150,31,87,31,55,31,174,31,17,31,253,31,91,31,91,30,113,31,113,30,87,31,31,31,31,30,229,31,67,31,157,31,195,31,195,30,180,31,246,31,137,31,137,30,189,31,56,31,56,30,79,31,214,31,88,31,81,31,113,31,113,30,169,31,169,31,54,31,158,31,158,30,73,31,252,31,83,31,44,31,115,31,91,31,135,31,135,30,168,31,76,31,254,31,98,31,174,31,122,31,122,30,66,31,197,31,170,31,140,31,126,31,149,31,250,31,250,30,93,31,26,31,149,31,247,31,247,30,247,29,70,31,73,31,97,31,209,31,129,31,177,31,26,31,246,31,196,31,35,31,190,31,234,31,214,31,73,31,155,31,82,31,44,31,159,31,228,31,174,31,3,31,3,30,205,31,223,31,134,31,253,31,74,31,60,31,10,31,6,31,197,31,213,31,213,30,155,31,53,31,193,31,88,31,14,31,235,31,153,31,135,31,81,31,123,31,167,31,217,31,145,31,246,31,140,31,107,31,107,30,230,31,249,31,237,31,59,31,60,31,3,31,23,31,199,31,199,30,254,31,39,31,215,31,215,30,146,31,246,31,69,31,102,31,102,31,112,31,197,31,21,31,90,31,90,30,213,31,180,31,182,31,25,31,137,31,120,31,223,31,116,31,159,31,195,31,23,31,23,30,192,31,151,31,136,31,101,31,198,31,194,31,194,30,28,31,121,31,128,31,164,31,36,31,157,31,112,31,112,30,73,31,73,30,217,31,253,31,246,31,161,31,161,30,106,31,106,30,185,31,75,31,34,31,153,31,70,31,223,31,221,31,238,31,116,31,116,30,248,31,47,31,72,31,43,31,18,31,134,31,114,31,114,30,224,31,131,31,83,31,83,30,174,31,82,31,119,31,119,30,248,31,253,31,253,30,253,29,253,28,94,31,67,31,67,30,22,31,191,31,224,31,235,31,141,31,48,31,48,30,48,29,97,31,237,31,188,31,48,31,48,30,15,31,156,31,9,31,210,31,249,31,249,30,119,31,119,30,54,31,54,30,54,29,179,31,203,31,24,31,251,31,107,31,231,31,231,30,129,31,106,31,106,30,224,31,77,31,77,30,201,31,130,31,28,31,16,31,79,31,79,30,79,29,188,31,141,31,221,31,221,30,214,31,80,31,80,30,135,31,232,31,221,31,221,30,58,31,244,31,128,31,128,30,26,31,193,31,112,31,75,31,23,31,67,31,67,30,119,31,119,31,152,31,128,31,4,31,215,31,83,31,83,30,179,31,41,31,41,30,110,31,156,31,159,31,138,31,2,31,241,31,241,30,181,31,172,31,128,31,112,31,230,31,210,31,94,31,94,30,165,31,164,31,51,31,51,30,186,31,205,31,205,30,205,29,205,28,100,31,40,31,143,31,230,31,165,31,251,31,108,31,137,31,137,30,217,31,129,31,189,31,20,31,14,31,14,30,255,31,186,31,36,31,113,31,145,31,124,31,80,31,106,31,235,31,151,31,121,31,155,31,202,31,162,31,59,31,26,31,26,30,182,31,27,31,27,30,158,31,179,31,236,31,122,31,122,30,155,31,114,31,6,31,132,31,131,31,131,30,131,29,131,28,247,31,71,31,71,30,71,29,3,31,70,31,31,31,31,30,59,31,155,31,1,31,167,31,76,31,198,31,145,31,145,30,95,31,230,31,96,31,67,31,101,31,211,31,80,31,223,31,69,31,162,31,162,31,152,31,15,31,15,30,248,31,248,30,220,31,167,31,93,31,83,31,194,31,75,31,224,31,23,31,157,31,91,31,29,31,57,31,87,31,224,31,238,31,167,31,212,31,212,30,11,31,198,31,185,31,185,30,6,31,6,30,145,31,108,31,255,31,18,31,40,31,70,31,111,31,124,31,73,31,77,31,44,31,73,31,245,31,51,31,51,30,49,31,210,31,1,31,155,31,155,30,194,31,229,31,229,30,229,29,172,31,118,31,49,31,39,31,143,31,116,31,250,31,246,31,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
