-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 270;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,116,0,202,0,35,0,184,0,75,0,6,0,226,0,190,0,51,0,0,0,197,0,0,0,125,0,0,0,105,0,0,0,90,0,16,0,139,0,215,0,206,0,1,0,101,0,241,0,32,0,76,0,181,0,156,0,0,0,91,0,74,0,164,0,58,0,162,0,5,0,0,0,209,0,0,0,42,0,4,0,55,0,189,0,166,0,201,0,203,0,0,0,63,0,0,0,101,0,0,0,91,0,77,0,151,0,145,0,156,0,237,0,0,0,17,0,0,0,0,0,243,0,44,0,89,0,46,0,88,0,149,0,56,0,133,0,99,0,0,0,28,0,0,0,175,0,202,0,0,0,0,0,228,0,45,0,0,0,192,0,143,0,53,0,200,0,201,0,239,0,243,0,174,0,49,0,190,0,104,0,149,0,224,0,68,0,110,0,253,0,232,0,163,0,122,0,38,0,178,0,0,0,28,0,230,0,0,0,214,0,135,0,0,0,232,0,102,0,6,0,105,0,51,0,96,0,12,0,252,0,49,0,116,0,237,0,0,0,226,0,164,0,0,0,158,0,0,0,69,0,90,0,120,0,122,0,250,0,116,0,9,0,211,0,0,0,162,0,93,0,66,0,174,0,125,0,48,0,8,0,134,0,166,0,191,0,64,0,220,0,100,0,0,0,227,0,178,0,56,0,136,0,26,0,9,0,63,0,229,0,58,0,0,0,13,0,9,0,54,0,184,0,240,0,0,0,46,0,82,0,153,0,237,0,0,0,112,0,0,0,0,0,244,0,72,0,0,0,36,0,71,0,128,0,251,0,0,0,114,0,26,0,213,0,45,0,0,0,230,0,216,0,216,0,30,0,233,0,143,0,0,0,0,0,35,0,0,0,243,0,163,0,236,0,129,0,0,0,146,0,183,0,0,0,249,0,137,0,110,0,208,0,59,0,189,0,172,0,67,0,132,0,24,0,0,0,33,0,0,0,157,0,83,0,244,0,24,0,120,0,46,0,157,0,147,0,90,0,117,0,246,0,88,0,0,0,109,0,66,0,82,0,213,0,70,0,0,0,152,0,205,0,0,0,175,0,199,0,211,0,0,0,152,0,17,0,0,0,125,0,0,0,41,0,0,0,46,0,56,0,164,0,0,0,13,0,99,0,0,0,26,0,119,0,0,0,42,0,0,0,16,0,0,0,65,0,68,0,0,0,232,0,139,0,236,0);
signal scenario_full  : scenario_type := (0,0,0,0,116,31,202,31,35,31,184,31,75,31,6,31,226,31,190,31,51,31,51,30,197,31,197,30,125,31,125,30,105,31,105,30,90,31,16,31,139,31,215,31,206,31,1,31,101,31,241,31,32,31,76,31,181,31,156,31,156,30,91,31,74,31,164,31,58,31,162,31,5,31,5,30,209,31,209,30,42,31,4,31,55,31,189,31,166,31,201,31,203,31,203,30,63,31,63,30,101,31,101,30,91,31,77,31,151,31,145,31,156,31,237,31,237,30,17,31,17,30,17,29,243,31,44,31,89,31,46,31,88,31,149,31,56,31,133,31,99,31,99,30,28,31,28,30,175,31,202,31,202,30,202,29,228,31,45,31,45,30,192,31,143,31,53,31,200,31,201,31,239,31,243,31,174,31,49,31,190,31,104,31,149,31,224,31,68,31,110,31,253,31,232,31,163,31,122,31,38,31,178,31,178,30,28,31,230,31,230,30,214,31,135,31,135,30,232,31,102,31,6,31,105,31,51,31,96,31,12,31,252,31,49,31,116,31,237,31,237,30,226,31,164,31,164,30,158,31,158,30,69,31,90,31,120,31,122,31,250,31,116,31,9,31,211,31,211,30,162,31,93,31,66,31,174,31,125,31,48,31,8,31,134,31,166,31,191,31,64,31,220,31,100,31,100,30,227,31,178,31,56,31,136,31,26,31,9,31,63,31,229,31,58,31,58,30,13,31,9,31,54,31,184,31,240,31,240,30,46,31,82,31,153,31,237,31,237,30,112,31,112,30,112,29,244,31,72,31,72,30,36,31,71,31,128,31,251,31,251,30,114,31,26,31,213,31,45,31,45,30,230,31,216,31,216,31,30,31,233,31,143,31,143,30,143,29,35,31,35,30,243,31,163,31,236,31,129,31,129,30,146,31,183,31,183,30,249,31,137,31,110,31,208,31,59,31,189,31,172,31,67,31,132,31,24,31,24,30,33,31,33,30,157,31,83,31,244,31,24,31,120,31,46,31,157,31,147,31,90,31,117,31,246,31,88,31,88,30,109,31,66,31,82,31,213,31,70,31,70,30,152,31,205,31,205,30,175,31,199,31,211,31,211,30,152,31,17,31,17,30,125,31,125,30,41,31,41,30,46,31,56,31,164,31,164,30,13,31,99,31,99,30,26,31,119,31,119,30,42,31,42,30,16,31,16,30,65,31,68,31,68,30,232,31,139,31,236,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
