-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 740;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,190,0,0,0,245,0,121,0,171,0,0,0,23,0,208,0,10,0,227,0,57,0,0,0,203,0,253,0,248,0,44,0,211,0,53,0,0,0,133,0,222,0,171,0,222,0,30,0,153,0,237,0,255,0,32,0,160,0,58,0,0,0,0,0,0,0,248,0,91,0,0,0,233,0,150,0,1,0,0,0,17,0,0,0,243,0,63,0,232,0,255,0,0,0,0,0,82,0,19,0,148,0,236,0,120,0,0,0,171,0,0,0,189,0,51,0,112,0,0,0,137,0,254,0,11,0,106,0,207,0,0,0,32,0,103,0,197,0,0,0,46,0,0,0,225,0,0,0,245,0,82,0,28,0,156,0,95,0,144,0,0,0,0,0,229,0,135,0,0,0,20,0,174,0,173,0,0,0,210,0,0,0,179,0,0,0,211,0,95,0,45,0,212,0,0,0,0,0,61,0,196,0,30,0,163,0,221,0,84,0,0,0,47,0,175,0,33,0,217,0,128,0,176,0,227,0,250,0,71,0,61,0,219,0,73,0,0,0,150,0,34,0,0,0,0,0,153,0,40,0,18,0,0,0,220,0,152,0,0,0,255,0,172,0,65,0,0,0,110,0,165,0,0,0,0,0,0,0,18,0,176,0,183,0,30,0,222,0,4,0,41,0,191,0,47,0,8,0,172,0,0,0,202,0,252,0,248,0,157,0,81,0,142,0,128,0,218,0,95,0,109,0,48,0,127,0,214,0,238,0,190,0,0,0,142,0,182,0,177,0,44,0,236,0,0,0,0,0,157,0,159,0,0,0,49,0,86,0,61,0,49,0,22,0,231,0,64,0,243,0,79,0,60,0,181,0,111,0,97,0,238,0,64,0,0,0,0,0,187,0,165,0,182,0,165,0,82,0,0,0,183,0,0,0,23,0,0,0,57,0,252,0,0,0,0,0,207,0,0,0,51,0,0,0,54,0,137,0,191,0,37,0,51,0,185,0,13,0,138,0,187,0,55,0,61,0,0,0,184,0,12,0,226,0,0,0,0,0,179,0,79,0,0,0,0,0,51,0,170,0,0,0,64,0,221,0,202,0,255,0,84,0,187,0,31,0,160,0,11,0,0,0,150,0,19,0,228,0,23,0,0,0,205,0,174,0,121,0,56,0,157,0,181,0,103,0,105,0,195,0,216,0,0,0,0,0,237,0,25,0,205,0,0,0,51,0,14,0,138,0,0,0,200,0,0,0,2,0,33,0,101,0,203,0,0,0,67,0,224,0,0,0,158,0,112,0,9,0,186,0,201,0,147,0,71,0,47,0,170,0,174,0,220,0,21,0,202,0,226,0,27,0,138,0,35,0,0,0,33,0,61,0,178,0,243,0,14,0,109,0,95,0,148,0,0,0,239,0,0,0,50,0,140,0,23,0,0,0,111,0,165,0,124,0,112,0,182,0,175,0,0,0,87,0,28,0,62,0,195,0,130,0,0,0,84,0,141,0,0,0,0,0,32,0,0,0,0,0,68,0,0,0,0,0,33,0,0,0,0,0,89,0,50,0,0,0,0,0,209,0,199,0,70,0,130,0,217,0,223,0,167,0,255,0,0,0,13,0,20,0,0,0,18,0,3,0,239,0,181,0,151,0,160,0,0,0,124,0,179,0,88,0,241,0,39,0,124,0,86,0,167,0,23,0,46,0,102,0,46,0,148,0,125,0,0,0,0,0,120,0,31,0,2,0,235,0,0,0,50,0,46,0,26,0,0,0,0,0,47,0,59,0,130,0,134,0,0,0,0,0,31,0,135,0,197,0,84,0,155,0,91,0,96,0,0,0,193,0,214,0,120,0,205,0,226,0,80,0,150,0,133,0,252,0,242,0,87,0,253,0,175,0,100,0,242,0,44,0,0,0,26,0,127,0,32,0,85,0,226,0,0,0,137,0,0,0,0,0,244,0,239,0,236,0,250,0,174,0,0,0,165,0,105,0,70,0,67,0,133,0,148,0,0,0,64,0,180,0,81,0,23,0,160,0,18,0,107,0,54,0,141,0,0,0,88,0,0,0,213,0,0,0,0,0,0,0,0,0,57,0,206,0,12,0,148,0,113,0,0,0,10,0,138,0,122,0,188,0,7,0,109,0,0,0,170,0,255,0,0,0,58,0,166,0,13,0,15,0,121,0,67,0,0,0,179,0,0,0,26,0,199,0,0,0,43,0,52,0,0,0,133,0,239,0,0,0,70,0,151,0,80,0,65,0,10,0,187,0,249,0,0,0,0,0,10,0,21,0,153,0,0,0,179,0,156,0,16,0,213,0,79,0,0,0,13,0,26,0,0,0,90,0,143,0,23,0,110,0,54,0,132,0,0,0,225,0,150,0,0,0,124,0,0,0,244,0,239,0,111,0,0,0,246,0,230,0,141,0,167,0,0,0,106,0,0,0,205,0,0,0,0,0,37,0,14,0,16,0,252,0,157,0,0,0,21,0,204,0,189,0,241,0,0,0,252,0,0,0,131,0,158,0,64,0,212,0,178,0,65,0,180,0,239,0,86,0,0,0,44,0,119,0,129,0,0,0,29,0,83,0,0,0,217,0,24,0,201,0,26,0,0,0,103,0,0,0,0,0,214,0,245,0,48,0,113,0,12,0,144,0,79,0,0,0,217,0,32,0,83,0,22,0,49,0,44,0,55,0,63,0,17,0,112,0,82,0,197,0,46,0,86,0,0,0,0,0,197,0,188,0,210,0,155,0,121,0,177,0,197,0,41,0,238,0,197,0,251,0,88,0,233,0,233,0,244,0,230,0,250,0,0,0,0,0,141,0,193,0,9,0,102,0,37,0,207,0,143,0,36,0,177,0,64,0,150,0,43,0,43,0,111,0,63,0,116,0,11,0,210,0,0,0,70,0,225,0,248,0,142,0,246,0,182,0,0,0,227,0,87,0,189,0,39,0,62,0,0,0,128,0,55,0,93,0,0,0,63,0,85,0,71,0,0,0,22,0,210,0,125,0,107,0,0,0,0,0,0,0,236,0,96,0,0,0,0,0,0,0,0,0,176,0,52,0,166,0,85,0,84,0,81,0,0,0,222,0,108,0,0,0,33,0,75,0,179,0,230,0,163,0,118,0,0,0,237,0,0,0,0,0,82,0,175,0,139,0,0,0,0,0,117,0,130,0,104,0,45,0,47,0,72,0,69,0,162,0,0,0,0,0,176,0,165,0,148,0,228,0,102,0,145,0,112,0,0,0,158,0,203,0,239,0,74,0,195,0,0,0,62,0,221,0,139,0,156,0,0,0,172,0,0,0,156,0,234,0,2,0,248,0,40,0,144,0,92,0,163,0);
signal scenario_full  : scenario_type := (181,31,190,31,190,30,245,31,121,31,171,31,171,30,23,31,208,31,10,31,227,31,57,31,57,30,203,31,253,31,248,31,44,31,211,31,53,31,53,30,133,31,222,31,171,31,222,31,30,31,153,31,237,31,255,31,32,31,160,31,58,31,58,30,58,29,58,28,248,31,91,31,91,30,233,31,150,31,1,31,1,30,17,31,17,30,243,31,63,31,232,31,255,31,255,30,255,29,82,31,19,31,148,31,236,31,120,31,120,30,171,31,171,30,189,31,51,31,112,31,112,30,137,31,254,31,11,31,106,31,207,31,207,30,32,31,103,31,197,31,197,30,46,31,46,30,225,31,225,30,245,31,82,31,28,31,156,31,95,31,144,31,144,30,144,29,229,31,135,31,135,30,20,31,174,31,173,31,173,30,210,31,210,30,179,31,179,30,211,31,95,31,45,31,212,31,212,30,212,29,61,31,196,31,30,31,163,31,221,31,84,31,84,30,47,31,175,31,33,31,217,31,128,31,176,31,227,31,250,31,71,31,61,31,219,31,73,31,73,30,150,31,34,31,34,30,34,29,153,31,40,31,18,31,18,30,220,31,152,31,152,30,255,31,172,31,65,31,65,30,110,31,165,31,165,30,165,29,165,28,18,31,176,31,183,31,30,31,222,31,4,31,41,31,191,31,47,31,8,31,172,31,172,30,202,31,252,31,248,31,157,31,81,31,142,31,128,31,218,31,95,31,109,31,48,31,127,31,214,31,238,31,190,31,190,30,142,31,182,31,177,31,44,31,236,31,236,30,236,29,157,31,159,31,159,30,49,31,86,31,61,31,49,31,22,31,231,31,64,31,243,31,79,31,60,31,181,31,111,31,97,31,238,31,64,31,64,30,64,29,187,31,165,31,182,31,165,31,82,31,82,30,183,31,183,30,23,31,23,30,57,31,252,31,252,30,252,29,207,31,207,30,51,31,51,30,54,31,137,31,191,31,37,31,51,31,185,31,13,31,138,31,187,31,55,31,61,31,61,30,184,31,12,31,226,31,226,30,226,29,179,31,79,31,79,30,79,29,51,31,170,31,170,30,64,31,221,31,202,31,255,31,84,31,187,31,31,31,160,31,11,31,11,30,150,31,19,31,228,31,23,31,23,30,205,31,174,31,121,31,56,31,157,31,181,31,103,31,105,31,195,31,216,31,216,30,216,29,237,31,25,31,205,31,205,30,51,31,14,31,138,31,138,30,200,31,200,30,2,31,33,31,101,31,203,31,203,30,67,31,224,31,224,30,158,31,112,31,9,31,186,31,201,31,147,31,71,31,47,31,170,31,174,31,220,31,21,31,202,31,226,31,27,31,138,31,35,31,35,30,33,31,61,31,178,31,243,31,14,31,109,31,95,31,148,31,148,30,239,31,239,30,50,31,140,31,23,31,23,30,111,31,165,31,124,31,112,31,182,31,175,31,175,30,87,31,28,31,62,31,195,31,130,31,130,30,84,31,141,31,141,30,141,29,32,31,32,30,32,29,68,31,68,30,68,29,33,31,33,30,33,29,89,31,50,31,50,30,50,29,209,31,199,31,70,31,130,31,217,31,223,31,167,31,255,31,255,30,13,31,20,31,20,30,18,31,3,31,239,31,181,31,151,31,160,31,160,30,124,31,179,31,88,31,241,31,39,31,124,31,86,31,167,31,23,31,46,31,102,31,46,31,148,31,125,31,125,30,125,29,120,31,31,31,2,31,235,31,235,30,50,31,46,31,26,31,26,30,26,29,47,31,59,31,130,31,134,31,134,30,134,29,31,31,135,31,197,31,84,31,155,31,91,31,96,31,96,30,193,31,214,31,120,31,205,31,226,31,80,31,150,31,133,31,252,31,242,31,87,31,253,31,175,31,100,31,242,31,44,31,44,30,26,31,127,31,32,31,85,31,226,31,226,30,137,31,137,30,137,29,244,31,239,31,236,31,250,31,174,31,174,30,165,31,105,31,70,31,67,31,133,31,148,31,148,30,64,31,180,31,81,31,23,31,160,31,18,31,107,31,54,31,141,31,141,30,88,31,88,30,213,31,213,30,213,29,213,28,213,27,57,31,206,31,12,31,148,31,113,31,113,30,10,31,138,31,122,31,188,31,7,31,109,31,109,30,170,31,255,31,255,30,58,31,166,31,13,31,15,31,121,31,67,31,67,30,179,31,179,30,26,31,199,31,199,30,43,31,52,31,52,30,133,31,239,31,239,30,70,31,151,31,80,31,65,31,10,31,187,31,249,31,249,30,249,29,10,31,21,31,153,31,153,30,179,31,156,31,16,31,213,31,79,31,79,30,13,31,26,31,26,30,90,31,143,31,23,31,110,31,54,31,132,31,132,30,225,31,150,31,150,30,124,31,124,30,244,31,239,31,111,31,111,30,246,31,230,31,141,31,167,31,167,30,106,31,106,30,205,31,205,30,205,29,37,31,14,31,16,31,252,31,157,31,157,30,21,31,204,31,189,31,241,31,241,30,252,31,252,30,131,31,158,31,64,31,212,31,178,31,65,31,180,31,239,31,86,31,86,30,44,31,119,31,129,31,129,30,29,31,83,31,83,30,217,31,24,31,201,31,26,31,26,30,103,31,103,30,103,29,214,31,245,31,48,31,113,31,12,31,144,31,79,31,79,30,217,31,32,31,83,31,22,31,49,31,44,31,55,31,63,31,17,31,112,31,82,31,197,31,46,31,86,31,86,30,86,29,197,31,188,31,210,31,155,31,121,31,177,31,197,31,41,31,238,31,197,31,251,31,88,31,233,31,233,31,244,31,230,31,250,31,250,30,250,29,141,31,193,31,9,31,102,31,37,31,207,31,143,31,36,31,177,31,64,31,150,31,43,31,43,31,111,31,63,31,116,31,11,31,210,31,210,30,70,31,225,31,248,31,142,31,246,31,182,31,182,30,227,31,87,31,189,31,39,31,62,31,62,30,128,31,55,31,93,31,93,30,63,31,85,31,71,31,71,30,22,31,210,31,125,31,107,31,107,30,107,29,107,28,236,31,96,31,96,30,96,29,96,28,96,27,176,31,52,31,166,31,85,31,84,31,81,31,81,30,222,31,108,31,108,30,33,31,75,31,179,31,230,31,163,31,118,31,118,30,237,31,237,30,237,29,82,31,175,31,139,31,139,30,139,29,117,31,130,31,104,31,45,31,47,31,72,31,69,31,162,31,162,30,162,29,176,31,165,31,148,31,228,31,102,31,145,31,112,31,112,30,158,31,203,31,239,31,74,31,195,31,195,30,62,31,221,31,139,31,156,31,156,30,172,31,172,30,156,31,234,31,2,31,248,31,40,31,144,31,92,31,163,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
