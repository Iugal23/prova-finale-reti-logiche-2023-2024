-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 908;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,230,0,0,0,117,0,0,0,21,0,0,0,131,0,56,0,172,0,193,0,215,0,15,0,237,0,29,0,228,0,0,0,231,0,163,0,245,0,71,0,96,0,165,0,94,0,72,0,0,0,226,0,0,0,34,0,146,0,238,0,139,0,156,0,168,0,2,0,173,0,81,0,53,0,0,0,30,0,156,0,0,0,0,0,122,0,247,0,0,0,0,0,0,0,211,0,25,0,243,0,0,0,118,0,199,0,71,0,131,0,196,0,152,0,53,0,52,0,24,0,41,0,203,0,0,0,219,0,97,0,40,0,240,0,231,0,161,0,121,0,0,0,0,0,0,0,53,0,182,0,206,0,23,0,62,0,211,0,67,0,43,0,19,0,28,0,194,0,31,0,219,0,26,0,0,0,0,0,99,0,85,0,197,0,221,0,242,0,0,0,236,0,0,0,9,0,85,0,17,0,127,0,109,0,208,0,73,0,0,0,17,0,74,0,149,0,11,0,93,0,0,0,161,0,21,0,238,0,255,0,92,0,204,0,27,0,233,0,4,0,141,0,0,0,223,0,27,0,109,0,176,0,111,0,101,0,187,0,102,0,26,0,0,0,87,0,127,0,171,0,162,0,38,0,175,0,159,0,221,0,58,0,0,0,0,0,131,0,55,0,0,0,0,0,186,0,104,0,102,0,0,0,0,0,156,0,218,0,0,0,176,0,50,0,27,0,255,0,148,0,63,0,79,0,0,0,0,0,202,0,11,0,0,0,112,0,193,0,4,0,0,0,0,0,61,0,0,0,120,0,194,0,82,0,53,0,63,0,99,0,0,0,141,0,18,0,235,0,163,0,80,0,241,0,12,0,207,0,140,0,131,0,156,0,52,0,0,0,127,0,190,0,176,0,247,0,251,0,227,0,142,0,166,0,120,0,95,0,218,0,50,0,131,0,136,0,15,0,216,0,0,0,51,0,59,0,63,0,0,0,108,0,2,0,26,0,152,0,100,0,243,0,0,0,68,0,68,0,154,0,121,0,0,0,36,0,0,0,0,0,175,0,240,0,140,0,0,0,0,0,0,0,125,0,110,0,0,0,207,0,183,0,5,0,220,0,9,0,197,0,122,0,32,0,220,0,218,0,0,0,29,0,66,0,237,0,119,0,122,0,99,0,132,0,155,0,0,0,0,0,219,0,215,0,211,0,80,0,47,0,20,0,188,0,13,0,174,0,226,0,0,0,90,0,253,0,135,0,144,0,62,0,0,0,24,0,53,0,0,0,8,0,182,0,78,0,167,0,30,0,123,0,0,0,51,0,178,0,18,0,113,0,43,0,0,0,115,0,197,0,203,0,95,0,0,0,203,0,118,0,174,0,200,0,0,0,126,0,126,0,112,0,206,0,147,0,237,0,127,0,134,0,27,0,0,0,55,0,42,0,246,0,230,0,20,0,161,0,184,0,60,0,45,0,193,0,178,0,0,0,164,0,133,0,24,0,81,0,197,0,199,0,222,0,26,0,57,0,0,0,159,0,182,0,63,0,168,0,120,0,72,0,221,0,48,0,6,0,47,0,86,0,89,0,14,0,0,0,0,0,135,0,43,0,176,0,135,0,227,0,125,0,0,0,122,0,0,0,236,0,172,0,73,0,251,0,33,0,141,0,142,0,189,0,179,0,109,0,83,0,118,0,0,0,120,0,180,0,154,0,41,0,160,0,43,0,157,0,239,0,124,0,139,0,184,0,228,0,0,0,179,0,252,0,0,0,0,0,226,0,13,0,0,0,120,0,94,0,247,0,33,0,221,0,114,0,0,0,170,0,53,0,2,0,132,0,233,0,242,0,215,0,195,0,0,0,187,0,251,0,81,0,53,0,85,0,229,0,241,0,0,0,177,0,210,0,207,0,194,0,225,0,15,0,122,0,233,0,0,0,41,0,0,0,112,0,1,0,92,0,145,0,213,0,168,0,254,0,0,0,0,0,127,0,0,0,224,0,0,0,209,0,0,0,68,0,93,0,0,0,212,0,241,0,91,0,223,0,225,0,228,0,106,0,232,0,89,0,128,0,0,0,57,0,42,0,144,0,201,0,150,0,147,0,0,0,206,0,84,0,0,0,0,0,244,0,55,0,16,0,245,0,188,0,217,0,197,0,250,0,165,0,249,0,49,0,189,0,136,0,137,0,243,0,203,0,130,0,130,0,0,0,232,0,40,0,57,0,137,0,26,0,43,0,145,0,248,0,142,0,255,0,182,0,192,0,228,0,169,0,170,0,188,0,205,0,20,0,250,0,189,0,86,0,79,0,211,0,166,0,160,0,0,0,101,0,35,0,0,0,38,0,120,0,50,0,179,0,140,0,0,0,188,0,130,0,7,0,247,0,210,0,50,0,239,0,161,0,72,0,0,0,225,0,73,0,42,0,0,0,103,0,142,0,0,0,158,0,155,0,223,0,84,0,111,0,196,0,139,0,0,0,31,0,140,0,155,0,105,0,0,0,63,0,51,0,0,0,17,0,0,0,165,0,61,0,23,0,238,0,130,0,0,0,159,0,1,0,255,0,145,0,0,0,0,0,0,0,26,0,111,0,119,0,195,0,218,0,207,0,72,0,13,0,83,0,110,0,173,0,188,0,246,0,101,0,231,0,168,0,0,0,113,0,169,0,164,0,57,0,153,0,0,0,102,0,0,0,207,0,183,0,234,0,122,0,0,0,229,0,66,0,201,0,252,0,83,0,187,0,0,0,200,0,0,0,192,0,0,0,0,0,102,0,92,0,178,0,189,0,44,0,0,0,225,0,235,0,249,0,90,0,190,0,18,0,231,0,156,0,0,0,73,0,0,0,237,0,65,0,26,0,0,0,123,0,120,0,173,0,0,0,0,0,106,0,12,0,79,0,0,0,0,0,11,0,0,0,12,0,48,0,171,0,77,0,0,0,164,0,93,0,0,0,152,0,99,0,0,0,165,0,90,0,242,0,71,0,151,0,40,0,105,0,226,0,115,0,0,0,232,0,219,0,193,0,207,0,36,0,180,0,145,0,8,0,10,0,0,0,0,0,0,0,47,0,3,0,65,0,62,0,0,0,134,0,0,0,249,0,139,0,178,0,142,0,144,0,44,0,235,0,61,0,0,0,41,0,0,0,46,0,152,0,179,0,199,0,16,0,212,0,0,0,111,0,108,0,91,0,0,0,32,0,0,0,87,0,4,0,172,0,242,0,31,0,191,0,111,0,76,0,160,0,62,0,0,0,250,0,65,0,211,0,106,0,142,0,71,0,171,0,5,0,99,0,66,0,0,0,0,0,0,0,58,0,190,0,63,0,176,0,182,0,211,0,0,0,200,0,67,0,166,0,164,0,0,0,3,0,83,0,43,0,193,0,194,0,125,0,115,0,215,0,195,0,31,0,49,0,111,0,27,0,134,0,135,0,85,0,31,0,0,0,81,0,173,0,241,0,130,0,146,0,218,0,0,0,0,0,97,0,241,0,45,0,195,0,130,0,0,0,124,0,0,0,109,0,3,0,15,0,120,0,120,0,4,0,0,0,115,0,0,0,237,0,0,0,0,0,237,0,93,0,12,0,137,0,0,0,169,0,49,0,221,0,199,0,0,0,11,0,126,0,48,0,167,0,20,0,171,0,22,0,246,0,40,0,76,0,189,0,127,0,0,0,0,0,0,0,203,0,132,0,96,0,169,0,216,0,0,0,116,0,199,0,43,0,230,0,25,0,210,0,90,0,44,0,3,0,19,0,158,0,64,0,203,0,20,0,168,0,0,0,152,0,42,0,96,0,246,0,39,0,0,0,84,0,230,0,252,0,142,0,87,0,170,0,0,0,0,0,64,0,0,0,213,0,0,0,70,0,189,0,0,0,3,0,28,0,215,0,253,0,0,0,197,0,48,0,225,0,125,0,149,0,5,0,224,0,21,0,193,0,232,0,148,0,138,0,118,0,20,0,0,0,123,0,161,0,68,0,215,0,252,0,178,0,23,0,51,0,0,0,70,0,199,0,133,0,6,0,164,0,17,0,207,0,254,0,204,0,41,0,0,0,191,0,34,0,29,0,200,0,185,0,83,0,243,0,120,0,0,0);
signal scenario_full  : scenario_type := (6,31,230,31,230,30,117,31,117,30,21,31,21,30,131,31,56,31,172,31,193,31,215,31,15,31,237,31,29,31,228,31,228,30,231,31,163,31,245,31,71,31,96,31,165,31,94,31,72,31,72,30,226,31,226,30,34,31,146,31,238,31,139,31,156,31,168,31,2,31,173,31,81,31,53,31,53,30,30,31,156,31,156,30,156,29,122,31,247,31,247,30,247,29,247,28,211,31,25,31,243,31,243,30,118,31,199,31,71,31,131,31,196,31,152,31,53,31,52,31,24,31,41,31,203,31,203,30,219,31,97,31,40,31,240,31,231,31,161,31,121,31,121,30,121,29,121,28,53,31,182,31,206,31,23,31,62,31,211,31,67,31,43,31,19,31,28,31,194,31,31,31,219,31,26,31,26,30,26,29,99,31,85,31,197,31,221,31,242,31,242,30,236,31,236,30,9,31,85,31,17,31,127,31,109,31,208,31,73,31,73,30,17,31,74,31,149,31,11,31,93,31,93,30,161,31,21,31,238,31,255,31,92,31,204,31,27,31,233,31,4,31,141,31,141,30,223,31,27,31,109,31,176,31,111,31,101,31,187,31,102,31,26,31,26,30,87,31,127,31,171,31,162,31,38,31,175,31,159,31,221,31,58,31,58,30,58,29,131,31,55,31,55,30,55,29,186,31,104,31,102,31,102,30,102,29,156,31,218,31,218,30,176,31,50,31,27,31,255,31,148,31,63,31,79,31,79,30,79,29,202,31,11,31,11,30,112,31,193,31,4,31,4,30,4,29,61,31,61,30,120,31,194,31,82,31,53,31,63,31,99,31,99,30,141,31,18,31,235,31,163,31,80,31,241,31,12,31,207,31,140,31,131,31,156,31,52,31,52,30,127,31,190,31,176,31,247,31,251,31,227,31,142,31,166,31,120,31,95,31,218,31,50,31,131,31,136,31,15,31,216,31,216,30,51,31,59,31,63,31,63,30,108,31,2,31,26,31,152,31,100,31,243,31,243,30,68,31,68,31,154,31,121,31,121,30,36,31,36,30,36,29,175,31,240,31,140,31,140,30,140,29,140,28,125,31,110,31,110,30,207,31,183,31,5,31,220,31,9,31,197,31,122,31,32,31,220,31,218,31,218,30,29,31,66,31,237,31,119,31,122,31,99,31,132,31,155,31,155,30,155,29,219,31,215,31,211,31,80,31,47,31,20,31,188,31,13,31,174,31,226,31,226,30,90,31,253,31,135,31,144,31,62,31,62,30,24,31,53,31,53,30,8,31,182,31,78,31,167,31,30,31,123,31,123,30,51,31,178,31,18,31,113,31,43,31,43,30,115,31,197,31,203,31,95,31,95,30,203,31,118,31,174,31,200,31,200,30,126,31,126,31,112,31,206,31,147,31,237,31,127,31,134,31,27,31,27,30,55,31,42,31,246,31,230,31,20,31,161,31,184,31,60,31,45,31,193,31,178,31,178,30,164,31,133,31,24,31,81,31,197,31,199,31,222,31,26,31,57,31,57,30,159,31,182,31,63,31,168,31,120,31,72,31,221,31,48,31,6,31,47,31,86,31,89,31,14,31,14,30,14,29,135,31,43,31,176,31,135,31,227,31,125,31,125,30,122,31,122,30,236,31,172,31,73,31,251,31,33,31,141,31,142,31,189,31,179,31,109,31,83,31,118,31,118,30,120,31,180,31,154,31,41,31,160,31,43,31,157,31,239,31,124,31,139,31,184,31,228,31,228,30,179,31,252,31,252,30,252,29,226,31,13,31,13,30,120,31,94,31,247,31,33,31,221,31,114,31,114,30,170,31,53,31,2,31,132,31,233,31,242,31,215,31,195,31,195,30,187,31,251,31,81,31,53,31,85,31,229,31,241,31,241,30,177,31,210,31,207,31,194,31,225,31,15,31,122,31,233,31,233,30,41,31,41,30,112,31,1,31,92,31,145,31,213,31,168,31,254,31,254,30,254,29,127,31,127,30,224,31,224,30,209,31,209,30,68,31,93,31,93,30,212,31,241,31,91,31,223,31,225,31,228,31,106,31,232,31,89,31,128,31,128,30,57,31,42,31,144,31,201,31,150,31,147,31,147,30,206,31,84,31,84,30,84,29,244,31,55,31,16,31,245,31,188,31,217,31,197,31,250,31,165,31,249,31,49,31,189,31,136,31,137,31,243,31,203,31,130,31,130,31,130,30,232,31,40,31,57,31,137,31,26,31,43,31,145,31,248,31,142,31,255,31,182,31,192,31,228,31,169,31,170,31,188,31,205,31,20,31,250,31,189,31,86,31,79,31,211,31,166,31,160,31,160,30,101,31,35,31,35,30,38,31,120,31,50,31,179,31,140,31,140,30,188,31,130,31,7,31,247,31,210,31,50,31,239,31,161,31,72,31,72,30,225,31,73,31,42,31,42,30,103,31,142,31,142,30,158,31,155,31,223,31,84,31,111,31,196,31,139,31,139,30,31,31,140,31,155,31,105,31,105,30,63,31,51,31,51,30,17,31,17,30,165,31,61,31,23,31,238,31,130,31,130,30,159,31,1,31,255,31,145,31,145,30,145,29,145,28,26,31,111,31,119,31,195,31,218,31,207,31,72,31,13,31,83,31,110,31,173,31,188,31,246,31,101,31,231,31,168,31,168,30,113,31,169,31,164,31,57,31,153,31,153,30,102,31,102,30,207,31,183,31,234,31,122,31,122,30,229,31,66,31,201,31,252,31,83,31,187,31,187,30,200,31,200,30,192,31,192,30,192,29,102,31,92,31,178,31,189,31,44,31,44,30,225,31,235,31,249,31,90,31,190,31,18,31,231,31,156,31,156,30,73,31,73,30,237,31,65,31,26,31,26,30,123,31,120,31,173,31,173,30,173,29,106,31,12,31,79,31,79,30,79,29,11,31,11,30,12,31,48,31,171,31,77,31,77,30,164,31,93,31,93,30,152,31,99,31,99,30,165,31,90,31,242,31,71,31,151,31,40,31,105,31,226,31,115,31,115,30,232,31,219,31,193,31,207,31,36,31,180,31,145,31,8,31,10,31,10,30,10,29,10,28,47,31,3,31,65,31,62,31,62,30,134,31,134,30,249,31,139,31,178,31,142,31,144,31,44,31,235,31,61,31,61,30,41,31,41,30,46,31,152,31,179,31,199,31,16,31,212,31,212,30,111,31,108,31,91,31,91,30,32,31,32,30,87,31,4,31,172,31,242,31,31,31,191,31,111,31,76,31,160,31,62,31,62,30,250,31,65,31,211,31,106,31,142,31,71,31,171,31,5,31,99,31,66,31,66,30,66,29,66,28,58,31,190,31,63,31,176,31,182,31,211,31,211,30,200,31,67,31,166,31,164,31,164,30,3,31,83,31,43,31,193,31,194,31,125,31,115,31,215,31,195,31,31,31,49,31,111,31,27,31,134,31,135,31,85,31,31,31,31,30,81,31,173,31,241,31,130,31,146,31,218,31,218,30,218,29,97,31,241,31,45,31,195,31,130,31,130,30,124,31,124,30,109,31,3,31,15,31,120,31,120,31,4,31,4,30,115,31,115,30,237,31,237,30,237,29,237,31,93,31,12,31,137,31,137,30,169,31,49,31,221,31,199,31,199,30,11,31,126,31,48,31,167,31,20,31,171,31,22,31,246,31,40,31,76,31,189,31,127,31,127,30,127,29,127,28,203,31,132,31,96,31,169,31,216,31,216,30,116,31,199,31,43,31,230,31,25,31,210,31,90,31,44,31,3,31,19,31,158,31,64,31,203,31,20,31,168,31,168,30,152,31,42,31,96,31,246,31,39,31,39,30,84,31,230,31,252,31,142,31,87,31,170,31,170,30,170,29,64,31,64,30,213,31,213,30,70,31,189,31,189,30,3,31,28,31,215,31,253,31,253,30,197,31,48,31,225,31,125,31,149,31,5,31,224,31,21,31,193,31,232,31,148,31,138,31,118,31,20,31,20,30,123,31,161,31,68,31,215,31,252,31,178,31,23,31,51,31,51,30,70,31,199,31,133,31,6,31,164,31,17,31,207,31,254,31,204,31,41,31,41,30,191,31,34,31,29,31,200,31,185,31,83,31,243,31,120,31,120,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
