-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 420;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,196,0,141,0,140,0,193,0,152,0,36,0,166,0,0,0,154,0,93,0,255,0,89,0,106,0,116,0,43,0,86,0,10,0,73,0,183,0,167,0,205,0,27,0,10,0,113,0,0,0,87,0,19,0,247,0,161,0,79,0,35,0,77,0,17,0,195,0,14,0,51,0,43,0,0,0,0,0,57,0,27,0,184,0,53,0,162,0,186,0,0,0,0,0,0,0,212,0,0,0,54,0,76,0,215,0,200,0,230,0,233,0,3,0,49,0,51,0,0,0,98,0,192,0,69,0,10,0,179,0,48,0,236,0,34,0,86,0,246,0,117,0,224,0,168,0,232,0,199,0,0,0,218,0,162,0,244,0,230,0,92,0,0,0,104,0,106,0,0,0,235,0,226,0,186,0,38,0,210,0,33,0,0,0,177,0,141,0,72,0,187,0,170,0,221,0,130,0,0,0,218,0,202,0,252,0,124,0,227,0,0,0,166,0,71,0,70,0,22,0,39,0,139,0,92,0,188,0,0,0,46,0,102,0,145,0,101,0,140,0,0,0,15,0,27,0,0,0,80,0,89,0,84,0,0,0,83,0,0,0,125,0,139,0,17,0,0,0,86,0,204,0,160,0,255,0,69,0,146,0,228,0,206,0,47,0,226,0,64,0,0,0,48,0,208,0,50,0,89,0,94,0,34,0,113,0,8,0,0,0,0,0,228,0,250,0,0,0,49,0,79,0,101,0,79,0,25,0,178,0,232,0,144,0,0,0,174,0,0,0,106,0,133,0,237,0,100,0,191,0,190,0,0,0,0,0,0,0,0,0,10,0,0,0,220,0,251,0,0,0,33,0,167,0,116,0,67,0,0,0,44,0,131,0,70,0,18,0,216,0,0,0,46,0,174,0,254,0,176,0,76,0,50,0,132,0,0,0,31,0,0,0,251,0,38,0,99,0,90,0,86,0,171,0,89,0,131,0,0,0,97,0,0,0,141,0,135,0,0,0,97,0,229,0,11,0,201,0,207,0,0,0,150,0,163,0,89,0,39,0,157,0,189,0,57,0,24,0,24,0,62,0,0,0,158,0,168,0,90,0,135,0,218,0,116,0,50,0,32,0,229,0,130,0,0,0,36,0,143,0,100,0,155,0,247,0,157,0,93,0,83,0,205,0,181,0,57,0,146,0,169,0,0,0,33,0,228,0,7,0,45,0,41,0,227,0,74,0,26,0,47,0,143,0,0,0,0,0,0,0,0,0,74,0,0,0,170,0,125,0,241,0,247,0,161,0,0,0,210,0,153,0,232,0,111,0,19,0,40,0,0,0,252,0,0,0,37,0,243,0,19,0,162,0,104,0,139,0,75,0,1,0,8,0,76,0,161,0,248,0,87,0,0,0,36,0,50,0,193,0,0,0,247,0,75,0,165,0,81,0,34,0,155,0,116,0,140,0,144,0,75,0,187,0,41,0,0,0,0,0,72,0,253,0,0,0,239,0,236,0,158,0,0,0,99,0,249,0,90,0,81,0,132,0,107,0,126,0,0,0,197,0,115,0,49,0,0,0,229,0,74,0,66,0,0,0,136,0,47,0,233,0,243,0,70,0,0,0,206,0,150,0,67,0,212,0,32,0,29,0,78,0,0,0,44,0,14,0,0,0,85,0,158,0,17,0,0,0,193,0,157,0,0,0,160,0,87,0,16,0,168,0,159,0,0,0,160,0,92,0,92,0,96,0,235,0,0,0,14,0,105,0,141,0,0,0,0,0,0,0,162,0,69,0,157,0,29,0,188,0,222,0,219,0,71,0,212,0,0,0,115,0,159,0,23,0,194,0,210,0,35,0,249,0,68,0,96,0,0,0,82,0,50,0,139,0,107,0,63,0,178,0,0,0,0,0,214,0);
signal scenario_full  : scenario_type := (0,0,196,31,141,31,140,31,193,31,152,31,36,31,166,31,166,30,154,31,93,31,255,31,89,31,106,31,116,31,43,31,86,31,10,31,73,31,183,31,167,31,205,31,27,31,10,31,113,31,113,30,87,31,19,31,247,31,161,31,79,31,35,31,77,31,17,31,195,31,14,31,51,31,43,31,43,30,43,29,57,31,27,31,184,31,53,31,162,31,186,31,186,30,186,29,186,28,212,31,212,30,54,31,76,31,215,31,200,31,230,31,233,31,3,31,49,31,51,31,51,30,98,31,192,31,69,31,10,31,179,31,48,31,236,31,34,31,86,31,246,31,117,31,224,31,168,31,232,31,199,31,199,30,218,31,162,31,244,31,230,31,92,31,92,30,104,31,106,31,106,30,235,31,226,31,186,31,38,31,210,31,33,31,33,30,177,31,141,31,72,31,187,31,170,31,221,31,130,31,130,30,218,31,202,31,252,31,124,31,227,31,227,30,166,31,71,31,70,31,22,31,39,31,139,31,92,31,188,31,188,30,46,31,102,31,145,31,101,31,140,31,140,30,15,31,27,31,27,30,80,31,89,31,84,31,84,30,83,31,83,30,125,31,139,31,17,31,17,30,86,31,204,31,160,31,255,31,69,31,146,31,228,31,206,31,47,31,226,31,64,31,64,30,48,31,208,31,50,31,89,31,94,31,34,31,113,31,8,31,8,30,8,29,228,31,250,31,250,30,49,31,79,31,101,31,79,31,25,31,178,31,232,31,144,31,144,30,174,31,174,30,106,31,133,31,237,31,100,31,191,31,190,31,190,30,190,29,190,28,190,27,10,31,10,30,220,31,251,31,251,30,33,31,167,31,116,31,67,31,67,30,44,31,131,31,70,31,18,31,216,31,216,30,46,31,174,31,254,31,176,31,76,31,50,31,132,31,132,30,31,31,31,30,251,31,38,31,99,31,90,31,86,31,171,31,89,31,131,31,131,30,97,31,97,30,141,31,135,31,135,30,97,31,229,31,11,31,201,31,207,31,207,30,150,31,163,31,89,31,39,31,157,31,189,31,57,31,24,31,24,31,62,31,62,30,158,31,168,31,90,31,135,31,218,31,116,31,50,31,32,31,229,31,130,31,130,30,36,31,143,31,100,31,155,31,247,31,157,31,93,31,83,31,205,31,181,31,57,31,146,31,169,31,169,30,33,31,228,31,7,31,45,31,41,31,227,31,74,31,26,31,47,31,143,31,143,30,143,29,143,28,143,27,74,31,74,30,170,31,125,31,241,31,247,31,161,31,161,30,210,31,153,31,232,31,111,31,19,31,40,31,40,30,252,31,252,30,37,31,243,31,19,31,162,31,104,31,139,31,75,31,1,31,8,31,76,31,161,31,248,31,87,31,87,30,36,31,50,31,193,31,193,30,247,31,75,31,165,31,81,31,34,31,155,31,116,31,140,31,144,31,75,31,187,31,41,31,41,30,41,29,72,31,253,31,253,30,239,31,236,31,158,31,158,30,99,31,249,31,90,31,81,31,132,31,107,31,126,31,126,30,197,31,115,31,49,31,49,30,229,31,74,31,66,31,66,30,136,31,47,31,233,31,243,31,70,31,70,30,206,31,150,31,67,31,212,31,32,31,29,31,78,31,78,30,44,31,14,31,14,30,85,31,158,31,17,31,17,30,193,31,157,31,157,30,160,31,87,31,16,31,168,31,159,31,159,30,160,31,92,31,92,31,96,31,235,31,235,30,14,31,105,31,141,31,141,30,141,29,141,28,162,31,69,31,157,31,29,31,188,31,222,31,219,31,71,31,212,31,212,30,115,31,159,31,23,31,194,31,210,31,35,31,249,31,68,31,96,31,96,30,82,31,50,31,139,31,107,31,63,31,178,31,178,30,178,29,214,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
