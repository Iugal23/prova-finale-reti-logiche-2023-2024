-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 674;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,30,0,15,0,57,0,138,0,105,0,0,0,140,0,104,0,109,0,57,0,74,0,110,0,187,0,107,0,24,0,35,0,17,0,240,0,0,0,219,0,83,0,70,0,0,0,47,0,155,0,115,0,0,0,79,0,0,0,19,0,210,0,219,0,63,0,136,0,122,0,164,0,137,0,108,0,37,0,0,0,194,0,27,0,129,0,0,0,239,0,30,0,0,0,251,0,250,0,134,0,47,0,165,0,243,0,0,0,153,0,43,0,36,0,0,0,77,0,157,0,170,0,33,0,38,0,149,0,83,0,72,0,42,0,126,0,119,0,0,0,168,0,0,0,0,0,190,0,226,0,185,0,198,0,147,0,153,0,25,0,0,0,100,0,0,0,185,0,12,0,44,0,226,0,126,0,0,0,236,0,117,0,203,0,109,0,156,0,75,0,0,0,0,0,135,0,83,0,106,0,178,0,199,0,0,0,0,0,193,0,60,0,249,0,83,0,60,0,56,0,154,0,0,0,0,0,68,0,159,0,203,0,102,0,232,0,27,0,43,0,213,0,156,0,54,0,4,0,46,0,65,0,231,0,150,0,14,0,0,0,158,0,224,0,91,0,139,0,132,0,0,0,74,0,66,0,0,0,126,0,21,0,209,0,194,0,244,0,0,0,0,0,0,0,0,0,243,0,0,0,242,0,0,0,29,0,1,0,31,0,181,0,236,0,70,0,15,0,0,0,190,0,2,0,237,0,124,0,0,0,118,0,29,0,15,0,17,0,183,0,15,0,210,0,190,0,129,0,111,0,0,0,50,0,11,0,117,0,182,0,93,0,245,0,0,0,0,0,75,0,0,0,104,0,0,0,143,0,145,0,117,0,230,0,0,0,248,0,213,0,234,0,240,0,251,0,115,0,59,0,0,0,89,0,206,0,77,0,11,0,88,0,66,0,0,0,228,0,0,0,198,0,0,0,126,0,197,0,175,0,143,0,132,0,0,0,222,0,245,0,79,0,163,0,107,0,188,0,213,0,49,0,17,0,146,0,197,0,3,0,107,0,91,0,86,0,240,0,156,0,0,0,246,0,0,0,0,0,118,0,0,0,18,0,221,0,0,0,244,0,0,0,142,0,230,0,228,0,147,0,218,0,248,0,0,0,239,0,116,0,127,0,0,0,213,0,103,0,28,0,0,0,55,0,155,0,84,0,192,0,88,0,82,0,162,0,3,0,87,0,0,0,0,0,130,0,16,0,61,0,218,0,0,0,143,0,224,0,15,0,0,0,25,0,155,0,63,0,113,0,113,0,94,0,253,0,244,0,219,0,139,0,222,0,102,0,2,0,241,0,94,0,110,0,244,0,0,0,56,0,95,0,0,0,41,0,0,0,114,0,162,0,137,0,101,0,0,0,49,0,0,0,187,0,134,0,0,0,14,0,130,0,219,0,29,0,237,0,120,0,181,0,0,0,203,0,13,0,174,0,201,0,78,0,0,0,1,0,158,0,91,0,0,0,215,0,0,0,239,0,191,0,139,0,133,0,0,0,50,0,156,0,110,0,233,0,241,0,182,0,55,0,122,0,0,0,0,0,167,0,107,0,188,0,0,0,116,0,201,0,0,0,96,0,28,0,83,0,156,0,105,0,96,0,0,0,114,0,0,0,91,0,103,0,0,0,0,0,245,0,0,0,214,0,228,0,25,0,242,0,212,0,97,0,155,0,95,0,213,0,45,0,217,0,126,0,245,0,195,0,4,0,223,0,98,0,100,0,183,0,12,0,181,0,55,0,58,0,75,0,80,0,0,0,182,0,161,0,29,0,125,0,140,0,0,0,0,0,83,0,183,0,114,0,236,0,54,0,156,0,0,0,17,0,175,0,0,0,0,0,190,0,182,0,228,0,214,0,244,0,0,0,117,0,219,0,81,0,232,0,64,0,205,0,105,0,163,0,71,0,0,0,14,0,216,0,145,0,103,0,220,0,205,0,56,0,141,0,199,0,30,0,0,0,104,0,0,0,15,0,62,0,189,0,186,0,151,0,68,0,130,0,64,0,175,0,206,0,71,0,164,0,86,0,23,0,0,0,82,0,0,0,199,0,244,0,83,0,245,0,0,0,101,0,213,0,148,0,223,0,169,0,37,0,0,0,230,0,198,0,41,0,16,0,176,0,144,0,216,0,168,0,124,0,93,0,59,0,107,0,251,0,8,0,95,0,112,0,160,0,6,0,177,0,28,0,239,0,31,0,32,0,232,0,0,0,145,0,16,0,102,0,177,0,19,0,216,0,119,0,26,0,177,0,0,0,171,0,202,0,57,0,0,0,134,0,73,0,72,0,138,0,166,0,0,0,182,0,112,0,211,0,38,0,181,0,0,0,244,0,16,0,58,0,0,0,157,0,73,0,199,0,67,0,108,0,243,0,34,0,31,0,117,0,163,0,196,0,31,0,0,0,147,0,194,0,175,0,224,0,12,0,93,0,152,0,25,0,228,0,255,0,77,0,231,0,26,0,245,0,10,0,207,0,0,0,35,0,124,0,146,0,25,0,191,0,154,0,0,0,241,0,196,0,243,0,0,0,7,0,232,0,208,0,15,0,230,0,190,0,176,0,207,0,6,0,67,0,0,0,139,0,251,0,78,0,205,0,64,0,74,0,73,0,0,0,0,0,0,0,236,0,44,0,0,0,141,0,33,0,106,0,0,0,20,0,29,0,210,0,48,0,133,0,6,0,23,0,67,0,89,0,196,0,47,0,13,0,158,0,75,0,213,0,19,0,207,0,27,0,187,0,85,0,91,0,168,0,149,0,92,0,30,0,0,0,255,0,116,0,231,0,92,0,137,0,123,0,114,0,27,0,0,0,225,0,60,0,112,0,205,0,124,0,225,0,6,0,0,0,0,0,250,0,118,0,0,0,141,0,4,0,251,0,114,0,29,0,187,0,44,0,45,0,157,0,6,0,61,0,0,0,187,0,18,0,18,0,23,0,74,0,95,0,73,0,0,0,253,0,138,0,39,0,235,0,38,0,250,0,22,0,137,0,40,0);
signal scenario_full  : scenario_type := (0,0,30,31,15,31,57,31,138,31,105,31,105,30,140,31,104,31,109,31,57,31,74,31,110,31,187,31,107,31,24,31,35,31,17,31,240,31,240,30,219,31,83,31,70,31,70,30,47,31,155,31,115,31,115,30,79,31,79,30,19,31,210,31,219,31,63,31,136,31,122,31,164,31,137,31,108,31,37,31,37,30,194,31,27,31,129,31,129,30,239,31,30,31,30,30,251,31,250,31,134,31,47,31,165,31,243,31,243,30,153,31,43,31,36,31,36,30,77,31,157,31,170,31,33,31,38,31,149,31,83,31,72,31,42,31,126,31,119,31,119,30,168,31,168,30,168,29,190,31,226,31,185,31,198,31,147,31,153,31,25,31,25,30,100,31,100,30,185,31,12,31,44,31,226,31,126,31,126,30,236,31,117,31,203,31,109,31,156,31,75,31,75,30,75,29,135,31,83,31,106,31,178,31,199,31,199,30,199,29,193,31,60,31,249,31,83,31,60,31,56,31,154,31,154,30,154,29,68,31,159,31,203,31,102,31,232,31,27,31,43,31,213,31,156,31,54,31,4,31,46,31,65,31,231,31,150,31,14,31,14,30,158,31,224,31,91,31,139,31,132,31,132,30,74,31,66,31,66,30,126,31,21,31,209,31,194,31,244,31,244,30,244,29,244,28,244,27,243,31,243,30,242,31,242,30,29,31,1,31,31,31,181,31,236,31,70,31,15,31,15,30,190,31,2,31,237,31,124,31,124,30,118,31,29,31,15,31,17,31,183,31,15,31,210,31,190,31,129,31,111,31,111,30,50,31,11,31,117,31,182,31,93,31,245,31,245,30,245,29,75,31,75,30,104,31,104,30,143,31,145,31,117,31,230,31,230,30,248,31,213,31,234,31,240,31,251,31,115,31,59,31,59,30,89,31,206,31,77,31,11,31,88,31,66,31,66,30,228,31,228,30,198,31,198,30,126,31,197,31,175,31,143,31,132,31,132,30,222,31,245,31,79,31,163,31,107,31,188,31,213,31,49,31,17,31,146,31,197,31,3,31,107,31,91,31,86,31,240,31,156,31,156,30,246,31,246,30,246,29,118,31,118,30,18,31,221,31,221,30,244,31,244,30,142,31,230,31,228,31,147,31,218,31,248,31,248,30,239,31,116,31,127,31,127,30,213,31,103,31,28,31,28,30,55,31,155,31,84,31,192,31,88,31,82,31,162,31,3,31,87,31,87,30,87,29,130,31,16,31,61,31,218,31,218,30,143,31,224,31,15,31,15,30,25,31,155,31,63,31,113,31,113,31,94,31,253,31,244,31,219,31,139,31,222,31,102,31,2,31,241,31,94,31,110,31,244,31,244,30,56,31,95,31,95,30,41,31,41,30,114,31,162,31,137,31,101,31,101,30,49,31,49,30,187,31,134,31,134,30,14,31,130,31,219,31,29,31,237,31,120,31,181,31,181,30,203,31,13,31,174,31,201,31,78,31,78,30,1,31,158,31,91,31,91,30,215,31,215,30,239,31,191,31,139,31,133,31,133,30,50,31,156,31,110,31,233,31,241,31,182,31,55,31,122,31,122,30,122,29,167,31,107,31,188,31,188,30,116,31,201,31,201,30,96,31,28,31,83,31,156,31,105,31,96,31,96,30,114,31,114,30,91,31,103,31,103,30,103,29,245,31,245,30,214,31,228,31,25,31,242,31,212,31,97,31,155,31,95,31,213,31,45,31,217,31,126,31,245,31,195,31,4,31,223,31,98,31,100,31,183,31,12,31,181,31,55,31,58,31,75,31,80,31,80,30,182,31,161,31,29,31,125,31,140,31,140,30,140,29,83,31,183,31,114,31,236,31,54,31,156,31,156,30,17,31,175,31,175,30,175,29,190,31,182,31,228,31,214,31,244,31,244,30,117,31,219,31,81,31,232,31,64,31,205,31,105,31,163,31,71,31,71,30,14,31,216,31,145,31,103,31,220,31,205,31,56,31,141,31,199,31,30,31,30,30,104,31,104,30,15,31,62,31,189,31,186,31,151,31,68,31,130,31,64,31,175,31,206,31,71,31,164,31,86,31,23,31,23,30,82,31,82,30,199,31,244,31,83,31,245,31,245,30,101,31,213,31,148,31,223,31,169,31,37,31,37,30,230,31,198,31,41,31,16,31,176,31,144,31,216,31,168,31,124,31,93,31,59,31,107,31,251,31,8,31,95,31,112,31,160,31,6,31,177,31,28,31,239,31,31,31,32,31,232,31,232,30,145,31,16,31,102,31,177,31,19,31,216,31,119,31,26,31,177,31,177,30,171,31,202,31,57,31,57,30,134,31,73,31,72,31,138,31,166,31,166,30,182,31,112,31,211,31,38,31,181,31,181,30,244,31,16,31,58,31,58,30,157,31,73,31,199,31,67,31,108,31,243,31,34,31,31,31,117,31,163,31,196,31,31,31,31,30,147,31,194,31,175,31,224,31,12,31,93,31,152,31,25,31,228,31,255,31,77,31,231,31,26,31,245,31,10,31,207,31,207,30,35,31,124,31,146,31,25,31,191,31,154,31,154,30,241,31,196,31,243,31,243,30,7,31,232,31,208,31,15,31,230,31,190,31,176,31,207,31,6,31,67,31,67,30,139,31,251,31,78,31,205,31,64,31,74,31,73,31,73,30,73,29,73,28,236,31,44,31,44,30,141,31,33,31,106,31,106,30,20,31,29,31,210,31,48,31,133,31,6,31,23,31,67,31,89,31,196,31,47,31,13,31,158,31,75,31,213,31,19,31,207,31,27,31,187,31,85,31,91,31,168,31,149,31,92,31,30,31,30,30,255,31,116,31,231,31,92,31,137,31,123,31,114,31,27,31,27,30,225,31,60,31,112,31,205,31,124,31,225,31,6,31,6,30,6,29,250,31,118,31,118,30,141,31,4,31,251,31,114,31,29,31,187,31,44,31,45,31,157,31,6,31,61,31,61,30,187,31,18,31,18,31,23,31,74,31,95,31,73,31,73,30,253,31,138,31,39,31,235,31,38,31,250,31,22,31,137,31,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
