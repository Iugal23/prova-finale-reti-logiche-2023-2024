-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_207 is
end project_tb_207;

architecture project_tb_arch_207 of project_tb_207 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 314;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,24,0,22,0,17,0,26,0,41,0,104,0,203,0,254,0,219,0,41,0,237,0,0,0,104,0,173,0,16,0,237,0,10,0,89,0,0,0,93,0,201,0,187,0,245,0,0,0,0,0,29,0,169,0,29,0,0,0,0,0,69,0,163,0,45,0,234,0,0,0,251,0,172,0,114,0,127,0,240,0,131,0,107,0,131,0,44,0,170,0,28,0,190,0,152,0,135,0,101,0,0,0,51,0,239,0,133,0,0,0,195,0,65,0,153,0,100,0,127,0,227,0,176,0,246,0,4,0,180,0,98,0,104,0,65,0,0,0,62,0,40,0,0,0,0,0,106,0,4,0,0,0,236,0,152,0,140,0,139,0,73,0,115,0,208,0,70,0,110,0,206,0,155,0,14,0,179,0,176,0,109,0,0,0,132,0,162,0,165,0,0,0,228,0,62,0,0,0,164,0,227,0,103,0,219,0,120,0,179,0,102,0,127,0,202,0,188,0,84,0,0,0,23,0,194,0,20,0,217,0,228,0,239,0,206,0,0,0,0,0,0,0,140,0,81,0,138,0,114,0,221,0,215,0,121,0,0,0,253,0,80,0,199,0,245,0,0,0,226,0,21,0,46,0,155,0,41,0,246,0,59,0,96,0,144,0,35,0,134,0,0,0,196,0,63,0,105,0,212,0,100,0,84,0,41,0,78,0,110,0,38,0,60,0,59,0,30,0,161,0,189,0,96,0,225,0,223,0,0,0,79,0,229,0,233,0,54,0,183,0,33,0,57,0,85,0,226,0,70,0,135,0,219,0,0,0,147,0,0,0,202,0,145,0,132,0,0,0,118,0,67,0,140,0,87,0,179,0,91,0,251,0,94,0,179,0,152,0,247,0,135,0,78,0,0,0,81,0,255,0,0,0,70,0,177,0,141,0,254,0,53,0,200,0,140,0,117,0,8,0,22,0,209,0,162,0,0,0,0,0,14,0,107,0,0,0,247,0,242,0,123,0,115,0,244,0,18,0,48,0,120,0,206,0,205,0,0,0,28,0,105,0,130,0,0,0,221,0,168,0,16,0,213,0,0,0,89,0,119,0,239,0,104,0,233,0,0,0,222,0,88,0,18,0,0,0,73,0,226,0,98,0,0,0,37,0,252,0,239,0,171,0,64,0,188,0,83,0,45,0,0,0,2,0,87,0,201,0,0,0,135,0,170,0,180,0,170,0,187,0,0,0,0,0,0,0,47,0,143,0,235,0,178,0,0,0,105,0,46,0,142,0,79,0,170,0,57,0,164,0,212,0,168,0,0,0,73,0,205,0,97,0,196,0,179,0,232,0,0,0,61,0,0,0,101,0,25,0,195,0,48,0,0,0,0,0,155,0,65,0,91,0,117,0,131,0,0,0,66,0,134,0,37,0,187,0);
signal scenario_full  : scenario_type := (68,31,24,31,22,31,17,31,26,31,41,31,104,31,203,31,254,31,219,31,41,31,237,31,237,30,104,31,173,31,16,31,237,31,10,31,89,31,89,30,93,31,201,31,187,31,245,31,245,30,245,29,29,31,169,31,29,31,29,30,29,29,69,31,163,31,45,31,234,31,234,30,251,31,172,31,114,31,127,31,240,31,131,31,107,31,131,31,44,31,170,31,28,31,190,31,152,31,135,31,101,31,101,30,51,31,239,31,133,31,133,30,195,31,65,31,153,31,100,31,127,31,227,31,176,31,246,31,4,31,180,31,98,31,104,31,65,31,65,30,62,31,40,31,40,30,40,29,106,31,4,31,4,30,236,31,152,31,140,31,139,31,73,31,115,31,208,31,70,31,110,31,206,31,155,31,14,31,179,31,176,31,109,31,109,30,132,31,162,31,165,31,165,30,228,31,62,31,62,30,164,31,227,31,103,31,219,31,120,31,179,31,102,31,127,31,202,31,188,31,84,31,84,30,23,31,194,31,20,31,217,31,228,31,239,31,206,31,206,30,206,29,206,28,140,31,81,31,138,31,114,31,221,31,215,31,121,31,121,30,253,31,80,31,199,31,245,31,245,30,226,31,21,31,46,31,155,31,41,31,246,31,59,31,96,31,144,31,35,31,134,31,134,30,196,31,63,31,105,31,212,31,100,31,84,31,41,31,78,31,110,31,38,31,60,31,59,31,30,31,161,31,189,31,96,31,225,31,223,31,223,30,79,31,229,31,233,31,54,31,183,31,33,31,57,31,85,31,226,31,70,31,135,31,219,31,219,30,147,31,147,30,202,31,145,31,132,31,132,30,118,31,67,31,140,31,87,31,179,31,91,31,251,31,94,31,179,31,152,31,247,31,135,31,78,31,78,30,81,31,255,31,255,30,70,31,177,31,141,31,254,31,53,31,200,31,140,31,117,31,8,31,22,31,209,31,162,31,162,30,162,29,14,31,107,31,107,30,247,31,242,31,123,31,115,31,244,31,18,31,48,31,120,31,206,31,205,31,205,30,28,31,105,31,130,31,130,30,221,31,168,31,16,31,213,31,213,30,89,31,119,31,239,31,104,31,233,31,233,30,222,31,88,31,18,31,18,30,73,31,226,31,98,31,98,30,37,31,252,31,239,31,171,31,64,31,188,31,83,31,45,31,45,30,2,31,87,31,201,31,201,30,135,31,170,31,180,31,170,31,187,31,187,30,187,29,187,28,47,31,143,31,235,31,178,31,178,30,105,31,46,31,142,31,79,31,170,31,57,31,164,31,212,31,168,31,168,30,73,31,205,31,97,31,196,31,179,31,232,31,232,30,61,31,61,30,101,31,25,31,195,31,48,31,48,30,48,29,155,31,65,31,91,31,117,31,131,31,131,30,66,31,134,31,37,31,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
