-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 247;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,112,0,40,0,81,0,139,0,0,0,76,0,74,0,53,0,19,0,0,0,244,0,247,0,100,0,79,0,6,0,163,0,0,0,83,0,191,0,0,0,144,0,222,0,201,0,0,0,245,0,180,0,152,0,66,0,0,0,46,0,81,0,64,0,27,0,168,0,0,0,251,0,146,0,19,0,0,0,94,0,228,0,100,0,240,0,0,0,81,0,68,0,230,0,55,0,54,0,115,0,178,0,25,0,171,0,8,0,171,0,233,0,0,0,0,0,159,0,65,0,0,0,244,0,93,0,0,0,73,0,182,0,170,0,173,0,0,0,118,0,235,0,208,0,126,0,194,0,0,0,74,0,254,0,177,0,11,0,160,0,34,0,188,0,20,0,93,0,237,0,164,0,46,0,0,0,117,0,252,0,0,0,221,0,80,0,234,0,21,0,54,0,102,0,0,0,0,0,84,0,203,0,88,0,23,0,104,0,219,0,251,0,118,0,205,0,53,0,0,0,196,0,225,0,194,0,221,0,35,0,195,0,32,0,0,0,64,0,227,0,165,0,0,0,143,0,143,0,29,0,55,0,207,0,0,0,126,0,5,0,110,0,210,0,149,0,167,0,186,0,54,0,45,0,226,0,115,0,73,0,0,0,10,0,132,0,134,0,0,0,5,0,119,0,172,0,0,0,134,0,0,0,167,0,245,0,5,0,0,0,30,0,4,0,55,0,0,0,0,0,215,0,5,0,0,0,146,0,168,0,201,0,241,0,8,0,138,0,0,0,0,0,73,0,143,0,152,0,44,0,69,0,107,0,189,0,11,0,189,0,225,0,0,0,17,0,168,0,107,0,90,0,18,0,9,0,163,0,238,0,6,0,239,0,212,0,24,0,27,0,0,0,229,0,0,0,224,0,234,0,86,0,244,0,0,0,81,0,0,0,152,0,0,0,222,0,73,0,168,0,58,0,48,0,224,0,141,0,0,0,0,0,0,0,21,0,42,0,82,0,0,0,188,0,168,0,51,0,116,0,122,0,33,0,0,0,130,0,0,0,204,0,0,0,0,0,128,0,159,0,0,0,227,0,15,0,0,0,74,0,0,0,226,0,0,0,97,0,214,0,0,0);
signal scenario_full  : scenario_type := (0,0,112,31,40,31,81,31,139,31,139,30,76,31,74,31,53,31,19,31,19,30,244,31,247,31,100,31,79,31,6,31,163,31,163,30,83,31,191,31,191,30,144,31,222,31,201,31,201,30,245,31,180,31,152,31,66,31,66,30,46,31,81,31,64,31,27,31,168,31,168,30,251,31,146,31,19,31,19,30,94,31,228,31,100,31,240,31,240,30,81,31,68,31,230,31,55,31,54,31,115,31,178,31,25,31,171,31,8,31,171,31,233,31,233,30,233,29,159,31,65,31,65,30,244,31,93,31,93,30,73,31,182,31,170,31,173,31,173,30,118,31,235,31,208,31,126,31,194,31,194,30,74,31,254,31,177,31,11,31,160,31,34,31,188,31,20,31,93,31,237,31,164,31,46,31,46,30,117,31,252,31,252,30,221,31,80,31,234,31,21,31,54,31,102,31,102,30,102,29,84,31,203,31,88,31,23,31,104,31,219,31,251,31,118,31,205,31,53,31,53,30,196,31,225,31,194,31,221,31,35,31,195,31,32,31,32,30,64,31,227,31,165,31,165,30,143,31,143,31,29,31,55,31,207,31,207,30,126,31,5,31,110,31,210,31,149,31,167,31,186,31,54,31,45,31,226,31,115,31,73,31,73,30,10,31,132,31,134,31,134,30,5,31,119,31,172,31,172,30,134,31,134,30,167,31,245,31,5,31,5,30,30,31,4,31,55,31,55,30,55,29,215,31,5,31,5,30,146,31,168,31,201,31,241,31,8,31,138,31,138,30,138,29,73,31,143,31,152,31,44,31,69,31,107,31,189,31,11,31,189,31,225,31,225,30,17,31,168,31,107,31,90,31,18,31,9,31,163,31,238,31,6,31,239,31,212,31,24,31,27,31,27,30,229,31,229,30,224,31,234,31,86,31,244,31,244,30,81,31,81,30,152,31,152,30,222,31,73,31,168,31,58,31,48,31,224,31,141,31,141,30,141,29,141,28,21,31,42,31,82,31,82,30,188,31,168,31,51,31,116,31,122,31,33,31,33,30,130,31,130,30,204,31,204,30,204,29,128,31,159,31,159,30,227,31,15,31,15,30,74,31,74,30,226,31,226,30,97,31,214,31,214,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
