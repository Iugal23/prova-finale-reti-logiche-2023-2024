-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 860;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,95,0,110,0,33,0,71,0,219,0,119,0,107,0,43,0,138,0,149,0,236,0,0,0,0,0,160,0,0,0,0,0,194,0,206,0,229,0,99,0,0,0,0,0,44,0,147,0,72,0,41,0,0,0,0,0,210,0,11,0,0,0,167,0,13,0,16,0,86,0,108,0,149,0,155,0,178,0,0,0,137,0,233,0,125,0,112,0,53,0,0,0,34,0,58,0,195,0,1,0,90,0,0,0,80,0,0,0,0,0,8,0,115,0,129,0,26,0,113,0,0,0,12,0,69,0,148,0,170,0,76,0,0,0,60,0,164,0,89,0,194,0,175,0,252,0,212,0,179,0,14,0,160,0,131,0,0,0,68,0,29,0,200,0,0,0,109,0,135,0,114,0,178,0,213,0,81,0,199,0,4,0,120,0,228,0,86,0,89,0,165,0,235,0,162,0,110,0,91,0,49,0,106,0,64,0,217,0,6,0,44,0,228,0,85,0,0,0,55,0,234,0,60,0,226,0,64,0,0,0,80,0,49,0,58,0,233,0,19,0,161,0,0,0,226,0,154,0,250,0,0,0,32,0,0,0,249,0,177,0,0,0,198,0,176,0,245,0,0,0,158,0,60,0,186,0,60,0,138,0,223,0,49,0,80,0,26,0,247,0,137,0,142,0,25,0,116,0,243,0,214,0,229,0,207,0,84,0,204,0,149,0,38,0,244,0,100,0,0,0,0,0,0,0,178,0,157,0,0,0,0,0,155,0,196,0,145,0,36,0,234,0,0,0,76,0,73,0,74,0,238,0,121,0,145,0,242,0,201,0,195,0,41,0,146,0,87,0,238,0,43,0,0,0,130,0,105,0,64,0,142,0,219,0,74,0,101,0,159,0,73,0,91,0,190,0,0,0,183,0,0,0,161,0,251,0,141,0,158,0,39,0,234,0,81,0,112,0,135,0,151,0,0,0,69,0,155,0,0,0,224,0,88,0,0,0,236,0,0,0,0,0,127,0,78,0,188,0,197,0,249,0,195,0,254,0,0,0,114,0,184,0,250,0,0,0,100,0,0,0,185,0,34,0,59,0,0,0,0,0,0,0,241,0,142,0,192,0,239,0,147,0,76,0,54,0,0,0,0,0,76,0,161,0,237,0,241,0,190,0,196,0,5,0,245,0,156,0,26,0,0,0,172,0,244,0,180,0,165,0,159,0,226,0,145,0,0,0,0,0,56,0,130,0,148,0,167,0,178,0,17,0,189,0,152,0,54,0,0,0,0,0,0,0,230,0,31,0,0,0,211,0,82,0,224,0,91,0,10,0,0,0,82,0,0,0,102,0,90,0,253,0,176,0,43,0,109,0,221,0,146,0,0,0,184,0,44,0,0,0,33,0,23,0,0,0,0,0,51,0,207,0,53,0,149,0,15,0,0,0,77,0,114,0,0,0,78,0,9,0,164,0,232,0,174,0,9,0,216,0,203,0,61,0,0,0,250,0,131,0,83,0,252,0,21,0,30,0,0,0,181,0,0,0,0,0,2,0,140,0,103,0,122,0,162,0,144,0,241,0,0,0,107,0,90,0,108,0,86,0,17,0,199,0,116,0,163,0,189,0,28,0,140,0,216,0,104,0,161,0,232,0,81,0,0,0,205,0,61,0,0,0,132,0,207,0,143,0,28,0,91,0,0,0,173,0,0,0,100,0,44,0,33,0,134,0,232,0,219,0,0,0,155,0,196,0,0,0,245,0,250,0,0,0,138,0,37,0,226,0,233,0,246,0,169,0,38,0,0,0,237,0,187,0,109,0,0,0,4,0,24,0,0,0,126,0,200,0,0,0,164,0,0,0,42,0,206,0,117,0,0,0,0,0,152,0,132,0,142,0,255,0,52,0,61,0,0,0,154,0,212,0,167,0,118,0,85,0,0,0,73,0,172,0,106,0,100,0,105,0,208,0,61,0,176,0,214,0,240,0,59,0,153,0,39,0,247,0,113,0,152,0,32,0,252,0,169,0,44,0,0,0,219,0,138,0,248,0,108,0,94,0,149,0,73,0,129,0,69,0,0,0,213,0,0,0,89,0,181,0,103,0,240,0,241,0,128,0,124,0,219,0,130,0,130,0,26,0,22,0,228,0,234,0,148,0,155,0,121,0,36,0,74,0,57,0,137,0,162,0,182,0,192,0,93,0,41,0,75,0,70,0,195,0,86,0,112,0,163,0,70,0,209,0,38,0,144,0,181,0,131,0,240,0,0,0,3,0,207,0,196,0,39,0,164,0,188,0,103,0,58,0,212,0,99,0,0,0,246,0,174,0,0,0,0,0,0,0,37,0,84,0,63,0,123,0,108,0,160,0,180,0,134,0,252,0,219,0,70,0,0,0,44,0,199,0,97,0,182,0,14,0,0,0,176,0,129,0,175,0,242,0,219,0,133,0,0,0,11,0,0,0,170,0,164,0,28,0,105,0,132,0,0,0,0,0,24,0,0,0,55,0,228,0,25,0,167,0,131,0,18,0,166,0,154,0,244,0,187,0,0,0,164,0,247,0,44,0,53,0,205,0,177,0,103,0,94,0,188,0,0,0,0,0,33,0,42,0,102,0,227,0,216,0,0,0,0,0,235,0,222,0,56,0,0,0,0,0,0,0,0,0,222,0,54,0,106,0,236,0,100,0,129,0,148,0,12,0,100,0,114,0,164,0,185,0,0,0,239,0,81,0,52,0,49,0,112,0,252,0,232,0,234,0,214,0,117,0,56,0,166,0,82,0,46,0,154,0,71,0,64,0,49,0,0,0,141,0,152,0,225,0,6,0,244,0,22,0,252,0,106,0,185,0,0,0,139,0,169,0,213,0,38,0,86,0,173,0,0,0,159,0,6,0,49,0,181,0,0,0,172,0,134,0,247,0,146,0,0,0,0,0,68,0,2,0,219,0,0,0,154,0,58,0,11,0,242,0,243,0,219,0,124,0,146,0,17,0,180,0,32,0,240,0,103,0,177,0,200,0,251,0,29,0,0,0,114,0,81,0,5,0,39,0,244,0,253,0,0,0,38,0,0,0,0,0,135,0,65,0,194,0,95,0,177,0,252,0,254,0,135,0,96,0,0,0,57,0,108,0,71,0,116,0,186,0,133,0,143,0,162,0,0,0,51,0,24,0,70,0,31,0,0,0,150,0,215,0,185,0,197,0,10,0,0,0,192,0,252,0,231,0,0,0,208,0,217,0,123,0,156,0,83,0,181,0,2,0,202,0,26,0,0,0,128,0,238,0,255,0,152,0,150,0,188,0,111,0,173,0,154,0,87,0,236,0,0,0,63,0,135,0,69,0,212,0,10,0,87,0,0,0,111,0,254,0,0,0,169,0,75,0,97,0,250,0,22,0,142,0,43,0,0,0,107,0,248,0,176,0,44,0,184,0,5,0,141,0,242,0,180,0,145,0,19,0,239,0,194,0,0,0,167,0,146,0,191,0,242,0,213,0,166,0,96,0,54,0,5,0,202,0,4,0,0,0,105,0,28,0,158,0,184,0,0,0,0,0,0,0,86,0,55,0,178,0,134,0,15,0,237,0,16,0,150,0,197,0,143,0,30,0,0,0,196,0,92,0,0,0,76,0,0,0,85,0,133,0,104,0,14,0,238,0,0,0,114,0,139,0,218,0,225,0,178,0,111,0,0,0,254,0,3,0,32,0,0,0,0,0,112,0,233,0,255,0,6,0,0,0,51,0,74,0,87,0,51,0,21,0,149,0,0,0,197,0,188,0,0,0,10,0,90,0,123,0,155,0,53,0,219,0,103,0,203,0,0,0,0,0,69,0,99,0,243,0,255,0,155,0,221,0,163,0,90,0,0,0,0,0,236,0,178,0,147,0,60,0);
signal scenario_full  : scenario_type := (71,31,95,31,110,31,33,31,71,31,219,31,119,31,107,31,43,31,138,31,149,31,236,31,236,30,236,29,160,31,160,30,160,29,194,31,206,31,229,31,99,31,99,30,99,29,44,31,147,31,72,31,41,31,41,30,41,29,210,31,11,31,11,30,167,31,13,31,16,31,86,31,108,31,149,31,155,31,178,31,178,30,137,31,233,31,125,31,112,31,53,31,53,30,34,31,58,31,195,31,1,31,90,31,90,30,80,31,80,30,80,29,8,31,115,31,129,31,26,31,113,31,113,30,12,31,69,31,148,31,170,31,76,31,76,30,60,31,164,31,89,31,194,31,175,31,252,31,212,31,179,31,14,31,160,31,131,31,131,30,68,31,29,31,200,31,200,30,109,31,135,31,114,31,178,31,213,31,81,31,199,31,4,31,120,31,228,31,86,31,89,31,165,31,235,31,162,31,110,31,91,31,49,31,106,31,64,31,217,31,6,31,44,31,228,31,85,31,85,30,55,31,234,31,60,31,226,31,64,31,64,30,80,31,49,31,58,31,233,31,19,31,161,31,161,30,226,31,154,31,250,31,250,30,32,31,32,30,249,31,177,31,177,30,198,31,176,31,245,31,245,30,158,31,60,31,186,31,60,31,138,31,223,31,49,31,80,31,26,31,247,31,137,31,142,31,25,31,116,31,243,31,214,31,229,31,207,31,84,31,204,31,149,31,38,31,244,31,100,31,100,30,100,29,100,28,178,31,157,31,157,30,157,29,155,31,196,31,145,31,36,31,234,31,234,30,76,31,73,31,74,31,238,31,121,31,145,31,242,31,201,31,195,31,41,31,146,31,87,31,238,31,43,31,43,30,130,31,105,31,64,31,142,31,219,31,74,31,101,31,159,31,73,31,91,31,190,31,190,30,183,31,183,30,161,31,251,31,141,31,158,31,39,31,234,31,81,31,112,31,135,31,151,31,151,30,69,31,155,31,155,30,224,31,88,31,88,30,236,31,236,30,236,29,127,31,78,31,188,31,197,31,249,31,195,31,254,31,254,30,114,31,184,31,250,31,250,30,100,31,100,30,185,31,34,31,59,31,59,30,59,29,59,28,241,31,142,31,192,31,239,31,147,31,76,31,54,31,54,30,54,29,76,31,161,31,237,31,241,31,190,31,196,31,5,31,245,31,156,31,26,31,26,30,172,31,244,31,180,31,165,31,159,31,226,31,145,31,145,30,145,29,56,31,130,31,148,31,167,31,178,31,17,31,189,31,152,31,54,31,54,30,54,29,54,28,230,31,31,31,31,30,211,31,82,31,224,31,91,31,10,31,10,30,82,31,82,30,102,31,90,31,253,31,176,31,43,31,109,31,221,31,146,31,146,30,184,31,44,31,44,30,33,31,23,31,23,30,23,29,51,31,207,31,53,31,149,31,15,31,15,30,77,31,114,31,114,30,78,31,9,31,164,31,232,31,174,31,9,31,216,31,203,31,61,31,61,30,250,31,131,31,83,31,252,31,21,31,30,31,30,30,181,31,181,30,181,29,2,31,140,31,103,31,122,31,162,31,144,31,241,31,241,30,107,31,90,31,108,31,86,31,17,31,199,31,116,31,163,31,189,31,28,31,140,31,216,31,104,31,161,31,232,31,81,31,81,30,205,31,61,31,61,30,132,31,207,31,143,31,28,31,91,31,91,30,173,31,173,30,100,31,44,31,33,31,134,31,232,31,219,31,219,30,155,31,196,31,196,30,245,31,250,31,250,30,138,31,37,31,226,31,233,31,246,31,169,31,38,31,38,30,237,31,187,31,109,31,109,30,4,31,24,31,24,30,126,31,200,31,200,30,164,31,164,30,42,31,206,31,117,31,117,30,117,29,152,31,132,31,142,31,255,31,52,31,61,31,61,30,154,31,212,31,167,31,118,31,85,31,85,30,73,31,172,31,106,31,100,31,105,31,208,31,61,31,176,31,214,31,240,31,59,31,153,31,39,31,247,31,113,31,152,31,32,31,252,31,169,31,44,31,44,30,219,31,138,31,248,31,108,31,94,31,149,31,73,31,129,31,69,31,69,30,213,31,213,30,89,31,181,31,103,31,240,31,241,31,128,31,124,31,219,31,130,31,130,31,26,31,22,31,228,31,234,31,148,31,155,31,121,31,36,31,74,31,57,31,137,31,162,31,182,31,192,31,93,31,41,31,75,31,70,31,195,31,86,31,112,31,163,31,70,31,209,31,38,31,144,31,181,31,131,31,240,31,240,30,3,31,207,31,196,31,39,31,164,31,188,31,103,31,58,31,212,31,99,31,99,30,246,31,174,31,174,30,174,29,174,28,37,31,84,31,63,31,123,31,108,31,160,31,180,31,134,31,252,31,219,31,70,31,70,30,44,31,199,31,97,31,182,31,14,31,14,30,176,31,129,31,175,31,242,31,219,31,133,31,133,30,11,31,11,30,170,31,164,31,28,31,105,31,132,31,132,30,132,29,24,31,24,30,55,31,228,31,25,31,167,31,131,31,18,31,166,31,154,31,244,31,187,31,187,30,164,31,247,31,44,31,53,31,205,31,177,31,103,31,94,31,188,31,188,30,188,29,33,31,42,31,102,31,227,31,216,31,216,30,216,29,235,31,222,31,56,31,56,30,56,29,56,28,56,27,222,31,54,31,106,31,236,31,100,31,129,31,148,31,12,31,100,31,114,31,164,31,185,31,185,30,239,31,81,31,52,31,49,31,112,31,252,31,232,31,234,31,214,31,117,31,56,31,166,31,82,31,46,31,154,31,71,31,64,31,49,31,49,30,141,31,152,31,225,31,6,31,244,31,22,31,252,31,106,31,185,31,185,30,139,31,169,31,213,31,38,31,86,31,173,31,173,30,159,31,6,31,49,31,181,31,181,30,172,31,134,31,247,31,146,31,146,30,146,29,68,31,2,31,219,31,219,30,154,31,58,31,11,31,242,31,243,31,219,31,124,31,146,31,17,31,180,31,32,31,240,31,103,31,177,31,200,31,251,31,29,31,29,30,114,31,81,31,5,31,39,31,244,31,253,31,253,30,38,31,38,30,38,29,135,31,65,31,194,31,95,31,177,31,252,31,254,31,135,31,96,31,96,30,57,31,108,31,71,31,116,31,186,31,133,31,143,31,162,31,162,30,51,31,24,31,70,31,31,31,31,30,150,31,215,31,185,31,197,31,10,31,10,30,192,31,252,31,231,31,231,30,208,31,217,31,123,31,156,31,83,31,181,31,2,31,202,31,26,31,26,30,128,31,238,31,255,31,152,31,150,31,188,31,111,31,173,31,154,31,87,31,236,31,236,30,63,31,135,31,69,31,212,31,10,31,87,31,87,30,111,31,254,31,254,30,169,31,75,31,97,31,250,31,22,31,142,31,43,31,43,30,107,31,248,31,176,31,44,31,184,31,5,31,141,31,242,31,180,31,145,31,19,31,239,31,194,31,194,30,167,31,146,31,191,31,242,31,213,31,166,31,96,31,54,31,5,31,202,31,4,31,4,30,105,31,28,31,158,31,184,31,184,30,184,29,184,28,86,31,55,31,178,31,134,31,15,31,237,31,16,31,150,31,197,31,143,31,30,31,30,30,196,31,92,31,92,30,76,31,76,30,85,31,133,31,104,31,14,31,238,31,238,30,114,31,139,31,218,31,225,31,178,31,111,31,111,30,254,31,3,31,32,31,32,30,32,29,112,31,233,31,255,31,6,31,6,30,51,31,74,31,87,31,51,31,21,31,149,31,149,30,197,31,188,31,188,30,10,31,90,31,123,31,155,31,53,31,219,31,103,31,203,31,203,30,203,29,69,31,99,31,243,31,255,31,155,31,221,31,163,31,90,31,90,30,90,29,236,31,178,31,147,31,60,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
