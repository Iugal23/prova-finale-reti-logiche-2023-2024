-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 180;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,205,0,2,0,51,0,169,0,56,0,106,0,255,0,48,0,23,0,247,0,77,0,236,0,166,0,27,0,92,0,48,0,0,0,185,0,240,0,238,0,200,0,36,0,214,0,192,0,0,0,207,0,251,0,250,0,137,0,83,0,7,0,54,0,21,0,146,0,0,0,144,0,135,0,50,0,190,0,150,0,0,0,24,0,234,0,221,0,119,0,208,0,137,0,227,0,135,0,221,0,168,0,97,0,48,0,143,0,4,0,0,0,249,0,0,0,32,0,0,0,62,0,39,0,0,0,157,0,193,0,201,0,5,0,201,0,6,0,223,0,12,0,0,0,165,0,97,0,176,0,8,0,154,0,41,0,77,0,191,0,185,0,34,0,136,0,236,0,56,0,0,0,133,0,131,0,42,0,229,0,190,0,0,0,2,0,3,0,221,0,69,0,139,0,30,0,56,0,0,0,41,0,59,0,145,0,234,0,75,0,38,0,163,0,0,0,233,0,230,0,4,0,0,0,155,0,88,0,159,0,0,0,119,0,0,0,0,0,2,0,142,0,193,0,7,0,77,0,221,0,0,0,3,0,181,0,141,0,0,0,0,0,154,0,159,0,115,0,26,0,110,0,0,0,102,0,118,0,0,0,30,0,0,0,194,0,0,0,28,0,0,0,184,0,0,0,175,0,0,0,50,0,96,0,179,0,74,0,93,0,241,0,0,0,0,0,217,0,0,0,105,0,135,0,0,0,107,0,10,0,157,0,74,0,0,0,158,0,155,0,221,0,0,0,237,0,116,0,20,0,136,0,86,0,0,0,193,0);
signal scenario_full  : scenario_type := (109,31,205,31,2,31,51,31,169,31,56,31,106,31,255,31,48,31,23,31,247,31,77,31,236,31,166,31,27,31,92,31,48,31,48,30,185,31,240,31,238,31,200,31,36,31,214,31,192,31,192,30,207,31,251,31,250,31,137,31,83,31,7,31,54,31,21,31,146,31,146,30,144,31,135,31,50,31,190,31,150,31,150,30,24,31,234,31,221,31,119,31,208,31,137,31,227,31,135,31,221,31,168,31,97,31,48,31,143,31,4,31,4,30,249,31,249,30,32,31,32,30,62,31,39,31,39,30,157,31,193,31,201,31,5,31,201,31,6,31,223,31,12,31,12,30,165,31,97,31,176,31,8,31,154,31,41,31,77,31,191,31,185,31,34,31,136,31,236,31,56,31,56,30,133,31,131,31,42,31,229,31,190,31,190,30,2,31,3,31,221,31,69,31,139,31,30,31,56,31,56,30,41,31,59,31,145,31,234,31,75,31,38,31,163,31,163,30,233,31,230,31,4,31,4,30,155,31,88,31,159,31,159,30,119,31,119,30,119,29,2,31,142,31,193,31,7,31,77,31,221,31,221,30,3,31,181,31,141,31,141,30,141,29,154,31,159,31,115,31,26,31,110,31,110,30,102,31,118,31,118,30,30,31,30,30,194,31,194,30,28,31,28,30,184,31,184,30,175,31,175,30,50,31,96,31,179,31,74,31,93,31,241,31,241,30,241,29,217,31,217,30,105,31,135,31,135,30,107,31,10,31,157,31,74,31,74,30,158,31,155,31,221,31,221,30,237,31,116,31,20,31,136,31,86,31,86,30,193,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
