-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 235;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (90,0,0,0,71,0,149,0,0,0,134,0,26,0,110,0,14,0,0,0,11,0,92,0,163,0,122,0,241,0,234,0,0,0,70,0,25,0,173,0,184,0,0,0,162,0,56,0,86,0,157,0,20,0,188,0,36,0,97,0,0,0,250,0,56,0,0,0,0,0,154,0,48,0,21,0,0,0,56,0,12,0,12,0,40,0,229,0,0,0,76,0,57,0,103,0,18,0,112,0,83,0,215,0,181,0,61,0,219,0,0,0,60,0,200,0,0,0,231,0,26,0,217,0,37,0,165,0,158,0,46,0,102,0,0,0,0,0,140,0,10,0,169,0,0,0,225,0,54,0,246,0,0,0,142,0,180,0,164,0,138,0,163,0,237,0,13,0,219,0,236,0,22,0,59,0,0,0,90,0,12,0,255,0,206,0,173,0,0,0,16,0,62,0,0,0,76,0,0,0,203,0,0,0,217,0,0,0,116,0,56,0,255,0,59,0,234,0,237,0,108,0,153,0,0,0,0,0,216,0,121,0,0,0,0,0,7,0,73,0,109,0,64,0,33,0,83,0,59,0,124,0,0,0,99,0,233,0,65,0,0,0,0,0,21,0,0,0,137,0,113,0,154,0,0,0,4,0,152,0,189,0,244,0,114,0,60,0,92,0,142,0,131,0,53,0,157,0,56,0,226,0,236,0,63,0,133,0,145,0,230,0,200,0,170,0,148,0,203,0,148,0,10,0,240,0,208,0,147,0,103,0,162,0,244,0,204,0,9,0,70,0,212,0,109,0,103,0,0,0,58,0,200,0,254,0,4,0,158,0,48,0,132,0,95,0,60,0,5,0,162,0,121,0,211,0,251,0,214,0,10,0,3,0,211,0,5,0,113,0,56,0,0,0,80,0,0,0,0,0,0,0,70,0,222,0,218,0,187,0,34,0,2,0,32,0,222,0,15,0,0,0,223,0,63,0,6,0,56,0,144,0,241,0,90,0,246,0,43,0,150,0,0,0,51,0,191,0,202,0,90,0,117,0,147,0,134,0,0,0,51,0,37,0,0,0,70,0,40,0);
signal scenario_full  : scenario_type := (90,31,90,30,71,31,149,31,149,30,134,31,26,31,110,31,14,31,14,30,11,31,92,31,163,31,122,31,241,31,234,31,234,30,70,31,25,31,173,31,184,31,184,30,162,31,56,31,86,31,157,31,20,31,188,31,36,31,97,31,97,30,250,31,56,31,56,30,56,29,154,31,48,31,21,31,21,30,56,31,12,31,12,31,40,31,229,31,229,30,76,31,57,31,103,31,18,31,112,31,83,31,215,31,181,31,61,31,219,31,219,30,60,31,200,31,200,30,231,31,26,31,217,31,37,31,165,31,158,31,46,31,102,31,102,30,102,29,140,31,10,31,169,31,169,30,225,31,54,31,246,31,246,30,142,31,180,31,164,31,138,31,163,31,237,31,13,31,219,31,236,31,22,31,59,31,59,30,90,31,12,31,255,31,206,31,173,31,173,30,16,31,62,31,62,30,76,31,76,30,203,31,203,30,217,31,217,30,116,31,56,31,255,31,59,31,234,31,237,31,108,31,153,31,153,30,153,29,216,31,121,31,121,30,121,29,7,31,73,31,109,31,64,31,33,31,83,31,59,31,124,31,124,30,99,31,233,31,65,31,65,30,65,29,21,31,21,30,137,31,113,31,154,31,154,30,4,31,152,31,189,31,244,31,114,31,60,31,92,31,142,31,131,31,53,31,157,31,56,31,226,31,236,31,63,31,133,31,145,31,230,31,200,31,170,31,148,31,203,31,148,31,10,31,240,31,208,31,147,31,103,31,162,31,244,31,204,31,9,31,70,31,212,31,109,31,103,31,103,30,58,31,200,31,254,31,4,31,158,31,48,31,132,31,95,31,60,31,5,31,162,31,121,31,211,31,251,31,214,31,10,31,3,31,211,31,5,31,113,31,56,31,56,30,80,31,80,30,80,29,80,28,70,31,222,31,218,31,187,31,34,31,2,31,32,31,222,31,15,31,15,30,223,31,63,31,6,31,56,31,144,31,241,31,90,31,246,31,43,31,150,31,150,30,51,31,191,31,202,31,90,31,117,31,147,31,134,31,134,30,51,31,37,31,37,30,70,31,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
