-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 389;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (237,0,108,0,119,0,95,0,0,0,0,0,119,0,209,0,0,0,10,0,173,0,192,0,2,0,143,0,51,0,169,0,202,0,0,0,28,0,0,0,187,0,114,0,0,0,235,0,29,0,176,0,215,0,162,0,33,0,8,0,162,0,163,0,239,0,185,0,85,0,200,0,11,0,172,0,192,0,253,0,87,0,225,0,0,0,207,0,12,0,0,0,165,0,224,0,0,0,13,0,6,0,0,0,215,0,135,0,94,0,118,0,14,0,131,0,0,0,193,0,255,0,166,0,77,0,72,0,7,0,20,0,19,0,0,0,255,0,120,0,0,0,105,0,0,0,0,0,164,0,232,0,72,0,57,0,0,0,141,0,0,0,0,0,50,0,176,0,31,0,176,0,202,0,201,0,21,0,181,0,38,0,0,0,8,0,208,0,161,0,0,0,250,0,134,0,0,0,12,0,58,0,121,0,0,0,0,0,82,0,0,0,0,0,242,0,144,0,188,0,142,0,84,0,159,0,150,0,0,0,104,0,166,0,193,0,0,0,0,0,0,0,115,0,128,0,101,0,188,0,14,0,234,0,143,0,176,0,0,0,23,0,120,0,163,0,154,0,0,0,49,0,39,0,194,0,183,0,0,0,0,0,0,0,237,0,0,0,0,0,68,0,0,0,181,0,145,0,6,0,160,0,0,0,47,0,228,0,39,0,0,0,215,0,0,0,252,0,31,0,0,0,113,0,202,0,0,0,234,0,165,0,0,0,201,0,230,0,0,0,0,0,149,0,0,0,154,0,183,0,30,0,116,0,177,0,248,0,223,0,0,0,195,0,96,0,1,0,0,0,61,0,246,0,45,0,96,0,58,0,71,0,63,0,0,0,0,0,58,0,43,0,0,0,0,0,179,0,105,0,109,0,130,0,0,0,253,0,106,0,0,0,112,0,61,0,46,0,56,0,0,0,190,0,205,0,207,0,0,0,159,0,116,0,0,0,78,0,86,0,0,0,39,0,69,0,111,0,0,0,147,0,62,0,238,0,42,0,0,0,0,0,0,0,207,0,0,0,104,0,71,0,0,0,84,0,141,0,83,0,228,0,116,0,136,0,0,0,174,0,141,0,184,0,0,0,174,0,0,0,3,0,0,0,0,0,88,0,34,0,0,0,0,0,0,0,35,0,241,0,227,0,174,0,140,0,199,0,21,0,166,0,13,0,29,0,0,0,81,0,48,0,85,0,0,0,96,0,5,0,105,0,0,0,23,0,143,0,80,0,153,0,239,0,89,0,141,0,12,0,72,0,22,0,61,0,79,0,105,0,201,0,140,0,0,0,0,0,0,0,43,0,109,0,35,0,83,0,99,0,121,0,205,0,36,0,105,0,5,0,7,0,98,0,241,0,218,0,0,0,187,0,230,0,0,0,176,0,197,0,138,0,141,0,62,0,0,0,220,0,36,0,236,0,61,0,41,0,206,0,1,0,42,0,72,0,81,0,62,0,141,0,128,0,170,0,0,0,54,0,40,0,248,0,92,0,15,0,60,0,173,0,249,0,26,0,187,0,246,0,0,0,7,0,113,0,142,0,60,0,87,0,94,0,129,0,73,0,32,0,186,0,255,0,178,0,77,0,170,0,232,0,139,0,122,0,0,0,85,0,67,0,242,0,157,0,41,0,0,0,16,0,109,0,18,0,0,0,157,0,79,0,170,0,65,0,0,0,203,0,81,0,202,0,43,0,28,0,147,0,196,0,80,0,244,0,129,0);
signal scenario_full  : scenario_type := (237,31,108,31,119,31,95,31,95,30,95,29,119,31,209,31,209,30,10,31,173,31,192,31,2,31,143,31,51,31,169,31,202,31,202,30,28,31,28,30,187,31,114,31,114,30,235,31,29,31,176,31,215,31,162,31,33,31,8,31,162,31,163,31,239,31,185,31,85,31,200,31,11,31,172,31,192,31,253,31,87,31,225,31,225,30,207,31,12,31,12,30,165,31,224,31,224,30,13,31,6,31,6,30,215,31,135,31,94,31,118,31,14,31,131,31,131,30,193,31,255,31,166,31,77,31,72,31,7,31,20,31,19,31,19,30,255,31,120,31,120,30,105,31,105,30,105,29,164,31,232,31,72,31,57,31,57,30,141,31,141,30,141,29,50,31,176,31,31,31,176,31,202,31,201,31,21,31,181,31,38,31,38,30,8,31,208,31,161,31,161,30,250,31,134,31,134,30,12,31,58,31,121,31,121,30,121,29,82,31,82,30,82,29,242,31,144,31,188,31,142,31,84,31,159,31,150,31,150,30,104,31,166,31,193,31,193,30,193,29,193,28,115,31,128,31,101,31,188,31,14,31,234,31,143,31,176,31,176,30,23,31,120,31,163,31,154,31,154,30,49,31,39,31,194,31,183,31,183,30,183,29,183,28,237,31,237,30,237,29,68,31,68,30,181,31,145,31,6,31,160,31,160,30,47,31,228,31,39,31,39,30,215,31,215,30,252,31,31,31,31,30,113,31,202,31,202,30,234,31,165,31,165,30,201,31,230,31,230,30,230,29,149,31,149,30,154,31,183,31,30,31,116,31,177,31,248,31,223,31,223,30,195,31,96,31,1,31,1,30,61,31,246,31,45,31,96,31,58,31,71,31,63,31,63,30,63,29,58,31,43,31,43,30,43,29,179,31,105,31,109,31,130,31,130,30,253,31,106,31,106,30,112,31,61,31,46,31,56,31,56,30,190,31,205,31,207,31,207,30,159,31,116,31,116,30,78,31,86,31,86,30,39,31,69,31,111,31,111,30,147,31,62,31,238,31,42,31,42,30,42,29,42,28,207,31,207,30,104,31,71,31,71,30,84,31,141,31,83,31,228,31,116,31,136,31,136,30,174,31,141,31,184,31,184,30,174,31,174,30,3,31,3,30,3,29,88,31,34,31,34,30,34,29,34,28,35,31,241,31,227,31,174,31,140,31,199,31,21,31,166,31,13,31,29,31,29,30,81,31,48,31,85,31,85,30,96,31,5,31,105,31,105,30,23,31,143,31,80,31,153,31,239,31,89,31,141,31,12,31,72,31,22,31,61,31,79,31,105,31,201,31,140,31,140,30,140,29,140,28,43,31,109,31,35,31,83,31,99,31,121,31,205,31,36,31,105,31,5,31,7,31,98,31,241,31,218,31,218,30,187,31,230,31,230,30,176,31,197,31,138,31,141,31,62,31,62,30,220,31,36,31,236,31,61,31,41,31,206,31,1,31,42,31,72,31,81,31,62,31,141,31,128,31,170,31,170,30,54,31,40,31,248,31,92,31,15,31,60,31,173,31,249,31,26,31,187,31,246,31,246,30,7,31,113,31,142,31,60,31,87,31,94,31,129,31,73,31,32,31,186,31,255,31,178,31,77,31,170,31,232,31,139,31,122,31,122,30,85,31,67,31,242,31,157,31,41,31,41,30,16,31,109,31,18,31,18,30,157,31,79,31,170,31,65,31,65,30,203,31,81,31,202,31,43,31,28,31,147,31,196,31,80,31,244,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
