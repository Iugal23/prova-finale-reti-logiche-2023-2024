-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_773 is
end project_tb_773;

architecture project_tb_arch_773 of project_tb_773 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 973;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (132,0,78,0,122,0,173,0,0,0,177,0,0,0,0,0,0,0,0,0,0,0,52,0,0,0,0,0,0,0,0,0,83,0,195,0,138,0,223,0,91,0,160,0,159,0,253,0,145,0,78,0,0,0,0,0,238,0,37,0,80,0,0,0,200,0,254,0,93,0,53,0,0,0,242,0,0,0,35,0,143,0,0,0,17,0,27,0,230,0,131,0,33,0,67,0,161,0,19,0,212,0,28,0,12,0,205,0,146,0,191,0,153,0,139,0,0,0,0,0,223,0,138,0,52,0,56,0,67,0,4,0,0,0,0,0,192,0,32,0,34,0,42,0,0,0,86,0,237,0,234,0,147,0,188,0,39,0,30,0,1,0,69,0,252,0,210,0,121,0,0,0,52,0,0,0,129,0,58,0,21,0,226,0,159,0,209,0,56,0,160,0,235,0,50,0,199,0,125,0,140,0,48,0,0,0,39,0,0,0,246,0,254,0,0,0,0,0,111,0,0,0,2,0,225,0,167,0,0,0,158,0,158,0,166,0,152,0,6,0,169,0,175,0,69,0,141,0,206,0,159,0,0,0,173,0,81,0,0,0,0,0,179,0,210,0,23,0,0,0,52,0,0,0,0,0,0,0,99,0,94,0,231,0,215,0,155,0,131,0,203,0,0,0,0,0,8,0,161,0,164,0,0,0,111,0,176,0,171,0,0,0,190,0,225,0,39,0,0,0,0,0,22,0,190,0,219,0,0,0,95,0,0,0,0,0,0,0,112,0,113,0,0,0,114,0,120,0,44,0,255,0,137,0,1,0,0,0,78,0,76,0,175,0,0,0,208,0,182,0,177,0,166,0,0,0,221,0,81,0,5,0,190,0,163,0,23,0,126,0,41,0,251,0,53,0,0,0,67,0,156,0,53,0,18,0,0,0,37,0,247,0,93,0,219,0,177,0,44,0,0,0,2,0,49,0,51,0,31,0,62,0,245,0,164,0,54,0,185,0,54,0,11,0,0,0,0,0,167,0,77,0,66,0,112,0,214,0,7,0,214,0,41,0,0,0,249,0,183,0,93,0,118,0,135,0,184,0,131,0,15,0,207,0,0,0,94,0,36,0,136,0,95,0,0,0,174,0,186,0,160,0,75,0,16,0,0,0,46,0,176,0,0,0,23,0,156,0,189,0,105,0,203,0,173,0,201,0,65,0,148,0,220,0,107,0,183,0,75,0,16,0,0,0,96,0,7,0,107,0,0,0,239,0,175,0,0,0,113,0,154,0,0,0,245,0,48,0,251,0,95,0,0,0,242,0,53,0,124,0,0,0,0,0,9,0,0,0,0,0,0,0,254,0,232,0,204,0,168,0,109,0,0,0,226,0,70,0,244,0,177,0,0,0,152,0,208,0,178,0,127,0,213,0,47,0,58,0,173,0,0,0,191,0,0,0,65,0,137,0,0,0,144,0,30,0,0,0,102,0,173,0,200,0,167,0,0,0,147,0,92,0,1,0,35,0,78,0,43,0,85,0,226,0,89,0,0,0,0,0,62,0,79,0,1,0,223,0,126,0,96,0,4,0,145,0,9,0,0,0,134,0,171,0,9,0,130,0,163,0,68,0,0,0,0,0,38,0,0,0,96,0,229,0,158,0,50,0,105,0,172,0,175,0,213,0,145,0,246,0,152,0,251,0,112,0,0,0,213,0,193,0,0,0,224,0,52,0,192,0,199,0,200,0,33,0,0,0,225,0,107,0,27,0,243,0,63,0,240,0,0,0,0,0,0,0,0,0,93,0,114,0,247,0,0,0,89,0,188,0,100,0,36,0,248,0,67,0,0,0,74,0,0,0,89,0,200,0,25,0,239,0,161,0,169,0,0,0,0,0,162,0,23,0,95,0,128,0,0,0,12,0,69,0,0,0,220,0,31,0,135,0,0,0,249,0,151,0,227,0,79,0,184,0,94,0,55,0,11,0,168,0,82,0,145,0,0,0,141,0,56,0,99,0,123,0,73,0,175,0,171,0,178,0,67,0,107,0,132,0,196,0,185,0,29,0,121,0,115,0,11,0,0,0,254,0,140,0,0,0,43,0,216,0,0,0,226,0,18,0,0,0,252,0,143,0,47,0,4,0,19,0,199,0,0,0,171,0,22,0,41,0,9,0,146,0,0,0,234,0,96,0,0,0,0,0,14,0,237,0,194,0,121,0,70,0,161,0,211,0,2,0,78,0,7,0,168,0,0,0,0,0,0,0,0,0,187,0,183,0,118,0,234,0,19,0,0,0,0,0,211,0,100,0,4,0,72,0,193,0,240,0,201,0,138,0,22,0,97,0,198,0,142,0,222,0,0,0,134,0,103,0,98,0,239,0,213,0,207,0,91,0,0,0,61,0,233,0,0,0,67,0,113,0,158,0,0,0,0,0,193,0,23,0,238,0,229,0,0,0,15,0,182,0,0,0,51,0,3,0,233,0,0,0,58,0,0,0,111,0,0,0,0,0,130,0,112,0,178,0,40,0,85,0,149,0,152,0,174,0,119,0,0,0,207,0,107,0,97,0,235,0,57,0,156,0,66,0,10,0,56,0,11,0,197,0,54,0,145,0,110,0,87,0,50,0,46,0,0,0,124,0,0,0,116,0,92,0,175,0,68,0,17,0,0,0,5,0,211,0,0,0,168,0,14,0,121,0,32,0,5,0,214,0,2,0,120,0,162,0,0,0,183,0,181,0,0,0,236,0,200,0,0,0,139,0,182,0,235,0,51,0,0,0,51,0,109,0,220,0,50,0,237,0,49,0,11,0,135,0,157,0,0,0,142,0,64,0,157,0,210,0,94,0,109,0,201,0,122,0,15,0,0,0,69,0,49,0,82,0,186,0,212,0,183,0,224,0,5,0,28,0,91,0,31,0,0,0,71,0,105,0,74,0,175,0,62,0,210,0,0,0,249,0,192,0,171,0,0,0,85,0,0,0,229,0,0,0,228,0,2,0,90,0,238,0,113,0,0,0,30,0,75,0,253,0,250,0,126,0,206,0,0,0,84,0,219,0,201,0,125,0,229,0,243,0,28,0,181,0,0,0,124,0,158,0,49,0,90,0,0,0,3,0,35,0,142,0,236,0,190,0,30,0,59,0,48,0,25,0,180,0,185,0,248,0,83,0,0,0,0,0,133,0,104,0,217,0,77,0,163,0,139,0,9,0,3,0,113,0,26,0,124,0,142,0,0,0,0,0,0,0,191,0,201,0,27,0,142,0,145,0,99,0,78,0,33,0,40,0,19,0,241,0,0,0,0,0,155,0,0,0,179,0,45,0,100,0,6,0,20,0,0,0,157,0,0,0,20,0,139,0,169,0,133,0,73,0,94,0,195,0,36,0,0,0,208,0,175,0,18,0,93,0,81,0,48,0,231,0,102,0,231,0,43,0,170,0,61,0,0,0,55,0,0,0,62,0,252,0,197,0,125,0,11,0,142,0,185,0,245,0,158,0,216,0,46,0,0,0,18,0,200,0,71,0,223,0,188,0,42,0,60,0,156,0,104,0,224,0,0,0,46,0,100,0,218,0,170,0,171,0,55,0,229,0,90,0,102,0,203,0,111,0,0,0,50,0,217,0,18,0,210,0,155,0,90,0,0,0,15,0,177,0,254,0,107,0,0,0,40,0,211,0,0,0,104,0,0,0,96,0,114,0,118,0,15,0,0,0,123,0,230,0,0,0,0,0,106,0,0,0,0,0,0,0,137,0,51,0,244,0,97,0,0,0,124,0,16,0,42,0,111,0,0,0,146,0,215,0,196,0,0,0,163,0,46,0,143,0,129,0,155,0,8,0,0,0,142,0,116,0,98,0,114,0,112,0,84,0,177,0,95,0,144,0,118,0,0,0,244,0,154,0,25,0,45,0,210,0,215,0,42,0,0,0,32,0,3,0,0,0,125,0,61,0,32,0,90,0,0,0,164,0,0,0,216,0,196,0,68,0,0,0,158,0,0,0,90,0,32,0,43,0,99,0,132,0,160,0,2,0,86,0,38,0,108,0,178,0,0,0,177,0,179,0,87,0,0,0,89,0,253,0,35,0,208,0,0,0,4,0,141,0,93,0,46,0,229,0,236,0,243,0,198,0,176,0,31,0,98,0,0,0,148,0,111,0,186,0,159,0,242,0,0,0,0,0,178,0,29,0,240,0,94,0,108,0,37,0,211,0,0,0,0,0,59,0,255,0,220,0,187,0,0,0,52,0,60,0,0,0,86,0,0,0,73,0,131,0,11,0,0,0,0,0,40,0,177,0,9,0,96,0,0,0,84,0,0,0,220,0,244,0,208,0,185,0,0,0,27,0,0,0,65,0,61,0,168,0,219,0,181,0,194,0,240,0,44,0,28,0,99,0,90,0);
signal scenario_full  : scenario_type := (132,31,78,31,122,31,173,31,173,30,177,31,177,30,177,29,177,28,177,27,177,26,52,31,52,30,52,29,52,28,52,27,83,31,195,31,138,31,223,31,91,31,160,31,159,31,253,31,145,31,78,31,78,30,78,29,238,31,37,31,80,31,80,30,200,31,254,31,93,31,53,31,53,30,242,31,242,30,35,31,143,31,143,30,17,31,27,31,230,31,131,31,33,31,67,31,161,31,19,31,212,31,28,31,12,31,205,31,146,31,191,31,153,31,139,31,139,30,139,29,223,31,138,31,52,31,56,31,67,31,4,31,4,30,4,29,192,31,32,31,34,31,42,31,42,30,86,31,237,31,234,31,147,31,188,31,39,31,30,31,1,31,69,31,252,31,210,31,121,31,121,30,52,31,52,30,129,31,58,31,21,31,226,31,159,31,209,31,56,31,160,31,235,31,50,31,199,31,125,31,140,31,48,31,48,30,39,31,39,30,246,31,254,31,254,30,254,29,111,31,111,30,2,31,225,31,167,31,167,30,158,31,158,31,166,31,152,31,6,31,169,31,175,31,69,31,141,31,206,31,159,31,159,30,173,31,81,31,81,30,81,29,179,31,210,31,23,31,23,30,52,31,52,30,52,29,52,28,99,31,94,31,231,31,215,31,155,31,131,31,203,31,203,30,203,29,8,31,161,31,164,31,164,30,111,31,176,31,171,31,171,30,190,31,225,31,39,31,39,30,39,29,22,31,190,31,219,31,219,30,95,31,95,30,95,29,95,28,112,31,113,31,113,30,114,31,120,31,44,31,255,31,137,31,1,31,1,30,78,31,76,31,175,31,175,30,208,31,182,31,177,31,166,31,166,30,221,31,81,31,5,31,190,31,163,31,23,31,126,31,41,31,251,31,53,31,53,30,67,31,156,31,53,31,18,31,18,30,37,31,247,31,93,31,219,31,177,31,44,31,44,30,2,31,49,31,51,31,31,31,62,31,245,31,164,31,54,31,185,31,54,31,11,31,11,30,11,29,167,31,77,31,66,31,112,31,214,31,7,31,214,31,41,31,41,30,249,31,183,31,93,31,118,31,135,31,184,31,131,31,15,31,207,31,207,30,94,31,36,31,136,31,95,31,95,30,174,31,186,31,160,31,75,31,16,31,16,30,46,31,176,31,176,30,23,31,156,31,189,31,105,31,203,31,173,31,201,31,65,31,148,31,220,31,107,31,183,31,75,31,16,31,16,30,96,31,7,31,107,31,107,30,239,31,175,31,175,30,113,31,154,31,154,30,245,31,48,31,251,31,95,31,95,30,242,31,53,31,124,31,124,30,124,29,9,31,9,30,9,29,9,28,254,31,232,31,204,31,168,31,109,31,109,30,226,31,70,31,244,31,177,31,177,30,152,31,208,31,178,31,127,31,213,31,47,31,58,31,173,31,173,30,191,31,191,30,65,31,137,31,137,30,144,31,30,31,30,30,102,31,173,31,200,31,167,31,167,30,147,31,92,31,1,31,35,31,78,31,43,31,85,31,226,31,89,31,89,30,89,29,62,31,79,31,1,31,223,31,126,31,96,31,4,31,145,31,9,31,9,30,134,31,171,31,9,31,130,31,163,31,68,31,68,30,68,29,38,31,38,30,96,31,229,31,158,31,50,31,105,31,172,31,175,31,213,31,145,31,246,31,152,31,251,31,112,31,112,30,213,31,193,31,193,30,224,31,52,31,192,31,199,31,200,31,33,31,33,30,225,31,107,31,27,31,243,31,63,31,240,31,240,30,240,29,240,28,240,27,93,31,114,31,247,31,247,30,89,31,188,31,100,31,36,31,248,31,67,31,67,30,74,31,74,30,89,31,200,31,25,31,239,31,161,31,169,31,169,30,169,29,162,31,23,31,95,31,128,31,128,30,12,31,69,31,69,30,220,31,31,31,135,31,135,30,249,31,151,31,227,31,79,31,184,31,94,31,55,31,11,31,168,31,82,31,145,31,145,30,141,31,56,31,99,31,123,31,73,31,175,31,171,31,178,31,67,31,107,31,132,31,196,31,185,31,29,31,121,31,115,31,11,31,11,30,254,31,140,31,140,30,43,31,216,31,216,30,226,31,18,31,18,30,252,31,143,31,47,31,4,31,19,31,199,31,199,30,171,31,22,31,41,31,9,31,146,31,146,30,234,31,96,31,96,30,96,29,14,31,237,31,194,31,121,31,70,31,161,31,211,31,2,31,78,31,7,31,168,31,168,30,168,29,168,28,168,27,187,31,183,31,118,31,234,31,19,31,19,30,19,29,211,31,100,31,4,31,72,31,193,31,240,31,201,31,138,31,22,31,97,31,198,31,142,31,222,31,222,30,134,31,103,31,98,31,239,31,213,31,207,31,91,31,91,30,61,31,233,31,233,30,67,31,113,31,158,31,158,30,158,29,193,31,23,31,238,31,229,31,229,30,15,31,182,31,182,30,51,31,3,31,233,31,233,30,58,31,58,30,111,31,111,30,111,29,130,31,112,31,178,31,40,31,85,31,149,31,152,31,174,31,119,31,119,30,207,31,107,31,97,31,235,31,57,31,156,31,66,31,10,31,56,31,11,31,197,31,54,31,145,31,110,31,87,31,50,31,46,31,46,30,124,31,124,30,116,31,92,31,175,31,68,31,17,31,17,30,5,31,211,31,211,30,168,31,14,31,121,31,32,31,5,31,214,31,2,31,120,31,162,31,162,30,183,31,181,31,181,30,236,31,200,31,200,30,139,31,182,31,235,31,51,31,51,30,51,31,109,31,220,31,50,31,237,31,49,31,11,31,135,31,157,31,157,30,142,31,64,31,157,31,210,31,94,31,109,31,201,31,122,31,15,31,15,30,69,31,49,31,82,31,186,31,212,31,183,31,224,31,5,31,28,31,91,31,31,31,31,30,71,31,105,31,74,31,175,31,62,31,210,31,210,30,249,31,192,31,171,31,171,30,85,31,85,30,229,31,229,30,228,31,2,31,90,31,238,31,113,31,113,30,30,31,75,31,253,31,250,31,126,31,206,31,206,30,84,31,219,31,201,31,125,31,229,31,243,31,28,31,181,31,181,30,124,31,158,31,49,31,90,31,90,30,3,31,35,31,142,31,236,31,190,31,30,31,59,31,48,31,25,31,180,31,185,31,248,31,83,31,83,30,83,29,133,31,104,31,217,31,77,31,163,31,139,31,9,31,3,31,113,31,26,31,124,31,142,31,142,30,142,29,142,28,191,31,201,31,27,31,142,31,145,31,99,31,78,31,33,31,40,31,19,31,241,31,241,30,241,29,155,31,155,30,179,31,45,31,100,31,6,31,20,31,20,30,157,31,157,30,20,31,139,31,169,31,133,31,73,31,94,31,195,31,36,31,36,30,208,31,175,31,18,31,93,31,81,31,48,31,231,31,102,31,231,31,43,31,170,31,61,31,61,30,55,31,55,30,62,31,252,31,197,31,125,31,11,31,142,31,185,31,245,31,158,31,216,31,46,31,46,30,18,31,200,31,71,31,223,31,188,31,42,31,60,31,156,31,104,31,224,31,224,30,46,31,100,31,218,31,170,31,171,31,55,31,229,31,90,31,102,31,203,31,111,31,111,30,50,31,217,31,18,31,210,31,155,31,90,31,90,30,15,31,177,31,254,31,107,31,107,30,40,31,211,31,211,30,104,31,104,30,96,31,114,31,118,31,15,31,15,30,123,31,230,31,230,30,230,29,106,31,106,30,106,29,106,28,137,31,51,31,244,31,97,31,97,30,124,31,16,31,42,31,111,31,111,30,146,31,215,31,196,31,196,30,163,31,46,31,143,31,129,31,155,31,8,31,8,30,142,31,116,31,98,31,114,31,112,31,84,31,177,31,95,31,144,31,118,31,118,30,244,31,154,31,25,31,45,31,210,31,215,31,42,31,42,30,32,31,3,31,3,30,125,31,61,31,32,31,90,31,90,30,164,31,164,30,216,31,196,31,68,31,68,30,158,31,158,30,90,31,32,31,43,31,99,31,132,31,160,31,2,31,86,31,38,31,108,31,178,31,178,30,177,31,179,31,87,31,87,30,89,31,253,31,35,31,208,31,208,30,4,31,141,31,93,31,46,31,229,31,236,31,243,31,198,31,176,31,31,31,98,31,98,30,148,31,111,31,186,31,159,31,242,31,242,30,242,29,178,31,29,31,240,31,94,31,108,31,37,31,211,31,211,30,211,29,59,31,255,31,220,31,187,31,187,30,52,31,60,31,60,30,86,31,86,30,73,31,131,31,11,31,11,30,11,29,40,31,177,31,9,31,96,31,96,30,84,31,84,30,220,31,244,31,208,31,185,31,185,30,27,31,27,30,65,31,61,31,168,31,219,31,181,31,194,31,240,31,44,31,28,31,99,31,90,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
