-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 931;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,37,0,17,0,212,0,255,0,99,0,0,0,173,0,159,0,98,0,61,0,0,0,216,0,0,0,141,0,37,0,162,0,226,0,206,0,156,0,235,0,224,0,237,0,136,0,190,0,191,0,152,0,103,0,62,0,14,0,161,0,209,0,213,0,63,0,182,0,236,0,0,0,66,0,102,0,254,0,174,0,245,0,155,0,249,0,0,0,83,0,13,0,79,0,88,0,46,0,249,0,0,0,215,0,191,0,13,0,0,0,254,0,0,0,228,0,236,0,235,0,234,0,230,0,49,0,217,0,197,0,158,0,52,0,53,0,210,0,205,0,248,0,77,0,183,0,0,0,12,0,18,0,126,0,0,0,181,0,0,0,12,0,0,0,119,0,76,0,191,0,204,0,0,0,78,0,244,0,115,0,0,0,108,0,77,0,72,0,5,0,151,0,163,0,232,0,87,0,62,0,82,0,181,0,178,0,97,0,232,0,3,0,65,0,0,0,16,0,0,0,208,0,0,0,198,0,0,0,0,0,0,0,187,0,254,0,0,0,145,0,0,0,39,0,166,0,194,0,93,0,78,0,184,0,145,0,94,0,0,0,0,0,0,0,187,0,49,0,116,0,196,0,40,0,73,0,206,0,126,0,201,0,15,0,0,0,44,0,0,0,117,0,179,0,224,0,241,0,71,0,198,0,63,0,31,0,53,0,71,0,0,0,11,0,255,0,198,0,0,0,64,0,245,0,234,0,216,0,169,0,89,0,0,0,47,0,159,0,240,0,52,0,227,0,0,0,78,0,131,0,60,0,230,0,60,0,154,0,0,0,0,0,173,0,214,0,230,0,227,0,156,0,42,0,176,0,112,0,207,0,140,0,49,0,77,0,205,0,59,0,0,0,165,0,223,0,185,0,0,0,0,0,0,0,14,0,147,0,0,0,92,0,220,0,123,0,0,0,41,0,0,0,176,0,245,0,168,0,76,0,0,0,14,0,210,0,167,0,0,0,182,0,4,0,42,0,255,0,28,0,180,0,159,0,103,0,218,0,0,0,189,0,0,0,104,0,0,0,157,0,216,0,0,0,136,0,101,0,210,0,52,0,0,0,60,0,160,0,151,0,165,0,210,0,0,0,210,0,66,0,0,0,47,0,26,0,199,0,160,0,5,0,186,0,0,0,236,0,0,0,178,0,97,0,0,0,10,0,95,0,155,0,37,0,235,0,94,0,0,0,151,0,233,0,185,0,0,0,10,0,158,0,170,0,180,0,0,0,5,0,215,0,2,0,77,0,0,0,198,0,0,0,177,0,59,0,149,0,73,0,74,0,30,0,225,0,222,0,220,0,235,0,19,0,62,0,146,0,250,0,56,0,0,0,37,0,125,0,0,0,63,0,32,0,0,0,30,0,0,0,0,0,0,0,11,0,0,0,27,0,43,0,76,0,68,0,236,0,63,0,15,0,21,0,0,0,254,0,219,0,0,0,201,0,65,0,0,0,108,0,1,0,48,0,0,0,137,0,252,0,86,0,57,0,249,0,57,0,141,0,115,0,196,0,180,0,121,0,249,0,67,0,235,0,22,0,90,0,73,0,240,0,86,0,0,0,222,0,3,0,0,0,202,0,161,0,0,0,4,0,33,0,122,0,219,0,0,0,0,0,232,0,6,0,240,0,141,0,14,0,90,0,0,0,8,0,0,0,120,0,157,0,144,0,0,0,0,0,83,0,0,0,0,0,178,0,70,0,179,0,8,0,0,0,238,0,125,0,104,0,53,0,189,0,82,0,9,0,111,0,0,0,21,0,91,0,110,0,0,0,89,0,0,0,232,0,122,0,233,0,130,0,243,0,38,0,67,0,48,0,168,0,210,0,141,0,113,0,102,0,102,0,0,0,187,0,124,0,130,0,1,0,0,0,105,0,234,0,108,0,89,0,0,0,227,0,72,0,197,0,0,0,0,0,0,0,128,0,124,0,196,0,164,0,232,0,136,0,64,0,0,0,102,0,30,0,110,0,130,0,205,0,142,0,139,0,81,0,0,0,0,0,93,0,178,0,124,0,53,0,230,0,0,0,243,0,10,0,130,0,195,0,177,0,64,0,86,0,70,0,243,0,85,0,0,0,250,0,194,0,184,0,0,0,121,0,50,0,200,0,82,0,102,0,120,0,217,0,216,0,184,0,221,0,184,0,4,0,144,0,202,0,230,0,161,0,83,0,28,0,37,0,116,0,0,0,224,0,0,0,62,0,63,0,72,0,127,0,236,0,109,0,0,0,32,0,50,0,152,0,0,0,133,0,228,0,133,0,204,0,26,0,125,0,0,0,0,0,100,0,62,0,0,0,138,0,126,0,25,0,191,0,23,0,234,0,67,0,216,0,202,0,0,0,213,0,131,0,219,0,0,0,157,0,8,0,229,0,249,0,69,0,34,0,0,0,249,0,26,0,0,0,24,0,0,0,25,0,169,0,74,0,228,0,0,0,133,0,0,0,32,0,0,0,229,0,138,0,49,0,110,0,0,0,43,0,156,0,13,0,249,0,29,0,243,0,231,0,233,0,0,0,139,0,254,0,0,0,221,0,142,0,0,0,0,0,236,0,202,0,137,0,0,0,103,0,18,0,161,0,254,0,204,0,201,0,179,0,210,0,0,0,63,0,58,0,197,0,0,0,149,0,0,0,0,0,177,0,25,0,18,0,193,0,141,0,0,0,79,0,251,0,111,0,223,0,8,0,0,0,120,0,202,0,208,0,208,0,83,0,63,0,199,0,13,0,5,0,143,0,244,0,243,0,0,0,17,0,58,0,93,0,41,0,204,0,154,0,21,0,20,0,254,0,11,0,38,0,144,0,31,0,155,0,0,0,0,0,30,0,139,0,0,0,0,0,2,0,105,0,7,0,70,0,153,0,175,0,0,0,209,0,227,0,129,0,0,0,27,0,78,0,0,0,71,0,25,0,0,0,108,0,65,0,38,0,0,0,206,0,107,0,40,0,54,0,0,0,231,0,168,0,0,0,254,0,98,0,151,0,170,0,122,0,144,0,238,0,208,0,95,0,69,0,72,0,0,0,88,0,54,0,0,0,0,0,0,0,27,0,215,0,22,0,160,0,78,0,242,0,1,0,197,0,0,0,39,0,101,0,97,0,0,0,29,0,215,0,72,0,167,0,218,0,15,0,12,0,187,0,0,0,143,0,79,0,0,0,113,0,0,0,0,0,87,0,104,0,115,0,110,0,8,0,0,0,149,0,0,0,147,0,177,0,191,0,79,0,0,0,0,0,205,0,93,0,246,0,46,0,134,0,149,0,105,0,80,0,208,0,10,0,0,0,168,0,148,0,0,0,10,0,63,0,200,0,83,0,76,0,185,0,157,0,149,0,0,0,212,0,249,0,106,0,0,0,149,0,245,0,47,0,0,0,117,0,0,0,230,0,248,0,0,0,70,0,212,0,140,0,112,0,67,0,56,0,150,0,97,0,0,0,34,0,235,0,132,0,76,0,0,0,130,0,253,0,123,0,24,0,195,0,51,0,50,0,0,0,0,0,189,0,140,0,121,0,30,0,210,0,241,0,54,0,220,0,2,0,0,0,0,0,74,0,119,0,113,0,90,0,34,0,0,0,179,0,2,0,25,0,78,0,210,0,100,0,0,0,229,0,55,0,0,0,255,0,185,0,0,0,35,0,204,0,126,0,116,0,0,0,112,0,0,0,44,0,0,0,148,0,48,0,26,0,0,0,39,0,33,0,119,0,109,0,218,0,79,0,106,0,64,0,65,0,138,0,0,0,60,0,133,0,25,0,116,0,104,0,0,0,237,0,144,0,0,0,54,0,10,0,71,0,0,0,0,0,73,0,58,0,0,0,184,0,253,0,88,0,0,0,93,0,3,0,97,0,0,0,7,0,0,0,15,0,73,0,0,0,116,0,126,0,0,0,90,0,21,0,32,0,120,0,0,0,48,0,180,0,117,0,107,0,98,0,18,0,139,0,73,0,141,0,37,0,0,0,0,0,134,0,247,0,16,0,249,0,245,0,181,0,56,0,177,0,246,0,0,0,114,0,201,0,74,0,178,0,164,0,115,0,0,0,0,0,0,0,0,0,212,0,13,0,17,0,0,0,182,0,0,0,15,0,116,0,11,0,72,0,95,0,132,0,232,0,0,0,209,0,0,0,147,0,23,0,0,0,223,0,26,0);
signal scenario_full  : scenario_type := (49,31,37,31,17,31,212,31,255,31,99,31,99,30,173,31,159,31,98,31,61,31,61,30,216,31,216,30,141,31,37,31,162,31,226,31,206,31,156,31,235,31,224,31,237,31,136,31,190,31,191,31,152,31,103,31,62,31,14,31,161,31,209,31,213,31,63,31,182,31,236,31,236,30,66,31,102,31,254,31,174,31,245,31,155,31,249,31,249,30,83,31,13,31,79,31,88,31,46,31,249,31,249,30,215,31,191,31,13,31,13,30,254,31,254,30,228,31,236,31,235,31,234,31,230,31,49,31,217,31,197,31,158,31,52,31,53,31,210,31,205,31,248,31,77,31,183,31,183,30,12,31,18,31,126,31,126,30,181,31,181,30,12,31,12,30,119,31,76,31,191,31,204,31,204,30,78,31,244,31,115,31,115,30,108,31,77,31,72,31,5,31,151,31,163,31,232,31,87,31,62,31,82,31,181,31,178,31,97,31,232,31,3,31,65,31,65,30,16,31,16,30,208,31,208,30,198,31,198,30,198,29,198,28,187,31,254,31,254,30,145,31,145,30,39,31,166,31,194,31,93,31,78,31,184,31,145,31,94,31,94,30,94,29,94,28,187,31,49,31,116,31,196,31,40,31,73,31,206,31,126,31,201,31,15,31,15,30,44,31,44,30,117,31,179,31,224,31,241,31,71,31,198,31,63,31,31,31,53,31,71,31,71,30,11,31,255,31,198,31,198,30,64,31,245,31,234,31,216,31,169,31,89,31,89,30,47,31,159,31,240,31,52,31,227,31,227,30,78,31,131,31,60,31,230,31,60,31,154,31,154,30,154,29,173,31,214,31,230,31,227,31,156,31,42,31,176,31,112,31,207,31,140,31,49,31,77,31,205,31,59,31,59,30,165,31,223,31,185,31,185,30,185,29,185,28,14,31,147,31,147,30,92,31,220,31,123,31,123,30,41,31,41,30,176,31,245,31,168,31,76,31,76,30,14,31,210,31,167,31,167,30,182,31,4,31,42,31,255,31,28,31,180,31,159,31,103,31,218,31,218,30,189,31,189,30,104,31,104,30,157,31,216,31,216,30,136,31,101,31,210,31,52,31,52,30,60,31,160,31,151,31,165,31,210,31,210,30,210,31,66,31,66,30,47,31,26,31,199,31,160,31,5,31,186,31,186,30,236,31,236,30,178,31,97,31,97,30,10,31,95,31,155,31,37,31,235,31,94,31,94,30,151,31,233,31,185,31,185,30,10,31,158,31,170,31,180,31,180,30,5,31,215,31,2,31,77,31,77,30,198,31,198,30,177,31,59,31,149,31,73,31,74,31,30,31,225,31,222,31,220,31,235,31,19,31,62,31,146,31,250,31,56,31,56,30,37,31,125,31,125,30,63,31,32,31,32,30,30,31,30,30,30,29,30,28,11,31,11,30,27,31,43,31,76,31,68,31,236,31,63,31,15,31,21,31,21,30,254,31,219,31,219,30,201,31,65,31,65,30,108,31,1,31,48,31,48,30,137,31,252,31,86,31,57,31,249,31,57,31,141,31,115,31,196,31,180,31,121,31,249,31,67,31,235,31,22,31,90,31,73,31,240,31,86,31,86,30,222,31,3,31,3,30,202,31,161,31,161,30,4,31,33,31,122,31,219,31,219,30,219,29,232,31,6,31,240,31,141,31,14,31,90,31,90,30,8,31,8,30,120,31,157,31,144,31,144,30,144,29,83,31,83,30,83,29,178,31,70,31,179,31,8,31,8,30,238,31,125,31,104,31,53,31,189,31,82,31,9,31,111,31,111,30,21,31,91,31,110,31,110,30,89,31,89,30,232,31,122,31,233,31,130,31,243,31,38,31,67,31,48,31,168,31,210,31,141,31,113,31,102,31,102,31,102,30,187,31,124,31,130,31,1,31,1,30,105,31,234,31,108,31,89,31,89,30,227,31,72,31,197,31,197,30,197,29,197,28,128,31,124,31,196,31,164,31,232,31,136,31,64,31,64,30,102,31,30,31,110,31,130,31,205,31,142,31,139,31,81,31,81,30,81,29,93,31,178,31,124,31,53,31,230,31,230,30,243,31,10,31,130,31,195,31,177,31,64,31,86,31,70,31,243,31,85,31,85,30,250,31,194,31,184,31,184,30,121,31,50,31,200,31,82,31,102,31,120,31,217,31,216,31,184,31,221,31,184,31,4,31,144,31,202,31,230,31,161,31,83,31,28,31,37,31,116,31,116,30,224,31,224,30,62,31,63,31,72,31,127,31,236,31,109,31,109,30,32,31,50,31,152,31,152,30,133,31,228,31,133,31,204,31,26,31,125,31,125,30,125,29,100,31,62,31,62,30,138,31,126,31,25,31,191,31,23,31,234,31,67,31,216,31,202,31,202,30,213,31,131,31,219,31,219,30,157,31,8,31,229,31,249,31,69,31,34,31,34,30,249,31,26,31,26,30,24,31,24,30,25,31,169,31,74,31,228,31,228,30,133,31,133,30,32,31,32,30,229,31,138,31,49,31,110,31,110,30,43,31,156,31,13,31,249,31,29,31,243,31,231,31,233,31,233,30,139,31,254,31,254,30,221,31,142,31,142,30,142,29,236,31,202,31,137,31,137,30,103,31,18,31,161,31,254,31,204,31,201,31,179,31,210,31,210,30,63,31,58,31,197,31,197,30,149,31,149,30,149,29,177,31,25,31,18,31,193,31,141,31,141,30,79,31,251,31,111,31,223,31,8,31,8,30,120,31,202,31,208,31,208,31,83,31,63,31,199,31,13,31,5,31,143,31,244,31,243,31,243,30,17,31,58,31,93,31,41,31,204,31,154,31,21,31,20,31,254,31,11,31,38,31,144,31,31,31,155,31,155,30,155,29,30,31,139,31,139,30,139,29,2,31,105,31,7,31,70,31,153,31,175,31,175,30,209,31,227,31,129,31,129,30,27,31,78,31,78,30,71,31,25,31,25,30,108,31,65,31,38,31,38,30,206,31,107,31,40,31,54,31,54,30,231,31,168,31,168,30,254,31,98,31,151,31,170,31,122,31,144,31,238,31,208,31,95,31,69,31,72,31,72,30,88,31,54,31,54,30,54,29,54,28,27,31,215,31,22,31,160,31,78,31,242,31,1,31,197,31,197,30,39,31,101,31,97,31,97,30,29,31,215,31,72,31,167,31,218,31,15,31,12,31,187,31,187,30,143,31,79,31,79,30,113,31,113,30,113,29,87,31,104,31,115,31,110,31,8,31,8,30,149,31,149,30,147,31,177,31,191,31,79,31,79,30,79,29,205,31,93,31,246,31,46,31,134,31,149,31,105,31,80,31,208,31,10,31,10,30,168,31,148,31,148,30,10,31,63,31,200,31,83,31,76,31,185,31,157,31,149,31,149,30,212,31,249,31,106,31,106,30,149,31,245,31,47,31,47,30,117,31,117,30,230,31,248,31,248,30,70,31,212,31,140,31,112,31,67,31,56,31,150,31,97,31,97,30,34,31,235,31,132,31,76,31,76,30,130,31,253,31,123,31,24,31,195,31,51,31,50,31,50,30,50,29,189,31,140,31,121,31,30,31,210,31,241,31,54,31,220,31,2,31,2,30,2,29,74,31,119,31,113,31,90,31,34,31,34,30,179,31,2,31,25,31,78,31,210,31,100,31,100,30,229,31,55,31,55,30,255,31,185,31,185,30,35,31,204,31,126,31,116,31,116,30,112,31,112,30,44,31,44,30,148,31,48,31,26,31,26,30,39,31,33,31,119,31,109,31,218,31,79,31,106,31,64,31,65,31,138,31,138,30,60,31,133,31,25,31,116,31,104,31,104,30,237,31,144,31,144,30,54,31,10,31,71,31,71,30,71,29,73,31,58,31,58,30,184,31,253,31,88,31,88,30,93,31,3,31,97,31,97,30,7,31,7,30,15,31,73,31,73,30,116,31,126,31,126,30,90,31,21,31,32,31,120,31,120,30,48,31,180,31,117,31,107,31,98,31,18,31,139,31,73,31,141,31,37,31,37,30,37,29,134,31,247,31,16,31,249,31,245,31,181,31,56,31,177,31,246,31,246,30,114,31,201,31,74,31,178,31,164,31,115,31,115,30,115,29,115,28,115,27,212,31,13,31,17,31,17,30,182,31,182,30,15,31,116,31,11,31,72,31,95,31,132,31,232,31,232,30,209,31,209,30,147,31,23,31,23,30,223,31,26,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
