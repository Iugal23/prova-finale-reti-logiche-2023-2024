-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 673;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,88,0,128,0,136,0,254,0,0,0,0,0,0,0,0,0,147,0,161,0,57,0,0,0,237,0,32,0,199,0,190,0,38,0,192,0,0,0,221,0,157,0,250,0,68,0,0,0,0,0,239,0,202,0,169,0,153,0,219,0,242,0,24,0,9,0,206,0,245,0,0,0,249,0,185,0,72,0,212,0,95,0,124,0,145,0,184,0,200,0,126,0,59,0,36,0,12,0,248,0,20,0,85,0,176,0,0,0,0,0,92,0,7,0,204,0,65,0,227,0,97,0,238,0,202,0,168,0,117,0,192,0,0,0,12,0,209,0,208,0,80,0,213,0,239,0,92,0,0,0,186,0,141,0,0,0,218,0,207,0,43,0,0,0,128,0,205,0,0,0,50,0,141,0,206,0,18,0,0,0,58,0,146,0,75,0,140,0,159,0,232,0,173,0,0,0,199,0,134,0,57,0,95,0,61,0,0,0,144,0,77,0,70,0,86,0,209,0,0,0,0,0,209,0,87,0,226,0,193,0,217,0,7,0,0,0,26,0,0,0,84,0,0,0,171,0,89,0,16,0,244,0,115,0,70,0,249,0,222,0,64,0,0,0,182,0,129,0,207,0,9,0,217,0,199,0,246,0,62,0,188,0,0,0,217,0,133,0,9,0,98,0,213,0,55,0,121,0,100,0,46,0,125,0,2,0,115,0,0,0,250,0,111,0,79,0,0,0,95,0,166,0,0,0,0,0,0,0,0,0,186,0,0,0,165,0,0,0,72,0,105,0,176,0,79,0,0,0,185,0,12,0,8,0,206,0,74,0,241,0,202,0,168,0,149,0,98,0,0,0,0,0,160,0,0,0,0,0,194,0,159,0,219,0,106,0,234,0,0,0,199,0,48,0,249,0,119,0,145,0,75,0,156,0,70,0,164,0,147,0,47,0,1,0,64,0,255,0,156,0,150,0,0,0,184,0,223,0,4,0,0,0,43,0,195,0,73,0,0,0,81,0,154,0,255,0,0,0,242,0,119,0,89,0,135,0,78,0,0,0,156,0,221,0,5,0,129,0,218,0,119,0,32,0,94,0,230,0,0,0,0,0,239,0,190,0,140,0,0,0,0,0,0,0,246,0,0,0,48,0,0,0,0,0,225,0,88,0,0,0,0,0,75,0,0,0,94,0,35,0,131,0,38,0,57,0,142,0,220,0,0,0,221,0,82,0,40,0,4,0,174,0,89,0,227,0,9,0,180,0,0,0,74,0,9,0,2,0,0,0,24,0,0,0,0,0,101,0,0,0,25,0,231,0,195,0,34,0,224,0,69,0,171,0,0,0,147,0,21,0,6,0,242,0,183,0,208,0,126,0,0,0,162,0,98,0,0,0,118,0,0,0,0,0,45,0,127,0,143,0,117,0,50,0,70,0,208,0,60,0,8,0,217,0,173,0,82,0,208,0,0,0,129,0,248,0,154,0,112,0,203,0,224,0,0,0,135,0,183,0,82,0,72,0,147,0,22,0,184,0,4,0,119,0,79,0,35,0,253,0,192,0,0,0,0,0,229,0,4,0,57,0,143,0,0,0,52,0,0,0,171,0,117,0,174,0,100,0,0,0,213,0,178,0,200,0,0,0,233,0,94,0,247,0,99,0,71,0,61,0,0,0,0,0,156,0,197,0,233,0,52,0,188,0,0,0,51,0,214,0,0,0,184,0,238,0,203,0,124,0,0,0,242,0,78,0,65,0,82,0,0,0,246,0,8,0,0,0,0,0,82,0,97,0,0,0,0,0,37,0,9,0,0,0,79,0,230,0,47,0,187,0,0,0,226,0,4,0,0,0,196,0,0,0,73,0,5,0,45,0,38,0,170,0,207,0,0,0,0,0,187,0,0,0,84,0,200,0,0,0,2,0,0,0,0,0,87,0,0,0,18,0,245,0,35,0,0,0,232,0,161,0,176,0,181,0,44,0,15,0,29,0,157,0,195,0,73,0,0,0,26,0,215,0,100,0,121,0,129,0,134,0,64,0,0,0,162,0,202,0,95,0,52,0,30,0,0,0,29,0,54,0,220,0,69,0,232,0,147,0,77,0,7,0,233,0,176,0,38,0,195,0,0,0,116,0,18,0,204,0,4,0,0,0,150,0,26,0,247,0,94,0,215,0,0,0,0,0,168,0,13,0,61,0,0,0,186,0,37,0,62,0,57,0,203,0,15,0,80,0,0,0,97,0,0,0,0,0,75,0,0,0,78,0,0,0,0,0,0,0,0,0,8,0,98,0,58,0,8,0,171,0,118,0,238,0,0,0,47,0,90,0,210,0,114,0,0,0,227,0,190,0,56,0,101,0,94,0,79,0,0,0,185,0,217,0,198,0,239,0,69,0,188,0,169,0,0,0,54,0,83,0,0,0,0,0,184,0,0,0,133,0,158,0,163,0,187,0,207,0,64,0,240,0,79,0,223,0,44,0,22,0,187,0,216,0,85,0,75,0,128,0,49,0,0,0,247,0,0,0,18,0,82,0,89,0,252,0,0,0,77,0,67,0,38,0,205,0,151,0,0,0,29,0,146,0,169,0,14,0,45,0,232,0,118,0,62,0,209,0,174,0,99,0,3,0,242,0,191,0,169,0,23,0,74,0,101,0,26,0,128,0,161,0,236,0,142,0,0,0,0,0,0,0,49,0,24,0,15,0,63,0,66,0,1,0,183,0,73,0,91,0,253,0,19,0,174,0,41,0,0,0,25,0,86,0,247,0,151,0,0,0,41,0,173,0,90,0,60,0,81,0,58,0,51,0,210,0,244,0,249,0,183,0,0,0,144,0,0,0,68,0,0,0,0,0,143,0,179,0,253,0,251,0,255,0,138,0,102,0,0,0,106,0,120,0,0,0,59,0,66,0,196,0,0,0,23,0,145,0,0,0,201,0,19,0,0,0,0,0,47,0,247,0,164,0,35,0,16,0,0,0,113,0,77,0,54,0,0,0,60,0,86,0,124,0,222,0,0,0,0,0,235,0,112,0,143,0,126,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,88,31,128,31,136,31,254,31,254,30,254,29,254,28,254,27,147,31,161,31,57,31,57,30,237,31,32,31,199,31,190,31,38,31,192,31,192,30,221,31,157,31,250,31,68,31,68,30,68,29,239,31,202,31,169,31,153,31,219,31,242,31,24,31,9,31,206,31,245,31,245,30,249,31,185,31,72,31,212,31,95,31,124,31,145,31,184,31,200,31,126,31,59,31,36,31,12,31,248,31,20,31,85,31,176,31,176,30,176,29,92,31,7,31,204,31,65,31,227,31,97,31,238,31,202,31,168,31,117,31,192,31,192,30,12,31,209,31,208,31,80,31,213,31,239,31,92,31,92,30,186,31,141,31,141,30,218,31,207,31,43,31,43,30,128,31,205,31,205,30,50,31,141,31,206,31,18,31,18,30,58,31,146,31,75,31,140,31,159,31,232,31,173,31,173,30,199,31,134,31,57,31,95,31,61,31,61,30,144,31,77,31,70,31,86,31,209,31,209,30,209,29,209,31,87,31,226,31,193,31,217,31,7,31,7,30,26,31,26,30,84,31,84,30,171,31,89,31,16,31,244,31,115,31,70,31,249,31,222,31,64,31,64,30,182,31,129,31,207,31,9,31,217,31,199,31,246,31,62,31,188,31,188,30,217,31,133,31,9,31,98,31,213,31,55,31,121,31,100,31,46,31,125,31,2,31,115,31,115,30,250,31,111,31,79,31,79,30,95,31,166,31,166,30,166,29,166,28,166,27,186,31,186,30,165,31,165,30,72,31,105,31,176,31,79,31,79,30,185,31,12,31,8,31,206,31,74,31,241,31,202,31,168,31,149,31,98,31,98,30,98,29,160,31,160,30,160,29,194,31,159,31,219,31,106,31,234,31,234,30,199,31,48,31,249,31,119,31,145,31,75,31,156,31,70,31,164,31,147,31,47,31,1,31,64,31,255,31,156,31,150,31,150,30,184,31,223,31,4,31,4,30,43,31,195,31,73,31,73,30,81,31,154,31,255,31,255,30,242,31,119,31,89,31,135,31,78,31,78,30,156,31,221,31,5,31,129,31,218,31,119,31,32,31,94,31,230,31,230,30,230,29,239,31,190,31,140,31,140,30,140,29,140,28,246,31,246,30,48,31,48,30,48,29,225,31,88,31,88,30,88,29,75,31,75,30,94,31,35,31,131,31,38,31,57,31,142,31,220,31,220,30,221,31,82,31,40,31,4,31,174,31,89,31,227,31,9,31,180,31,180,30,74,31,9,31,2,31,2,30,24,31,24,30,24,29,101,31,101,30,25,31,231,31,195,31,34,31,224,31,69,31,171,31,171,30,147,31,21,31,6,31,242,31,183,31,208,31,126,31,126,30,162,31,98,31,98,30,118,31,118,30,118,29,45,31,127,31,143,31,117,31,50,31,70,31,208,31,60,31,8,31,217,31,173,31,82,31,208,31,208,30,129,31,248,31,154,31,112,31,203,31,224,31,224,30,135,31,183,31,82,31,72,31,147,31,22,31,184,31,4,31,119,31,79,31,35,31,253,31,192,31,192,30,192,29,229,31,4,31,57,31,143,31,143,30,52,31,52,30,171,31,117,31,174,31,100,31,100,30,213,31,178,31,200,31,200,30,233,31,94,31,247,31,99,31,71,31,61,31,61,30,61,29,156,31,197,31,233,31,52,31,188,31,188,30,51,31,214,31,214,30,184,31,238,31,203,31,124,31,124,30,242,31,78,31,65,31,82,31,82,30,246,31,8,31,8,30,8,29,82,31,97,31,97,30,97,29,37,31,9,31,9,30,79,31,230,31,47,31,187,31,187,30,226,31,4,31,4,30,196,31,196,30,73,31,5,31,45,31,38,31,170,31,207,31,207,30,207,29,187,31,187,30,84,31,200,31,200,30,2,31,2,30,2,29,87,31,87,30,18,31,245,31,35,31,35,30,232,31,161,31,176,31,181,31,44,31,15,31,29,31,157,31,195,31,73,31,73,30,26,31,215,31,100,31,121,31,129,31,134,31,64,31,64,30,162,31,202,31,95,31,52,31,30,31,30,30,29,31,54,31,220,31,69,31,232,31,147,31,77,31,7,31,233,31,176,31,38,31,195,31,195,30,116,31,18,31,204,31,4,31,4,30,150,31,26,31,247,31,94,31,215,31,215,30,215,29,168,31,13,31,61,31,61,30,186,31,37,31,62,31,57,31,203,31,15,31,80,31,80,30,97,31,97,30,97,29,75,31,75,30,78,31,78,30,78,29,78,28,78,27,8,31,98,31,58,31,8,31,171,31,118,31,238,31,238,30,47,31,90,31,210,31,114,31,114,30,227,31,190,31,56,31,101,31,94,31,79,31,79,30,185,31,217,31,198,31,239,31,69,31,188,31,169,31,169,30,54,31,83,31,83,30,83,29,184,31,184,30,133,31,158,31,163,31,187,31,207,31,64,31,240,31,79,31,223,31,44,31,22,31,187,31,216,31,85,31,75,31,128,31,49,31,49,30,247,31,247,30,18,31,82,31,89,31,252,31,252,30,77,31,67,31,38,31,205,31,151,31,151,30,29,31,146,31,169,31,14,31,45,31,232,31,118,31,62,31,209,31,174,31,99,31,3,31,242,31,191,31,169,31,23,31,74,31,101,31,26,31,128,31,161,31,236,31,142,31,142,30,142,29,142,28,49,31,24,31,15,31,63,31,66,31,1,31,183,31,73,31,91,31,253,31,19,31,174,31,41,31,41,30,25,31,86,31,247,31,151,31,151,30,41,31,173,31,90,31,60,31,81,31,58,31,51,31,210,31,244,31,249,31,183,31,183,30,144,31,144,30,68,31,68,30,68,29,143,31,179,31,253,31,251,31,255,31,138,31,102,31,102,30,106,31,120,31,120,30,59,31,66,31,196,31,196,30,23,31,145,31,145,30,201,31,19,31,19,30,19,29,47,31,247,31,164,31,35,31,16,31,16,30,113,31,77,31,54,31,54,30,60,31,86,31,124,31,222,31,222,30,222,29,235,31,112,31,143,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
