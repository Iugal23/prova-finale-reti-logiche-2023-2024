-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_278 is
end project_tb_278;

architecture project_tb_arch_278 of project_tb_278 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 276;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,197,0,170,0,144,0,212,0,245,0,0,0,7,0,26,0,199,0,88,0,253,0,69,0,177,0,196,0,116,0,0,0,15,0,238,0,195,0,228,0,0,0,0,0,201,0,0,0,225,0,36,0,71,0,233,0,83,0,0,0,183,0,108,0,203,0,184,0,1,0,233,0,237,0,99,0,209,0,32,0,194,0,5,0,163,0,0,0,0,0,18,0,0,0,58,0,121,0,19,0,132,0,110,0,220,0,0,0,9,0,188,0,247,0,74,0,187,0,57,0,251,0,29,0,25,0,44,0,115,0,127,0,58,0,122,0,17,0,14,0,0,0,43,0,246,0,125,0,137,0,230,0,169,0,61,0,0,0,0,0,24,0,251,0,238,0,242,0,209,0,82,0,197,0,101,0,21,0,98,0,18,0,188,0,0,0,242,0,0,0,0,0,145,0,194,0,255,0,60,0,136,0,17,0,210,0,120,0,207,0,0,0,237,0,15,0,0,0,72,0,125,0,100,0,48,0,0,0,144,0,167,0,46,0,49,0,207,0,0,0,0,0,215,0,47,0,18,0,9,0,37,0,236,0,139,0,0,0,115,0,0,0,0,0,0,0,0,0,152,0,29,0,146,0,57,0,3,0,58,0,89,0,0,0,241,0,0,0,172,0,246,0,0,0,216,0,177,0,0,0,184,0,0,0,130,0,19,0,251,0,162,0,0,0,200,0,0,0,211,0,0,0,4,0,208,0,247,0,2,0,25,0,103,0,0,0,255,0,50,0,121,0,129,0,14,0,42,0,0,0,0,0,126,0,231,0,106,0,69,0,0,0,167,0,174,0,32,0,201,0,213,0,47,0,204,0,252,0,79,0,0,0,0,0,206,0,43,0,176,0,0,0,85,0,194,0,215,0,196,0,194,0,0,0,0,0,247,0,3,0,231,0,195,0,139,0,40,0,49,0,65,0,168,0,29,0,237,0,114,0,142,0,31,0,98,0,130,0,129,0,24,0,124,0,146,0,104,0,0,0,184,0,15,0,52,0,0,0,54,0,108,0,172,0,0,0,94,0,205,0,26,0,222,0,134,0,247,0,0,0,222,0,65,0,143,0,22,0,171,0,191,0,172,0,0,0,189,0,0,0,104,0,5,0,0,0,0,0,108,0,0,0,225,0,146,0,217,0,241,0,211,0,33,0,0,0,241,0,0,0,102,0,138,0,107,0,95,0,184,0,203,0,23,0,57,0,132,0,164,0);
signal scenario_full  : scenario_type := (133,31,197,31,170,31,144,31,212,31,245,31,245,30,7,31,26,31,199,31,88,31,253,31,69,31,177,31,196,31,116,31,116,30,15,31,238,31,195,31,228,31,228,30,228,29,201,31,201,30,225,31,36,31,71,31,233,31,83,31,83,30,183,31,108,31,203,31,184,31,1,31,233,31,237,31,99,31,209,31,32,31,194,31,5,31,163,31,163,30,163,29,18,31,18,30,58,31,121,31,19,31,132,31,110,31,220,31,220,30,9,31,188,31,247,31,74,31,187,31,57,31,251,31,29,31,25,31,44,31,115,31,127,31,58,31,122,31,17,31,14,31,14,30,43,31,246,31,125,31,137,31,230,31,169,31,61,31,61,30,61,29,24,31,251,31,238,31,242,31,209,31,82,31,197,31,101,31,21,31,98,31,18,31,188,31,188,30,242,31,242,30,242,29,145,31,194,31,255,31,60,31,136,31,17,31,210,31,120,31,207,31,207,30,237,31,15,31,15,30,72,31,125,31,100,31,48,31,48,30,144,31,167,31,46,31,49,31,207,31,207,30,207,29,215,31,47,31,18,31,9,31,37,31,236,31,139,31,139,30,115,31,115,30,115,29,115,28,115,27,152,31,29,31,146,31,57,31,3,31,58,31,89,31,89,30,241,31,241,30,172,31,246,31,246,30,216,31,177,31,177,30,184,31,184,30,130,31,19,31,251,31,162,31,162,30,200,31,200,30,211,31,211,30,4,31,208,31,247,31,2,31,25,31,103,31,103,30,255,31,50,31,121,31,129,31,14,31,42,31,42,30,42,29,126,31,231,31,106,31,69,31,69,30,167,31,174,31,32,31,201,31,213,31,47,31,204,31,252,31,79,31,79,30,79,29,206,31,43,31,176,31,176,30,85,31,194,31,215,31,196,31,194,31,194,30,194,29,247,31,3,31,231,31,195,31,139,31,40,31,49,31,65,31,168,31,29,31,237,31,114,31,142,31,31,31,98,31,130,31,129,31,24,31,124,31,146,31,104,31,104,30,184,31,15,31,52,31,52,30,54,31,108,31,172,31,172,30,94,31,205,31,26,31,222,31,134,31,247,31,247,30,222,31,65,31,143,31,22,31,171,31,191,31,172,31,172,30,189,31,189,30,104,31,5,31,5,30,5,29,108,31,108,30,225,31,146,31,217,31,241,31,211,31,33,31,33,30,241,31,241,30,102,31,138,31,107,31,95,31,184,31,203,31,23,31,57,31,132,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
