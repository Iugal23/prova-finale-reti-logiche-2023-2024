-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_311 is
end project_tb_311;

architecture project_tb_arch_311 of project_tb_311 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 939;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,0,0,112,0,9,0,0,0,229,0,40,0,181,0,150,0,0,0,0,0,244,0,82,0,163,0,57,0,158,0,0,0,199,0,10,0,145,0,58,0,0,0,118,0,73,0,103,0,0,0,197,0,13,0,183,0,0,0,0,0,32,0,0,0,21,0,103,0,248,0,0,0,11,0,196,0,154,0,206,0,239,0,34,0,154,0,60,0,85,0,0,0,89,0,73,0,43,0,0,0,0,0,26,0,29,0,55,0,106,0,143,0,0,0,111,0,170,0,98,0,0,0,194,0,0,0,141,0,133,0,0,0,230,0,186,0,104,0,0,0,98,0,84,0,53,0,202,0,107,0,0,0,0,0,0,0,207,0,219,0,32,0,187,0,234,0,72,0,254,0,109,0,149,0,75,0,21,0,171,0,182,0,0,0,135,0,114,0,86,0,6,0,188,0,0,0,0,0,71,0,34,0,64,0,148,0,19,0,177,0,0,0,90,0,58,0,161,0,25,0,79,0,195,0,148,0,74,0,224,0,15,0,177,0,67,0,164,0,15,0,203,0,106,0,0,0,0,0,61,0,89,0,241,0,152,0,0,0,228,0,177,0,144,0,67,0,152,0,218,0,121,0,248,0,219,0,6,0,125,0,53,0,15,0,0,0,204,0,113,0,25,0,97,0,187,0,27,0,5,0,212,0,92,0,162,0,49,0,228,0,0,0,10,0,129,0,0,0,162,0,210,0,0,0,0,0,227,0,56,0,0,0,161,0,231,0,218,0,216,0,61,0,0,0,0,0,140,0,77,0,20,0,30,0,25,0,128,0,154,0,147,0,97,0,109,0,225,0,229,0,138,0,0,0,11,0,57,0,0,0,127,0,168,0,121,0,191,0,0,0,71,0,38,0,221,0,48,0,9,0,198,0,177,0,177,0,138,0,0,0,117,0,181,0,245,0,168,0,0,0,158,0,139,0,18,0,22,0,148,0,16,0,0,0,212,0,57,0,142,0,44,0,83,0,42,0,107,0,83,0,58,0,213,0,30,0,217,0,190,0,108,0,221,0,175,0,0,0,0,0,197,0,0,0,166,0,102,0,0,0,228,0,72,0,0,0,141,0,231,0,0,0,26,0,0,0,85,0,52,0,0,0,100,0,86,0,101,0,0,0,218,0,0,0,87,0,218,0,230,0,100,0,161,0,0,0,74,0,109,0,135,0,53,0,0,0,108,0,0,0,75,0,122,0,169,0,0,0,136,0,67,0,196,0,183,0,0,0,253,0,22,0,88,0,200,0,5,0,253,0,185,0,77,0,0,0,236,0,0,0,0,0,0,0,98,0,141,0,0,0,132,0,196,0,243,0,158,0,0,0,246,0,0,0,80,0,0,0,45,0,77,0,104,0,132,0,199,0,77,0,6,0,90,0,13,0,253,0,145,0,62,0,240,0,235,0,169,0,118,0,88,0,46,0,100,0,176,0,0,0,200,0,0,0,0,0,12,0,58,0,0,0,0,0,59,0,130,0,60,0,122,0,0,0,61,0,0,0,14,0,197,0,9,0,53,0,39,0,34,0,161,0,89,0,170,0,215,0,27,0,78,0,202,0,204,0,0,0,92,0,18,0,0,0,223,0,207,0,175,0,239,0,61,0,3,0,131,0,146,0,12,0,123,0,0,0,182,0,210,0,0,0,51,0,28,0,241,0,0,0,64,0,0,0,86,0,69,0,229,0,199,0,111,0,85,0,21,0,0,0,7,0,220,0,0,0,183,0,167,0,243,0,0,0,11,0,184,0,0,0,79,0,164,0,0,0,210,0,200,0,251,0,0,0,2,0,133,0,0,0,213,0,134,0,0,0,254,0,46,0,8,0,20,0,47,0,183,0,81,0,0,0,191,0,109,0,184,0,0,0,122,0,96,0,76,0,0,0,115,0,0,0,12,0,93,0,24,0,160,0,57,0,16,0,250,0,137,0,66,0,234,0,132,0,86,0,2,0,242,0,112,0,138,0,0,0,129,0,65,0,41,0,42,0,0,0,224,0,214,0,198,0,200,0,220,0,249,0,11,0,226,0,161,0,0,0,21,0,197,0,43,0,62,0,12,0,94,0,103,0,199,0,189,0,186,0,32,0,186,0,224,0,240,0,94,0,80,0,52,0,14,0,231,0,237,0,0,0,0,0,0,0,186,0,127,0,249,0,98,0,0,0,23,0,133,0,0,0,194,0,51,0,205,0,0,0,3,0,10,0,66,0,221,0,151,0,192,0,250,0,106,0,32,0,142,0,190,0,58,0,137,0,254,0,31,0,163,0,87,0,36,0,0,0,104,0,220,0,255,0,245,0,0,0,11,0,102,0,0,0,0,0,0,0,233,0,130,0,109,0,83,0,4,0,11,0,9,0,198,0,105,0,0,0,133,0,163,0,198,0,203,0,22,0,60,0,0,0,137,0,173,0,0,0,0,0,154,0,36,0,85,0,222,0,198,0,191,0,169,0,216,0,11,0,35,0,0,0,137,0,0,0,0,0,184,0,187,0,0,0,91,0,23,0,130,0,158,0,0,0,0,0,125,0,0,0,191,0,229,0,170,0,126,0,209,0,172,0,0,0,67,0,0,0,0,0,133,0,179,0,64,0,168,0,166,0,0,0,131,0,248,0,177,0,0,0,0,0,0,0,0,0,230,0,72,0,192,0,228,0,149,0,42,0,103,0,50,0,148,0,221,0,73,0,49,0,133,0,91,0,5,0,184,0,108,0,191,0,191,0,150,0,34,0,37,0,200,0,144,0,44,0,74,0,0,0,187,0,0,0,107,0,45,0,189,0,200,0,127,0,212,0,189,0,197,0,73,0,233,0,0,0,0,0,163,0,84,0,67,0,87,0,67,0,229,0,7,0,145,0,174,0,108,0,0,0,148,0,62,0,183,0,0,0,191,0,238,0,50,0,110,0,74,0,131,0,165,0,177,0,0,0,134,0,95,0,0,0,166,0,64,0,57,0,0,0,0,0,100,0,28,0,249,0,39,0,149,0,154,0,151,0,63,0,200,0,31,0,0,0,111,0,111,0,0,0,87,0,226,0,250,0,59,0,197,0,172,0,165,0,0,0,245,0,0,0,228,0,135,0,0,0,204,0,201,0,84,0,95,0,0,0,181,0,224,0,214,0,108,0,205,0,0,0,164,0,146,0,51,0,122,0,191,0,0,0,0,0,196,0,222,0,170,0,22,0,252,0,232,0,81,0,103,0,152,0,196,0,51,0,2,0,207,0,0,0,57,0,189,0,28,0,203,0,83,0,0,0,238,0,214,0,81,0,21,0,212,0,236,0,58,0,66,0,142,0,0,0,45,0,0,0,206,0,29,0,166,0,0,0,140,0,130,0,141,0,121,0,40,0,0,0,99,0,33,0,35,0,0,0,6,0,168,0,90,0,122,0,137,0,37,0,0,0,220,0,17,0,52,0,0,0,143,0,0,0,55,0,152,0,0,0,0,0,252,0,128,0,227,0,44,0,0,0,126,0,176,0,18,0,40,0,187,0,88,0,201,0,189,0,240,0,18,0,119,0,0,0,234,0,7,0,194,0,101,0,48,0,134,0,134,0,0,0,9,0,44,0,216,0,210,0,0,0,192,0,0,0,222,0,50,0,208,0,0,0,183,0,125,0,184,0,160,0,56,0,0,0,0,0,0,0,62,0,0,0,157,0,23,0,95,0,155,0,121,0,223,0,191,0,26,0,187,0,0,0,9,0,26,0,173,0,120,0,140,0,0,0,128,0,220,0,54,0,66,0,252,0,9,0,73,0,172,0,139,0,38,0,232,0,109,0,185,0,0,0,0,0,81,0,169,0,157,0,0,0,145,0,39,0,241,0,235,0,179,0,0,0,0,0,142,0,57,0,43,0,61,0,161,0,58,0,47,0,250,0,0,0,113,0,29,0,3,0,0,0,67,0,0,0,1,0,150,0,76,0,217,0,209,0,0,0,171,0,208,0,0,0,122,0,45,0,108,0,66,0,19,0,253,0,125,0,138,0,102,0,109,0,101,0,0,0,238,0,176,0,114,0,246,0,47,0,196,0,225,0,218,0,103,0,49,0,0,0,0,0,0,0,9,0,252,0,42,0,220,0,162,0,48,0,0,0,44,0,0,0,173,0,255,0,139,0,18,0,188,0,148,0,127,0,221,0,0,0,217,0,137,0,38,0,49,0,152,0,24,0,176,0,54,0,0,0,91,0,116,0);
signal scenario_full  : scenario_type := (105,31,105,30,112,31,9,31,9,30,229,31,40,31,181,31,150,31,150,30,150,29,244,31,82,31,163,31,57,31,158,31,158,30,199,31,10,31,145,31,58,31,58,30,118,31,73,31,103,31,103,30,197,31,13,31,183,31,183,30,183,29,32,31,32,30,21,31,103,31,248,31,248,30,11,31,196,31,154,31,206,31,239,31,34,31,154,31,60,31,85,31,85,30,89,31,73,31,43,31,43,30,43,29,26,31,29,31,55,31,106,31,143,31,143,30,111,31,170,31,98,31,98,30,194,31,194,30,141,31,133,31,133,30,230,31,186,31,104,31,104,30,98,31,84,31,53,31,202,31,107,31,107,30,107,29,107,28,207,31,219,31,32,31,187,31,234,31,72,31,254,31,109,31,149,31,75,31,21,31,171,31,182,31,182,30,135,31,114,31,86,31,6,31,188,31,188,30,188,29,71,31,34,31,64,31,148,31,19,31,177,31,177,30,90,31,58,31,161,31,25,31,79,31,195,31,148,31,74,31,224,31,15,31,177,31,67,31,164,31,15,31,203,31,106,31,106,30,106,29,61,31,89,31,241,31,152,31,152,30,228,31,177,31,144,31,67,31,152,31,218,31,121,31,248,31,219,31,6,31,125,31,53,31,15,31,15,30,204,31,113,31,25,31,97,31,187,31,27,31,5,31,212,31,92,31,162,31,49,31,228,31,228,30,10,31,129,31,129,30,162,31,210,31,210,30,210,29,227,31,56,31,56,30,161,31,231,31,218,31,216,31,61,31,61,30,61,29,140,31,77,31,20,31,30,31,25,31,128,31,154,31,147,31,97,31,109,31,225,31,229,31,138,31,138,30,11,31,57,31,57,30,127,31,168,31,121,31,191,31,191,30,71,31,38,31,221,31,48,31,9,31,198,31,177,31,177,31,138,31,138,30,117,31,181,31,245,31,168,31,168,30,158,31,139,31,18,31,22,31,148,31,16,31,16,30,212,31,57,31,142,31,44,31,83,31,42,31,107,31,83,31,58,31,213,31,30,31,217,31,190,31,108,31,221,31,175,31,175,30,175,29,197,31,197,30,166,31,102,31,102,30,228,31,72,31,72,30,141,31,231,31,231,30,26,31,26,30,85,31,52,31,52,30,100,31,86,31,101,31,101,30,218,31,218,30,87,31,218,31,230,31,100,31,161,31,161,30,74,31,109,31,135,31,53,31,53,30,108,31,108,30,75,31,122,31,169,31,169,30,136,31,67,31,196,31,183,31,183,30,253,31,22,31,88,31,200,31,5,31,253,31,185,31,77,31,77,30,236,31,236,30,236,29,236,28,98,31,141,31,141,30,132,31,196,31,243,31,158,31,158,30,246,31,246,30,80,31,80,30,45,31,77,31,104,31,132,31,199,31,77,31,6,31,90,31,13,31,253,31,145,31,62,31,240,31,235,31,169,31,118,31,88,31,46,31,100,31,176,31,176,30,200,31,200,30,200,29,12,31,58,31,58,30,58,29,59,31,130,31,60,31,122,31,122,30,61,31,61,30,14,31,197,31,9,31,53,31,39,31,34,31,161,31,89,31,170,31,215,31,27,31,78,31,202,31,204,31,204,30,92,31,18,31,18,30,223,31,207,31,175,31,239,31,61,31,3,31,131,31,146,31,12,31,123,31,123,30,182,31,210,31,210,30,51,31,28,31,241,31,241,30,64,31,64,30,86,31,69,31,229,31,199,31,111,31,85,31,21,31,21,30,7,31,220,31,220,30,183,31,167,31,243,31,243,30,11,31,184,31,184,30,79,31,164,31,164,30,210,31,200,31,251,31,251,30,2,31,133,31,133,30,213,31,134,31,134,30,254,31,46,31,8,31,20,31,47,31,183,31,81,31,81,30,191,31,109,31,184,31,184,30,122,31,96,31,76,31,76,30,115,31,115,30,12,31,93,31,24,31,160,31,57,31,16,31,250,31,137,31,66,31,234,31,132,31,86,31,2,31,242,31,112,31,138,31,138,30,129,31,65,31,41,31,42,31,42,30,224,31,214,31,198,31,200,31,220,31,249,31,11,31,226,31,161,31,161,30,21,31,197,31,43,31,62,31,12,31,94,31,103,31,199,31,189,31,186,31,32,31,186,31,224,31,240,31,94,31,80,31,52,31,14,31,231,31,237,31,237,30,237,29,237,28,186,31,127,31,249,31,98,31,98,30,23,31,133,31,133,30,194,31,51,31,205,31,205,30,3,31,10,31,66,31,221,31,151,31,192,31,250,31,106,31,32,31,142,31,190,31,58,31,137,31,254,31,31,31,163,31,87,31,36,31,36,30,104,31,220,31,255,31,245,31,245,30,11,31,102,31,102,30,102,29,102,28,233,31,130,31,109,31,83,31,4,31,11,31,9,31,198,31,105,31,105,30,133,31,163,31,198,31,203,31,22,31,60,31,60,30,137,31,173,31,173,30,173,29,154,31,36,31,85,31,222,31,198,31,191,31,169,31,216,31,11,31,35,31,35,30,137,31,137,30,137,29,184,31,187,31,187,30,91,31,23,31,130,31,158,31,158,30,158,29,125,31,125,30,191,31,229,31,170,31,126,31,209,31,172,31,172,30,67,31,67,30,67,29,133,31,179,31,64,31,168,31,166,31,166,30,131,31,248,31,177,31,177,30,177,29,177,28,177,27,230,31,72,31,192,31,228,31,149,31,42,31,103,31,50,31,148,31,221,31,73,31,49,31,133,31,91,31,5,31,184,31,108,31,191,31,191,31,150,31,34,31,37,31,200,31,144,31,44,31,74,31,74,30,187,31,187,30,107,31,45,31,189,31,200,31,127,31,212,31,189,31,197,31,73,31,233,31,233,30,233,29,163,31,84,31,67,31,87,31,67,31,229,31,7,31,145,31,174,31,108,31,108,30,148,31,62,31,183,31,183,30,191,31,238,31,50,31,110,31,74,31,131,31,165,31,177,31,177,30,134,31,95,31,95,30,166,31,64,31,57,31,57,30,57,29,100,31,28,31,249,31,39,31,149,31,154,31,151,31,63,31,200,31,31,31,31,30,111,31,111,31,111,30,87,31,226,31,250,31,59,31,197,31,172,31,165,31,165,30,245,31,245,30,228,31,135,31,135,30,204,31,201,31,84,31,95,31,95,30,181,31,224,31,214,31,108,31,205,31,205,30,164,31,146,31,51,31,122,31,191,31,191,30,191,29,196,31,222,31,170,31,22,31,252,31,232,31,81,31,103,31,152,31,196,31,51,31,2,31,207,31,207,30,57,31,189,31,28,31,203,31,83,31,83,30,238,31,214,31,81,31,21,31,212,31,236,31,58,31,66,31,142,31,142,30,45,31,45,30,206,31,29,31,166,31,166,30,140,31,130,31,141,31,121,31,40,31,40,30,99,31,33,31,35,31,35,30,6,31,168,31,90,31,122,31,137,31,37,31,37,30,220,31,17,31,52,31,52,30,143,31,143,30,55,31,152,31,152,30,152,29,252,31,128,31,227,31,44,31,44,30,126,31,176,31,18,31,40,31,187,31,88,31,201,31,189,31,240,31,18,31,119,31,119,30,234,31,7,31,194,31,101,31,48,31,134,31,134,31,134,30,9,31,44,31,216,31,210,31,210,30,192,31,192,30,222,31,50,31,208,31,208,30,183,31,125,31,184,31,160,31,56,31,56,30,56,29,56,28,62,31,62,30,157,31,23,31,95,31,155,31,121,31,223,31,191,31,26,31,187,31,187,30,9,31,26,31,173,31,120,31,140,31,140,30,128,31,220,31,54,31,66,31,252,31,9,31,73,31,172,31,139,31,38,31,232,31,109,31,185,31,185,30,185,29,81,31,169,31,157,31,157,30,145,31,39,31,241,31,235,31,179,31,179,30,179,29,142,31,57,31,43,31,61,31,161,31,58,31,47,31,250,31,250,30,113,31,29,31,3,31,3,30,67,31,67,30,1,31,150,31,76,31,217,31,209,31,209,30,171,31,208,31,208,30,122,31,45,31,108,31,66,31,19,31,253,31,125,31,138,31,102,31,109,31,101,31,101,30,238,31,176,31,114,31,246,31,47,31,196,31,225,31,218,31,103,31,49,31,49,30,49,29,49,28,9,31,252,31,42,31,220,31,162,31,48,31,48,30,44,31,44,30,173,31,255,31,139,31,18,31,188,31,148,31,127,31,221,31,221,30,217,31,137,31,38,31,49,31,152,31,24,31,176,31,54,31,54,30,91,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
