-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 768;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (3,0,82,0,194,0,213,0,0,0,70,0,228,0,37,0,0,0,0,0,1,0,0,0,137,0,72,0,201,0,61,0,62,0,146,0,131,0,70,0,86,0,132,0,76,0,43,0,49,0,107,0,238,0,32,0,68,0,0,0,32,0,21,0,101,0,110,0,89,0,0,0,4,0,109,0,190,0,15,0,215,0,164,0,55,0,181,0,187,0,0,0,13,0,0,0,76,0,117,0,23,0,245,0,45,0,140,0,201,0,49,0,84,0,62,0,119,0,118,0,252,0,140,0,162,0,117,0,2,0,182,0,0,0,0,0,190,0,0,0,0,0,92,0,239,0,72,0,37,0,0,0,46,0,236,0,173,0,234,0,249,0,34,0,225,0,88,0,172,0,0,0,134,0,38,0,76,0,247,0,169,0,0,0,0,0,137,0,48,0,15,0,7,0,183,0,80,0,0,0,136,0,167,0,40,0,0,0,143,0,3,0,224,0,0,0,180,0,0,0,52,0,198,0,193,0,239,0,0,0,66,0,6,0,17,0,236,0,127,0,65,0,194,0,48,0,212,0,172,0,120,0,253,0,244,0,197,0,109,0,18,0,0,0,72,0,191,0,1,0,0,0,0,0,155,0,203,0,0,0,206,0,90,0,0,0,0,0,28,0,230,0,159,0,174,0,236,0,37,0,19,0,157,0,145,0,0,0,131,0,0,0,0,0,197,0,198,0,255,0,0,0,35,0,10,0,0,0,6,0,177,0,83,0,244,0,0,0,68,0,17,0,98,0,231,0,22,0,0,0,183,0,255,0,138,0,0,0,139,0,213,0,113,0,144,0,28,0,213,0,152,0,73,0,118,0,78,0,154,0,41,0,0,0,207,0,0,0,2,0,24,0,106,0,217,0,0,0,62,0,224,0,0,0,24,0,227,0,211,0,243,0,159,0,91,0,163,0,149,0,54,0,0,0,37,0,12,0,62,0,0,0,216,0,179,0,0,0,0,0,255,0,159,0,25,0,140,0,235,0,238,0,51,0,16,0,166,0,188,0,9,0,0,0,242,0,31,0,0,0,72,0,97,0,30,0,0,0,94,0,0,0,44,0,64,0,42,0,0,0,23,0,71,0,44,0,188,0,181,0,153,0,0,0,0,0,74,0,135,0,0,0,0,0,227,0,74,0,232,0,71,0,0,0,185,0,20,0,235,0,118,0,0,0,0,0,246,0,16,0,181,0,75,0,32,0,0,0,120,0,100,0,0,0,146,0,63,0,72,0,79,0,0,0,13,0,114,0,33,0,44,0,125,0,179,0,81,0,123,0,117,0,0,0,177,0,0,0,239,0,169,0,0,0,186,0,222,0,0,0,120,0,188,0,201,0,181,0,20,0,207,0,152,0,0,0,103,0,12,0,0,0,38,0,23,0,9,0,0,0,0,0,0,0,20,0,166,0,74,0,158,0,7,0,44,0,241,0,215,0,57,0,141,0,0,0,131,0,0,0,47,0,215,0,50,0,2,0,0,0,0,0,210,0,232,0,151,0,218,0,185,0,78,0,4,0,154,0,0,0,0,0,198,0,18,0,0,0,5,0,0,0,210,0,87,0,0,0,172,0,61,0,0,0,181,0,176,0,26,0,20,0,188,0,112,0,0,0,15,0,49,0,115,0,209,0,150,0,20,0,126,0,180,0,138,0,71,0,206,0,240,0,65,0,249,0,152,0,0,0,111,0,0,0,7,0,10,0,192,0,56,0,0,0,168,0,136,0,223,0,129,0,247,0,6,0,226,0,93,0,125,0,165,0,13,0,0,0,0,0,57,0,243,0,157,0,91,0,145,0,129,0,49,0,15,0,225,0,69,0,27,0,0,0,0,0,0,0,141,0,0,0,193,0,0,0,171,0,144,0,131,0,142,0,151,0,106,0,30,0,0,0,228,0,98,0,223,0,221,0,45,0,121,0,117,0,107,0,24,0,203,0,0,0,242,0,107,0,0,0,67,0,63,0,0,0,67,0,176,0,28,0,0,0,88,0,210,0,121,0,175,0,246,0,190,0,92,0,6,0,81,0,132,0,164,0,93,0,183,0,35,0,0,0,117,0,136,0,123,0,120,0,206,0,248,0,0,0,224,0,198,0,102,0,0,0,0,0,222,0,0,0,0,0,159,0,97,0,237,0,0,0,138,0,112,0,0,0,129,0,249,0,83,0,252,0,73,0,235,0,21,0,93,0,0,0,83,0,186,0,0,0,0,0,246,0,0,0,0,0,91,0,0,0,0,0,0,0,1,0,96,0,142,0,240,0,145,0,41,0,10,0,199,0,206,0,0,0,243,0,231,0,54,0,210,0,210,0,60,0,12,0,28,0,1,0,103,0,136,0,0,0,2,0,0,0,93,0,205,0,225,0,109,0,0,0,14,0,0,0,0,0,92,0,0,0,0,0,98,0,17,0,121,0,224,0,62,0,64,0,190,0,202,0,181,0,126,0,99,0,133,0,7,0,146,0,194,0,0,0,207,0,0,0,0,0,40,0,207,0,191,0,26,0,126,0,108,0,180,0,0,0,0,0,5,0,135,0,0,0,56,0,66,0,64,0,92,0,0,0,139,0,98,0,47,0,0,0,79,0,0,0,217,0,131,0,129,0,53,0,164,0,0,0,12,0,224,0,191,0,2,0,40,0,124,0,59,0,166,0,173,0,71,0,139,0,240,0,107,0,229,0,212,0,23,0,108,0,0,0,93,0,63,0,0,0,222,0,69,0,255,0,117,0,0,0,32,0,145,0,120,0,128,0,141,0,99,0,103,0,232,0,57,0,49,0,158,0,189,0,42,0,159,0,82,0,0,0,0,0,11,0,199,0,182,0,216,0,0,0,158,0,230,0,199,0,22,0,0,0,120,0,235,0,217,0,146,0,37,0,248,0,18,0,248,0,152,0,134,0,46,0,0,0,0,0,75,0,47,0,250,0,90,0,0,0,45,0,132,0,0,0,66,0,108,0,216,0,0,0,195,0,36,0,6,0,0,0,41,0,34,0,36,0,0,0,224,0,0,0,0,0,35,0,40,0,22,0,42,0,108,0,101,0,16,0,182,0,230,0,0,0,186,0,98,0,0,0,76,0,123,0,221,0,128,0,145,0,219,0,82,0,139,0,0,0,80,0,140,0,0,0,191,0,82,0,161,0,49,0,0,0,195,0,86,0,0,0,7,0,0,0,0,0,107,0,203,0,164,0,127,0,51,0,68,0,68,0,205,0,115,0,251,0,23,0,130,0,40,0,143,0,72,0,142,0,47,0,0,0,123,0,175,0,0,0,120,0,98,0,0,0,145,0,173,0,218,0,72,0,131,0,242,0,0,0,0,0,157,0,5,0,65,0,139,0,0,0,73,0,114,0,181,0,214,0,103,0,221,0,205,0,134,0,217,0,4,0,60,0,58,0,235,0,208,0,206,0,93,0,224,0,72,0,115,0);
signal scenario_full  : scenario_type := (3,31,82,31,194,31,213,31,213,30,70,31,228,31,37,31,37,30,37,29,1,31,1,30,137,31,72,31,201,31,61,31,62,31,146,31,131,31,70,31,86,31,132,31,76,31,43,31,49,31,107,31,238,31,32,31,68,31,68,30,32,31,21,31,101,31,110,31,89,31,89,30,4,31,109,31,190,31,15,31,215,31,164,31,55,31,181,31,187,31,187,30,13,31,13,30,76,31,117,31,23,31,245,31,45,31,140,31,201,31,49,31,84,31,62,31,119,31,118,31,252,31,140,31,162,31,117,31,2,31,182,31,182,30,182,29,190,31,190,30,190,29,92,31,239,31,72,31,37,31,37,30,46,31,236,31,173,31,234,31,249,31,34,31,225,31,88,31,172,31,172,30,134,31,38,31,76,31,247,31,169,31,169,30,169,29,137,31,48,31,15,31,7,31,183,31,80,31,80,30,136,31,167,31,40,31,40,30,143,31,3,31,224,31,224,30,180,31,180,30,52,31,198,31,193,31,239,31,239,30,66,31,6,31,17,31,236,31,127,31,65,31,194,31,48,31,212,31,172,31,120,31,253,31,244,31,197,31,109,31,18,31,18,30,72,31,191,31,1,31,1,30,1,29,155,31,203,31,203,30,206,31,90,31,90,30,90,29,28,31,230,31,159,31,174,31,236,31,37,31,19,31,157,31,145,31,145,30,131,31,131,30,131,29,197,31,198,31,255,31,255,30,35,31,10,31,10,30,6,31,177,31,83,31,244,31,244,30,68,31,17,31,98,31,231,31,22,31,22,30,183,31,255,31,138,31,138,30,139,31,213,31,113,31,144,31,28,31,213,31,152,31,73,31,118,31,78,31,154,31,41,31,41,30,207,31,207,30,2,31,24,31,106,31,217,31,217,30,62,31,224,31,224,30,24,31,227,31,211,31,243,31,159,31,91,31,163,31,149,31,54,31,54,30,37,31,12,31,62,31,62,30,216,31,179,31,179,30,179,29,255,31,159,31,25,31,140,31,235,31,238,31,51,31,16,31,166,31,188,31,9,31,9,30,242,31,31,31,31,30,72,31,97,31,30,31,30,30,94,31,94,30,44,31,64,31,42,31,42,30,23,31,71,31,44,31,188,31,181,31,153,31,153,30,153,29,74,31,135,31,135,30,135,29,227,31,74,31,232,31,71,31,71,30,185,31,20,31,235,31,118,31,118,30,118,29,246,31,16,31,181,31,75,31,32,31,32,30,120,31,100,31,100,30,146,31,63,31,72,31,79,31,79,30,13,31,114,31,33,31,44,31,125,31,179,31,81,31,123,31,117,31,117,30,177,31,177,30,239,31,169,31,169,30,186,31,222,31,222,30,120,31,188,31,201,31,181,31,20,31,207,31,152,31,152,30,103,31,12,31,12,30,38,31,23,31,9,31,9,30,9,29,9,28,20,31,166,31,74,31,158,31,7,31,44,31,241,31,215,31,57,31,141,31,141,30,131,31,131,30,47,31,215,31,50,31,2,31,2,30,2,29,210,31,232,31,151,31,218,31,185,31,78,31,4,31,154,31,154,30,154,29,198,31,18,31,18,30,5,31,5,30,210,31,87,31,87,30,172,31,61,31,61,30,181,31,176,31,26,31,20,31,188,31,112,31,112,30,15,31,49,31,115,31,209,31,150,31,20,31,126,31,180,31,138,31,71,31,206,31,240,31,65,31,249,31,152,31,152,30,111,31,111,30,7,31,10,31,192,31,56,31,56,30,168,31,136,31,223,31,129,31,247,31,6,31,226,31,93,31,125,31,165,31,13,31,13,30,13,29,57,31,243,31,157,31,91,31,145,31,129,31,49,31,15,31,225,31,69,31,27,31,27,30,27,29,27,28,141,31,141,30,193,31,193,30,171,31,144,31,131,31,142,31,151,31,106,31,30,31,30,30,228,31,98,31,223,31,221,31,45,31,121,31,117,31,107,31,24,31,203,31,203,30,242,31,107,31,107,30,67,31,63,31,63,30,67,31,176,31,28,31,28,30,88,31,210,31,121,31,175,31,246,31,190,31,92,31,6,31,81,31,132,31,164,31,93,31,183,31,35,31,35,30,117,31,136,31,123,31,120,31,206,31,248,31,248,30,224,31,198,31,102,31,102,30,102,29,222,31,222,30,222,29,159,31,97,31,237,31,237,30,138,31,112,31,112,30,129,31,249,31,83,31,252,31,73,31,235,31,21,31,93,31,93,30,83,31,186,31,186,30,186,29,246,31,246,30,246,29,91,31,91,30,91,29,91,28,1,31,96,31,142,31,240,31,145,31,41,31,10,31,199,31,206,31,206,30,243,31,231,31,54,31,210,31,210,31,60,31,12,31,28,31,1,31,103,31,136,31,136,30,2,31,2,30,93,31,205,31,225,31,109,31,109,30,14,31,14,30,14,29,92,31,92,30,92,29,98,31,17,31,121,31,224,31,62,31,64,31,190,31,202,31,181,31,126,31,99,31,133,31,7,31,146,31,194,31,194,30,207,31,207,30,207,29,40,31,207,31,191,31,26,31,126,31,108,31,180,31,180,30,180,29,5,31,135,31,135,30,56,31,66,31,64,31,92,31,92,30,139,31,98,31,47,31,47,30,79,31,79,30,217,31,131,31,129,31,53,31,164,31,164,30,12,31,224,31,191,31,2,31,40,31,124,31,59,31,166,31,173,31,71,31,139,31,240,31,107,31,229,31,212,31,23,31,108,31,108,30,93,31,63,31,63,30,222,31,69,31,255,31,117,31,117,30,32,31,145,31,120,31,128,31,141,31,99,31,103,31,232,31,57,31,49,31,158,31,189,31,42,31,159,31,82,31,82,30,82,29,11,31,199,31,182,31,216,31,216,30,158,31,230,31,199,31,22,31,22,30,120,31,235,31,217,31,146,31,37,31,248,31,18,31,248,31,152,31,134,31,46,31,46,30,46,29,75,31,47,31,250,31,90,31,90,30,45,31,132,31,132,30,66,31,108,31,216,31,216,30,195,31,36,31,6,31,6,30,41,31,34,31,36,31,36,30,224,31,224,30,224,29,35,31,40,31,22,31,42,31,108,31,101,31,16,31,182,31,230,31,230,30,186,31,98,31,98,30,76,31,123,31,221,31,128,31,145,31,219,31,82,31,139,31,139,30,80,31,140,31,140,30,191,31,82,31,161,31,49,31,49,30,195,31,86,31,86,30,7,31,7,30,7,29,107,31,203,31,164,31,127,31,51,31,68,31,68,31,205,31,115,31,251,31,23,31,130,31,40,31,143,31,72,31,142,31,47,31,47,30,123,31,175,31,175,30,120,31,98,31,98,30,145,31,173,31,218,31,72,31,131,31,242,31,242,30,242,29,157,31,5,31,65,31,139,31,139,30,73,31,114,31,181,31,214,31,103,31,221,31,205,31,134,31,217,31,4,31,60,31,58,31,235,31,208,31,206,31,93,31,224,31,72,31,115,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
