-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1019;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (16,0,0,0,110,0,0,0,222,0,48,0,47,0,34,0,20,0,237,0,208,0,0,0,41,0,0,0,183,0,210,0,0,0,0,0,132,0,169,0,81,0,104,0,188,0,119,0,184,0,0,0,0,0,0,0,82,0,0,0,181,0,0,0,0,0,21,0,183,0,155,0,0,0,0,0,122,0,0,0,77,0,0,0,0,0,243,0,36,0,156,0,34,0,150,0,77,0,247,0,132,0,125,0,9,0,134,0,133,0,51,0,226,0,242,0,163,0,23,0,0,0,193,0,177,0,61,0,0,0,118,0,17,0,0,0,0,0,200,0,90,0,0,0,0,0,92,0,255,0,26,0,0,0,153,0,86,0,145,0,0,0,43,0,210,0,0,0,42,0,206,0,203,0,78,0,124,0,0,0,205,0,173,0,58,0,31,0,249,0,0,0,0,0,102,0,0,0,62,0,115,0,2,0,23,0,234,0,249,0,5,0,54,0,0,0,0,0,129,0,0,0,173,0,0,0,212,0,10,0,0,0,219,0,23,0,237,0,44,0,0,0,0,0,117,0,156,0,50,0,111,0,55,0,200,0,100,0,48,0,52,0,60,0,184,0,229,0,0,0,203,0,183,0,108,0,70,0,99,0,15,0,0,0,90,0,150,0,226,0,0,0,62,0,7,0,0,0,226,0,83,0,58,0,196,0,191,0,0,0,109,0,165,0,105,0,223,0,65,0,175,0,109,0,24,0,0,0,211,0,245,0,148,0,0,0,94,0,12,0,114,0,0,0,250,0,58,0,40,0,232,0,0,0,0,0,123,0,219,0,108,0,0,0,226,0,0,0,225,0,239,0,0,0,118,0,11,0,86,0,221,0,241,0,0,0,83,0,81,0,0,0,0,0,92,0,81,0,229,0,185,0,218,0,22,0,32,0,0,0,196,0,122,0,71,0,247,0,0,0,4,0,192,0,19,0,250,0,221,0,158,0,157,0,245,0,0,0,200,0,205,0,15,0,125,0,79,0,10,0,164,0,231,0,0,0,97,0,137,0,0,0,144,0,193,0,49,0,154,0,173,0,0,0,0,0,96,0,141,0,20,0,239,0,23,0,73,0,254,0,0,0,106,0,6,0,220,0,30,0,140,0,96,0,139,0,50,0,0,0,41,0,119,0,204,0,135,0,0,0,0,0,0,0,221,0,177,0,121,0,113,0,24,0,146,0,0,0,210,0,50,0,202,0,157,0,159,0,93,0,68,0,137,0,124,0,243,0,83,0,30,0,0,0,91,0,193,0,39,0,225,0,60,0,65,0,249,0,0,0,88,0,63,0,215,0,174,0,0,0,0,0,102,0,36,0,0,0,0,0,61,0,134,0,0,0,0,0,40,0,217,0,212,0,0,0,251,0,193,0,100,0,124,0,44,0,31,0,0,0,13,0,165,0,169,0,33,0,0,0,46,0,88,0,32,0,83,0,245,0,110,0,80,0,237,0,56,0,174,0,0,0,0,0,85,0,117,0,171,0,19,0,177,0,246,0,255,0,95,0,111,0,97,0,0,0,1,0,177,0,224,0,150,0,149,0,118,0,166,0,0,0,0,0,79,0,120,0,39,0,0,0,158,0,0,0,67,0,239,0,211,0,10,0,231,0,177,0,210,0,0,0,140,0,129,0,214,0,104,0,108,0,155,0,166,0,97,0,28,0,0,0,108,0,181,0,112,0,0,0,243,0,204,0,186,0,0,0,0,0,51,0,38,0,115,0,0,0,149,0,0,0,0,0,36,0,86,0,22,0,179,0,192,0,49,0,0,0,0,0,27,0,0,0,229,0,0,0,16,0,210,0,232,0,64,0,97,0,66,0,0,0,173,0,87,0,146,0,100,0,211,0,185,0,0,0,188,0,222,0,114,0,4,0,122,0,29,0,37,0,113,0,226,0,58,0,86,0,14,0,183,0,189,0,0,0,120,0,85,0,165,0,75,0,129,0,214,0,63,0,252,0,94,0,164,0,86,0,48,0,140,0,240,0,244,0,48,0,157,0,176,0,166,0,0,0,238,0,114,0,161,0,0,0,73,0,158,0,201,0,0,0,176,0,0,0,76,0,143,0,249,0,0,0,0,0,222,0,212,0,0,0,60,0,0,0,7,0,0,0,0,0,0,0,129,0,3,0,28,0,41,0,99,0,70,0,101,0,68,0,0,0,43,0,223,0,6,0,17,0,220,0,0,0,80,0,37,0,110,0,0,0,229,0,217,0,0,0,177,0,4,0,205,0,224,0,31,0,225,0,171,0,252,0,51,0,148,0,213,0,124,0,62,0,0,0,106,0,62,0,240,0,167,0,5,0,190,0,44,0,209,0,184,0,94,0,0,0,161,0,237,0,0,0,184,0,171,0,149,0,123,0,0,0,63,0,188,0,45,0,6,0,77,0,0,0,61,0,178,0,0,0,180,0,214,0,69,0,61,0,192,0,198,0,46,0,236,0,160,0,0,0,202,0,39,0,99,0,202,0,0,0,106,0,120,0,99,0,151,0,185,0,66,0,0,0,55,0,0,0,12,0,237,0,78,0,58,0,54,0,32,0,131,0,149,0,114,0,78,0,55,0,178,0,130,0,176,0,5,0,192,0,192,0,247,0,0,0,180,0,153,0,242,0,151,0,0,0,228,0,164,0,219,0,145,0,39,0,169,0,204,0,35,0,58,0,0,0,222,0,201,0,238,0,183,0,245,0,0,0,30,0,0,0,166,0,120,0,0,0,0,0,0,0,97,0,154,0,12,0,189,0,90,0,0,0,7,0,0,0,0,0,34,0,0,0,151,0,61,0,79,0,33,0,154,0,157,0,137,0,0,0,163,0,182,0,185,0,130,0,63,0,243,0,96,0,36,0,131,0,188,0,169,0,32,0,100,0,0,0,237,0,78,0,71,0,53,0,252,0,0,0,173,0,255,0,52,0,15,0,69,0,95,0,83,0,198,0,97,0,125,0,0,0,97,0,113,0,0,0,0,0,21,0,99,0,120,0,44,0,0,0,19,0,0,0,48,0,9,0,193,0,234,0,141,0,243,0,62,0,243,0,98,0,229,0,193,0,238,0,48,0,196,0,0,0,229,0,205,0,191,0,191,0,121,0,0,0,124,0,0,0,47,0,42,0,67,0,68,0,27,0,209,0,0,0,194,0,58,0,37,0,113,0,195,0,0,0,206,0,106,0,0,0,70,0,160,0,39,0,62,0,200,0,17,0,0,0,147,0,37,0,64,0,38,0,108,0,238,0,0,0,30,0,50,0,0,0,63,0,137,0,246,0,214,0,40,0,68,0,0,0,225,0,143,0,10,0,193,0,31,0,94,0,24,0,217,0,135,0,70,0,223,0,45,0,0,0,237,0,233,0,0,0,62,0,165,0,0,0,68,0,235,0,0,0,67,0,145,0,0,0,248,0,38,0,147,0,0,0,90,0,11,0,62,0,154,0,205,0,224,0,45,0,105,0,0,0,149,0,225,0,147,0,174,0,0,0,0,0,165,0,85,0,0,0,204,0,234,0,0,0,35,0,0,0,0,0,185,0,126,0,0,0,2,0,93,0,48,0,162,0,204,0,147,0,235,0,117,0,0,0,204,0,149,0,189,0,0,0,48,0,164,0,0,0,0,0,83,0,0,0,9,0,96,0,113,0,77,0,70,0,96,0,157,0,35,0,137,0,0,0,219,0,223,0,186,0,78,0,167,0,27,0,139,0,252,0,214,0,0,0,3,0,199,0,159,0,206,0,0,0,227,0,92,0,15,0,180,0,211,0,175,0,1,0,108,0,178,0,205,0,231,0,136,0,118,0,207,0,157,0,156,0,0,0,86,0,196,0,204,0,242,0,154,0,194,0,145,0,221,0,21,0,173,0,171,0,85,0,2,0,69,0,40,0,189,0,224,0,59,0,151,0,249,0,101,0,0,0,0,0,58,0,0,0,253,0,170,0,123,0,246,0,124,0,234,0,0,0,170,0,30,0,178,0,82,0,91,0,27,0,107,0,182,0,0,0,149,0,0,0,2,0,0,0,125,0,131,0,202,0,112,0,216,0,47,0,152,0,249,0,171,0,185,0,176,0,120,0,0,0,204,0,86,0,253,0,188,0,192,0,32,0,0,0,175,0,255,0,133,0,76,0,16,0,0,0,131,0,0,0,0,0,238,0,89,0,248,0,191,0,174,0,26,0,0,0,27,0,26,0,144,0,160,0,0,0,114,0,0,0,87,0,77,0,0,0,146,0,0,0,154,0,6,0,229,0,107,0,241,0,151,0,57,0,247,0,224,0,0,0,0,0,145,0,78,0,0,0,0,0,75,0,157,0,247,0,76,0,6,0,29,0,164,0,235,0,235,0,162,0,186,0,159,0,61,0,0,0,220,0,0,0,144,0,80,0,0,0,0,0,211,0,100,0,106,0,112,0,0,0,0,0,5,0,252,0,138,0,69,0,224,0,96,0,80,0,0,0,45,0,21,0,159,0,0,0,0,0,38,0,18,0,91,0,27,0,165,0,168,0,231,0,52,0,195,0,29,0,0,0,108,0,168,0,0,0,0,0,3,0,184,0,223,0,80,0);
signal scenario_full  : scenario_type := (16,31,16,30,110,31,110,30,222,31,48,31,47,31,34,31,20,31,237,31,208,31,208,30,41,31,41,30,183,31,210,31,210,30,210,29,132,31,169,31,81,31,104,31,188,31,119,31,184,31,184,30,184,29,184,28,82,31,82,30,181,31,181,30,181,29,21,31,183,31,155,31,155,30,155,29,122,31,122,30,77,31,77,30,77,29,243,31,36,31,156,31,34,31,150,31,77,31,247,31,132,31,125,31,9,31,134,31,133,31,51,31,226,31,242,31,163,31,23,31,23,30,193,31,177,31,61,31,61,30,118,31,17,31,17,30,17,29,200,31,90,31,90,30,90,29,92,31,255,31,26,31,26,30,153,31,86,31,145,31,145,30,43,31,210,31,210,30,42,31,206,31,203,31,78,31,124,31,124,30,205,31,173,31,58,31,31,31,249,31,249,30,249,29,102,31,102,30,62,31,115,31,2,31,23,31,234,31,249,31,5,31,54,31,54,30,54,29,129,31,129,30,173,31,173,30,212,31,10,31,10,30,219,31,23,31,237,31,44,31,44,30,44,29,117,31,156,31,50,31,111,31,55,31,200,31,100,31,48,31,52,31,60,31,184,31,229,31,229,30,203,31,183,31,108,31,70,31,99,31,15,31,15,30,90,31,150,31,226,31,226,30,62,31,7,31,7,30,226,31,83,31,58,31,196,31,191,31,191,30,109,31,165,31,105,31,223,31,65,31,175,31,109,31,24,31,24,30,211,31,245,31,148,31,148,30,94,31,12,31,114,31,114,30,250,31,58,31,40,31,232,31,232,30,232,29,123,31,219,31,108,31,108,30,226,31,226,30,225,31,239,31,239,30,118,31,11,31,86,31,221,31,241,31,241,30,83,31,81,31,81,30,81,29,92,31,81,31,229,31,185,31,218,31,22,31,32,31,32,30,196,31,122,31,71,31,247,31,247,30,4,31,192,31,19,31,250,31,221,31,158,31,157,31,245,31,245,30,200,31,205,31,15,31,125,31,79,31,10,31,164,31,231,31,231,30,97,31,137,31,137,30,144,31,193,31,49,31,154,31,173,31,173,30,173,29,96,31,141,31,20,31,239,31,23,31,73,31,254,31,254,30,106,31,6,31,220,31,30,31,140,31,96,31,139,31,50,31,50,30,41,31,119,31,204,31,135,31,135,30,135,29,135,28,221,31,177,31,121,31,113,31,24,31,146,31,146,30,210,31,50,31,202,31,157,31,159,31,93,31,68,31,137,31,124,31,243,31,83,31,30,31,30,30,91,31,193,31,39,31,225,31,60,31,65,31,249,31,249,30,88,31,63,31,215,31,174,31,174,30,174,29,102,31,36,31,36,30,36,29,61,31,134,31,134,30,134,29,40,31,217,31,212,31,212,30,251,31,193,31,100,31,124,31,44,31,31,31,31,30,13,31,165,31,169,31,33,31,33,30,46,31,88,31,32,31,83,31,245,31,110,31,80,31,237,31,56,31,174,31,174,30,174,29,85,31,117,31,171,31,19,31,177,31,246,31,255,31,95,31,111,31,97,31,97,30,1,31,177,31,224,31,150,31,149,31,118,31,166,31,166,30,166,29,79,31,120,31,39,31,39,30,158,31,158,30,67,31,239,31,211,31,10,31,231,31,177,31,210,31,210,30,140,31,129,31,214,31,104,31,108,31,155,31,166,31,97,31,28,31,28,30,108,31,181,31,112,31,112,30,243,31,204,31,186,31,186,30,186,29,51,31,38,31,115,31,115,30,149,31,149,30,149,29,36,31,86,31,22,31,179,31,192,31,49,31,49,30,49,29,27,31,27,30,229,31,229,30,16,31,210,31,232,31,64,31,97,31,66,31,66,30,173,31,87,31,146,31,100,31,211,31,185,31,185,30,188,31,222,31,114,31,4,31,122,31,29,31,37,31,113,31,226,31,58,31,86,31,14,31,183,31,189,31,189,30,120,31,85,31,165,31,75,31,129,31,214,31,63,31,252,31,94,31,164,31,86,31,48,31,140,31,240,31,244,31,48,31,157,31,176,31,166,31,166,30,238,31,114,31,161,31,161,30,73,31,158,31,201,31,201,30,176,31,176,30,76,31,143,31,249,31,249,30,249,29,222,31,212,31,212,30,60,31,60,30,7,31,7,30,7,29,7,28,129,31,3,31,28,31,41,31,99,31,70,31,101,31,68,31,68,30,43,31,223,31,6,31,17,31,220,31,220,30,80,31,37,31,110,31,110,30,229,31,217,31,217,30,177,31,4,31,205,31,224,31,31,31,225,31,171,31,252,31,51,31,148,31,213,31,124,31,62,31,62,30,106,31,62,31,240,31,167,31,5,31,190,31,44,31,209,31,184,31,94,31,94,30,161,31,237,31,237,30,184,31,171,31,149,31,123,31,123,30,63,31,188,31,45,31,6,31,77,31,77,30,61,31,178,31,178,30,180,31,214,31,69,31,61,31,192,31,198,31,46,31,236,31,160,31,160,30,202,31,39,31,99,31,202,31,202,30,106,31,120,31,99,31,151,31,185,31,66,31,66,30,55,31,55,30,12,31,237,31,78,31,58,31,54,31,32,31,131,31,149,31,114,31,78,31,55,31,178,31,130,31,176,31,5,31,192,31,192,31,247,31,247,30,180,31,153,31,242,31,151,31,151,30,228,31,164,31,219,31,145,31,39,31,169,31,204,31,35,31,58,31,58,30,222,31,201,31,238,31,183,31,245,31,245,30,30,31,30,30,166,31,120,31,120,30,120,29,120,28,97,31,154,31,12,31,189,31,90,31,90,30,7,31,7,30,7,29,34,31,34,30,151,31,61,31,79,31,33,31,154,31,157,31,137,31,137,30,163,31,182,31,185,31,130,31,63,31,243,31,96,31,36,31,131,31,188,31,169,31,32,31,100,31,100,30,237,31,78,31,71,31,53,31,252,31,252,30,173,31,255,31,52,31,15,31,69,31,95,31,83,31,198,31,97,31,125,31,125,30,97,31,113,31,113,30,113,29,21,31,99,31,120,31,44,31,44,30,19,31,19,30,48,31,9,31,193,31,234,31,141,31,243,31,62,31,243,31,98,31,229,31,193,31,238,31,48,31,196,31,196,30,229,31,205,31,191,31,191,31,121,31,121,30,124,31,124,30,47,31,42,31,67,31,68,31,27,31,209,31,209,30,194,31,58,31,37,31,113,31,195,31,195,30,206,31,106,31,106,30,70,31,160,31,39,31,62,31,200,31,17,31,17,30,147,31,37,31,64,31,38,31,108,31,238,31,238,30,30,31,50,31,50,30,63,31,137,31,246,31,214,31,40,31,68,31,68,30,225,31,143,31,10,31,193,31,31,31,94,31,24,31,217,31,135,31,70,31,223,31,45,31,45,30,237,31,233,31,233,30,62,31,165,31,165,30,68,31,235,31,235,30,67,31,145,31,145,30,248,31,38,31,147,31,147,30,90,31,11,31,62,31,154,31,205,31,224,31,45,31,105,31,105,30,149,31,225,31,147,31,174,31,174,30,174,29,165,31,85,31,85,30,204,31,234,31,234,30,35,31,35,30,35,29,185,31,126,31,126,30,2,31,93,31,48,31,162,31,204,31,147,31,235,31,117,31,117,30,204,31,149,31,189,31,189,30,48,31,164,31,164,30,164,29,83,31,83,30,9,31,96,31,113,31,77,31,70,31,96,31,157,31,35,31,137,31,137,30,219,31,223,31,186,31,78,31,167,31,27,31,139,31,252,31,214,31,214,30,3,31,199,31,159,31,206,31,206,30,227,31,92,31,15,31,180,31,211,31,175,31,1,31,108,31,178,31,205,31,231,31,136,31,118,31,207,31,157,31,156,31,156,30,86,31,196,31,204,31,242,31,154,31,194,31,145,31,221,31,21,31,173,31,171,31,85,31,2,31,69,31,40,31,189,31,224,31,59,31,151,31,249,31,101,31,101,30,101,29,58,31,58,30,253,31,170,31,123,31,246,31,124,31,234,31,234,30,170,31,30,31,178,31,82,31,91,31,27,31,107,31,182,31,182,30,149,31,149,30,2,31,2,30,125,31,131,31,202,31,112,31,216,31,47,31,152,31,249,31,171,31,185,31,176,31,120,31,120,30,204,31,86,31,253,31,188,31,192,31,32,31,32,30,175,31,255,31,133,31,76,31,16,31,16,30,131,31,131,30,131,29,238,31,89,31,248,31,191,31,174,31,26,31,26,30,27,31,26,31,144,31,160,31,160,30,114,31,114,30,87,31,77,31,77,30,146,31,146,30,154,31,6,31,229,31,107,31,241,31,151,31,57,31,247,31,224,31,224,30,224,29,145,31,78,31,78,30,78,29,75,31,157,31,247,31,76,31,6,31,29,31,164,31,235,31,235,31,162,31,186,31,159,31,61,31,61,30,220,31,220,30,144,31,80,31,80,30,80,29,211,31,100,31,106,31,112,31,112,30,112,29,5,31,252,31,138,31,69,31,224,31,96,31,80,31,80,30,45,31,21,31,159,31,159,30,159,29,38,31,18,31,91,31,27,31,165,31,168,31,231,31,52,31,195,31,29,31,29,30,108,31,168,31,168,30,168,29,3,31,184,31,223,31,80,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
