-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 974;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,223,0,185,0,0,0,105,0,22,0,208,0,0,0,170,0,107,0,153,0,200,0,6,0,185,0,147,0,17,0,0,0,106,0,199,0,198,0,39,0,0,0,172,0,31,0,71,0,11,0,237,0,86,0,56,0,31,0,88,0,166,0,0,0,219,0,172,0,0,0,7,0,0,0,0,0,186,0,0,0,112,0,99,0,245,0,30,0,0,0,72,0,106,0,214,0,206,0,221,0,70,0,78,0,246,0,51,0,234,0,182,0,0,0,146,0,55,0,0,0,97,0,241,0,190,0,0,0,0,0,0,0,89,0,0,0,71,0,142,0,180,0,102,0,119,0,147,0,242,0,86,0,183,0,18,0,160,0,161,0,179,0,0,0,14,0,0,0,218,0,134,0,0,0,0,0,99,0,0,0,107,0,200,0,15,0,1,0,155,0,39,0,53,0,72,0,209,0,231,0,232,0,69,0,0,0,202,0,0,0,133,0,23,0,85,0,8,0,153,0,96,0,0,0,21,0,43,0,107,0,0,0,0,0,57,0,251,0,168,0,183,0,181,0,224,0,0,0,131,0,230,0,252,0,137,0,82,0,68,0,132,0,0,0,209,0,32,0,0,0,204,0,84,0,114,0,23,0,161,0,236,0,54,0,11,0,0,0,19,0,0,0,228,0,37,0,147,0,240,0,211,0,0,0,140,0,0,0,68,0,255,0,17,0,0,0,171,0,251,0,237,0,140,0,0,0,150,0,20,0,163,0,0,0,192,0,16,0,0,0,252,0,0,0,117,0,105,0,0,0,247,0,0,0,9,0,31,0,0,0,0,0,20,0,202,0,0,0,40,0,243,0,136,0,252,0,232,0,103,0,22,0,40,0,19,0,252,0,0,0,0,0,129,0,121,0,43,0,139,0,159,0,154,0,197,0,195,0,147,0,52,0,240,0,121,0,218,0,176,0,190,0,32,0,0,0,32,0,101,0,29,0,0,0,14,0,159,0,0,0,84,0,217,0,0,0,119,0,188,0,23,0,0,0,89,0,0,0,233,0,194,0,170,0,155,0,0,0,60,0,161,0,24,0,225,0,79,0,202,0,0,0,205,0,11,0,139,0,0,0,0,0,231,0,196,0,17,0,72,0,0,0,0,0,0,0,186,0,254,0,73,0,101,0,171,0,0,0,0,0,113,0,163,0,198,0,168,0,252,0,0,0,160,0,46,0,143,0,228,0,0,0,113,0,25,0,0,0,37,0,153,0,33,0,0,0,82,0,211,0,56,0,0,0,54,0,0,0,30,0,0,0,0,0,179,0,0,0,0,0,139,0,165,0,127,0,134,0,37,0,50,0,0,0,0,0,0,0,100,0,66,0,42,0,199,0,205,0,0,0,130,0,0,0,55,0,0,0,0,0,116,0,61,0,253,0,218,0,150,0,0,0,108,0,92,0,0,0,69,0,224,0,0,0,244,0,180,0,36,0,195,0,0,0,19,0,176,0,0,0,122,0,91,0,73,0,66,0,250,0,194,0,255,0,74,0,183,0,0,0,6,0,52,0,194,0,120,0,28,0,237,0,161,0,0,0,45,0,11,0,113,0,76,0,125,0,115,0,211,0,152,0,119,0,0,0,247,0,173,0,157,0,253,0,164,0,16,0,152,0,12,0,51,0,3,0,225,0,185,0,211,0,132,0,222,0,225,0,213,0,247,0,168,0,1,0,237,0,0,0,77,0,60,0,13,0,122,0,66,0,52,0,221,0,169,0,237,0,230,0,58,0,210,0,100,0,103,0,177,0,38,0,249,0,139,0,0,0,179,0,140,0,199,0,126,0,168,0,0,0,91,0,250,0,213,0,139,0,209,0,196,0,0,0,182,0,174,0,33,0,13,0,17,0,50,0,242,0,41,0,194,0,71,0,22,0,92,0,110,0,82,0,0,0,43,0,108,0,0,0,218,0,222,0,190,0,0,0,170,0,0,0,29,0,15,0,162,0,82,0,126,0,222,0,95,0,126,0,26,0,166,0,62,0,0,0,174,0,225,0,207,0,0,0,202,0,236,0,59,0,134,0,0,0,0,0,0,0,0,0,137,0,50,0,0,0,167,0,0,0,248,0,44,0,0,0,188,0,161,0,143,0,243,0,232,0,0,0,0,0,151,0,174,0,20,0,151,0,0,0,0,0,209,0,202,0,252,0,0,0,92,0,183,0,0,0,119,0,164,0,204,0,111,0,239,0,190,0,0,0,139,0,239,0,215,0,0,0,33,0,222,0,181,0,214,0,0,0,56,0,0,0,128,0,203,0,152,0,13,0,176,0,243,0,155,0,111,0,0,0,0,0,239,0,0,0,210,0,65,0,234,0,202,0,0,0,165,0,1,0,177,0,2,0,141,0,191,0,102,0,242,0,56,0,35,0,70,0,111,0,239,0,145,0,40,0,188,0,5,0,151,0,196,0,0,0,16,0,2,0,86,0,0,0,64,0,186,0,166,0,0,0,239,0,254,0,23,0,116,0,168,0,183,0,12,0,28,0,128,0,209,0,17,0,200,0,150,0,126,0,238,0,236,0,105,0,166,0,207,0,61,0,212,0,125,0,0,0,124,0,14,0,9,0,52,0,28,0,138,0,0,0,33,0,69,0,0,0,30,0,194,0,79,0,248,0,0,0,46,0,119,0,184,0,84,0,78,0,186,0,32,0,109,0,220,0,207,0,25,0,0,0,253,0,126,0,216,0,45,0,0,0,211,0,224,0,0,0,230,0,193,0,6,0,11,0,244,0,186,0,235,0,229,0,244,0,121,0,0,0,137,0,159,0,76,0,91,0,25,0,0,0,27,0,42,0,52,0,113,0,0,0,1,0,61,0,187,0,107,0,152,0,102,0,222,0,38,0,81,0,184,0,0,0,0,0,204,0,41,0,0,0,0,0,49,0,122,0,0,0,216,0,5,0,180,0,241,0,140,0,82,0,70,0,0,0,0,0,4,0,80,0,43,0,199,0,13,0,37,0,0,0,236,0,22,0,15,0,178,0,0,0,240,0,112,0,0,0,245,0,220,0,201,0,50,0,66,0,0,0,59,0,0,0,13,0,0,0,175,0,23,0,12,0,183,0,41,0,67,0,236,0,37,0,66,0,5,0,48,0,48,0,168,0,34,0,111,0,0,0,144,0,0,0,3,0,78,0,64,0,190,0,35,0,71,0,143,0,209,0,116,0,226,0,231,0,199,0,107,0,141,0,155,0,170,0,125,0,0,0,77,0,251,0,110,0,11,0,95,0,23,0,11,0,0,0,166,0,234,0,45,0,43,0,5,0,0,0,44,0,27,0,220,0,217,0,65,0,0,0,243,0,226,0,118,0,85,0,0,0,111,0,207,0,47,0,60,0,208,0,128,0,0,0,2,0,73,0,8,0,96,0,239,0,155,0,0,0,10,0,180,0,69,0,119,0,195,0,140,0,69,0,78,0,81,0,146,0,62,0,83,0,0,0,0,0,229,0,174,0,160,0,197,0,194,0,30,0,68,0,1,0,0,0,167,0,0,0,210,0,0,0,64,0,86,0,0,0,198,0,0,0,206,0,181,0,91,0,58,0,0,0,74,0,93,0,30,0,83,0,197,0,224,0,115,0,133,0,116,0,153,0,234,0,19,0,236,0,0,0,8,0,81,0,195,0,130,0,26,0,16,0,81,0,0,0,130,0,50,0,124,0,0,0,150,0,139,0,126,0,92,0,3,0,209,0,173,0,225,0,60,0,58,0,0,0,46,0,0,0,61,0,0,0,173,0,161,0,0,0,0,0,18,0,0,0,57,0,103,0,150,0,193,0,167,0,0,0,53,0,239,0,0,0,104,0,179,0,148,0,220,0,66,0,254,0,0,0,5,0,200,0,199,0,0,0,221,0,248,0,0,0,0,0,60,0,0,0,0,0,149,0,102,0,171,0,86,0,118,0,54,0,0,0,124,0,186,0,49,0,227,0,0,0,222,0,7,0,0,0,67,0,74,0,146,0,153,0,179,0,27,0,46,0,131,0,110,0,0,0,0,0,232,0,165,0,33,0,0,0,15,0,6,0,0,0,0,0,91,0,0,0,0,0,0,0,108,0,18,0,245,0,0,0,24,0,215,0,220,0,233,0,44,0,201,0,16,0,0,0,198,0,81,0,69,0,28,0,22,0,170,0,0,0,131,0,6,0,0,0,241,0,101,0,89,0,1,0,201,0,204,0,253,0,152,0,0,0,186,0,142,0,5,0,166,0,0,0,0,0,202,0,74,0,0,0,69,0,178,0,24,0,185,0,201,0,0,0,139,0,0,0,0,0,0,0,215,0,48,0,243,0,215,0,168,0,109,0,5,0,23,0,229,0,239,0,172,0,174,0,0,0,130,0,187,0);
signal scenario_full  : scenario_type := (105,31,223,31,185,31,185,30,105,31,22,31,208,31,208,30,170,31,107,31,153,31,200,31,6,31,185,31,147,31,17,31,17,30,106,31,199,31,198,31,39,31,39,30,172,31,31,31,71,31,11,31,237,31,86,31,56,31,31,31,88,31,166,31,166,30,219,31,172,31,172,30,7,31,7,30,7,29,186,31,186,30,112,31,99,31,245,31,30,31,30,30,72,31,106,31,214,31,206,31,221,31,70,31,78,31,246,31,51,31,234,31,182,31,182,30,146,31,55,31,55,30,97,31,241,31,190,31,190,30,190,29,190,28,89,31,89,30,71,31,142,31,180,31,102,31,119,31,147,31,242,31,86,31,183,31,18,31,160,31,161,31,179,31,179,30,14,31,14,30,218,31,134,31,134,30,134,29,99,31,99,30,107,31,200,31,15,31,1,31,155,31,39,31,53,31,72,31,209,31,231,31,232,31,69,31,69,30,202,31,202,30,133,31,23,31,85,31,8,31,153,31,96,31,96,30,21,31,43,31,107,31,107,30,107,29,57,31,251,31,168,31,183,31,181,31,224,31,224,30,131,31,230,31,252,31,137,31,82,31,68,31,132,31,132,30,209,31,32,31,32,30,204,31,84,31,114,31,23,31,161,31,236,31,54,31,11,31,11,30,19,31,19,30,228,31,37,31,147,31,240,31,211,31,211,30,140,31,140,30,68,31,255,31,17,31,17,30,171,31,251,31,237,31,140,31,140,30,150,31,20,31,163,31,163,30,192,31,16,31,16,30,252,31,252,30,117,31,105,31,105,30,247,31,247,30,9,31,31,31,31,30,31,29,20,31,202,31,202,30,40,31,243,31,136,31,252,31,232,31,103,31,22,31,40,31,19,31,252,31,252,30,252,29,129,31,121,31,43,31,139,31,159,31,154,31,197,31,195,31,147,31,52,31,240,31,121,31,218,31,176,31,190,31,32,31,32,30,32,31,101,31,29,31,29,30,14,31,159,31,159,30,84,31,217,31,217,30,119,31,188,31,23,31,23,30,89,31,89,30,233,31,194,31,170,31,155,31,155,30,60,31,161,31,24,31,225,31,79,31,202,31,202,30,205,31,11,31,139,31,139,30,139,29,231,31,196,31,17,31,72,31,72,30,72,29,72,28,186,31,254,31,73,31,101,31,171,31,171,30,171,29,113,31,163,31,198,31,168,31,252,31,252,30,160,31,46,31,143,31,228,31,228,30,113,31,25,31,25,30,37,31,153,31,33,31,33,30,82,31,211,31,56,31,56,30,54,31,54,30,30,31,30,30,30,29,179,31,179,30,179,29,139,31,165,31,127,31,134,31,37,31,50,31,50,30,50,29,50,28,100,31,66,31,42,31,199,31,205,31,205,30,130,31,130,30,55,31,55,30,55,29,116,31,61,31,253,31,218,31,150,31,150,30,108,31,92,31,92,30,69,31,224,31,224,30,244,31,180,31,36,31,195,31,195,30,19,31,176,31,176,30,122,31,91,31,73,31,66,31,250,31,194,31,255,31,74,31,183,31,183,30,6,31,52,31,194,31,120,31,28,31,237,31,161,31,161,30,45,31,11,31,113,31,76,31,125,31,115,31,211,31,152,31,119,31,119,30,247,31,173,31,157,31,253,31,164,31,16,31,152,31,12,31,51,31,3,31,225,31,185,31,211,31,132,31,222,31,225,31,213,31,247,31,168,31,1,31,237,31,237,30,77,31,60,31,13,31,122,31,66,31,52,31,221,31,169,31,237,31,230,31,58,31,210,31,100,31,103,31,177,31,38,31,249,31,139,31,139,30,179,31,140,31,199,31,126,31,168,31,168,30,91,31,250,31,213,31,139,31,209,31,196,31,196,30,182,31,174,31,33,31,13,31,17,31,50,31,242,31,41,31,194,31,71,31,22,31,92,31,110,31,82,31,82,30,43,31,108,31,108,30,218,31,222,31,190,31,190,30,170,31,170,30,29,31,15,31,162,31,82,31,126,31,222,31,95,31,126,31,26,31,166,31,62,31,62,30,174,31,225,31,207,31,207,30,202,31,236,31,59,31,134,31,134,30,134,29,134,28,134,27,137,31,50,31,50,30,167,31,167,30,248,31,44,31,44,30,188,31,161,31,143,31,243,31,232,31,232,30,232,29,151,31,174,31,20,31,151,31,151,30,151,29,209,31,202,31,252,31,252,30,92,31,183,31,183,30,119,31,164,31,204,31,111,31,239,31,190,31,190,30,139,31,239,31,215,31,215,30,33,31,222,31,181,31,214,31,214,30,56,31,56,30,128,31,203,31,152,31,13,31,176,31,243,31,155,31,111,31,111,30,111,29,239,31,239,30,210,31,65,31,234,31,202,31,202,30,165,31,1,31,177,31,2,31,141,31,191,31,102,31,242,31,56,31,35,31,70,31,111,31,239,31,145,31,40,31,188,31,5,31,151,31,196,31,196,30,16,31,2,31,86,31,86,30,64,31,186,31,166,31,166,30,239,31,254,31,23,31,116,31,168,31,183,31,12,31,28,31,128,31,209,31,17,31,200,31,150,31,126,31,238,31,236,31,105,31,166,31,207,31,61,31,212,31,125,31,125,30,124,31,14,31,9,31,52,31,28,31,138,31,138,30,33,31,69,31,69,30,30,31,194,31,79,31,248,31,248,30,46,31,119,31,184,31,84,31,78,31,186,31,32,31,109,31,220,31,207,31,25,31,25,30,253,31,126,31,216,31,45,31,45,30,211,31,224,31,224,30,230,31,193,31,6,31,11,31,244,31,186,31,235,31,229,31,244,31,121,31,121,30,137,31,159,31,76,31,91,31,25,31,25,30,27,31,42,31,52,31,113,31,113,30,1,31,61,31,187,31,107,31,152,31,102,31,222,31,38,31,81,31,184,31,184,30,184,29,204,31,41,31,41,30,41,29,49,31,122,31,122,30,216,31,5,31,180,31,241,31,140,31,82,31,70,31,70,30,70,29,4,31,80,31,43,31,199,31,13,31,37,31,37,30,236,31,22,31,15,31,178,31,178,30,240,31,112,31,112,30,245,31,220,31,201,31,50,31,66,31,66,30,59,31,59,30,13,31,13,30,175,31,23,31,12,31,183,31,41,31,67,31,236,31,37,31,66,31,5,31,48,31,48,31,168,31,34,31,111,31,111,30,144,31,144,30,3,31,78,31,64,31,190,31,35,31,71,31,143,31,209,31,116,31,226,31,231,31,199,31,107,31,141,31,155,31,170,31,125,31,125,30,77,31,251,31,110,31,11,31,95,31,23,31,11,31,11,30,166,31,234,31,45,31,43,31,5,31,5,30,44,31,27,31,220,31,217,31,65,31,65,30,243,31,226,31,118,31,85,31,85,30,111,31,207,31,47,31,60,31,208,31,128,31,128,30,2,31,73,31,8,31,96,31,239,31,155,31,155,30,10,31,180,31,69,31,119,31,195,31,140,31,69,31,78,31,81,31,146,31,62,31,83,31,83,30,83,29,229,31,174,31,160,31,197,31,194,31,30,31,68,31,1,31,1,30,167,31,167,30,210,31,210,30,64,31,86,31,86,30,198,31,198,30,206,31,181,31,91,31,58,31,58,30,74,31,93,31,30,31,83,31,197,31,224,31,115,31,133,31,116,31,153,31,234,31,19,31,236,31,236,30,8,31,81,31,195,31,130,31,26,31,16,31,81,31,81,30,130,31,50,31,124,31,124,30,150,31,139,31,126,31,92,31,3,31,209,31,173,31,225,31,60,31,58,31,58,30,46,31,46,30,61,31,61,30,173,31,161,31,161,30,161,29,18,31,18,30,57,31,103,31,150,31,193,31,167,31,167,30,53,31,239,31,239,30,104,31,179,31,148,31,220,31,66,31,254,31,254,30,5,31,200,31,199,31,199,30,221,31,248,31,248,30,248,29,60,31,60,30,60,29,149,31,102,31,171,31,86,31,118,31,54,31,54,30,124,31,186,31,49,31,227,31,227,30,222,31,7,31,7,30,67,31,74,31,146,31,153,31,179,31,27,31,46,31,131,31,110,31,110,30,110,29,232,31,165,31,33,31,33,30,15,31,6,31,6,30,6,29,91,31,91,30,91,29,91,28,108,31,18,31,245,31,245,30,24,31,215,31,220,31,233,31,44,31,201,31,16,31,16,30,198,31,81,31,69,31,28,31,22,31,170,31,170,30,131,31,6,31,6,30,241,31,101,31,89,31,1,31,201,31,204,31,253,31,152,31,152,30,186,31,142,31,5,31,166,31,166,30,166,29,202,31,74,31,74,30,69,31,178,31,24,31,185,31,201,31,201,30,139,31,139,30,139,29,139,28,215,31,48,31,243,31,215,31,168,31,109,31,5,31,23,31,229,31,239,31,172,31,174,31,174,30,130,31,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
