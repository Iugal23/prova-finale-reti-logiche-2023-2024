-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 740;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,113,0,135,0,91,0,120,0,231,0,0,0,22,0,0,0,82,0,22,0,210,0,41,0,14,0,62,0,158,0,0,0,115,0,2,0,248,0,87,0,0,0,230,0,71,0,29,0,172,0,172,0,117,0,0,0,161,0,0,0,121,0,124,0,87,0,0,0,167,0,152,0,92,0,55,0,0,0,0,0,7,0,193,0,231,0,0,0,251,0,0,0,236,0,176,0,63,0,221,0,122,0,53,0,245,0,0,0,226,0,184,0,0,0,0,0,146,0,94,0,0,0,31,0,243,0,22,0,222,0,0,0,228,0,0,0,138,0,90,0,174,0,103,0,56,0,0,0,0,0,85,0,249,0,55,0,126,0,250,0,174,0,6,0,162,0,27,0,222,0,9,0,79,0,51,0,56,0,10,0,94,0,0,0,21,0,0,0,255,0,37,0,129,0,88,0,182,0,194,0,222,0,39,0,171,0,196,0,31,0,116,0,19,0,0,0,197,0,0,0,0,0,83,0,113,0,26,0,225,0,0,0,125,0,175,0,210,0,45,0,64,0,0,0,251,0,11,0,207,0,76,0,76,0,167,0,0,0,173,0,201,0,233,0,0,0,0,0,91,0,49,0,43,0,249,0,0,0,23,0,0,0,150,0,29,0,249,0,0,0,0,0,134,0,75,0,240,0,139,0,118,0,205,0,0,0,4,0,0,0,0,0,0,0,232,0,0,0,194,0,153,0,178,0,192,0,0,0,0,0,0,0,148,0,190,0,103,0,183,0,127,0,0,0,3,0,51,0,234,0,0,0,17,0,5,0,162,0,122,0,36,0,130,0,153,0,218,0,46,0,0,0,213,0,177,0,0,0,0,0,137,0,212,0,144,0,249,0,59,0,80,0,220,0,0,0,172,0,169,0,157,0,117,0,159,0,13,0,0,0,228,0,213,0,66,0,163,0,174,0,0,0,180,0,60,0,44,0,126,0,0,0,35,0,183,0,0,0,186,0,24,0,89,0,32,0,6,0,110,0,0,0,217,0,0,0,0,0,0,0,134,0,156,0,252,0,86,0,142,0,137,0,173,0,180,0,119,0,127,0,99,0,0,0,251,0,79,0,89,0,48,0,217,0,38,0,52,0,229,0,0,0,69,0,16,0,78,0,51,0,22,0,50,0,138,0,0,0,0,0,0,0,73,0,0,0,51,0,0,0,241,0,20,0,23,0,73,0,40,0,21,0,234,0,196,0,214,0,173,0,162,0,4,0,131,0,34,0,66,0,0,0,246,0,229,0,0,0,239,0,0,0,93,0,218,0,86,0,254,0,0,0,104,0,252,0,0,0,102,0,48,0,128,0,11,0,243,0,0,0,109,0,150,0,102,0,75,0,0,0,125,0,0,0,103,0,76,0,125,0,210,0,221,0,0,0,0,0,146,0,254,0,80,0,57,0,100,0,0,0,237,0,0,0,81,0,226,0,198,0,0,0,157,0,32,0,162,0,12,0,0,0,166,0,47,0,97,0,0,0,1,0,151,0,8,0,69,0,223,0,74,0,0,0,122,0,103,0,217,0,146,0,10,0,75,0,126,0,0,0,21,0,195,0,89,0,185,0,134,0,7,0,158,0,209,0,132,0,21,0,14,0,53,0,81,0,68,0,174,0,0,0,129,0,43,0,72,0,0,0,55,0,41,0,14,0,248,0,0,0,162,0,180,0,228,0,0,0,13,0,155,0,202,0,87,0,3,0,40,0,0,0,0,0,235,0,47,0,76,0,236,0,77,0,159,0,0,0,112,0,248,0,0,0,192,0,0,0,0,0,97,0,195,0,202,0,0,0,55,0,64,0,0,0,0,0,197,0,206,0,203,0,232,0,71,0,0,0,0,0,167,0,235,0,149,0,110,0,207,0,46,0,0,0,96,0,34,0,175,0,186,0,40,0,118,0,0,0,112,0,11,0,0,0,230,0,20,0,168,0,212,0,158,0,8,0,46,0,220,0,0,0,37,0,92,0,0,0,0,0,168,0,156,0,128,0,4,0,124,0,58,0,0,0,28,0,150,0,82,0,0,0,40,0,54,0,115,0,89,0,174,0,0,0,35,0,132,0,0,0,76,0,181,0,169,0,126,0,170,0,0,0,0,0,202,0,46,0,250,0,0,0,0,0,38,0,254,0,52,0,0,0,96,0,151,0,103,0,0,0,58,0,244,0,0,0,0,0,188,0,0,0,239,0,187,0,0,0,112,0,192,0,190,0,61,0,0,0,240,0,104,0,57,0,0,0,4,0,118,0,7,0,173,0,160,0,0,0,210,0,0,0,77,0,45,0,0,0,29,0,156,0,0,0,196,0,125,0,182,0,232,0,121,0,0,0,129,0,33,0,202,0,2,0,142,0,126,0,14,0,145,0,60,0,116,0,131,0,90,0,63,0,55,0,130,0,95,0,23,0,82,0,149,0,166,0,34,0,0,0,30,0,214,0,0,0,143,0,20,0,213,0,163,0,156,0,119,0,47,0,114,0,187,0,0,0,80,0,103,0,203,0,226,0,162,0,0,0,240,0,0,0,0,0,141,0,102,0,0,0,0,0,60,0,0,0,126,0,0,0,126,0,120,0,244,0,8,0,3,0,207,0,108,0,0,0,127,0,9,0,0,0,208,0,161,0,148,0,11,0,0,0,184,0,126,0,193,0,0,0,0,0,181,0,187,0,28,0,113,0,173,0,210,0,92,0,156,0,0,0,102,0,62,0,120,0,78,0,44,0,0,0,0,0,185,0,0,0,185,0,144,0,251,0,117,0,0,0,191,0,15,0,248,0,67,0,225,0,65,0,22,0,70,0,207,0,206,0,199,0,92,0,75,0,175,0,222,0,42,0,218,0,82,0,241,0,40,0,17,0,51,0,180,0,120,0,174,0,73,0,131,0,249,0,249,0,192,0,219,0,193,0,239,0,25,0,0,0,83,0,180,0,153,0,206,0,0,0,219,0,39,0,52,0,0,0,0,0,177,0,58,0,0,0,62,0,22,0,0,0,170,0,0,0,150,0,166,0,12,0,244,0,25,0,0,0,0,0,13,0,250,0,205,0,34,0,237,0,145,0,197,0,63,0,0,0,241,0,71,0,91,0,65,0,185,0,198,0,0,0,234,0,139,0,0,0,45,0,143,0,233,0,198,0,82,0,79,0,168,0,0,0,6,0,0,0,68,0,39,0,0,0,175,0,185,0,0,0,231,0,177,0,0,0,98,0,239,0,0,0,182,0,0,0,88,0,138,0,0,0,107,0,63,0,201,0,0,0,162,0,0,0,249,0,143,0,110,0,178,0,52,0,140,0,196,0,208,0);
signal scenario_full  : scenario_type := (0,0,113,31,135,31,91,31,120,31,231,31,231,30,22,31,22,30,82,31,22,31,210,31,41,31,14,31,62,31,158,31,158,30,115,31,2,31,248,31,87,31,87,30,230,31,71,31,29,31,172,31,172,31,117,31,117,30,161,31,161,30,121,31,124,31,87,31,87,30,167,31,152,31,92,31,55,31,55,30,55,29,7,31,193,31,231,31,231,30,251,31,251,30,236,31,176,31,63,31,221,31,122,31,53,31,245,31,245,30,226,31,184,31,184,30,184,29,146,31,94,31,94,30,31,31,243,31,22,31,222,31,222,30,228,31,228,30,138,31,90,31,174,31,103,31,56,31,56,30,56,29,85,31,249,31,55,31,126,31,250,31,174,31,6,31,162,31,27,31,222,31,9,31,79,31,51,31,56,31,10,31,94,31,94,30,21,31,21,30,255,31,37,31,129,31,88,31,182,31,194,31,222,31,39,31,171,31,196,31,31,31,116,31,19,31,19,30,197,31,197,30,197,29,83,31,113,31,26,31,225,31,225,30,125,31,175,31,210,31,45,31,64,31,64,30,251,31,11,31,207,31,76,31,76,31,167,31,167,30,173,31,201,31,233,31,233,30,233,29,91,31,49,31,43,31,249,31,249,30,23,31,23,30,150,31,29,31,249,31,249,30,249,29,134,31,75,31,240,31,139,31,118,31,205,31,205,30,4,31,4,30,4,29,4,28,232,31,232,30,194,31,153,31,178,31,192,31,192,30,192,29,192,28,148,31,190,31,103,31,183,31,127,31,127,30,3,31,51,31,234,31,234,30,17,31,5,31,162,31,122,31,36,31,130,31,153,31,218,31,46,31,46,30,213,31,177,31,177,30,177,29,137,31,212,31,144,31,249,31,59,31,80,31,220,31,220,30,172,31,169,31,157,31,117,31,159,31,13,31,13,30,228,31,213,31,66,31,163,31,174,31,174,30,180,31,60,31,44,31,126,31,126,30,35,31,183,31,183,30,186,31,24,31,89,31,32,31,6,31,110,31,110,30,217,31,217,30,217,29,217,28,134,31,156,31,252,31,86,31,142,31,137,31,173,31,180,31,119,31,127,31,99,31,99,30,251,31,79,31,89,31,48,31,217,31,38,31,52,31,229,31,229,30,69,31,16,31,78,31,51,31,22,31,50,31,138,31,138,30,138,29,138,28,73,31,73,30,51,31,51,30,241,31,20,31,23,31,73,31,40,31,21,31,234,31,196,31,214,31,173,31,162,31,4,31,131,31,34,31,66,31,66,30,246,31,229,31,229,30,239,31,239,30,93,31,218,31,86,31,254,31,254,30,104,31,252,31,252,30,102,31,48,31,128,31,11,31,243,31,243,30,109,31,150,31,102,31,75,31,75,30,125,31,125,30,103,31,76,31,125,31,210,31,221,31,221,30,221,29,146,31,254,31,80,31,57,31,100,31,100,30,237,31,237,30,81,31,226,31,198,31,198,30,157,31,32,31,162,31,12,31,12,30,166,31,47,31,97,31,97,30,1,31,151,31,8,31,69,31,223,31,74,31,74,30,122,31,103,31,217,31,146,31,10,31,75,31,126,31,126,30,21,31,195,31,89,31,185,31,134,31,7,31,158,31,209,31,132,31,21,31,14,31,53,31,81,31,68,31,174,31,174,30,129,31,43,31,72,31,72,30,55,31,41,31,14,31,248,31,248,30,162,31,180,31,228,31,228,30,13,31,155,31,202,31,87,31,3,31,40,31,40,30,40,29,235,31,47,31,76,31,236,31,77,31,159,31,159,30,112,31,248,31,248,30,192,31,192,30,192,29,97,31,195,31,202,31,202,30,55,31,64,31,64,30,64,29,197,31,206,31,203,31,232,31,71,31,71,30,71,29,167,31,235,31,149,31,110,31,207,31,46,31,46,30,96,31,34,31,175,31,186,31,40,31,118,31,118,30,112,31,11,31,11,30,230,31,20,31,168,31,212,31,158,31,8,31,46,31,220,31,220,30,37,31,92,31,92,30,92,29,168,31,156,31,128,31,4,31,124,31,58,31,58,30,28,31,150,31,82,31,82,30,40,31,54,31,115,31,89,31,174,31,174,30,35,31,132,31,132,30,76,31,181,31,169,31,126,31,170,31,170,30,170,29,202,31,46,31,250,31,250,30,250,29,38,31,254,31,52,31,52,30,96,31,151,31,103,31,103,30,58,31,244,31,244,30,244,29,188,31,188,30,239,31,187,31,187,30,112,31,192,31,190,31,61,31,61,30,240,31,104,31,57,31,57,30,4,31,118,31,7,31,173,31,160,31,160,30,210,31,210,30,77,31,45,31,45,30,29,31,156,31,156,30,196,31,125,31,182,31,232,31,121,31,121,30,129,31,33,31,202,31,2,31,142,31,126,31,14,31,145,31,60,31,116,31,131,31,90,31,63,31,55,31,130,31,95,31,23,31,82,31,149,31,166,31,34,31,34,30,30,31,214,31,214,30,143,31,20,31,213,31,163,31,156,31,119,31,47,31,114,31,187,31,187,30,80,31,103,31,203,31,226,31,162,31,162,30,240,31,240,30,240,29,141,31,102,31,102,30,102,29,60,31,60,30,126,31,126,30,126,31,120,31,244,31,8,31,3,31,207,31,108,31,108,30,127,31,9,31,9,30,208,31,161,31,148,31,11,31,11,30,184,31,126,31,193,31,193,30,193,29,181,31,187,31,28,31,113,31,173,31,210,31,92,31,156,31,156,30,102,31,62,31,120,31,78,31,44,31,44,30,44,29,185,31,185,30,185,31,144,31,251,31,117,31,117,30,191,31,15,31,248,31,67,31,225,31,65,31,22,31,70,31,207,31,206,31,199,31,92,31,75,31,175,31,222,31,42,31,218,31,82,31,241,31,40,31,17,31,51,31,180,31,120,31,174,31,73,31,131,31,249,31,249,31,192,31,219,31,193,31,239,31,25,31,25,30,83,31,180,31,153,31,206,31,206,30,219,31,39,31,52,31,52,30,52,29,177,31,58,31,58,30,62,31,22,31,22,30,170,31,170,30,150,31,166,31,12,31,244,31,25,31,25,30,25,29,13,31,250,31,205,31,34,31,237,31,145,31,197,31,63,31,63,30,241,31,71,31,91,31,65,31,185,31,198,31,198,30,234,31,139,31,139,30,45,31,143,31,233,31,198,31,82,31,79,31,168,31,168,30,6,31,6,30,68,31,39,31,39,30,175,31,185,31,185,30,231,31,177,31,177,30,98,31,239,31,239,30,182,31,182,30,88,31,138,31,138,30,107,31,63,31,201,31,201,30,162,31,162,30,249,31,143,31,110,31,178,31,52,31,140,31,196,31,208,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
