-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 333;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (183,0,163,0,0,0,0,0,58,0,0,0,43,0,7,0,211,0,142,0,52,0,140,0,48,0,174,0,0,0,177,0,0,0,0,0,138,0,226,0,94,0,121,0,211,0,5,0,0,0,52,0,163,0,229,0,165,0,189,0,145,0,103,0,69,0,0,0,137,0,246,0,190,0,7,0,0,0,0,0,192,0,80,0,108,0,197,0,155,0,84,0,0,0,117,0,74,0,0,0,120,0,45,0,180,0,0,0,15,0,224,0,47,0,203,0,0,0,131,0,44,0,0,0,176,0,237,0,105,0,126,0,149,0,35,0,211,0,231,0,171,0,138,0,93,0,0,0,42,0,0,0,216,0,19,0,97,0,220,0,225,0,67,0,98,0,228,0,193,0,92,0,32,0,249,0,14,0,42,0,75,0,0,0,203,0,0,0,0,0,8,0,0,0,44,0,236,0,156,0,72,0,67,0,194,0,0,0,252,0,77,0,42,0,74,0,57,0,43,0,4,0,23,0,80,0,203,0,82,0,159,0,62,0,123,0,188,0,237,0,59,0,0,0,148,0,140,0,78,0,157,0,32,0,242,0,136,0,100,0,0,0,124,0,0,0,42,0,96,0,128,0,78,0,187,0,116,0,38,0,148,0,0,0,0,0,221,0,211,0,237,0,39,0,188,0,0,0,232,0,0,0,95,0,0,0,39,0,222,0,0,0,101,0,249,0,21,0,125,0,0,0,92,0,71,0,207,0,19,0,200,0,224,0,0,0,0,0,74,0,0,0,26,0,212,0,63,0,174,0,194,0,187,0,164,0,81,0,0,0,239,0,0,0,0,0,0,0,0,0,29,0,189,0,12,0,0,0,197,0,222,0,110,0,0,0,65,0,174,0,60,0,44,0,221,0,234,0,182,0,0,0,115,0,0,0,182,0,47,0,0,0,0,0,0,0,218,0,196,0,0,0,187,0,85,0,211,0,1,0,169,0,118,0,114,0,19,0,28,0,0,0,10,0,245,0,224,0,91,0,249,0,58,0,121,0,0,0,74,0,0,0,25,0,0,0,80,0,0,0,41,0,0,0,234,0,0,0,97,0,225,0,92,0,25,0,167,0,4,0,139,0,38,0,31,0,0,0,0,0,182,0,0,0,0,0,163,0,27,0,8,0,0,0,0,0,1,0,231,0,169,0,220,0,77,0,125,0,0,0,0,0,0,0,90,0,0,0,108,0,0,0,14,0,105,0,91,0,76,0,7,0,0,0,41,0,83,0,0,0,176,0,110,0,3,0,37,0,0,0,0,0,113,0,0,0,53,0,205,0,0,0,203,0,0,0,0,0,98,0,49,0,18,0,242,0,0,0,0,0,15,0,54,0,58,0,5,0,72,0,81,0,237,0,223,0,46,0,173,0,221,0,0,0,98,0,97,0,0,0,124,0,114,0,199,0,176,0,0,0,0,0,0,0,46,0,54,0,224,0,37,0,0,0,83,0,0,0,143,0,217,0,73,0,163,0);
signal scenario_full  : scenario_type := (183,31,163,31,163,30,163,29,58,31,58,30,43,31,7,31,211,31,142,31,52,31,140,31,48,31,174,31,174,30,177,31,177,30,177,29,138,31,226,31,94,31,121,31,211,31,5,31,5,30,52,31,163,31,229,31,165,31,189,31,145,31,103,31,69,31,69,30,137,31,246,31,190,31,7,31,7,30,7,29,192,31,80,31,108,31,197,31,155,31,84,31,84,30,117,31,74,31,74,30,120,31,45,31,180,31,180,30,15,31,224,31,47,31,203,31,203,30,131,31,44,31,44,30,176,31,237,31,105,31,126,31,149,31,35,31,211,31,231,31,171,31,138,31,93,31,93,30,42,31,42,30,216,31,19,31,97,31,220,31,225,31,67,31,98,31,228,31,193,31,92,31,32,31,249,31,14,31,42,31,75,31,75,30,203,31,203,30,203,29,8,31,8,30,44,31,236,31,156,31,72,31,67,31,194,31,194,30,252,31,77,31,42,31,74,31,57,31,43,31,4,31,23,31,80,31,203,31,82,31,159,31,62,31,123,31,188,31,237,31,59,31,59,30,148,31,140,31,78,31,157,31,32,31,242,31,136,31,100,31,100,30,124,31,124,30,42,31,96,31,128,31,78,31,187,31,116,31,38,31,148,31,148,30,148,29,221,31,211,31,237,31,39,31,188,31,188,30,232,31,232,30,95,31,95,30,39,31,222,31,222,30,101,31,249,31,21,31,125,31,125,30,92,31,71,31,207,31,19,31,200,31,224,31,224,30,224,29,74,31,74,30,26,31,212,31,63,31,174,31,194,31,187,31,164,31,81,31,81,30,239,31,239,30,239,29,239,28,239,27,29,31,189,31,12,31,12,30,197,31,222,31,110,31,110,30,65,31,174,31,60,31,44,31,221,31,234,31,182,31,182,30,115,31,115,30,182,31,47,31,47,30,47,29,47,28,218,31,196,31,196,30,187,31,85,31,211,31,1,31,169,31,118,31,114,31,19,31,28,31,28,30,10,31,245,31,224,31,91,31,249,31,58,31,121,31,121,30,74,31,74,30,25,31,25,30,80,31,80,30,41,31,41,30,234,31,234,30,97,31,225,31,92,31,25,31,167,31,4,31,139,31,38,31,31,31,31,30,31,29,182,31,182,30,182,29,163,31,27,31,8,31,8,30,8,29,1,31,231,31,169,31,220,31,77,31,125,31,125,30,125,29,125,28,90,31,90,30,108,31,108,30,14,31,105,31,91,31,76,31,7,31,7,30,41,31,83,31,83,30,176,31,110,31,3,31,37,31,37,30,37,29,113,31,113,30,53,31,205,31,205,30,203,31,203,30,203,29,98,31,49,31,18,31,242,31,242,30,242,29,15,31,54,31,58,31,5,31,72,31,81,31,237,31,223,31,46,31,173,31,221,31,221,30,98,31,97,31,97,30,124,31,114,31,199,31,176,31,176,30,176,29,176,28,46,31,54,31,224,31,37,31,37,30,83,31,83,30,143,31,217,31,73,31,163,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
