-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 539;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,53,0,37,0,159,0,180,0,141,0,127,0,75,0,241,0,25,0,120,0,240,0,204,0,250,0,0,0,0,0,157,0,228,0,91,0,2,0,176,0,133,0,44,0,181,0,16,0,40,0,254,0,0,0,0,0,39,0,253,0,0,0,250,0,49,0,64,0,0,0,251,0,78,0,0,0,156,0,181,0,135,0,2,0,194,0,89,0,55,0,0,0,196,0,150,0,220,0,158,0,201,0,64,0,69,0,66,0,126,0,62,0,229,0,0,0,0,0,237,0,44,0,167,0,144,0,206,0,161,0,150,0,0,0,204,0,154,0,41,0,215,0,189,0,186,0,102,0,210,0,229,0,51,0,29,0,114,0,0,0,160,0,0,0,21,0,54,0,0,0,83,0,0,0,165,0,211,0,157,0,0,0,252,0,235,0,115,0,134,0,196,0,0,0,0,0,124,0,162,0,128,0,0,0,0,0,195,0,130,0,194,0,15,0,86,0,229,0,133,0,188,0,255,0,127,0,180,0,114,0,216,0,16,0,62,0,246,0,0,0,223,0,239,0,166,0,142,0,0,0,215,0,214,0,124,0,147,0,100,0,169,0,60,0,216,0,172,0,0,0,228,0,0,0,212,0,253,0,211,0,236,0,59,0,102,0,0,0,223,0,228,0,0,0,0,0,0,0,247,0,236,0,111,0,77,0,64,0,133,0,152,0,88,0,227,0,164,0,138,0,248,0,13,0,41,0,82,0,0,0,0,0,120,0,0,0,246,0,169,0,177,0,205,0,224,0,63,0,0,0,126,0,145,0,228,0,73,0,32,0,125,0,0,0,227,0,41,0,255,0,0,0,163,0,3,0,108,0,199,0,188,0,0,0,28,0,208,0,12,0,247,0,0,0,0,0,0,0,243,0,219,0,126,0,249,0,0,0,34,0,96,0,33,0,181,0,194,0,214,0,208,0,0,0,195,0,134,0,114,0,235,0,91,0,253,0,228,0,106,0,0,0,132,0,224,0,0,0,43,0,199,0,227,0,91,0,0,0,4,0,226,0,243,0,217,0,0,0,0,0,172,0,80,0,0,0,192,0,0,0,57,0,146,0,220,0,70,0,145,0,160,0,208,0,83,0,164,0,140,0,0,0,236,0,57,0,0,0,63,0,195,0,42,0,114,0,0,0,141,0,86,0,0,0,129,0,166,0,0,0,156,0,4,0,224,0,135,0,181,0,116,0,251,0,134,0,5,0,226,0,15,0,126,0,0,0,206,0,104,0,213,0,192,0,104,0,0,0,0,0,0,0,196,0,22,0,108,0,217,0,211,0,133,0,25,0,0,0,225,0,141,0,229,0,14,0,229,0,217,0,22,0,31,0,226,0,188,0,0,0,245,0,227,0,37,0,208,0,210,0,0,0,17,0,146,0,141,0,172,0,21,0,236,0,0,0,225,0,118,0,199,0,126,0,0,0,0,0,47,0,0,0,0,0,19,0,110,0,0,0,65,0,19,0,98,0,0,0,238,0,35,0,0,0,189,0,168,0,237,0,64,0,38,0,233,0,143,0,170,0,0,0,49,0,2,0,0,0,205,0,70,0,202,0,22,0,93,0,59,0,0,0,74,0,0,0,107,0,88,0,118,0,83,0,37,0,0,0,0,0,2,0,53,0,0,0,0,0,239,0,0,0,1,0,59,0,166,0,55,0,0,0,108,0,27,0,0,0,0,0,222,0,202,0,133,0,124,0,0,0,72,0,81,0,92,0,198,0,53,0,0,0,254,0,0,0,23,0,186,0,189,0,104,0,104,0,87,0,196,0,6,0,135,0,172,0,0,0,74,0,187,0,177,0,0,0,111,0,254,0,199,0,243,0,200,0,218,0,76,0,49,0,5,0,56,0,0,0,0,0,248,0,0,0,0,0,53,0,0,0,77,0,58,0,0,0,34,0,2,0,42,0,151,0,58,0,180,0,222,0,0,0,48,0,142,0,208,0,197,0,219,0,0,0,152,0,0,0,15,0,63,0,40,0,0,0,103,0,190,0,0,0,0,0,74,0,180,0,0,0,0,0,0,0,218,0,179,0,186,0,0,0,155,0,161,0,0,0,137,0,0,0,217,0,237,0,229,0,254,0,52,0,108,0,149,0,0,0,0,0,234,0,0,0,83,0,224,0,88,0,0,0,95,0,46,0,91,0,161,0,0,0,20,0,218,0,0,0,162,0,205,0,124,0,152,0,3,0,102,0,49,0,182,0,0,0,99,0,241,0,191,0,69,0,166,0,0,0,0,0,0,0,40,0,250,0,129,0,126,0,69,0,159,0,105,0,3,0,80,0,45,0,46,0,0,0,0,0,214,0,51,0,38,0,72,0,0,0,19,0,0,0,242,0,167,0,10,0,242,0,217,0,82,0,173,0,20,0,250,0,95,0,119,0,111,0);
signal scenario_full  : scenario_type := (0,0,53,31,37,31,159,31,180,31,141,31,127,31,75,31,241,31,25,31,120,31,240,31,204,31,250,31,250,30,250,29,157,31,228,31,91,31,2,31,176,31,133,31,44,31,181,31,16,31,40,31,254,31,254,30,254,29,39,31,253,31,253,30,250,31,49,31,64,31,64,30,251,31,78,31,78,30,156,31,181,31,135,31,2,31,194,31,89,31,55,31,55,30,196,31,150,31,220,31,158,31,201,31,64,31,69,31,66,31,126,31,62,31,229,31,229,30,229,29,237,31,44,31,167,31,144,31,206,31,161,31,150,31,150,30,204,31,154,31,41,31,215,31,189,31,186,31,102,31,210,31,229,31,51,31,29,31,114,31,114,30,160,31,160,30,21,31,54,31,54,30,83,31,83,30,165,31,211,31,157,31,157,30,252,31,235,31,115,31,134,31,196,31,196,30,196,29,124,31,162,31,128,31,128,30,128,29,195,31,130,31,194,31,15,31,86,31,229,31,133,31,188,31,255,31,127,31,180,31,114,31,216,31,16,31,62,31,246,31,246,30,223,31,239,31,166,31,142,31,142,30,215,31,214,31,124,31,147,31,100,31,169,31,60,31,216,31,172,31,172,30,228,31,228,30,212,31,253,31,211,31,236,31,59,31,102,31,102,30,223,31,228,31,228,30,228,29,228,28,247,31,236,31,111,31,77,31,64,31,133,31,152,31,88,31,227,31,164,31,138,31,248,31,13,31,41,31,82,31,82,30,82,29,120,31,120,30,246,31,169,31,177,31,205,31,224,31,63,31,63,30,126,31,145,31,228,31,73,31,32,31,125,31,125,30,227,31,41,31,255,31,255,30,163,31,3,31,108,31,199,31,188,31,188,30,28,31,208,31,12,31,247,31,247,30,247,29,247,28,243,31,219,31,126,31,249,31,249,30,34,31,96,31,33,31,181,31,194,31,214,31,208,31,208,30,195,31,134,31,114,31,235,31,91,31,253,31,228,31,106,31,106,30,132,31,224,31,224,30,43,31,199,31,227,31,91,31,91,30,4,31,226,31,243,31,217,31,217,30,217,29,172,31,80,31,80,30,192,31,192,30,57,31,146,31,220,31,70,31,145,31,160,31,208,31,83,31,164,31,140,31,140,30,236,31,57,31,57,30,63,31,195,31,42,31,114,31,114,30,141,31,86,31,86,30,129,31,166,31,166,30,156,31,4,31,224,31,135,31,181,31,116,31,251,31,134,31,5,31,226,31,15,31,126,31,126,30,206,31,104,31,213,31,192,31,104,31,104,30,104,29,104,28,196,31,22,31,108,31,217,31,211,31,133,31,25,31,25,30,225,31,141,31,229,31,14,31,229,31,217,31,22,31,31,31,226,31,188,31,188,30,245,31,227,31,37,31,208,31,210,31,210,30,17,31,146,31,141,31,172,31,21,31,236,31,236,30,225,31,118,31,199,31,126,31,126,30,126,29,47,31,47,30,47,29,19,31,110,31,110,30,65,31,19,31,98,31,98,30,238,31,35,31,35,30,189,31,168,31,237,31,64,31,38,31,233,31,143,31,170,31,170,30,49,31,2,31,2,30,205,31,70,31,202,31,22,31,93,31,59,31,59,30,74,31,74,30,107,31,88,31,118,31,83,31,37,31,37,30,37,29,2,31,53,31,53,30,53,29,239,31,239,30,1,31,59,31,166,31,55,31,55,30,108,31,27,31,27,30,27,29,222,31,202,31,133,31,124,31,124,30,72,31,81,31,92,31,198,31,53,31,53,30,254,31,254,30,23,31,186,31,189,31,104,31,104,31,87,31,196,31,6,31,135,31,172,31,172,30,74,31,187,31,177,31,177,30,111,31,254,31,199,31,243,31,200,31,218,31,76,31,49,31,5,31,56,31,56,30,56,29,248,31,248,30,248,29,53,31,53,30,77,31,58,31,58,30,34,31,2,31,42,31,151,31,58,31,180,31,222,31,222,30,48,31,142,31,208,31,197,31,219,31,219,30,152,31,152,30,15,31,63,31,40,31,40,30,103,31,190,31,190,30,190,29,74,31,180,31,180,30,180,29,180,28,218,31,179,31,186,31,186,30,155,31,161,31,161,30,137,31,137,30,217,31,237,31,229,31,254,31,52,31,108,31,149,31,149,30,149,29,234,31,234,30,83,31,224,31,88,31,88,30,95,31,46,31,91,31,161,31,161,30,20,31,218,31,218,30,162,31,205,31,124,31,152,31,3,31,102,31,49,31,182,31,182,30,99,31,241,31,191,31,69,31,166,31,166,30,166,29,166,28,40,31,250,31,129,31,126,31,69,31,159,31,105,31,3,31,80,31,45,31,46,31,46,30,46,29,214,31,51,31,38,31,72,31,72,30,19,31,19,30,242,31,167,31,10,31,242,31,217,31,82,31,173,31,20,31,250,31,95,31,119,31,111,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
