-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 868;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (73,0,111,0,138,0,141,0,73,0,107,0,213,0,0,0,153,0,34,0,107,0,45,0,0,0,57,0,69,0,0,0,158,0,217,0,0,0,153,0,21,0,219,0,123,0,222,0,9,0,0,0,67,0,214,0,0,0,81,0,218,0,52,0,110,0,30,0,0,0,211,0,0,0,0,0,66,0,74,0,233,0,67,0,139,0,84,0,5,0,165,0,161,0,54,0,0,0,102,0,69,0,91,0,0,0,0,0,245,0,254,0,62,0,208,0,43,0,214,0,0,0,249,0,82,0,230,0,0,0,165,0,92,0,100,0,228,0,0,0,0,0,63,0,198,0,253,0,3,0,0,0,41,0,72,0,0,0,80,0,133,0,165,0,157,0,19,0,26,0,30,0,205,0,225,0,0,0,127,0,0,0,243,0,0,0,200,0,81,0,244,0,224,0,0,0,34,0,255,0,48,0,0,0,0,0,117,0,213,0,66,0,0,0,131,0,54,0,126,0,70,0,195,0,223,0,0,0,214,0,233,0,0,0,164,0,0,0,236,0,0,0,48,0,0,0,52,0,207,0,249,0,115,0,0,0,76,0,217,0,85,0,187,0,0,0,15,0,4,0,113,0,219,0,0,0,22,0,0,0,51,0,212,0,122,0,0,0,8,0,0,0,0,0,136,0,136,0,0,0,19,0,212,0,0,0,182,0,253,0,26,0,162,0,129,0,0,0,133,0,224,0,218,0,196,0,238,0,215,0,0,0,170,0,28,0,195,0,220,0,0,0,70,0,202,0,153,0,0,0,208,0,201,0,0,0,194,0,0,0,10,0,77,0,15,0,115,0,0,0,173,0,0,0,0,0,176,0,107,0,225,0,0,0,52,0,235,0,8,0,117,0,222,0,163,0,26,0,85,0,183,0,234,0,51,0,87,0,226,0,0,0,88,0,0,0,13,0,0,0,0,0,138,0,16,0,144,0,137,0,109,0,246,0,0,0,190,0,178,0,0,0,228,0,28,0,0,0,0,0,132,0,102,0,143,0,165,0,110,0,253,0,141,0,0,0,171,0,0,0,0,0,81,0,0,0,80,0,0,0,34,0,134,0,128,0,70,0,168,0,132,0,216,0,103,0,192,0,61,0,99,0,52,0,188,0,166,0,0,0,247,0,46,0,0,0,94,0,194,0,226,0,19,0,43,0,193,0,62,0,241,0,0,0,116,0,169,0,41,0,0,0,163,0,20,0,138,0,250,0,2,0,0,0,94,0,120,0,30,0,107,0,0,0,0,0,137,0,0,0,0,0,58,0,185,0,161,0,141,0,167,0,73,0,211,0,82,0,207,0,234,0,185,0,97,0,42,0,241,0,97,0,0,0,0,0,77,0,0,0,38,0,172,0,0,0,176,0,107,0,0,0,34,0,180,0,0,0,22,0,63,0,209,0,247,0,217,0,191,0,0,0,91,0,0,0,234,0,167,0,0,0,95,0,0,0,234,0,186,0,85,0,138,0,8,0,250,0,144,0,124,0,159,0,35,0,204,0,255,0,0,0,219,0,66,0,68,0,201,0,46,0,130,0,94,0,63,0,107,0,65,0,152,0,76,0,0,0,92,0,0,0,36,0,0,0,66,0,40,0,112,0,225,0,186,0,13,0,213,0,0,0,0,0,103,0,174,0,90,0,210,0,0,0,0,0,87,0,17,0,236,0,0,0,183,0,121,0,127,0,0,0,123,0,134,0,130,0,5,0,7,0,127,0,252,0,0,0,0,0,0,0,0,0,57,0,233,0,169,0,236,0,78,0,0,0,160,0,234,0,19,0,18,0,175,0,180,0,3,0,130,0,154,0,119,0,143,0,0,0,201,0,0,0,20,0,143,0,36,0,0,0,0,0,163,0,226,0,52,0,196,0,43,0,25,0,47,0,37,0,0,0,236,0,192,0,73,0,170,0,0,0,253,0,0,0,30,0,238,0,0,0,241,0,156,0,54,0,0,0,0,0,23,0,135,0,196,0,150,0,3,0,169,0,76,0,60,0,0,0,216,0,237,0,140,0,195,0,0,0,165,0,139,0,0,0,231,0,139,0,0,0,162,0,116,0,79,0,103,0,0,0,0,0,0,0,0,0,251,0,0,0,0,0,188,0,0,0,71,0,213,0,11,0,5,0,180,0,151,0,1,0,5,0,0,0,248,0,184,0,246,0,22,0,0,0,193,0,0,0,67,0,0,0,171,0,0,0,0,0,199,0,132,0,29,0,0,0,127,0,235,0,206,0,0,0,177,0,106,0,0,0,0,0,59,0,217,0,0,0,113,0,159,0,219,0,16,0,94,0,99,0,189,0,0,0,203,0,113,0,0,0,61,0,253,0,189,0,214,0,103,0,157,0,66,0,147,0,44,0,203,0,112,0,29,0,69,0,163,0,125,0,86,0,149,0,0,0,188,0,228,0,132,0,0,0,0,0,130,0,55,0,148,0,88,0,187,0,190,0,114,0,0,0,181,0,76,0,0,0,0,0,101,0,186,0,225,0,176,0,181,0,146,0,208,0,236,0,121,0,22,0,0,0,23,0,247,0,166,0,191,0,188,0,165,0,237,0,0,0,227,0,249,0,134,0,38,0,0,0,0,0,255,0,149,0,0,0,213,0,125,0,149,0,118,0,118,0,27,0,139,0,159,0,0,0,253,0,254,0,28,0,90,0,86,0,209,0,192,0,180,0,0,0,52,0,229,0,223,0,101,0,121,0,93,0,223,0,113,0,47,0,161,0,190,0,140,0,180,0,174,0,15,0,233,0,0,0,72,0,9,0,0,0,27,0,219,0,216,0,34,0,227,0,212,0,69,0,87,0,190,0,192,0,150,0,91,0,0,0,0,0,57,0,157,0,0,0,24,0,121,0,65,0,144,0,38,0,14,0,0,0,43,0,0,0,122,0,187,0,166,0,0,0,72,0,200,0,21,0,135,0,0,0,11,0,97,0,95,0,35,0,61,0,0,0,44,0,156,0,7,0,215,0,176,0,210,0,85,0,0,0,186,0,0,0,20,0,189,0,207,0,215,0,51,0,0,0,143,0,0,0,157,0,132,0,191,0,11,0,83,0,73,0,141,0,0,0,242,0,0,0,247,0,34,0,110,0,110,0,108,0,150,0,160,0,84,0,197,0,93,0,169,0,14,0,182,0,0,0,199,0,0,0,94,0,97,0,0,0,0,0,175,0,54,0,132,0,6,0,131,0,45,0,37,0,38,0,149,0,159,0,80,0,202,0,157,0,98,0,172,0,39,0,48,0,0,0,144,0,91,0,39,0,237,0,94,0,0,0,131,0,0,0,0,0,115,0,63,0,0,0,251,0,207,0,37,0,191,0,72,0,183,0,173,0,41,0,170,0,124,0,0,0,187,0,0,0,251,0,178,0,0,0,115,0,80,0,0,0,237,0,72,0,31,0,216,0,119,0,249,0,156,0,0,0,0,0,30,0,0,0,0,0,126,0,0,0,59,0,0,0,0,0,165,0,189,0,0,0,0,0,0,0,254,0,196,0,0,0,0,0,117,0,0,0,49,0,0,0,56,0,224,0,58,0,151,0,155,0,0,0,121,0,92,0,0,0,0,0,43,0,0,0,0,0,0,0,14,0,0,0,74,0,101,0,71,0,244,0,28,0,102,0,89,0,192,0,200,0,229,0,0,0,0,0,225,0,162,0,102,0,0,0,180,0,0,0,89,0,181,0,246,0,140,0,187,0,154,0,77,0,64,0,187,0,203,0,161,0,175,0,104,0,0,0,68,0,131,0,172,0,73,0,96,0,164,0,216,0,107,0,198,0,121,0,255,0,251,0,177,0,0,0,32,0,154,0,161,0,252,0,0,0,143,0,51,0,38,0,81,0,12,0,0,0,160,0,87,0,0,0,162,0,213,0);
signal scenario_full  : scenario_type := (73,31,111,31,138,31,141,31,73,31,107,31,213,31,213,30,153,31,34,31,107,31,45,31,45,30,57,31,69,31,69,30,158,31,217,31,217,30,153,31,21,31,219,31,123,31,222,31,9,31,9,30,67,31,214,31,214,30,81,31,218,31,52,31,110,31,30,31,30,30,211,31,211,30,211,29,66,31,74,31,233,31,67,31,139,31,84,31,5,31,165,31,161,31,54,31,54,30,102,31,69,31,91,31,91,30,91,29,245,31,254,31,62,31,208,31,43,31,214,31,214,30,249,31,82,31,230,31,230,30,165,31,92,31,100,31,228,31,228,30,228,29,63,31,198,31,253,31,3,31,3,30,41,31,72,31,72,30,80,31,133,31,165,31,157,31,19,31,26,31,30,31,205,31,225,31,225,30,127,31,127,30,243,31,243,30,200,31,81,31,244,31,224,31,224,30,34,31,255,31,48,31,48,30,48,29,117,31,213,31,66,31,66,30,131,31,54,31,126,31,70,31,195,31,223,31,223,30,214,31,233,31,233,30,164,31,164,30,236,31,236,30,48,31,48,30,52,31,207,31,249,31,115,31,115,30,76,31,217,31,85,31,187,31,187,30,15,31,4,31,113,31,219,31,219,30,22,31,22,30,51,31,212,31,122,31,122,30,8,31,8,30,8,29,136,31,136,31,136,30,19,31,212,31,212,30,182,31,253,31,26,31,162,31,129,31,129,30,133,31,224,31,218,31,196,31,238,31,215,31,215,30,170,31,28,31,195,31,220,31,220,30,70,31,202,31,153,31,153,30,208,31,201,31,201,30,194,31,194,30,10,31,77,31,15,31,115,31,115,30,173,31,173,30,173,29,176,31,107,31,225,31,225,30,52,31,235,31,8,31,117,31,222,31,163,31,26,31,85,31,183,31,234,31,51,31,87,31,226,31,226,30,88,31,88,30,13,31,13,30,13,29,138,31,16,31,144,31,137,31,109,31,246,31,246,30,190,31,178,31,178,30,228,31,28,31,28,30,28,29,132,31,102,31,143,31,165,31,110,31,253,31,141,31,141,30,171,31,171,30,171,29,81,31,81,30,80,31,80,30,34,31,134,31,128,31,70,31,168,31,132,31,216,31,103,31,192,31,61,31,99,31,52,31,188,31,166,31,166,30,247,31,46,31,46,30,94,31,194,31,226,31,19,31,43,31,193,31,62,31,241,31,241,30,116,31,169,31,41,31,41,30,163,31,20,31,138,31,250,31,2,31,2,30,94,31,120,31,30,31,107,31,107,30,107,29,137,31,137,30,137,29,58,31,185,31,161,31,141,31,167,31,73,31,211,31,82,31,207,31,234,31,185,31,97,31,42,31,241,31,97,31,97,30,97,29,77,31,77,30,38,31,172,31,172,30,176,31,107,31,107,30,34,31,180,31,180,30,22,31,63,31,209,31,247,31,217,31,191,31,191,30,91,31,91,30,234,31,167,31,167,30,95,31,95,30,234,31,186,31,85,31,138,31,8,31,250,31,144,31,124,31,159,31,35,31,204,31,255,31,255,30,219,31,66,31,68,31,201,31,46,31,130,31,94,31,63,31,107,31,65,31,152,31,76,31,76,30,92,31,92,30,36,31,36,30,66,31,40,31,112,31,225,31,186,31,13,31,213,31,213,30,213,29,103,31,174,31,90,31,210,31,210,30,210,29,87,31,17,31,236,31,236,30,183,31,121,31,127,31,127,30,123,31,134,31,130,31,5,31,7,31,127,31,252,31,252,30,252,29,252,28,252,27,57,31,233,31,169,31,236,31,78,31,78,30,160,31,234,31,19,31,18,31,175,31,180,31,3,31,130,31,154,31,119,31,143,31,143,30,201,31,201,30,20,31,143,31,36,31,36,30,36,29,163,31,226,31,52,31,196,31,43,31,25,31,47,31,37,31,37,30,236,31,192,31,73,31,170,31,170,30,253,31,253,30,30,31,238,31,238,30,241,31,156,31,54,31,54,30,54,29,23,31,135,31,196,31,150,31,3,31,169,31,76,31,60,31,60,30,216,31,237,31,140,31,195,31,195,30,165,31,139,31,139,30,231,31,139,31,139,30,162,31,116,31,79,31,103,31,103,30,103,29,103,28,103,27,251,31,251,30,251,29,188,31,188,30,71,31,213,31,11,31,5,31,180,31,151,31,1,31,5,31,5,30,248,31,184,31,246,31,22,31,22,30,193,31,193,30,67,31,67,30,171,31,171,30,171,29,199,31,132,31,29,31,29,30,127,31,235,31,206,31,206,30,177,31,106,31,106,30,106,29,59,31,217,31,217,30,113,31,159,31,219,31,16,31,94,31,99,31,189,31,189,30,203,31,113,31,113,30,61,31,253,31,189,31,214,31,103,31,157,31,66,31,147,31,44,31,203,31,112,31,29,31,69,31,163,31,125,31,86,31,149,31,149,30,188,31,228,31,132,31,132,30,132,29,130,31,55,31,148,31,88,31,187,31,190,31,114,31,114,30,181,31,76,31,76,30,76,29,101,31,186,31,225,31,176,31,181,31,146,31,208,31,236,31,121,31,22,31,22,30,23,31,247,31,166,31,191,31,188,31,165,31,237,31,237,30,227,31,249,31,134,31,38,31,38,30,38,29,255,31,149,31,149,30,213,31,125,31,149,31,118,31,118,31,27,31,139,31,159,31,159,30,253,31,254,31,28,31,90,31,86,31,209,31,192,31,180,31,180,30,52,31,229,31,223,31,101,31,121,31,93,31,223,31,113,31,47,31,161,31,190,31,140,31,180,31,174,31,15,31,233,31,233,30,72,31,9,31,9,30,27,31,219,31,216,31,34,31,227,31,212,31,69,31,87,31,190,31,192,31,150,31,91,31,91,30,91,29,57,31,157,31,157,30,24,31,121,31,65,31,144,31,38,31,14,31,14,30,43,31,43,30,122,31,187,31,166,31,166,30,72,31,200,31,21,31,135,31,135,30,11,31,97,31,95,31,35,31,61,31,61,30,44,31,156,31,7,31,215,31,176,31,210,31,85,31,85,30,186,31,186,30,20,31,189,31,207,31,215,31,51,31,51,30,143,31,143,30,157,31,132,31,191,31,11,31,83,31,73,31,141,31,141,30,242,31,242,30,247,31,34,31,110,31,110,31,108,31,150,31,160,31,84,31,197,31,93,31,169,31,14,31,182,31,182,30,199,31,199,30,94,31,97,31,97,30,97,29,175,31,54,31,132,31,6,31,131,31,45,31,37,31,38,31,149,31,159,31,80,31,202,31,157,31,98,31,172,31,39,31,48,31,48,30,144,31,91,31,39,31,237,31,94,31,94,30,131,31,131,30,131,29,115,31,63,31,63,30,251,31,207,31,37,31,191,31,72,31,183,31,173,31,41,31,170,31,124,31,124,30,187,31,187,30,251,31,178,31,178,30,115,31,80,31,80,30,237,31,72,31,31,31,216,31,119,31,249,31,156,31,156,30,156,29,30,31,30,30,30,29,126,31,126,30,59,31,59,30,59,29,165,31,189,31,189,30,189,29,189,28,254,31,196,31,196,30,196,29,117,31,117,30,49,31,49,30,56,31,224,31,58,31,151,31,155,31,155,30,121,31,92,31,92,30,92,29,43,31,43,30,43,29,43,28,14,31,14,30,74,31,101,31,71,31,244,31,28,31,102,31,89,31,192,31,200,31,229,31,229,30,229,29,225,31,162,31,102,31,102,30,180,31,180,30,89,31,181,31,246,31,140,31,187,31,154,31,77,31,64,31,187,31,203,31,161,31,175,31,104,31,104,30,68,31,131,31,172,31,73,31,96,31,164,31,216,31,107,31,198,31,121,31,255,31,251,31,177,31,177,30,32,31,154,31,161,31,252,31,252,30,143,31,51,31,38,31,81,31,12,31,12,30,160,31,87,31,87,30,162,31,213,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
