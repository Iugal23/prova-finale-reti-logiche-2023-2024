-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 831;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (216,0,0,0,243,0,0,0,203,0,60,0,229,0,221,0,190,0,238,0,15,0,0,0,207,0,214,0,49,0,0,0,49,0,0,0,231,0,0,0,102,0,152,0,181,0,0,0,87,0,136,0,171,0,167,0,131,0,154,0,74,0,0,0,95,0,134,0,130,0,0,0,210,0,181,0,26,0,189,0,8,0,246,0,197,0,206,0,120,0,31,0,28,0,137,0,175,0,181,0,14,0,116,0,174,0,118,0,233,0,54,0,200,0,162,0,0,0,235,0,0,0,175,0,253,0,197,0,250,0,46,0,54,0,82,0,0,0,0,0,11,0,54,0,153,0,0,0,91,0,130,0,110,0,53,0,156,0,243,0,123,0,187,0,112,0,0,0,63,0,119,0,110,0,0,0,36,0,0,0,0,0,207,0,73,0,152,0,0,0,14,0,65,0,79,0,72,0,242,0,17,0,0,0,56,0,223,0,0,0,59,0,96,0,98,0,4,0,0,0,126,0,0,0,0,0,191,0,243,0,63,0,0,0,106,0,53,0,0,0,249,0,83,0,255,0,25,0,248,0,177,0,1,0,221,0,210,0,0,0,0,0,54,0,247,0,50,0,31,0,9,0,54,0,0,0,157,0,190,0,138,0,173,0,69,0,71,0,61,0,29,0,0,0,0,0,139,0,15,0,0,0,16,0,5,0,129,0,180,0,106,0,74,0,96,0,19,0,118,0,18,0,0,0,0,0,0,0,27,0,18,0,67,0,24,0,0,0,142,0,40,0,200,0,29,0,130,0,222,0,119,0,127,0,140,0,221,0,155,0,94,0,246,0,95,0,252,0,0,0,0,0,111,0,23,0,0,0,0,0,79,0,239,0,167,0,56,0,0,0,133,0,17,0,35,0,0,0,0,0,127,0,0,0,210,0,0,0,0,0,115,0,0,0,188,0,126,0,109,0,159,0,89,0,0,0,42,0,1,0,103,0,126,0,221,0,214,0,150,0,221,0,165,0,18,0,240,0,235,0,175,0,214,0,0,0,74,0,37,0,169,0,112,0,155,0,0,0,98,0,32,0,57,0,127,0,48,0,38,0,132,0,40,0,216,0,164,0,251,0,216,0,168,0,70,0,0,0,117,0,143,0,93,0,0,0,32,0,0,0,154,0,0,0,224,0,167,0,127,0,0,0,14,0,48,0,122,0,67,0,85,0,153,0,37,0,0,0,21,0,0,0,0,0,121,0,130,0,0,0,143,0,35,0,12,0,224,0,0,0,49,0,192,0,89,0,202,0,94,0,0,0,0,0,245,0,44,0,8,0,17,0,40,0,225,0,201,0,179,0,32,0,20,0,24,0,41,0,44,0,0,0,73,0,22,0,116,0,214,0,8,0,110,0,16,0,151,0,202,0,0,0,252,0,33,0,19,0,148,0,197,0,109,0,0,0,69,0,0,0,6,0,144,0,32,0,119,0,192,0,70,0,127,0,0,0,0,0,59,0,0,0,255,0,24,0,85,0,227,0,72,0,33,0,169,0,165,0,3,0,136,0,39,0,0,0,0,0,46,0,0,0,198,0,127,0,0,0,101,0,228,0,248,0,232,0,162,0,91,0,0,0,7,0,36,0,170,0,66,0,122,0,194,0,236,0,231,0,108,0,41,0,7,0,69,0,229,0,99,0,189,0,83,0,49,0,165,0,123,0,61,0,37,0,6,0,182,0,117,0,0,0,122,0,144,0,216,0,193,0,121,0,181,0,0,0,98,0,0,0,253,0,135,0,152,0,66,0,6,0,84,0,114,0,186,0,231,0,182,0,70,0,39,0,210,0,44,0,212,0,36,0,77,0,141,0,154,0,53,0,162,0,228,0,236,0,0,0,46,0,17,0,189,0,196,0,179,0,184,0,0,0,43,0,27,0,12,0,0,0,76,0,76,0,67,0,196,0,188,0,41,0,243,0,0,0,0,0,227,0,13,0,21,0,41,0,85,0,0,0,199,0,80,0,243,0,192,0,22,0,214,0,128,0,152,0,165,0,92,0,0,0,0,0,166,0,0,0,0,0,0,0,170,0,249,0,28,0,0,0,124,0,0,0,143,0,43,0,176,0,55,0,199,0,143,0,0,0,169,0,147,0,210,0,6,0,143,0,19,0,0,0,129,0,133,0,71,0,0,0,28,0,253,0,189,0,247,0,110,0,37,0,180,0,195,0,121,0,15,0,127,0,49,0,15,0,251,0,179,0,115,0,178,0,167,0,240,0,110,0,69,0,148,0,0,0,97,0,40,0,0,0,18,0,0,0,72,0,138,0,180,0,27,0,153,0,225,0,33,0,8,0,165,0,246,0,90,0,0,0,31,0,235,0,223,0,173,0,176,0,109,0,45,0,168,0,111,0,0,0,234,0,183,0,7,0,40,0,94,0,192,0,0,0,69,0,44,0,0,0,204,0,125,0,0,0,131,0,65,0,0,0,206,0,15,0,147,0,0,0,0,0,60,0,73,0,143,0,120,0,0,0,66,0,118,0,74,0,3,0,252,0,252,0,157,0,59,0,37,0,0,0,0,0,125,0,0,0,0,0,0,0,231,0,69,0,129,0,63,0,75,0,93,0,115,0,4,0,32,0,40,0,0,0,138,0,210,0,235,0,234,0,214,0,0,0,255,0,233,0,0,0,25,0,84,0,47,0,74,0,0,0,28,0,185,0,0,0,53,0,139,0,253,0,0,0,0,0,71,0,0,0,146,0,107,0,78,0,2,0,208,0,153,0,56,0,136,0,139,0,198,0,61,0,172,0,202,0,248,0,168,0,38,0,203,0,247,0,11,0,221,0,217,0,145,0,87,0,143,0,182,0,149,0,166,0,16,0,111,0,3,0,181,0,0,0,141,0,0,0,0,0,66,0,40,0,5,0,82,0,17,0,83,0,0,0,79,0,44,0,212,0,159,0,0,0,188,0,109,0,0,0,191,0,49,0,82,0,6,0,42,0,252,0,0,0,0,0,169,0,255,0,146,0,0,0,0,0,177,0,0,0,244,0,73,0,180,0,105,0,19,0,190,0,74,0,0,0,127,0,175,0,210,0,141,0,180,0,219,0,43,0,232,0,89,0,198,0,3,0,0,0,75,0,52,0,187,0,147,0,71,0,44,0,184,0,55,0,199,0,0,0,47,0,49,0,206,0,234,0,247,0,13,0,125,0,251,0,44,0,8,0,0,0,0,0,0,0,178,0,52,0,116,0,0,0,182,0,87,0,0,0,0,0,213,0,161,0,65,0,199,0,244,0,245,0,127,0,0,0,0,0,0,0,195,0,46,0,209,0,100,0,156,0,0,0,66,0,80,0,0,0,36,0,175,0,140,0,107,0,88,0,190,0,236,0,0,0,184,0,102,0,50,0,149,0,94,0,0,0,0,0,118,0,222,0,201,0,3,0,207,0,235,0,199,0,53,0,243,0,154,0,95,0,21,0,0,0,5,0,0,0,228,0,149,0,220,0,127,0,175,0,60,0,221,0,237,0,29,0,22,0,22,0,205,0,204,0,0,0,137,0,22,0,88,0,73,0,199,0,55,0,0,0,74,0,101,0,214,0,148,0,44,0,0,0,31,0,0,0,124,0,94,0,80,0,161,0,204,0,130,0,149,0,223,0,18,0,196,0,0,0,0,0,112,0,70,0,236,0,220,0,0,0,0,0,232,0,54,0,205,0,0,0,175,0,0,0,67,0,178,0,129,0,221,0,126,0,204,0,206,0);
signal scenario_full  : scenario_type := (216,31,216,30,243,31,243,30,203,31,60,31,229,31,221,31,190,31,238,31,15,31,15,30,207,31,214,31,49,31,49,30,49,31,49,30,231,31,231,30,102,31,152,31,181,31,181,30,87,31,136,31,171,31,167,31,131,31,154,31,74,31,74,30,95,31,134,31,130,31,130,30,210,31,181,31,26,31,189,31,8,31,246,31,197,31,206,31,120,31,31,31,28,31,137,31,175,31,181,31,14,31,116,31,174,31,118,31,233,31,54,31,200,31,162,31,162,30,235,31,235,30,175,31,253,31,197,31,250,31,46,31,54,31,82,31,82,30,82,29,11,31,54,31,153,31,153,30,91,31,130,31,110,31,53,31,156,31,243,31,123,31,187,31,112,31,112,30,63,31,119,31,110,31,110,30,36,31,36,30,36,29,207,31,73,31,152,31,152,30,14,31,65,31,79,31,72,31,242,31,17,31,17,30,56,31,223,31,223,30,59,31,96,31,98,31,4,31,4,30,126,31,126,30,126,29,191,31,243,31,63,31,63,30,106,31,53,31,53,30,249,31,83,31,255,31,25,31,248,31,177,31,1,31,221,31,210,31,210,30,210,29,54,31,247,31,50,31,31,31,9,31,54,31,54,30,157,31,190,31,138,31,173,31,69,31,71,31,61,31,29,31,29,30,29,29,139,31,15,31,15,30,16,31,5,31,129,31,180,31,106,31,74,31,96,31,19,31,118,31,18,31,18,30,18,29,18,28,27,31,18,31,67,31,24,31,24,30,142,31,40,31,200,31,29,31,130,31,222,31,119,31,127,31,140,31,221,31,155,31,94,31,246,31,95,31,252,31,252,30,252,29,111,31,23,31,23,30,23,29,79,31,239,31,167,31,56,31,56,30,133,31,17,31,35,31,35,30,35,29,127,31,127,30,210,31,210,30,210,29,115,31,115,30,188,31,126,31,109,31,159,31,89,31,89,30,42,31,1,31,103,31,126,31,221,31,214,31,150,31,221,31,165,31,18,31,240,31,235,31,175,31,214,31,214,30,74,31,37,31,169,31,112,31,155,31,155,30,98,31,32,31,57,31,127,31,48,31,38,31,132,31,40,31,216,31,164,31,251,31,216,31,168,31,70,31,70,30,117,31,143,31,93,31,93,30,32,31,32,30,154,31,154,30,224,31,167,31,127,31,127,30,14,31,48,31,122,31,67,31,85,31,153,31,37,31,37,30,21,31,21,30,21,29,121,31,130,31,130,30,143,31,35,31,12,31,224,31,224,30,49,31,192,31,89,31,202,31,94,31,94,30,94,29,245,31,44,31,8,31,17,31,40,31,225,31,201,31,179,31,32,31,20,31,24,31,41,31,44,31,44,30,73,31,22,31,116,31,214,31,8,31,110,31,16,31,151,31,202,31,202,30,252,31,33,31,19,31,148,31,197,31,109,31,109,30,69,31,69,30,6,31,144,31,32,31,119,31,192,31,70,31,127,31,127,30,127,29,59,31,59,30,255,31,24,31,85,31,227,31,72,31,33,31,169,31,165,31,3,31,136,31,39,31,39,30,39,29,46,31,46,30,198,31,127,31,127,30,101,31,228,31,248,31,232,31,162,31,91,31,91,30,7,31,36,31,170,31,66,31,122,31,194,31,236,31,231,31,108,31,41,31,7,31,69,31,229,31,99,31,189,31,83,31,49,31,165,31,123,31,61,31,37,31,6,31,182,31,117,31,117,30,122,31,144,31,216,31,193,31,121,31,181,31,181,30,98,31,98,30,253,31,135,31,152,31,66,31,6,31,84,31,114,31,186,31,231,31,182,31,70,31,39,31,210,31,44,31,212,31,36,31,77,31,141,31,154,31,53,31,162,31,228,31,236,31,236,30,46,31,17,31,189,31,196,31,179,31,184,31,184,30,43,31,27,31,12,31,12,30,76,31,76,31,67,31,196,31,188,31,41,31,243,31,243,30,243,29,227,31,13,31,21,31,41,31,85,31,85,30,199,31,80,31,243,31,192,31,22,31,214,31,128,31,152,31,165,31,92,31,92,30,92,29,166,31,166,30,166,29,166,28,170,31,249,31,28,31,28,30,124,31,124,30,143,31,43,31,176,31,55,31,199,31,143,31,143,30,169,31,147,31,210,31,6,31,143,31,19,31,19,30,129,31,133,31,71,31,71,30,28,31,253,31,189,31,247,31,110,31,37,31,180,31,195,31,121,31,15,31,127,31,49,31,15,31,251,31,179,31,115,31,178,31,167,31,240,31,110,31,69,31,148,31,148,30,97,31,40,31,40,30,18,31,18,30,72,31,138,31,180,31,27,31,153,31,225,31,33,31,8,31,165,31,246,31,90,31,90,30,31,31,235,31,223,31,173,31,176,31,109,31,45,31,168,31,111,31,111,30,234,31,183,31,7,31,40,31,94,31,192,31,192,30,69,31,44,31,44,30,204,31,125,31,125,30,131,31,65,31,65,30,206,31,15,31,147,31,147,30,147,29,60,31,73,31,143,31,120,31,120,30,66,31,118,31,74,31,3,31,252,31,252,31,157,31,59,31,37,31,37,30,37,29,125,31,125,30,125,29,125,28,231,31,69,31,129,31,63,31,75,31,93,31,115,31,4,31,32,31,40,31,40,30,138,31,210,31,235,31,234,31,214,31,214,30,255,31,233,31,233,30,25,31,84,31,47,31,74,31,74,30,28,31,185,31,185,30,53,31,139,31,253,31,253,30,253,29,71,31,71,30,146,31,107,31,78,31,2,31,208,31,153,31,56,31,136,31,139,31,198,31,61,31,172,31,202,31,248,31,168,31,38,31,203,31,247,31,11,31,221,31,217,31,145,31,87,31,143,31,182,31,149,31,166,31,16,31,111,31,3,31,181,31,181,30,141,31,141,30,141,29,66,31,40,31,5,31,82,31,17,31,83,31,83,30,79,31,44,31,212,31,159,31,159,30,188,31,109,31,109,30,191,31,49,31,82,31,6,31,42,31,252,31,252,30,252,29,169,31,255,31,146,31,146,30,146,29,177,31,177,30,244,31,73,31,180,31,105,31,19,31,190,31,74,31,74,30,127,31,175,31,210,31,141,31,180,31,219,31,43,31,232,31,89,31,198,31,3,31,3,30,75,31,52,31,187,31,147,31,71,31,44,31,184,31,55,31,199,31,199,30,47,31,49,31,206,31,234,31,247,31,13,31,125,31,251,31,44,31,8,31,8,30,8,29,8,28,178,31,52,31,116,31,116,30,182,31,87,31,87,30,87,29,213,31,161,31,65,31,199,31,244,31,245,31,127,31,127,30,127,29,127,28,195,31,46,31,209,31,100,31,156,31,156,30,66,31,80,31,80,30,36,31,175,31,140,31,107,31,88,31,190,31,236,31,236,30,184,31,102,31,50,31,149,31,94,31,94,30,94,29,118,31,222,31,201,31,3,31,207,31,235,31,199,31,53,31,243,31,154,31,95,31,21,31,21,30,5,31,5,30,228,31,149,31,220,31,127,31,175,31,60,31,221,31,237,31,29,31,22,31,22,31,205,31,204,31,204,30,137,31,22,31,88,31,73,31,199,31,55,31,55,30,74,31,101,31,214,31,148,31,44,31,44,30,31,31,31,30,124,31,94,31,80,31,161,31,204,31,130,31,149,31,223,31,18,31,196,31,196,30,196,29,112,31,70,31,236,31,220,31,220,30,220,29,232,31,54,31,205,31,205,30,175,31,175,30,67,31,178,31,129,31,221,31,126,31,204,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
