-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 897;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,133,0,84,0,61,0,111,0,190,0,18,0,193,0,129,0,97,0,0,0,180,0,98,0,115,0,116,0,163,0,20,0,0,0,7,0,113,0,0,0,138,0,25,0,93,0,65,0,200,0,156,0,0,0,171,0,116,0,54,0,0,0,22,0,43,0,254,0,188,0,235,0,215,0,166,0,152,0,156,0,73,0,45,0,194,0,133,0,19,0,86,0,32,0,74,0,214,0,93,0,209,0,223,0,144,0,55,0,0,0,0,0,162,0,32,0,129,0,141,0,46,0,240,0,0,0,231,0,73,0,20,0,0,0,117,0,222,0,0,0,0,0,16,0,38,0,0,0,0,0,223,0,113,0,177,0,29,0,115,0,85,0,236,0,154,0,0,0,162,0,205,0,162,0,225,0,132,0,0,0,0,0,0,0,89,0,4,0,245,0,88,0,213,0,57,0,145,0,23,0,0,0,0,0,16,0,0,0,0,0,251,0,192,0,232,0,20,0,41,0,144,0,142,0,32,0,177,0,79,0,0,0,33,0,6,0,77,0,35,0,0,0,184,0,23,0,162,0,41,0,228,0,224,0,243,0,57,0,52,0,0,0,0,0,129,0,97,0,90,0,98,0,0,0,80,0,125,0,182,0,59,0,206,0,64,0,146,0,90,0,159,0,89,0,243,0,45,0,242,0,0,0,70,0,0,0,76,0,160,0,24,0,46,0,37,0,51,0,139,0,157,0,99,0,200,0,0,0,83,0,223,0,78,0,80,0,166,0,64,0,138,0,113,0,254,0,162,0,0,0,188,0,151,0,20,0,0,0,129,0,8,0,16,0,255,0,91,0,0,0,178,0,64,0,196,0,9,0,121,0,0,0,130,0,173,0,50,0,247,0,16,0,174,0,97,0,215,0,0,0,82,0,0,0,134,0,62,0,0,0,101,0,0,0,162,0,175,0,140,0,243,0,246,0,91,0,222,0,116,0,62,0,79,0,176,0,60,0,135,0,86,0,180,0,0,0,220,0,49,0,135,0,212,0,110,0,96,0,150,0,166,0,0,0,255,0,113,0,246,0,252,0,32,0,125,0,240,0,241,0,163,0,205,0,248,0,193,0,203,0,163,0,6,0,144,0,42,0,5,0,165,0,59,0,14,0,123,0,69,0,14,0,15,0,156,0,212,0,0,0,243,0,0,0,0,0,0,0,28,0,17,0,150,0,200,0,243,0,0,0,224,0,183,0,223,0,95,0,158,0,0,0,0,0,0,0,99,0,86,0,242,0,71,0,0,0,210,0,64,0,131,0,246,0,237,0,220,0,0,0,243,0,0,0,73,0,146,0,25,0,239,0,117,0,40,0,196,0,120,0,234,0,208,0,73,0,0,0,138,0,119,0,82,0,109,0,114,0,215,0,226,0,0,0,0,0,215,0,9,0,10,0,74,0,0,0,10,0,232,0,128,0,230,0,123,0,57,0,226,0,170,0,193,0,92,0,223,0,227,0,232,0,184,0,0,0,0,0,238,0,234,0,48,0,0,0,225,0,207,0,111,0,233,0,109,0,150,0,254,0,219,0,80,0,0,0,55,0,74,0,159,0,0,0,9,0,109,0,226,0,242,0,31,0,239,0,0,0,107,0,185,0,0,0,148,0,22,0,0,0,108,0,158,0,212,0,0,0,48,0,119,0,117,0,0,0,90,0,0,0,0,0,85,0,22,0,3,0,197,0,0,0,85,0,63,0,207,0,33,0,0,0,71,0,233,0,213,0,0,0,89,0,143,0,8,0,48,0,98,0,122,0,127,0,249,0,140,0,57,0,125,0,23,0,112,0,51,0,191,0,205,0,97,0,37,0,1,0,78,0,0,0,244,0,28,0,97,0,148,0,54,0,196,0,120,0,142,0,179,0,158,0,0,0,158,0,0,0,119,0,103,0,4,0,218,0,124,0,221,0,39,0,0,0,107,0,0,0,195,0,127,0,0,0,0,0,230,0,130,0,224,0,167,0,0,0,119,0,185,0,191,0,72,0,156,0,78,0,129,0,218,0,0,0,230,0,241,0,20,0,0,0,198,0,203,0,143,0,0,0,248,0,0,0,231,0,106,0,0,0,219,0,151,0,175,0,240,0,85,0,120,0,47,0,136,0,72,0,0,0,146,0,139,0,72,0,143,0,86,0,86,0,0,0,85,0,179,0,9,0,0,0,215,0,240,0,19,0,93,0,196,0,76,0,4,0,71,0,247,0,0,0,0,0,100,0,175,0,83,0,160,0,180,0,0,0,226,0,52,0,220,0,39,0,28,0,154,0,0,0,131,0,202,0,128,0,57,0,85,0,198,0,99,0,160,0,88,0,0,0,30,0,85,0,148,0,54,0,183,0,0,0,238,0,250,0,193,0,113,0,0,0,3,0,10,0,63,0,137,0,0,0,0,0,208,0,205,0,17,0,213,0,64,0,0,0,168,0,39,0,0,0,149,0,229,0,109,0,187,0,132,0,0,0,30,0,201,0,124,0,231,0,0,0,252,0,221,0,70,0,180,0,217,0,0,0,85,0,0,0,0,0,152,0,112,0,0,0,170,0,3,0,181,0,0,0,245,0,34,0,151,0,149,0,175,0,254,0,229,0,223,0,18,0,40,0,0,0,194,0,85,0,39,0,0,0,0,0,226,0,8,0,49,0,0,0,62,0,0,0,122,0,28,0,244,0,232,0,159,0,110,0,0,0,33,0,163,0,0,0,0,0,180,0,205,0,176,0,206,0,164,0,46,0,0,0,204,0,52,0,249,0,106,0,119,0,151,0,95,0,37,0,0,0,155,0,68,0,136,0,119,0,202,0,0,0,38,0,112,0,148,0,77,0,153,0,0,0,0,0,31,0,0,0,36,0,113,0,97,0,10,0,127,0,6,0,0,0,218,0,0,0,0,0,90,0,0,0,61,0,94,0,127,0,234,0,107,0,110,0,36,0,0,0,121,0,67,0,0,0,109,0,68,0,230,0,0,0,76,0,217,0,134,0,141,0,82,0,220,0,232,0,0,0,186,0,38,0,46,0,0,0,35,0,0,0,5,0,0,0,26,0,230,0,5,0,0,0,163,0,199,0,0,0,246,0,35,0,234,0,0,0,202,0,182,0,0,0,204,0,233,0,42,0,168,0,20,0,187,0,42,0,213,0,187,0,168,0,35,0,59,0,124,0,189,0,165,0,65,0,203,0,229,0,0,0,119,0,91,0,251,0,51,0,141,0,32,0,100,0,163,0,0,0,119,0,0,0,142,0,104,0,206,0,172,0,81,0,100,0,28,0,0,0,0,0,0,0,160,0,95,0,36,0,150,0,199,0,49,0,122,0,116,0,230,0,218,0,123,0,225,0,0,0,241,0,140,0,166,0,0,0,37,0,215,0,147,0,145,0,112,0,111,0,0,0,0,0,243,0,243,0,254,0,179,0,231,0,188,0,0,0,113,0,31,0,193,0,213,0,159,0,222,0,142,0,24,0,76,0,203,0,192,0,65,0,222,0,0,0,105,0,223,0,77,0,58,0,0,0,218,0,252,0,0,0,101,0,0,0,0,0,0,0,40,0,189,0,196,0,139,0,238,0,0,0,163,0,45,0,58,0,254,0,0,0,119,0,158,0,0,0,136,0,0,0,187,0,254,0,198,0,45,0,223,0,38,0,217,0,193,0,42,0,0,0,0,0,241,0,33,0,175,0,158,0,79,0,104,0,105,0,222,0,132,0,63,0,111,0,185,0,0,0,226,0,171,0,245,0,0,0,28,0,248,0,0,0,0,0,0,0,182,0,120,0,55,0,0,0,0,0,251,0,44,0,78,0,189,0,95,0,234,0,235,0,68,0,111,0,0,0,135,0,113,0,0,0,23,0,244,0,142,0,194,0,24,0,135,0,0,0,89,0,47,0,0,0,106,0,0,0,239,0,181,0,236,0,105,0,0,0,250,0,0,0,205,0,189,0,198,0,148,0,96,0,142,0,239,0,51,0,0,0,0,0,172,0,11,0,33,0,34,0,87,0,1,0,180,0,121,0);
signal scenario_full  : scenario_type := (147,31,133,31,84,31,61,31,111,31,190,31,18,31,193,31,129,31,97,31,97,30,180,31,98,31,115,31,116,31,163,31,20,31,20,30,7,31,113,31,113,30,138,31,25,31,93,31,65,31,200,31,156,31,156,30,171,31,116,31,54,31,54,30,22,31,43,31,254,31,188,31,235,31,215,31,166,31,152,31,156,31,73,31,45,31,194,31,133,31,19,31,86,31,32,31,74,31,214,31,93,31,209,31,223,31,144,31,55,31,55,30,55,29,162,31,32,31,129,31,141,31,46,31,240,31,240,30,231,31,73,31,20,31,20,30,117,31,222,31,222,30,222,29,16,31,38,31,38,30,38,29,223,31,113,31,177,31,29,31,115,31,85,31,236,31,154,31,154,30,162,31,205,31,162,31,225,31,132,31,132,30,132,29,132,28,89,31,4,31,245,31,88,31,213,31,57,31,145,31,23,31,23,30,23,29,16,31,16,30,16,29,251,31,192,31,232,31,20,31,41,31,144,31,142,31,32,31,177,31,79,31,79,30,33,31,6,31,77,31,35,31,35,30,184,31,23,31,162,31,41,31,228,31,224,31,243,31,57,31,52,31,52,30,52,29,129,31,97,31,90,31,98,31,98,30,80,31,125,31,182,31,59,31,206,31,64,31,146,31,90,31,159,31,89,31,243,31,45,31,242,31,242,30,70,31,70,30,76,31,160,31,24,31,46,31,37,31,51,31,139,31,157,31,99,31,200,31,200,30,83,31,223,31,78,31,80,31,166,31,64,31,138,31,113,31,254,31,162,31,162,30,188,31,151,31,20,31,20,30,129,31,8,31,16,31,255,31,91,31,91,30,178,31,64,31,196,31,9,31,121,31,121,30,130,31,173,31,50,31,247,31,16,31,174,31,97,31,215,31,215,30,82,31,82,30,134,31,62,31,62,30,101,31,101,30,162,31,175,31,140,31,243,31,246,31,91,31,222,31,116,31,62,31,79,31,176,31,60,31,135,31,86,31,180,31,180,30,220,31,49,31,135,31,212,31,110,31,96,31,150,31,166,31,166,30,255,31,113,31,246,31,252,31,32,31,125,31,240,31,241,31,163,31,205,31,248,31,193,31,203,31,163,31,6,31,144,31,42,31,5,31,165,31,59,31,14,31,123,31,69,31,14,31,15,31,156,31,212,31,212,30,243,31,243,30,243,29,243,28,28,31,17,31,150,31,200,31,243,31,243,30,224,31,183,31,223,31,95,31,158,31,158,30,158,29,158,28,99,31,86,31,242,31,71,31,71,30,210,31,64,31,131,31,246,31,237,31,220,31,220,30,243,31,243,30,73,31,146,31,25,31,239,31,117,31,40,31,196,31,120,31,234,31,208,31,73,31,73,30,138,31,119,31,82,31,109,31,114,31,215,31,226,31,226,30,226,29,215,31,9,31,10,31,74,31,74,30,10,31,232,31,128,31,230,31,123,31,57,31,226,31,170,31,193,31,92,31,223,31,227,31,232,31,184,31,184,30,184,29,238,31,234,31,48,31,48,30,225,31,207,31,111,31,233,31,109,31,150,31,254,31,219,31,80,31,80,30,55,31,74,31,159,31,159,30,9,31,109,31,226,31,242,31,31,31,239,31,239,30,107,31,185,31,185,30,148,31,22,31,22,30,108,31,158,31,212,31,212,30,48,31,119,31,117,31,117,30,90,31,90,30,90,29,85,31,22,31,3,31,197,31,197,30,85,31,63,31,207,31,33,31,33,30,71,31,233,31,213,31,213,30,89,31,143,31,8,31,48,31,98,31,122,31,127,31,249,31,140,31,57,31,125,31,23,31,112,31,51,31,191,31,205,31,97,31,37,31,1,31,78,31,78,30,244,31,28,31,97,31,148,31,54,31,196,31,120,31,142,31,179,31,158,31,158,30,158,31,158,30,119,31,103,31,4,31,218,31,124,31,221,31,39,31,39,30,107,31,107,30,195,31,127,31,127,30,127,29,230,31,130,31,224,31,167,31,167,30,119,31,185,31,191,31,72,31,156,31,78,31,129,31,218,31,218,30,230,31,241,31,20,31,20,30,198,31,203,31,143,31,143,30,248,31,248,30,231,31,106,31,106,30,219,31,151,31,175,31,240,31,85,31,120,31,47,31,136,31,72,31,72,30,146,31,139,31,72,31,143,31,86,31,86,31,86,30,85,31,179,31,9,31,9,30,215,31,240,31,19,31,93,31,196,31,76,31,4,31,71,31,247,31,247,30,247,29,100,31,175,31,83,31,160,31,180,31,180,30,226,31,52,31,220,31,39,31,28,31,154,31,154,30,131,31,202,31,128,31,57,31,85,31,198,31,99,31,160,31,88,31,88,30,30,31,85,31,148,31,54,31,183,31,183,30,238,31,250,31,193,31,113,31,113,30,3,31,10,31,63,31,137,31,137,30,137,29,208,31,205,31,17,31,213,31,64,31,64,30,168,31,39,31,39,30,149,31,229,31,109,31,187,31,132,31,132,30,30,31,201,31,124,31,231,31,231,30,252,31,221,31,70,31,180,31,217,31,217,30,85,31,85,30,85,29,152,31,112,31,112,30,170,31,3,31,181,31,181,30,245,31,34,31,151,31,149,31,175,31,254,31,229,31,223,31,18,31,40,31,40,30,194,31,85,31,39,31,39,30,39,29,226,31,8,31,49,31,49,30,62,31,62,30,122,31,28,31,244,31,232,31,159,31,110,31,110,30,33,31,163,31,163,30,163,29,180,31,205,31,176,31,206,31,164,31,46,31,46,30,204,31,52,31,249,31,106,31,119,31,151,31,95,31,37,31,37,30,155,31,68,31,136,31,119,31,202,31,202,30,38,31,112,31,148,31,77,31,153,31,153,30,153,29,31,31,31,30,36,31,113,31,97,31,10,31,127,31,6,31,6,30,218,31,218,30,218,29,90,31,90,30,61,31,94,31,127,31,234,31,107,31,110,31,36,31,36,30,121,31,67,31,67,30,109,31,68,31,230,31,230,30,76,31,217,31,134,31,141,31,82,31,220,31,232,31,232,30,186,31,38,31,46,31,46,30,35,31,35,30,5,31,5,30,26,31,230,31,5,31,5,30,163,31,199,31,199,30,246,31,35,31,234,31,234,30,202,31,182,31,182,30,204,31,233,31,42,31,168,31,20,31,187,31,42,31,213,31,187,31,168,31,35,31,59,31,124,31,189,31,165,31,65,31,203,31,229,31,229,30,119,31,91,31,251,31,51,31,141,31,32,31,100,31,163,31,163,30,119,31,119,30,142,31,104,31,206,31,172,31,81,31,100,31,28,31,28,30,28,29,28,28,160,31,95,31,36,31,150,31,199,31,49,31,122,31,116,31,230,31,218,31,123,31,225,31,225,30,241,31,140,31,166,31,166,30,37,31,215,31,147,31,145,31,112,31,111,31,111,30,111,29,243,31,243,31,254,31,179,31,231,31,188,31,188,30,113,31,31,31,193,31,213,31,159,31,222,31,142,31,24,31,76,31,203,31,192,31,65,31,222,31,222,30,105,31,223,31,77,31,58,31,58,30,218,31,252,31,252,30,101,31,101,30,101,29,101,28,40,31,189,31,196,31,139,31,238,31,238,30,163,31,45,31,58,31,254,31,254,30,119,31,158,31,158,30,136,31,136,30,187,31,254,31,198,31,45,31,223,31,38,31,217,31,193,31,42,31,42,30,42,29,241,31,33,31,175,31,158,31,79,31,104,31,105,31,222,31,132,31,63,31,111,31,185,31,185,30,226,31,171,31,245,31,245,30,28,31,248,31,248,30,248,29,248,28,182,31,120,31,55,31,55,30,55,29,251,31,44,31,78,31,189,31,95,31,234,31,235,31,68,31,111,31,111,30,135,31,113,31,113,30,23,31,244,31,142,31,194,31,24,31,135,31,135,30,89,31,47,31,47,30,106,31,106,30,239,31,181,31,236,31,105,31,105,30,250,31,250,30,205,31,189,31,198,31,148,31,96,31,142,31,239,31,51,31,51,30,51,29,172,31,11,31,33,31,34,31,87,31,1,31,180,31,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
