-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_242 is
end project_tb_242;

architecture project_tb_arch_242 of project_tb_242 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 373;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (194,0,65,0,181,0,73,0,249,0,70,0,184,0,188,0,241,0,0,0,0,0,156,0,225,0,125,0,2,0,0,0,157,0,221,0,36,0,203,0,0,0,0,0,105,0,231,0,98,0,47,0,127,0,30,0,82,0,0,0,0,0,52,0,0,0,207,0,220,0,116,0,0,0,0,0,227,0,9,0,154,0,181,0,130,0,128,0,184,0,148,0,249,0,131,0,50,0,84,0,67,0,0,0,0,0,0,0,101,0,0,0,210,0,0,0,57,0,23,0,131,0,91,0,212,0,159,0,0,0,149,0,28,0,48,0,82,0,132,0,100,0,19,0,220,0,224,0,22,0,147,0,220,0,58,0,86,0,221,0,0,0,46,0,126,0,0,0,0,0,139,0,4,0,144,0,66,0,163,0,58,0,0,0,67,0,56,0,18,0,27,0,211,0,31,0,34,0,96,0,196,0,122,0,69,0,5,0,0,0,0,0,98,0,255,0,0,0,218,0,138,0,0,0,115,0,115,0,0,0,114,0,238,0,0,0,33,0,155,0,174,0,170,0,32,0,0,0,138,0,154,0,226,0,0,0,227,0,130,0,174,0,40,0,185,0,193,0,1,0,184,0,151,0,20,0,0,0,0,0,80,0,214,0,196,0,22,0,71,0,109,0,82,0,0,0,0,0,91,0,185,0,90,0,62,0,83,0,77,0,217,0,88,0,53,0,166,0,51,0,237,0,189,0,227,0,219,0,219,0,0,0,192,0,235,0,0,0,240,0,203,0,0,0,135,0,0,0,129,0,0,0,189,0,0,0,91,0,156,0,242,0,76,0,0,0,93,0,241,0,0,0,136,0,134,0,241,0,0,0,138,0,229,0,15,0,141,0,159,0,102,0,192,0,235,0,246,0,50,0,89,0,234,0,106,0,198,0,70,0,46,0,71,0,177,0,75,0,0,0,162,0,60,0,105,0,84,0,143,0,0,0,140,0,166,0,0,0,124,0,54,0,0,0,76,0,219,0,0,0,116,0,75,0,40,0,175,0,0,0,104,0,53,0,109,0,113,0,45,0,127,0,110,0,206,0,0,0,0,0,136,0,157,0,235,0,75,0,253,0,0,0,185,0,108,0,85,0,186,0,160,0,87,0,211,0,90,0,0,0,3,0,161,0,0,0,124,0,0,0,0,0,0,0,248,0,0,0,37,0,47,0,0,0,112,0,164,0,18,0,0,0,0,0,62,0,121,0,0,0,252,0,124,0,214,0,154,0,0,0,0,0,0,0,151,0,128,0,86,0,216,0,68,0,49,0,74,0,177,0,66,0,0,0,60,0,78,0,17,0,0,0,179,0,72,0,62,0,0,0,23,0,0,0,201,0,133,0,189,0,205,0,68,0,221,0,0,0,129,0,7,0,188,0,12,0,0,0,0,0,172,0,208,0,0,0,42,0,254,0,26,0,138,0,73,0,0,0,9,0,105,0,3,0,148,0,144,0,202,0,210,0,49,0,147,0,52,0,57,0,0,0,48,0,0,0,119,0,231,0,150,0,10,0,0,0,15,0,110,0,220,0,66,0,163,0,237,0,93,0,207,0,69,0,4,0,0,0,0,0,187,0,247,0,169,0,0,0,237,0,110,0,210,0,135,0,0,0,0,0,252,0,227,0,0,0,0,0,169,0,191,0,135,0,0,0);
signal scenario_full  : scenario_type := (194,31,65,31,181,31,73,31,249,31,70,31,184,31,188,31,241,31,241,30,241,29,156,31,225,31,125,31,2,31,2,30,157,31,221,31,36,31,203,31,203,30,203,29,105,31,231,31,98,31,47,31,127,31,30,31,82,31,82,30,82,29,52,31,52,30,207,31,220,31,116,31,116,30,116,29,227,31,9,31,154,31,181,31,130,31,128,31,184,31,148,31,249,31,131,31,50,31,84,31,67,31,67,30,67,29,67,28,101,31,101,30,210,31,210,30,57,31,23,31,131,31,91,31,212,31,159,31,159,30,149,31,28,31,48,31,82,31,132,31,100,31,19,31,220,31,224,31,22,31,147,31,220,31,58,31,86,31,221,31,221,30,46,31,126,31,126,30,126,29,139,31,4,31,144,31,66,31,163,31,58,31,58,30,67,31,56,31,18,31,27,31,211,31,31,31,34,31,96,31,196,31,122,31,69,31,5,31,5,30,5,29,98,31,255,31,255,30,218,31,138,31,138,30,115,31,115,31,115,30,114,31,238,31,238,30,33,31,155,31,174,31,170,31,32,31,32,30,138,31,154,31,226,31,226,30,227,31,130,31,174,31,40,31,185,31,193,31,1,31,184,31,151,31,20,31,20,30,20,29,80,31,214,31,196,31,22,31,71,31,109,31,82,31,82,30,82,29,91,31,185,31,90,31,62,31,83,31,77,31,217,31,88,31,53,31,166,31,51,31,237,31,189,31,227,31,219,31,219,31,219,30,192,31,235,31,235,30,240,31,203,31,203,30,135,31,135,30,129,31,129,30,189,31,189,30,91,31,156,31,242,31,76,31,76,30,93,31,241,31,241,30,136,31,134,31,241,31,241,30,138,31,229,31,15,31,141,31,159,31,102,31,192,31,235,31,246,31,50,31,89,31,234,31,106,31,198,31,70,31,46,31,71,31,177,31,75,31,75,30,162,31,60,31,105,31,84,31,143,31,143,30,140,31,166,31,166,30,124,31,54,31,54,30,76,31,219,31,219,30,116,31,75,31,40,31,175,31,175,30,104,31,53,31,109,31,113,31,45,31,127,31,110,31,206,31,206,30,206,29,136,31,157,31,235,31,75,31,253,31,253,30,185,31,108,31,85,31,186,31,160,31,87,31,211,31,90,31,90,30,3,31,161,31,161,30,124,31,124,30,124,29,124,28,248,31,248,30,37,31,47,31,47,30,112,31,164,31,18,31,18,30,18,29,62,31,121,31,121,30,252,31,124,31,214,31,154,31,154,30,154,29,154,28,151,31,128,31,86,31,216,31,68,31,49,31,74,31,177,31,66,31,66,30,60,31,78,31,17,31,17,30,179,31,72,31,62,31,62,30,23,31,23,30,201,31,133,31,189,31,205,31,68,31,221,31,221,30,129,31,7,31,188,31,12,31,12,30,12,29,172,31,208,31,208,30,42,31,254,31,26,31,138,31,73,31,73,30,9,31,105,31,3,31,148,31,144,31,202,31,210,31,49,31,147,31,52,31,57,31,57,30,48,31,48,30,119,31,231,31,150,31,10,31,10,30,15,31,110,31,220,31,66,31,163,31,237,31,93,31,207,31,69,31,4,31,4,30,4,29,187,31,247,31,169,31,169,30,237,31,110,31,210,31,135,31,135,30,135,29,252,31,227,31,227,30,227,29,169,31,191,31,135,31,135,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
