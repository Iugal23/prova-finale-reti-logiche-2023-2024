-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 982;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,178,0,129,0,190,0,119,0,4,0,0,0,76,0,156,0,112,0,26,0,218,0,249,0,122,0,50,0,89,0,16,0,243,0,182,0,0,0,0,0,0,0,220,0,0,0,0,0,60,0,111,0,131,0,157,0,60,0,63,0,212,0,100,0,59,0,174,0,75,0,1,0,19,0,0,0,27,0,203,0,74,0,245,0,246,0,73,0,244,0,113,0,0,0,85,0,14,0,0,0,25,0,205,0,108,0,14,0,66,0,229,0,185,0,241,0,0,0,206,0,30,0,103,0,83,0,54,0,189,0,0,0,237,0,28,0,84,0,30,0,134,0,46,0,249,0,0,0,67,0,248,0,101,0,131,0,224,0,40,0,0,0,237,0,175,0,89,0,213,0,153,0,139,0,205,0,44,0,14,0,24,0,0,0,0,0,246,0,245,0,186,0,209,0,107,0,0,0,0,0,0,0,227,0,139,0,186,0,65,0,0,0,200,0,61,0,106,0,0,0,71,0,0,0,68,0,0,0,58,0,0,0,105,0,0,0,25,0,255,0,249,0,72,0,89,0,147,0,170,0,24,0,157,0,64,0,196,0,19,0,145,0,0,0,214,0,149,0,3,0,92,0,72,0,115,0,200,0,208,0,0,0,227,0,147,0,43,0,201,0,148,0,120,0,60,0,20,0,135,0,55,0,0,0,21,0,106,0,60,0,0,0,44,0,22,0,36,0,61,0,248,0,8,0,26,0,104,0,227,0,0,0,20,0,150,0,139,0,209,0,126,0,0,0,78,0,227,0,0,0,0,0,0,0,8,0,80,0,198,0,189,0,215,0,0,0,208,0,138,0,46,0,36,0,0,0,0,0,0,0,214,0,205,0,39,0,219,0,0,0,0,0,0,0,85,0,203,0,2,0,132,0,81,0,0,0,112,0,218,0,77,0,177,0,76,0,40,0,252,0,133,0,61,0,253,0,119,0,101,0,169,0,61,0,0,0,0,0,0,0,132,0,196,0,174,0,48,0,170,0,192,0,71,0,239,0,57,0,120,0,89,0,145,0,0,0,0,0,250,0,145,0,137,0,66,0,74,0,0,0,225,0,99,0,241,0,235,0,159,0,0,0,34,0,104,0,48,0,45,0,3,0,58,0,75,0,0,0,4,0,236,0,105,0,128,0,144,0,174,0,0,0,228,0,16,0,31,0,62,0,43,0,11,0,0,0,28,0,5,0,200,0,211,0,234,0,0,0,44,0,245,0,116,0,46,0,102,0,215,0,198,0,233,0,112,0,0,0,35,0,27,0,0,0,86,0,244,0,0,0,18,0,240,0,168,0,83,0,79,0,222,0,9,0,93,0,107,0,0,0,0,0,0,0,0,0,0,0,89,0,39,0,195,0,0,0,109,0,90,0,245,0,230,0,0,0,246,0,114,0,46,0,183,0,203,0,100,0,92,0,0,0,92,0,217,0,123,0,0,0,0,0,240,0,30,0,84,0,172,0,107,0,196,0,199,0,22,0,0,0,59,0,0,0,105,0,0,0,173,0,0,0,147,0,133,0,175,0,106,0,63,0,176,0,230,0,94,0,88,0,249,0,144,0,0,0,143,0,41,0,199,0,158,0,142,0,176,0,132,0,237,0,0,0,200,0,43,0,133,0,179,0,98,0,209,0,197,0,0,0,45,0,109,0,166,0,201,0,169,0,115,0,0,0,16,0,176,0,122,0,181,0,72,0,71,0,89,0,0,0,141,0,0,0,232,0,216,0,102,0,49,0,88,0,24,0,220,0,163,0,209,0,200,0,0,0,82,0,0,0,0,0,0,0,0,0,145,0,132,0,85,0,0,0,0,0,21,0,182,0,219,0,50,0,110,0,66,0,226,0,25,0,129,0,0,0,181,0,248,0,122,0,221,0,200,0,58,0,0,0,89,0,0,0,28,0,68,0,0,0,0,0,149,0,16,0,0,0,170,0,133,0,238,0,164,0,194,0,197,0,178,0,0,0,0,0,83,0,32,0,83,0,243,0,138,0,10,0,64,0,0,0,0,0,247,0,167,0,78,0,68,0,82,0,203,0,252,0,219,0,0,0,0,0,0,0,114,0,0,0,239,0,0,0,0,0,0,0,123,0,0,0,215,0,227,0,25,0,0,0,169,0,114,0,110,0,0,0,0,0,89,0,54,0,60,0,25,0,0,0,91,0,0,0,152,0,165,0,0,0,183,0,182,0,96,0,120,0,128,0,0,0,202,0,0,0,75,0,170,0,236,0,108,0,123,0,39,0,144,0,221,0,235,0,81,0,222,0,212,0,169,0,29,0,0,0,9,0,152,0,187,0,120,0,0,0,0,0,186,0,0,0,13,0,125,0,0,0,0,0,226,0,244,0,236,0,0,0,99,0,0,0,253,0,158,0,249,0,13,0,219,0,139,0,0,0,0,0,52,0,40,0,65,0,29,0,83,0,231,0,59,0,0,0,98,0,7,0,0,0,59,0,131,0,13,0,0,0,112,0,69,0,183,0,246,0,16,0,152,0,56,0,0,0,198,0,18,0,114,0,249,0,99,0,0,0,168,0,212,0,204,0,253,0,0,0,41,0,0,0,238,0,128,0,114,0,91,0,30,0,134,0,20,0,0,0,0,0,228,0,39,0,71,0,15,0,150,0,0,0,33,0,0,0,120,0,0,0,0,0,19,0,132,0,100,0,106,0,74,0,78,0,1,0,33,0,107,0,45,0,253,0,0,0,23,0,207,0,112,0,245,0,199,0,113,0,0,0,125,0,40,0,30,0,251,0,26,0,23,0,0,0,174,0,109,0,100,0,65,0,130,0,200,0,129,0,113,0,19,0,37,0,170,0,93,0,137,0,209,0,64,0,28,0,102,0,131,0,17,0,151,0,31,0,242,0,13,0,122,0,24,0,234,0,113,0,121,0,144,0,11,0,219,0,14,0,137,0,67,0,115,0,0,0,169,0,248,0,93,0,0,0,77,0,106,0,76,0,128,0,0,0,160,0,118,0,221,0,246,0,0,0,220,0,0,0,16,0,0,0,223,0,13,0,0,0,48,0,247,0,51,0,104,0,217,0,169,0,163,0,0,0,0,0,218,0,130,0,0,0,119,0,0,0,0,0,30,0,146,0,248,0,221,0,87,0,36,0,145,0,147,0,21,0,198,0,113,0,24,0,0,0,235,0,52,0,145,0,24,0,250,0,209,0,144,0,32,0,70,0,170,0,164,0,206,0,0,0,44,0,0,0,230,0,64,0,102,0,27,0,238,0,115,0,0,0,199,0,41,0,46,0,119,0,123,0,139,0,0,0,0,0,73,0,0,0,59,0,204,0,37,0,0,0,210,0,33,0,63,0,100,0,165,0,0,0,187,0,233,0,215,0,1,0,0,0,226,0,183,0,54,0,92,0,0,0,0,0,101,0,14,0,120,0,48,0,0,0,189,0,77,0,146,0,116,0,248,0,8,0,185,0,0,0,63,0,204,0,116,0,123,0,0,0,42,0,197,0,0,0,165,0,201,0,166,0,0,0,56,0,246,0,98,0,212,0,92,0,240,0,187,0,122,0,0,0,73,0,28,0,117,0,199,0,130,0,113,0,0,0,5,0,152,0,91,0,109,0,197,0,0,0,97,0,215,0,19,0,173,0,225,0,245,0,0,0,60,0,162,0,186,0,180,0,91,0,92,0,153,0,6,0,195,0,29,0,65,0,250,0,0,0,86,0,15,0,77,0,226,0,0,0,12,0,153,0,155,0,203,0,0,0,227,0,127,0,30,0,89,0,66,0,7,0,31,0,201,0,19,0,74,0,198,0,208,0,110,0,0,0,73,0,56,0,67,0,107,0,234,0,81,0,166,0,111,0,17,0,161,0,0,0,209,0,18,0,132,0,56,0,119,0,132,0,198,0,243,0,25,0,189,0,180,0,84,0,0,0,111,0,240,0,5,0,197,0,52,0,136,0,0,0,71,0,78,0,0,0,54,0,143,0,162,0,198,0,182,0,206,0,245,0,217,0,0,0,85,0,204,0,42,0,200,0,159,0,195,0,189,0,248,0,251,0,232,0,213,0,209,0,212,0,170,0,147,0,115,0,34,0,130,0,210,0,225,0,0,0,48,0,0,0,112,0,0,0,197,0,89,0,141,0,82,0,92,0,113,0,33,0,75,0,213,0,57,0,49,0,96,0,190,0,236,0,23,0,0,0,199,0,0,0,199,0,0,0,64,0,0,0,0,0,38,0,109,0,74,0,0,0,3,0,180,0,192,0,7,0,92,0,52,0,147,0,93,0,12,0,125,0,133,0,60,0,217,0,118,0,0,0,77,0,0,0,0,0,95,0,129,0,0,0,65,0,0,0,132,0,16,0,207,0,39,0,135,0,150,0,120,0,109,0,21,0,0,0,66,0,168,0,194,0);
signal scenario_full  : scenario_type := (181,31,178,31,129,31,190,31,119,31,4,31,4,30,76,31,156,31,112,31,26,31,218,31,249,31,122,31,50,31,89,31,16,31,243,31,182,31,182,30,182,29,182,28,220,31,220,30,220,29,60,31,111,31,131,31,157,31,60,31,63,31,212,31,100,31,59,31,174,31,75,31,1,31,19,31,19,30,27,31,203,31,74,31,245,31,246,31,73,31,244,31,113,31,113,30,85,31,14,31,14,30,25,31,205,31,108,31,14,31,66,31,229,31,185,31,241,31,241,30,206,31,30,31,103,31,83,31,54,31,189,31,189,30,237,31,28,31,84,31,30,31,134,31,46,31,249,31,249,30,67,31,248,31,101,31,131,31,224,31,40,31,40,30,237,31,175,31,89,31,213,31,153,31,139,31,205,31,44,31,14,31,24,31,24,30,24,29,246,31,245,31,186,31,209,31,107,31,107,30,107,29,107,28,227,31,139,31,186,31,65,31,65,30,200,31,61,31,106,31,106,30,71,31,71,30,68,31,68,30,58,31,58,30,105,31,105,30,25,31,255,31,249,31,72,31,89,31,147,31,170,31,24,31,157,31,64,31,196,31,19,31,145,31,145,30,214,31,149,31,3,31,92,31,72,31,115,31,200,31,208,31,208,30,227,31,147,31,43,31,201,31,148,31,120,31,60,31,20,31,135,31,55,31,55,30,21,31,106,31,60,31,60,30,44,31,22,31,36,31,61,31,248,31,8,31,26,31,104,31,227,31,227,30,20,31,150,31,139,31,209,31,126,31,126,30,78,31,227,31,227,30,227,29,227,28,8,31,80,31,198,31,189,31,215,31,215,30,208,31,138,31,46,31,36,31,36,30,36,29,36,28,214,31,205,31,39,31,219,31,219,30,219,29,219,28,85,31,203,31,2,31,132,31,81,31,81,30,112,31,218,31,77,31,177,31,76,31,40,31,252,31,133,31,61,31,253,31,119,31,101,31,169,31,61,31,61,30,61,29,61,28,132,31,196,31,174,31,48,31,170,31,192,31,71,31,239,31,57,31,120,31,89,31,145,31,145,30,145,29,250,31,145,31,137,31,66,31,74,31,74,30,225,31,99,31,241,31,235,31,159,31,159,30,34,31,104,31,48,31,45,31,3,31,58,31,75,31,75,30,4,31,236,31,105,31,128,31,144,31,174,31,174,30,228,31,16,31,31,31,62,31,43,31,11,31,11,30,28,31,5,31,200,31,211,31,234,31,234,30,44,31,245,31,116,31,46,31,102,31,215,31,198,31,233,31,112,31,112,30,35,31,27,31,27,30,86,31,244,31,244,30,18,31,240,31,168,31,83,31,79,31,222,31,9,31,93,31,107,31,107,30,107,29,107,28,107,27,107,26,89,31,39,31,195,31,195,30,109,31,90,31,245,31,230,31,230,30,246,31,114,31,46,31,183,31,203,31,100,31,92,31,92,30,92,31,217,31,123,31,123,30,123,29,240,31,30,31,84,31,172,31,107,31,196,31,199,31,22,31,22,30,59,31,59,30,105,31,105,30,173,31,173,30,147,31,133,31,175,31,106,31,63,31,176,31,230,31,94,31,88,31,249,31,144,31,144,30,143,31,41,31,199,31,158,31,142,31,176,31,132,31,237,31,237,30,200,31,43,31,133,31,179,31,98,31,209,31,197,31,197,30,45,31,109,31,166,31,201,31,169,31,115,31,115,30,16,31,176,31,122,31,181,31,72,31,71,31,89,31,89,30,141,31,141,30,232,31,216,31,102,31,49,31,88,31,24,31,220,31,163,31,209,31,200,31,200,30,82,31,82,30,82,29,82,28,82,27,145,31,132,31,85,31,85,30,85,29,21,31,182,31,219,31,50,31,110,31,66,31,226,31,25,31,129,31,129,30,181,31,248,31,122,31,221,31,200,31,58,31,58,30,89,31,89,30,28,31,68,31,68,30,68,29,149,31,16,31,16,30,170,31,133,31,238,31,164,31,194,31,197,31,178,31,178,30,178,29,83,31,32,31,83,31,243,31,138,31,10,31,64,31,64,30,64,29,247,31,167,31,78,31,68,31,82,31,203,31,252,31,219,31,219,30,219,29,219,28,114,31,114,30,239,31,239,30,239,29,239,28,123,31,123,30,215,31,227,31,25,31,25,30,169,31,114,31,110,31,110,30,110,29,89,31,54,31,60,31,25,31,25,30,91,31,91,30,152,31,165,31,165,30,183,31,182,31,96,31,120,31,128,31,128,30,202,31,202,30,75,31,170,31,236,31,108,31,123,31,39,31,144,31,221,31,235,31,81,31,222,31,212,31,169,31,29,31,29,30,9,31,152,31,187,31,120,31,120,30,120,29,186,31,186,30,13,31,125,31,125,30,125,29,226,31,244,31,236,31,236,30,99,31,99,30,253,31,158,31,249,31,13,31,219,31,139,31,139,30,139,29,52,31,40,31,65,31,29,31,83,31,231,31,59,31,59,30,98,31,7,31,7,30,59,31,131,31,13,31,13,30,112,31,69,31,183,31,246,31,16,31,152,31,56,31,56,30,198,31,18,31,114,31,249,31,99,31,99,30,168,31,212,31,204,31,253,31,253,30,41,31,41,30,238,31,128,31,114,31,91,31,30,31,134,31,20,31,20,30,20,29,228,31,39,31,71,31,15,31,150,31,150,30,33,31,33,30,120,31,120,30,120,29,19,31,132,31,100,31,106,31,74,31,78,31,1,31,33,31,107,31,45,31,253,31,253,30,23,31,207,31,112,31,245,31,199,31,113,31,113,30,125,31,40,31,30,31,251,31,26,31,23,31,23,30,174,31,109,31,100,31,65,31,130,31,200,31,129,31,113,31,19,31,37,31,170,31,93,31,137,31,209,31,64,31,28,31,102,31,131,31,17,31,151,31,31,31,242,31,13,31,122,31,24,31,234,31,113,31,121,31,144,31,11,31,219,31,14,31,137,31,67,31,115,31,115,30,169,31,248,31,93,31,93,30,77,31,106,31,76,31,128,31,128,30,160,31,118,31,221,31,246,31,246,30,220,31,220,30,16,31,16,30,223,31,13,31,13,30,48,31,247,31,51,31,104,31,217,31,169,31,163,31,163,30,163,29,218,31,130,31,130,30,119,31,119,30,119,29,30,31,146,31,248,31,221,31,87,31,36,31,145,31,147,31,21,31,198,31,113,31,24,31,24,30,235,31,52,31,145,31,24,31,250,31,209,31,144,31,32,31,70,31,170,31,164,31,206,31,206,30,44,31,44,30,230,31,64,31,102,31,27,31,238,31,115,31,115,30,199,31,41,31,46,31,119,31,123,31,139,31,139,30,139,29,73,31,73,30,59,31,204,31,37,31,37,30,210,31,33,31,63,31,100,31,165,31,165,30,187,31,233,31,215,31,1,31,1,30,226,31,183,31,54,31,92,31,92,30,92,29,101,31,14,31,120,31,48,31,48,30,189,31,77,31,146,31,116,31,248,31,8,31,185,31,185,30,63,31,204,31,116,31,123,31,123,30,42,31,197,31,197,30,165,31,201,31,166,31,166,30,56,31,246,31,98,31,212,31,92,31,240,31,187,31,122,31,122,30,73,31,28,31,117,31,199,31,130,31,113,31,113,30,5,31,152,31,91,31,109,31,197,31,197,30,97,31,215,31,19,31,173,31,225,31,245,31,245,30,60,31,162,31,186,31,180,31,91,31,92,31,153,31,6,31,195,31,29,31,65,31,250,31,250,30,86,31,15,31,77,31,226,31,226,30,12,31,153,31,155,31,203,31,203,30,227,31,127,31,30,31,89,31,66,31,7,31,31,31,201,31,19,31,74,31,198,31,208,31,110,31,110,30,73,31,56,31,67,31,107,31,234,31,81,31,166,31,111,31,17,31,161,31,161,30,209,31,18,31,132,31,56,31,119,31,132,31,198,31,243,31,25,31,189,31,180,31,84,31,84,30,111,31,240,31,5,31,197,31,52,31,136,31,136,30,71,31,78,31,78,30,54,31,143,31,162,31,198,31,182,31,206,31,245,31,217,31,217,30,85,31,204,31,42,31,200,31,159,31,195,31,189,31,248,31,251,31,232,31,213,31,209,31,212,31,170,31,147,31,115,31,34,31,130,31,210,31,225,31,225,30,48,31,48,30,112,31,112,30,197,31,89,31,141,31,82,31,92,31,113,31,33,31,75,31,213,31,57,31,49,31,96,31,190,31,236,31,23,31,23,30,199,31,199,30,199,31,199,30,64,31,64,30,64,29,38,31,109,31,74,31,74,30,3,31,180,31,192,31,7,31,92,31,52,31,147,31,93,31,12,31,125,31,133,31,60,31,217,31,118,31,118,30,77,31,77,30,77,29,95,31,129,31,129,30,65,31,65,30,132,31,16,31,207,31,39,31,135,31,150,31,120,31,109,31,21,31,21,30,66,31,168,31,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
