-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 438;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (98,0,92,0,254,0,4,0,221,0,22,0,108,0,111,0,31,0,0,0,241,0,218,0,169,0,0,0,245,0,36,0,82,0,136,0,228,0,0,0,1,0,0,0,167,0,24,0,0,0,58,0,0,0,28,0,0,0,182,0,133,0,11,0,63,0,35,0,120,0,60,0,173,0,215,0,228,0,11,0,0,0,63,0,230,0,205,0,177,0,119,0,44,0,29,0,0,0,131,0,0,0,192,0,39,0,51,0,12,0,1,0,197,0,0,0,83,0,113,0,48,0,195,0,0,0,127,0,37,0,122,0,87,0,6,0,247,0,147,0,52,0,56,0,126,0,2,0,165,0,73,0,97,0,0,0,0,0,109,0,54,0,117,0,133,0,106,0,82,0,0,0,149,0,237,0,0,0,8,0,84,0,0,0,165,0,238,0,0,0,168,0,200,0,0,0,4,0,181,0,0,0,107,0,0,0,12,0,202,0,191,0,32,0,252,0,181,0,228,0,0,0,0,0,167,0,103,0,45,0,161,0,59,0,0,0,10,0,150,0,117,0,0,0,190,0,247,0,107,0,0,0,14,0,245,0,0,0,84,0,89,0,119,0,0,0,117,0,0,0,234,0,0,0,0,0,181,0,234,0,84,0,62,0,105,0,245,0,55,0,169,0,0,0,0,0,85,0,0,0,0,0,228,0,107,0,117,0,15,0,0,0,166,0,197,0,0,0,237,0,131,0,159,0,0,0,131,0,251,0,76,0,57,0,7,0,0,0,0,0,9,0,208,0,0,0,18,0,162,0,195,0,171,0,196,0,26,0,129,0,0,0,28,0,18,0,96,0,173,0,215,0,23,0,0,0,159,0,0,0,0,0,0,0,113,0,229,0,43,0,181,0,97,0,142,0,135,0,219,0,0,0,243,0,21,0,79,0,247,0,175,0,58,0,125,0,0,0,136,0,0,0,46,0,0,0,197,0,19,0,155,0,121,0,51,0,219,0,156,0,112,0,117,0,83,0,227,0,7,0,235,0,129,0,59,0,0,0,64,0,0,0,219,0,60,0,129,0,250,0,136,0,148,0,150,0,189,0,158,0,10,0,136,0,182,0,40,0,0,0,164,0,31,0,224,0,0,0,237,0,102,0,239,0,246,0,1,0,203,0,219,0,80,0,0,0,101,0,74,0,131,0,180,0,0,0,1,0,131,0,132,0,237,0,227,0,33,0,0,0,87,0,0,0,0,0,108,0,46,0,100,0,244,0,183,0,40,0,183,0,129,0,14,0,185,0,167,0,14,0,0,0,70,0,52,0,82,0,122,0,72,0,143,0,242,0,140,0,48,0,179,0,57,0,138,0,0,0,0,0,119,0,0,0,26,0,17,0,0,0,42,0,96,0,109,0,86,0,109,0,0,0,129,0,217,0,203,0,57,0,114,0,0,0,48,0,0,0,112,0,192,0,0,0,235,0,78,0,57,0,0,0,227,0,82,0,94,0,39,0,238,0,194,0,234,0,249,0,48,0,35,0,0,0,0,0,37,0,64,0,0,0,16,0,62,0,0,0,0,0,0,0,112,0,176,0,135,0,20,0,24,0,1,0,90,0,0,0,150,0,186,0,0,0,0,0,0,0,151,0,0,0,233,0,66,0,187,0,25,0,185,0,31,0,210,0,146,0,65,0,179,0,0,0,0,0,129,0,0,0,178,0,69,0,0,0,249,0,30,0,102,0,16,0,81,0,102,0,210,0,112,0,18,0,213,0,141,0,0,0,13,0,94,0,0,0,206,0,221,0,81,0,250,0,90,0,87,0,129,0,23,0,0,0,248,0,27,0,38,0,170,0,186,0,237,0,90,0,186,0,0,0,40,0,0,0,0,0,87,0,57,0,98,0,179,0,170,0,218,0,138,0,0,0,182,0,202,0,118,0,189,0,11,0,14,0,135,0,0,0,161,0,85,0,91,0,254,0,0,0,0,0,121,0,70,0);
signal scenario_full  : scenario_type := (98,31,92,31,254,31,4,31,221,31,22,31,108,31,111,31,31,31,31,30,241,31,218,31,169,31,169,30,245,31,36,31,82,31,136,31,228,31,228,30,1,31,1,30,167,31,24,31,24,30,58,31,58,30,28,31,28,30,182,31,133,31,11,31,63,31,35,31,120,31,60,31,173,31,215,31,228,31,11,31,11,30,63,31,230,31,205,31,177,31,119,31,44,31,29,31,29,30,131,31,131,30,192,31,39,31,51,31,12,31,1,31,197,31,197,30,83,31,113,31,48,31,195,31,195,30,127,31,37,31,122,31,87,31,6,31,247,31,147,31,52,31,56,31,126,31,2,31,165,31,73,31,97,31,97,30,97,29,109,31,54,31,117,31,133,31,106,31,82,31,82,30,149,31,237,31,237,30,8,31,84,31,84,30,165,31,238,31,238,30,168,31,200,31,200,30,4,31,181,31,181,30,107,31,107,30,12,31,202,31,191,31,32,31,252,31,181,31,228,31,228,30,228,29,167,31,103,31,45,31,161,31,59,31,59,30,10,31,150,31,117,31,117,30,190,31,247,31,107,31,107,30,14,31,245,31,245,30,84,31,89,31,119,31,119,30,117,31,117,30,234,31,234,30,234,29,181,31,234,31,84,31,62,31,105,31,245,31,55,31,169,31,169,30,169,29,85,31,85,30,85,29,228,31,107,31,117,31,15,31,15,30,166,31,197,31,197,30,237,31,131,31,159,31,159,30,131,31,251,31,76,31,57,31,7,31,7,30,7,29,9,31,208,31,208,30,18,31,162,31,195,31,171,31,196,31,26,31,129,31,129,30,28,31,18,31,96,31,173,31,215,31,23,31,23,30,159,31,159,30,159,29,159,28,113,31,229,31,43,31,181,31,97,31,142,31,135,31,219,31,219,30,243,31,21,31,79,31,247,31,175,31,58,31,125,31,125,30,136,31,136,30,46,31,46,30,197,31,19,31,155,31,121,31,51,31,219,31,156,31,112,31,117,31,83,31,227,31,7,31,235,31,129,31,59,31,59,30,64,31,64,30,219,31,60,31,129,31,250,31,136,31,148,31,150,31,189,31,158,31,10,31,136,31,182,31,40,31,40,30,164,31,31,31,224,31,224,30,237,31,102,31,239,31,246,31,1,31,203,31,219,31,80,31,80,30,101,31,74,31,131,31,180,31,180,30,1,31,131,31,132,31,237,31,227,31,33,31,33,30,87,31,87,30,87,29,108,31,46,31,100,31,244,31,183,31,40,31,183,31,129,31,14,31,185,31,167,31,14,31,14,30,70,31,52,31,82,31,122,31,72,31,143,31,242,31,140,31,48,31,179,31,57,31,138,31,138,30,138,29,119,31,119,30,26,31,17,31,17,30,42,31,96,31,109,31,86,31,109,31,109,30,129,31,217,31,203,31,57,31,114,31,114,30,48,31,48,30,112,31,192,31,192,30,235,31,78,31,57,31,57,30,227,31,82,31,94,31,39,31,238,31,194,31,234,31,249,31,48,31,35,31,35,30,35,29,37,31,64,31,64,30,16,31,62,31,62,30,62,29,62,28,112,31,176,31,135,31,20,31,24,31,1,31,90,31,90,30,150,31,186,31,186,30,186,29,186,28,151,31,151,30,233,31,66,31,187,31,25,31,185,31,31,31,210,31,146,31,65,31,179,31,179,30,179,29,129,31,129,30,178,31,69,31,69,30,249,31,30,31,102,31,16,31,81,31,102,31,210,31,112,31,18,31,213,31,141,31,141,30,13,31,94,31,94,30,206,31,221,31,81,31,250,31,90,31,87,31,129,31,23,31,23,30,248,31,27,31,38,31,170,31,186,31,237,31,90,31,186,31,186,30,40,31,40,30,40,29,87,31,57,31,98,31,179,31,170,31,218,31,138,31,138,30,182,31,202,31,118,31,189,31,11,31,14,31,135,31,135,30,161,31,85,31,91,31,254,31,254,30,254,29,121,31,70,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
