-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_256 is
end project_tb_256;

architecture project_tb_arch_256 of project_tb_256 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 837;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (254,0,221,0,57,0,244,0,62,0,0,0,229,0,89,0,0,0,0,0,0,0,249,0,223,0,184,0,185,0,231,0,145,0,97,0,190,0,116,0,0,0,194,0,0,0,178,0,64,0,191,0,114,0,3,0,140,0,141,0,113,0,43,0,90,0,55,0,49,0,171,0,147,0,67,0,38,0,249,0,95,0,5,0,99,0,244,0,129,0,173,0,235,0,0,0,30,0,224,0,0,0,0,0,162,0,0,0,150,0,20,0,52,0,224,0,44,0,5,0,201,0,70,0,166,0,222,0,230,0,199,0,0,0,179,0,0,0,28,0,79,0,78,0,86,0,72,0,6,0,180,0,0,0,146,0,44,0,48,0,93,0,249,0,56,0,102,0,89,0,0,0,227,0,184,0,23,0,202,0,55,0,94,0,232,0,160,0,70,0,115,0,113,0,72,0,211,0,87,0,1,0,145,0,242,0,0,0,8,0,0,0,0,0,62,0,102,0,173,0,0,0,4,0,178,0,0,0,0,0,0,0,67,0,117,0,119,0,127,0,182,0,49,0,142,0,0,0,67,0,0,0,20,0,246,0,135,0,142,0,187,0,41,0,3,0,9,0,253,0,145,0,68,0,144,0,63,0,192,0,19,0,104,0,28,0,0,0,0,0,0,0,232,0,235,0,0,0,0,0,178,0,84,0,73,0,111,0,146,0,7,0,138,0,102,0,0,0,11,0,49,0,255,0,127,0,61,0,222,0,209,0,0,0,74,0,11,0,7,0,0,0,245,0,29,0,193,0,9,0,28,0,185,0,194,0,49,0,147,0,134,0,239,0,203,0,83,0,42,0,215,0,50,0,218,0,9,0,214,0,0,0,216,0,115,0,35,0,180,0,0,0,66,0,181,0,78,0,99,0,112,0,35,0,88,0,0,0,3,0,46,0,187,0,0,0,101,0,90,0,0,0,177,0,2,0,120,0,161,0,0,0,75,0,183,0,84,0,232,0,46,0,155,0,179,0,170,0,210,0,204,0,191,0,54,0,25,0,9,0,44,0,137,0,58,0,59,0,116,0,106,0,0,0,216,0,0,0,125,0,137,0,44,0,163,0,161,0,123,0,216,0,244,0,130,0,87,0,89,0,139,0,146,0,202,0,0,0,131,0,197,0,130,0,79,0,63,0,229,0,239,0,125,0,0,0,0,0,156,0,0,0,203,0,250,0,207,0,145,0,214,0,218,0,175,0,86,0,208,0,120,0,114,0,0,0,167,0,95,0,196,0,0,0,120,0,54,0,148,0,92,0,47,0,34,0,92,0,95,0,0,0,0,0,226,0,162,0,79,0,66,0,227,0,217,0,160,0,6,0,162,0,0,0,102,0,0,0,230,0,92,0,21,0,111,0,206,0,123,0,49,0,247,0,243,0,99,0,0,0,192,0,111,0,77,0,15,0,182,0,200,0,183,0,255,0,0,0,231,0,214,0,26,0,0,0,118,0,159,0,199,0,47,0,252,0,216,0,179,0,190,0,0,0,94,0,0,0,6,0,4,0,137,0,103,0,29,0,212,0,223,0,0,0,0,0,0,0,30,0,65,0,252,0,65,0,36,0,241,0,129,0,0,0,0,0,46,0,128,0,93,0,180,0,179,0,44,0,194,0,0,0,11,0,36,0,0,0,111,0,0,0,114,0,159,0,180,0,33,0,0,0,0,0,75,0,0,0,0,0,109,0,131,0,39,0,91,0,52,0,204,0,0,0,0,0,252,0,0,0,71,0,243,0,86,0,75,0,34,0,205,0,215,0,0,0,231,0,108,0,80,0,0,0,206,0,69,0,60,0,177,0,8,0,179,0,172,0,159,0,64,0,77,0,158,0,152,0,3,0,211,0,175,0,1,0,0,0,36,0,0,0,96,0,6,0,115,0,236,0,0,0,214,0,0,0,200,0,254,0,0,0,189,0,0,0,111,0,124,0,79,0,48,0,12,0,50,0,141,0,138,0,6,0,174,0,176,0,0,0,0,0,250,0,200,0,174,0,51,0,0,0,18,0,170,0,0,0,0,0,214,0,106,0,125,0,40,0,113,0,21,0,155,0,0,0,0,0,141,0,9,0,244,0,0,0,238,0,120,0,143,0,4,0,63,0,150,0,66,0,22,0,99,0,249,0,52,0,207,0,52,0,134,0,236,0,145,0,225,0,100,0,183,0,65,0,74,0,150,0,0,0,202,0,0,0,18,0,153,0,0,0,45,0,181,0,178,0,102,0,86,0,0,0,73,0,159,0,177,0,138,0,149,0,0,0,186,0,0,0,229,0,240,0,96,0,154,0,39,0,7,0,75,0,238,0,98,0,122,0,230,0,226,0,76,0,59,0,241,0,116,0,30,0,174,0,50,0,244,0,0,0,226,0,114,0,126,0,121,0,241,0,58,0,154,0,0,0,202,0,242,0,138,0,31,0,0,0,0,0,241,0,0,0,0,0,172,0,0,0,0,0,149,0,46,0,188,0,163,0,46,0,237,0,99,0,100,0,194,0,0,0,0,0,182,0,159,0,238,0,131,0,0,0,0,0,141,0,0,0,98,0,136,0,48,0,138,0,131,0,57,0,189,0,217,0,77,0,0,0,217,0,133,0,0,0,196,0,49,0,0,0,139,0,68,0,0,0,55,0,31,0,0,0,204,0,152,0,231,0,160,0,0,0,157,0,213,0,43,0,94,0,223,0,21,0,216,0,71,0,0,0,18,0,166,0,81,0,245,0,170,0,131,0,127,0,0,0,132,0,215,0,251,0,121,0,157,0,23,0,124,0,46,0,205,0,128,0,180,0,227,0,0,0,79,0,79,0,228,0,245,0,0,0,211,0,167,0,0,0,64,0,128,0,160,0,178,0,130,0,82,0,174,0,199,0,9,0,118,0,78,0,0,0,40,0,38,0,235,0,252,0,241,0,227,0,55,0,0,0,0,0,230,0,51,0,36,0,0,0,25,0,0,0,174,0,83,0,23,0,60,0,167,0,255,0,43,0,0,0,116,0,101,0,2,0,157,0,0,0,0,0,224,0,52,0,115,0,82,0,0,0,0,0,218,0,6,0,93,0,42,0,254,0,254,0,7,0,175,0,0,0,17,0,72,0,165,0,0,0,225,0,175,0,83,0,69,0,234,0,165,0,148,0,41,0,0,0,233,0,55,0,0,0,201,0,132,0,189,0,0,0,116,0,184,0,141,0,109,0,59,0,84,0,243,0,240,0,40,0,37,0,35,0,29,0,221,0,84,0,92,0,109,0,0,0,0,0,99,0,0,0,90,0,82,0,18,0,202,0,0,0,182,0,8,0,103,0,0,0,0,0,114,0,76,0,0,0,36,0,26,0,120,0,0,0,33,0,0,0,252,0,191,0,61,0,96,0,0,0,224,0,85,0,40,0,0,0,188,0,0,0,95,0,0,0,96,0,3,0,117,0,140,0,46,0,239,0,0,0,160,0,206,0,204,0,237,0,48,0,175,0,85,0,222,0,64,0,0,0,133,0,78,0,131,0,56,0,40,0,0,0,0,0,93,0,5,0,0,0,21,0,217,0,126,0,0,0,0,0,229,0,200,0,39,0,63,0,0,0,211,0,0,0,11,0,0,0,97,0,118,0,89,0,188,0,109,0,247,0,224,0,72,0,56,0,18,0,190,0,48,0,47,0,0,0,0,0,253,0,52,0,96,0,84,0,170,0,192,0,137,0,227,0,87,0,0,0,104,0,0,0,187,0,34,0,114,0,0,0,244,0,240,0);
signal scenario_full  : scenario_type := (254,31,221,31,57,31,244,31,62,31,62,30,229,31,89,31,89,30,89,29,89,28,249,31,223,31,184,31,185,31,231,31,145,31,97,31,190,31,116,31,116,30,194,31,194,30,178,31,64,31,191,31,114,31,3,31,140,31,141,31,113,31,43,31,90,31,55,31,49,31,171,31,147,31,67,31,38,31,249,31,95,31,5,31,99,31,244,31,129,31,173,31,235,31,235,30,30,31,224,31,224,30,224,29,162,31,162,30,150,31,20,31,52,31,224,31,44,31,5,31,201,31,70,31,166,31,222,31,230,31,199,31,199,30,179,31,179,30,28,31,79,31,78,31,86,31,72,31,6,31,180,31,180,30,146,31,44,31,48,31,93,31,249,31,56,31,102,31,89,31,89,30,227,31,184,31,23,31,202,31,55,31,94,31,232,31,160,31,70,31,115,31,113,31,72,31,211,31,87,31,1,31,145,31,242,31,242,30,8,31,8,30,8,29,62,31,102,31,173,31,173,30,4,31,178,31,178,30,178,29,178,28,67,31,117,31,119,31,127,31,182,31,49,31,142,31,142,30,67,31,67,30,20,31,246,31,135,31,142,31,187,31,41,31,3,31,9,31,253,31,145,31,68,31,144,31,63,31,192,31,19,31,104,31,28,31,28,30,28,29,28,28,232,31,235,31,235,30,235,29,178,31,84,31,73,31,111,31,146,31,7,31,138,31,102,31,102,30,11,31,49,31,255,31,127,31,61,31,222,31,209,31,209,30,74,31,11,31,7,31,7,30,245,31,29,31,193,31,9,31,28,31,185,31,194,31,49,31,147,31,134,31,239,31,203,31,83,31,42,31,215,31,50,31,218,31,9,31,214,31,214,30,216,31,115,31,35,31,180,31,180,30,66,31,181,31,78,31,99,31,112,31,35,31,88,31,88,30,3,31,46,31,187,31,187,30,101,31,90,31,90,30,177,31,2,31,120,31,161,31,161,30,75,31,183,31,84,31,232,31,46,31,155,31,179,31,170,31,210,31,204,31,191,31,54,31,25,31,9,31,44,31,137,31,58,31,59,31,116,31,106,31,106,30,216,31,216,30,125,31,137,31,44,31,163,31,161,31,123,31,216,31,244,31,130,31,87,31,89,31,139,31,146,31,202,31,202,30,131,31,197,31,130,31,79,31,63,31,229,31,239,31,125,31,125,30,125,29,156,31,156,30,203,31,250,31,207,31,145,31,214,31,218,31,175,31,86,31,208,31,120,31,114,31,114,30,167,31,95,31,196,31,196,30,120,31,54,31,148,31,92,31,47,31,34,31,92,31,95,31,95,30,95,29,226,31,162,31,79,31,66,31,227,31,217,31,160,31,6,31,162,31,162,30,102,31,102,30,230,31,92,31,21,31,111,31,206,31,123,31,49,31,247,31,243,31,99,31,99,30,192,31,111,31,77,31,15,31,182,31,200,31,183,31,255,31,255,30,231,31,214,31,26,31,26,30,118,31,159,31,199,31,47,31,252,31,216,31,179,31,190,31,190,30,94,31,94,30,6,31,4,31,137,31,103,31,29,31,212,31,223,31,223,30,223,29,223,28,30,31,65,31,252,31,65,31,36,31,241,31,129,31,129,30,129,29,46,31,128,31,93,31,180,31,179,31,44,31,194,31,194,30,11,31,36,31,36,30,111,31,111,30,114,31,159,31,180,31,33,31,33,30,33,29,75,31,75,30,75,29,109,31,131,31,39,31,91,31,52,31,204,31,204,30,204,29,252,31,252,30,71,31,243,31,86,31,75,31,34,31,205,31,215,31,215,30,231,31,108,31,80,31,80,30,206,31,69,31,60,31,177,31,8,31,179,31,172,31,159,31,64,31,77,31,158,31,152,31,3,31,211,31,175,31,1,31,1,30,36,31,36,30,96,31,6,31,115,31,236,31,236,30,214,31,214,30,200,31,254,31,254,30,189,31,189,30,111,31,124,31,79,31,48,31,12,31,50,31,141,31,138,31,6,31,174,31,176,31,176,30,176,29,250,31,200,31,174,31,51,31,51,30,18,31,170,31,170,30,170,29,214,31,106,31,125,31,40,31,113,31,21,31,155,31,155,30,155,29,141,31,9,31,244,31,244,30,238,31,120,31,143,31,4,31,63,31,150,31,66,31,22,31,99,31,249,31,52,31,207,31,52,31,134,31,236,31,145,31,225,31,100,31,183,31,65,31,74,31,150,31,150,30,202,31,202,30,18,31,153,31,153,30,45,31,181,31,178,31,102,31,86,31,86,30,73,31,159,31,177,31,138,31,149,31,149,30,186,31,186,30,229,31,240,31,96,31,154,31,39,31,7,31,75,31,238,31,98,31,122,31,230,31,226,31,76,31,59,31,241,31,116,31,30,31,174,31,50,31,244,31,244,30,226,31,114,31,126,31,121,31,241,31,58,31,154,31,154,30,202,31,242,31,138,31,31,31,31,30,31,29,241,31,241,30,241,29,172,31,172,30,172,29,149,31,46,31,188,31,163,31,46,31,237,31,99,31,100,31,194,31,194,30,194,29,182,31,159,31,238,31,131,31,131,30,131,29,141,31,141,30,98,31,136,31,48,31,138,31,131,31,57,31,189,31,217,31,77,31,77,30,217,31,133,31,133,30,196,31,49,31,49,30,139,31,68,31,68,30,55,31,31,31,31,30,204,31,152,31,231,31,160,31,160,30,157,31,213,31,43,31,94,31,223,31,21,31,216,31,71,31,71,30,18,31,166,31,81,31,245,31,170,31,131,31,127,31,127,30,132,31,215,31,251,31,121,31,157,31,23,31,124,31,46,31,205,31,128,31,180,31,227,31,227,30,79,31,79,31,228,31,245,31,245,30,211,31,167,31,167,30,64,31,128,31,160,31,178,31,130,31,82,31,174,31,199,31,9,31,118,31,78,31,78,30,40,31,38,31,235,31,252,31,241,31,227,31,55,31,55,30,55,29,230,31,51,31,36,31,36,30,25,31,25,30,174,31,83,31,23,31,60,31,167,31,255,31,43,31,43,30,116,31,101,31,2,31,157,31,157,30,157,29,224,31,52,31,115,31,82,31,82,30,82,29,218,31,6,31,93,31,42,31,254,31,254,31,7,31,175,31,175,30,17,31,72,31,165,31,165,30,225,31,175,31,83,31,69,31,234,31,165,31,148,31,41,31,41,30,233,31,55,31,55,30,201,31,132,31,189,31,189,30,116,31,184,31,141,31,109,31,59,31,84,31,243,31,240,31,40,31,37,31,35,31,29,31,221,31,84,31,92,31,109,31,109,30,109,29,99,31,99,30,90,31,82,31,18,31,202,31,202,30,182,31,8,31,103,31,103,30,103,29,114,31,76,31,76,30,36,31,26,31,120,31,120,30,33,31,33,30,252,31,191,31,61,31,96,31,96,30,224,31,85,31,40,31,40,30,188,31,188,30,95,31,95,30,96,31,3,31,117,31,140,31,46,31,239,31,239,30,160,31,206,31,204,31,237,31,48,31,175,31,85,31,222,31,64,31,64,30,133,31,78,31,131,31,56,31,40,31,40,30,40,29,93,31,5,31,5,30,21,31,217,31,126,31,126,30,126,29,229,31,200,31,39,31,63,31,63,30,211,31,211,30,11,31,11,30,97,31,118,31,89,31,188,31,109,31,247,31,224,31,72,31,56,31,18,31,190,31,48,31,47,31,47,30,47,29,253,31,52,31,96,31,84,31,170,31,192,31,137,31,227,31,87,31,87,30,104,31,104,30,187,31,34,31,114,31,114,30,244,31,240,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
