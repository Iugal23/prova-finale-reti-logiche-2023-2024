-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 855;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (86,0,10,0,0,0,224,0,83,0,101,0,200,0,4,0,103,0,233,0,20,0,26,0,154,0,88,0,0,0,42,0,0,0,73,0,27,0,56,0,44,0,240,0,156,0,0,0,139,0,189,0,200,0,82,0,0,0,244,0,241,0,0,0,254,0,147,0,0,0,21,0,151,0,20,0,88,0,247,0,133,0,151,0,249,0,0,0,52,0,113,0,117,0,0,0,116,0,143,0,86,0,132,0,113,0,211,0,21,0,154,0,118,0,178,0,0,0,0,0,22,0,0,0,0,0,151,0,97,0,88,0,87,0,0,0,234,0,175,0,0,0,142,0,129,0,168,0,175,0,164,0,30,0,95,0,14,0,101,0,181,0,0,0,140,0,4,0,18,0,32,0,227,0,3,0,55,0,30,0,38,0,0,0,178,0,50,0,239,0,23,0,0,0,216,0,17,0,136,0,0,0,154,0,147,0,56,0,139,0,0,0,0,0,76,0,79,0,50,0,54,0,173,0,125,0,213,0,243,0,217,0,134,0,233,0,157,0,136,0,0,0,254,0,249,0,0,0,177,0,181,0,69,0,92,0,149,0,73,0,21,0,11,0,83,0,0,0,0,0,205,0,85,0,247,0,66,0,14,0,32,0,129,0,55,0,218,0,155,0,0,0,126,0,16,0,158,0,142,0,209,0,175,0,65,0,69,0,137,0,203,0,153,0,14,0,224,0,34,0,253,0,0,0,45,0,56,0,17,0,18,0,48,0,114,0,246,0,152,0,143,0,109,0,100,0,144,0,186,0,166,0,116,0,40,0,0,0,0,0,183,0,94,0,27,0,106,0,206,0,146,0,47,0,253,0,77,0,155,0,55,0,238,0,0,0,0,0,75,0,136,0,185,0,142,0,131,0,104,0,0,0,253,0,187,0,211,0,29,0,94,0,153,0,99,0,204,0,20,0,91,0,86,0,24,0,234,0,188,0,106,0,0,0,83,0,0,0,0,0,190,0,134,0,0,0,31,0,208,0,142,0,191,0,34,0,0,0,0,0,220,0,166,0,0,0,0,0,0,0,249,0,251,0,0,0,0,0,215,0,233,0,87,0,15,0,34,0,240,0,194,0,95,0,48,0,221,0,129,0,198,0,73,0,124,0,197,0,121,0,128,0,211,0,171,0,224,0,49,0,253,0,182,0,122,0,214,0,59,0,52,0,126,0,73,0,132,0,74,0,252,0,202,0,138,0,161,0,8,0,0,0,184,0,80,0,44,0,154,0,239,0,182,0,34,0,76,0,52,0,14,0,226,0,38,0,0,0,0,0,0,0,233,0,0,0,0,0,212,0,152,0,57,0,94,0,85,0,0,0,0,0,117,0,109,0,111,0,153,0,106,0,0,0,215,0,37,0,0,0,184,0,178,0,168,0,184,0,232,0,114,0,0,0,60,0,254,0,15,0,137,0,0,0,80,0,28,0,72,0,58,0,159,0,74,0,29,0,2,0,0,0,223,0,126,0,156,0,0,0,66,0,136,0,230,0,127,0,0,0,0,0,104,0,0,0,0,0,247,0,202,0,214,0,164,0,0,0,0,0,238,0,159,0,105,0,221,0,81,0,134,0,0,0,249,0,0,0,209,0,96,0,52,0,0,0,32,0,0,0,145,0,198,0,70,0,164,0,198,0,76,0,184,0,149,0,0,0,164,0,201,0,0,0,195,0,155,0,115,0,9,0,77,0,0,0,218,0,157,0,46,0,105,0,163,0,228,0,217,0,177,0,138,0,0,0,198,0,13,0,163,0,254,0,0,0,0,0,56,0,0,0,143,0,0,0,46,0,251,0,133,0,0,0,102,0,0,0,108,0,14,0,0,0,0,0,79,0,0,0,0,0,201,0,0,0,0,0,53,0,236,0,185,0,208,0,51,0,130,0,221,0,186,0,102,0,195,0,29,0,214,0,0,0,55,0,156,0,53,0,131,0,18,0,92,0,35,0,0,0,0,0,211,0,0,0,122,0,0,0,112,0,104,0,111,0,0,0,143,0,123,0,34,0,202,0,215,0,0,0,248,0,37,0,0,0,22,0,85,0,168,0,91,0,205,0,154,0,187,0,240,0,142,0,241,0,177,0,248,0,51,0,0,0,148,0,129,0,0,0,0,0,81,0,172,0,236,0,200,0,73,0,247,0,242,0,28,0,166,0,22,0,119,0,73,0,118,0,116,0,212,0,0,0,137,0,1,0,0,0,4,0,3,0,200,0,220,0,169,0,233,0,218,0,207,0,116,0,152,0,0,0,84,0,22,0,161,0,0,0,104,0,0,0,254,0,113,0,146,0,0,0,180,0,4,0,35,0,139,0,0,0,228,0,126,0,219,0,208,0,16,0,75,0,225,0,176,0,5,0,203,0,106,0,0,0,0,0,0,0,54,0,134,0,81,0,45,0,188,0,146,0,0,0,231,0,32,0,28,0,104,0,247,0,7,0,188,0,169,0,3,0,191,0,47,0,0,0,58,0,55,0,63,0,10,0,152,0,180,0,0,0,89,0,132,0,164,0,150,0,80,0,235,0,8,0,4,0,151,0,44,0,0,0,181,0,51,0,218,0,64,0,58,0,67,0,135,0,235,0,196,0,254,0,0,0,78,0,101,0,253,0,188,0,15,0,110,0,137,0,79,0,98,0,66,0,21,0,77,0,231,0,28,0,0,0,231,0,1,0,158,0,71,0,3,0,0,0,15,0,174,0,200,0,140,0,56,0,244,0,65,0,253,0,226,0,128,0,157,0,124,0,82,0,130,0,145,0,8,0,163,0,174,0,20,0,141,0,16,0,0,0,0,0,0,0,123,0,0,0,61,0,71,0,92,0,233,0,0,0,158,0,0,0,190,0,120,0,0,0,180,0,106,0,53,0,140,0,30,0,194,0,236,0,0,0,228,0,0,0,0,0,132,0,2,0,135,0,231,0,0,0,184,0,246,0,0,0,81,0,8,0,184,0,113,0,104,0,0,0,0,0,0,0,52,0,0,0,41,0,184,0,196,0,222,0,148,0,17,0,0,0,0,0,6,0,216,0,196,0,37,0,0,0,162,0,114,0,0,0,47,0,63,0,24,0,139,0,253,0,203,0,13,0,48,0,205,0,27,0,146,0,136,0,49,0,0,0,0,0,204,0,157,0,132,0,0,0,115,0,207,0,236,0,0,0,0,0,39,0,253,0,98,0,131,0,0,0,126,0,150,0,156,0,0,0,225,0,0,0,15,0,175,0,27,0,15,0,148,0,103,0,227,0,168,0,0,0,0,0,201,0,18,0,197,0,158,0,76,0,153,0,116,0,1,0,195,0,140,0,0,0,145,0,153,0,202,0,239,0,124,0,0,0,0,0,208,0,12,0,80,0,0,0,26,0,96,0,0,0,65,0,77,0,39,0,91,0,57,0,77,0,95,0,121,0,27,0,193,0,197,0,142,0,209,0,134,0,153,0,70,0,43,0,182,0,64,0,152,0,0,0,239,0,169,0,17,0,6,0,87,0,0,0,190,0,0,0,0,0,36,0,241,0,223,0,246,0,6,0,24,0,0,0,0,0,224,0,159,0,84,0,0,0,166,0,142,0,0,0,0,0,70,0,0,0,170,0,24,0,128,0,0,0,0,0,201,0,108,0,195,0,0,0,79,0,0,0,0,0,0,0,168,0,0,0,122,0,180,0,0,0,219,0,0,0,194,0,13,0,73,0,54,0,201,0,208,0,0,0,144,0,122,0,245,0,40,0,8,0,8,0,138,0,124,0,79,0,193,0,1,0,30,0,142,0,0,0,0,0,138,0,197,0,220,0,0,0,132,0,157,0,92,0,105,0,141,0,10,0);
signal scenario_full  : scenario_type := (86,31,10,31,10,30,224,31,83,31,101,31,200,31,4,31,103,31,233,31,20,31,26,31,154,31,88,31,88,30,42,31,42,30,73,31,27,31,56,31,44,31,240,31,156,31,156,30,139,31,189,31,200,31,82,31,82,30,244,31,241,31,241,30,254,31,147,31,147,30,21,31,151,31,20,31,88,31,247,31,133,31,151,31,249,31,249,30,52,31,113,31,117,31,117,30,116,31,143,31,86,31,132,31,113,31,211,31,21,31,154,31,118,31,178,31,178,30,178,29,22,31,22,30,22,29,151,31,97,31,88,31,87,31,87,30,234,31,175,31,175,30,142,31,129,31,168,31,175,31,164,31,30,31,95,31,14,31,101,31,181,31,181,30,140,31,4,31,18,31,32,31,227,31,3,31,55,31,30,31,38,31,38,30,178,31,50,31,239,31,23,31,23,30,216,31,17,31,136,31,136,30,154,31,147,31,56,31,139,31,139,30,139,29,76,31,79,31,50,31,54,31,173,31,125,31,213,31,243,31,217,31,134,31,233,31,157,31,136,31,136,30,254,31,249,31,249,30,177,31,181,31,69,31,92,31,149,31,73,31,21,31,11,31,83,31,83,30,83,29,205,31,85,31,247,31,66,31,14,31,32,31,129,31,55,31,218,31,155,31,155,30,126,31,16,31,158,31,142,31,209,31,175,31,65,31,69,31,137,31,203,31,153,31,14,31,224,31,34,31,253,31,253,30,45,31,56,31,17,31,18,31,48,31,114,31,246,31,152,31,143,31,109,31,100,31,144,31,186,31,166,31,116,31,40,31,40,30,40,29,183,31,94,31,27,31,106,31,206,31,146,31,47,31,253,31,77,31,155,31,55,31,238,31,238,30,238,29,75,31,136,31,185,31,142,31,131,31,104,31,104,30,253,31,187,31,211,31,29,31,94,31,153,31,99,31,204,31,20,31,91,31,86,31,24,31,234,31,188,31,106,31,106,30,83,31,83,30,83,29,190,31,134,31,134,30,31,31,208,31,142,31,191,31,34,31,34,30,34,29,220,31,166,31,166,30,166,29,166,28,249,31,251,31,251,30,251,29,215,31,233,31,87,31,15,31,34,31,240,31,194,31,95,31,48,31,221,31,129,31,198,31,73,31,124,31,197,31,121,31,128,31,211,31,171,31,224,31,49,31,253,31,182,31,122,31,214,31,59,31,52,31,126,31,73,31,132,31,74,31,252,31,202,31,138,31,161,31,8,31,8,30,184,31,80,31,44,31,154,31,239,31,182,31,34,31,76,31,52,31,14,31,226,31,38,31,38,30,38,29,38,28,233,31,233,30,233,29,212,31,152,31,57,31,94,31,85,31,85,30,85,29,117,31,109,31,111,31,153,31,106,31,106,30,215,31,37,31,37,30,184,31,178,31,168,31,184,31,232,31,114,31,114,30,60,31,254,31,15,31,137,31,137,30,80,31,28,31,72,31,58,31,159,31,74,31,29,31,2,31,2,30,223,31,126,31,156,31,156,30,66,31,136,31,230,31,127,31,127,30,127,29,104,31,104,30,104,29,247,31,202,31,214,31,164,31,164,30,164,29,238,31,159,31,105,31,221,31,81,31,134,31,134,30,249,31,249,30,209,31,96,31,52,31,52,30,32,31,32,30,145,31,198,31,70,31,164,31,198,31,76,31,184,31,149,31,149,30,164,31,201,31,201,30,195,31,155,31,115,31,9,31,77,31,77,30,218,31,157,31,46,31,105,31,163,31,228,31,217,31,177,31,138,31,138,30,198,31,13,31,163,31,254,31,254,30,254,29,56,31,56,30,143,31,143,30,46,31,251,31,133,31,133,30,102,31,102,30,108,31,14,31,14,30,14,29,79,31,79,30,79,29,201,31,201,30,201,29,53,31,236,31,185,31,208,31,51,31,130,31,221,31,186,31,102,31,195,31,29,31,214,31,214,30,55,31,156,31,53,31,131,31,18,31,92,31,35,31,35,30,35,29,211,31,211,30,122,31,122,30,112,31,104,31,111,31,111,30,143,31,123,31,34,31,202,31,215,31,215,30,248,31,37,31,37,30,22,31,85,31,168,31,91,31,205,31,154,31,187,31,240,31,142,31,241,31,177,31,248,31,51,31,51,30,148,31,129,31,129,30,129,29,81,31,172,31,236,31,200,31,73,31,247,31,242,31,28,31,166,31,22,31,119,31,73,31,118,31,116,31,212,31,212,30,137,31,1,31,1,30,4,31,3,31,200,31,220,31,169,31,233,31,218,31,207,31,116,31,152,31,152,30,84,31,22,31,161,31,161,30,104,31,104,30,254,31,113,31,146,31,146,30,180,31,4,31,35,31,139,31,139,30,228,31,126,31,219,31,208,31,16,31,75,31,225,31,176,31,5,31,203,31,106,31,106,30,106,29,106,28,54,31,134,31,81,31,45,31,188,31,146,31,146,30,231,31,32,31,28,31,104,31,247,31,7,31,188,31,169,31,3,31,191,31,47,31,47,30,58,31,55,31,63,31,10,31,152,31,180,31,180,30,89,31,132,31,164,31,150,31,80,31,235,31,8,31,4,31,151,31,44,31,44,30,181,31,51,31,218,31,64,31,58,31,67,31,135,31,235,31,196,31,254,31,254,30,78,31,101,31,253,31,188,31,15,31,110,31,137,31,79,31,98,31,66,31,21,31,77,31,231,31,28,31,28,30,231,31,1,31,158,31,71,31,3,31,3,30,15,31,174,31,200,31,140,31,56,31,244,31,65,31,253,31,226,31,128,31,157,31,124,31,82,31,130,31,145,31,8,31,163,31,174,31,20,31,141,31,16,31,16,30,16,29,16,28,123,31,123,30,61,31,71,31,92,31,233,31,233,30,158,31,158,30,190,31,120,31,120,30,180,31,106,31,53,31,140,31,30,31,194,31,236,31,236,30,228,31,228,30,228,29,132,31,2,31,135,31,231,31,231,30,184,31,246,31,246,30,81,31,8,31,184,31,113,31,104,31,104,30,104,29,104,28,52,31,52,30,41,31,184,31,196,31,222,31,148,31,17,31,17,30,17,29,6,31,216,31,196,31,37,31,37,30,162,31,114,31,114,30,47,31,63,31,24,31,139,31,253,31,203,31,13,31,48,31,205,31,27,31,146,31,136,31,49,31,49,30,49,29,204,31,157,31,132,31,132,30,115,31,207,31,236,31,236,30,236,29,39,31,253,31,98,31,131,31,131,30,126,31,150,31,156,31,156,30,225,31,225,30,15,31,175,31,27,31,15,31,148,31,103,31,227,31,168,31,168,30,168,29,201,31,18,31,197,31,158,31,76,31,153,31,116,31,1,31,195,31,140,31,140,30,145,31,153,31,202,31,239,31,124,31,124,30,124,29,208,31,12,31,80,31,80,30,26,31,96,31,96,30,65,31,77,31,39,31,91,31,57,31,77,31,95,31,121,31,27,31,193,31,197,31,142,31,209,31,134,31,153,31,70,31,43,31,182,31,64,31,152,31,152,30,239,31,169,31,17,31,6,31,87,31,87,30,190,31,190,30,190,29,36,31,241,31,223,31,246,31,6,31,24,31,24,30,24,29,224,31,159,31,84,31,84,30,166,31,142,31,142,30,142,29,70,31,70,30,170,31,24,31,128,31,128,30,128,29,201,31,108,31,195,31,195,30,79,31,79,30,79,29,79,28,168,31,168,30,122,31,180,31,180,30,219,31,219,30,194,31,13,31,73,31,54,31,201,31,208,31,208,30,144,31,122,31,245,31,40,31,8,31,8,31,138,31,124,31,79,31,193,31,1,31,30,31,142,31,142,30,142,29,138,31,197,31,220,31,220,30,132,31,157,31,92,31,105,31,141,31,10,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
