-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_379 is
end project_tb_379;

architecture project_tb_arch_379 of project_tb_379 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 551;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (4,0,0,0,74,0,113,0,103,0,68,0,169,0,9,0,188,0,209,0,0,0,228,0,66,0,141,0,169,0,0,0,0,0,0,0,148,0,107,0,0,0,36,0,152,0,178,0,244,0,200,0,0,0,194,0,96,0,178,0,217,0,0,0,36,0,0,0,52,0,239,0,234,0,106,0,200,0,0,0,122,0,21,0,0,0,130,0,80,0,0,0,27,0,214,0,2,0,159,0,192,0,0,0,62,0,242,0,192,0,108,0,38,0,3,0,103,0,151,0,223,0,0,0,134,0,96,0,8,0,62,0,162,0,196,0,178,0,36,0,24,0,131,0,13,0,177,0,0,0,0,0,250,0,241,0,187,0,228,0,86,0,0,0,174,0,60,0,23,0,232,0,31,0,60,0,75,0,0,0,230,0,207,0,160,0,59,0,156,0,0,0,49,0,78,0,2,0,71,0,66,0,32,0,231,0,0,0,166,0,70,0,228,0,87,0,152,0,61,0,212,0,5,0,0,0,63,0,97,0,0,0,66,0,47,0,0,0,24,0,150,0,0,0,181,0,151,0,165,0,0,0,189,0,0,0,0,0,0,0,4,0,0,0,205,0,100,0,33,0,0,0,10,0,124,0,150,0,172,0,188,0,114,0,55,0,134,0,0,0,123,0,242,0,66,0,131,0,194,0,156,0,92,0,174,0,225,0,247,0,20,0,15,0,19,0,245,0,68,0,123,0,0,0,9,0,154,0,93,0,0,0,0,0,167,0,0,0,0,0,150,0,15,0,141,0,73,0,230,0,227,0,184,0,73,0,7,0,195,0,143,0,127,0,119,0,116,0,160,0,45,0,241,0,110,0,74,0,185,0,132,0,18,0,242,0,115,0,187,0,171,0,138,0,0,0,231,0,24,0,0,0,23,0,102,0,243,0,0,0,213,0,0,0,41,0,10,0,0,0,0,0,41,0,36,0,179,0,199,0,152,0,87,0,0,0,108,0,118,0,204,0,186,0,192,0,230,0,161,0,255,0,4,0,6,0,241,0,41,0,17,0,7,0,209,0,0,0,0,0,154,0,195,0,190,0,179,0,0,0,127,0,37,0,182,0,0,0,197,0,87,0,189,0,48,0,64,0,211,0,167,0,157,0,90,0,0,0,0,0,110,0,82,0,0,0,228,0,229,0,255,0,174,0,16,0,104,0,233,0,0,0,71,0,182,0,162,0,128,0,57,0,40,0,204,0,199,0,0,0,181,0,237,0,209,0,211,0,181,0,247,0,146,0,0,0,158,0,14,0,59,0,0,0,154,0,248,0,103,0,86,0,0,0,247,0,147,0,95,0,13,0,0,0,187,0,190,0,38,0,60,0,0,0,170,0,132,0,0,0,23,0,162,0,175,0,56,0,207,0,43,0,0,0,181,0,152,0,0,0,159,0,0,0,229,0,205,0,24,0,239,0,0,0,217,0,131,0,0,0,0,0,195,0,231,0,124,0,211,0,92,0,0,0,135,0,29,0,137,0,41,0,16,0,195,0,239,0,37,0,0,0,147,0,170,0,129,0,21,0,0,0,85,0,127,0,203,0,145,0,67,0,21,0,5,0,238,0,58,0,0,0,1,0,38,0,0,0,0,0,163,0,172,0,174,0,50,0,130,0,174,0,199,0,180,0,25,0,96,0,25,0,15,0,123,0,78,0,239,0,12,0,91,0,116,0,40,0,100,0,207,0,220,0,162,0,124,0,50,0,0,0,240,0,141,0,97,0,188,0,247,0,195,0,46,0,41,0,0,0,185,0,135,0,86,0,0,0,137,0,0,0,30,0,7,0,77,0,16,0,252,0,253,0,196,0,0,0,111,0,18,0,166,0,0,0,0,0,183,0,229,0,134,0,67,0,5,0,16,0,157,0,192,0,0,0,246,0,243,0,0,0,123,0,153,0,167,0,156,0,143,0,0,0,109,0,0,0,225,0,123,0,95,0,23,0,102,0,225,0,0,0,16,0,0,0,0,0,208,0,100,0,88,0,186,0,0,0,205,0,96,0,107,0,39,0,30,0,16,0,187,0,44,0,247,0,0,0,0,0,167,0,82,0,49,0,0,0,10,0,89,0,83,0,204,0,0,0,70,0,128,0,87,0,116,0,142,0,92,0,111,0,241,0,114,0,223,0,0,0,88,0,97,0,0,0,0,0,224,0,4,0,125,0,0,0,248,0,242,0,75,0,139,0,0,0,0,0,197,0,0,0,177,0,125,0,135,0,166,0,27,0,0,0,0,0,22,0,148,0,0,0,52,0,133,0,62,0,151,0,0,0,95,0,0,0,55,0,67,0,175,0,77,0,115,0,0,0,0,0,145,0,239,0,0,0,142,0,25,0,126,0,28,0,0,0,90,0,24,0,178,0,43,0,202,0,246,0,27,0,157,0,0,0,231,0,0,0,180,0,88,0,0,0,106,0,44,0,18,0,85,0,57,0,127,0,72,0,24,0,0,0);
signal scenario_full  : scenario_type := (4,31,4,30,74,31,113,31,103,31,68,31,169,31,9,31,188,31,209,31,209,30,228,31,66,31,141,31,169,31,169,30,169,29,169,28,148,31,107,31,107,30,36,31,152,31,178,31,244,31,200,31,200,30,194,31,96,31,178,31,217,31,217,30,36,31,36,30,52,31,239,31,234,31,106,31,200,31,200,30,122,31,21,31,21,30,130,31,80,31,80,30,27,31,214,31,2,31,159,31,192,31,192,30,62,31,242,31,192,31,108,31,38,31,3,31,103,31,151,31,223,31,223,30,134,31,96,31,8,31,62,31,162,31,196,31,178,31,36,31,24,31,131,31,13,31,177,31,177,30,177,29,250,31,241,31,187,31,228,31,86,31,86,30,174,31,60,31,23,31,232,31,31,31,60,31,75,31,75,30,230,31,207,31,160,31,59,31,156,31,156,30,49,31,78,31,2,31,71,31,66,31,32,31,231,31,231,30,166,31,70,31,228,31,87,31,152,31,61,31,212,31,5,31,5,30,63,31,97,31,97,30,66,31,47,31,47,30,24,31,150,31,150,30,181,31,151,31,165,31,165,30,189,31,189,30,189,29,189,28,4,31,4,30,205,31,100,31,33,31,33,30,10,31,124,31,150,31,172,31,188,31,114,31,55,31,134,31,134,30,123,31,242,31,66,31,131,31,194,31,156,31,92,31,174,31,225,31,247,31,20,31,15,31,19,31,245,31,68,31,123,31,123,30,9,31,154,31,93,31,93,30,93,29,167,31,167,30,167,29,150,31,15,31,141,31,73,31,230,31,227,31,184,31,73,31,7,31,195,31,143,31,127,31,119,31,116,31,160,31,45,31,241,31,110,31,74,31,185,31,132,31,18,31,242,31,115,31,187,31,171,31,138,31,138,30,231,31,24,31,24,30,23,31,102,31,243,31,243,30,213,31,213,30,41,31,10,31,10,30,10,29,41,31,36,31,179,31,199,31,152,31,87,31,87,30,108,31,118,31,204,31,186,31,192,31,230,31,161,31,255,31,4,31,6,31,241,31,41,31,17,31,7,31,209,31,209,30,209,29,154,31,195,31,190,31,179,31,179,30,127,31,37,31,182,31,182,30,197,31,87,31,189,31,48,31,64,31,211,31,167,31,157,31,90,31,90,30,90,29,110,31,82,31,82,30,228,31,229,31,255,31,174,31,16,31,104,31,233,31,233,30,71,31,182,31,162,31,128,31,57,31,40,31,204,31,199,31,199,30,181,31,237,31,209,31,211,31,181,31,247,31,146,31,146,30,158,31,14,31,59,31,59,30,154,31,248,31,103,31,86,31,86,30,247,31,147,31,95,31,13,31,13,30,187,31,190,31,38,31,60,31,60,30,170,31,132,31,132,30,23,31,162,31,175,31,56,31,207,31,43,31,43,30,181,31,152,31,152,30,159,31,159,30,229,31,205,31,24,31,239,31,239,30,217,31,131,31,131,30,131,29,195,31,231,31,124,31,211,31,92,31,92,30,135,31,29,31,137,31,41,31,16,31,195,31,239,31,37,31,37,30,147,31,170,31,129,31,21,31,21,30,85,31,127,31,203,31,145,31,67,31,21,31,5,31,238,31,58,31,58,30,1,31,38,31,38,30,38,29,163,31,172,31,174,31,50,31,130,31,174,31,199,31,180,31,25,31,96,31,25,31,15,31,123,31,78,31,239,31,12,31,91,31,116,31,40,31,100,31,207,31,220,31,162,31,124,31,50,31,50,30,240,31,141,31,97,31,188,31,247,31,195,31,46,31,41,31,41,30,185,31,135,31,86,31,86,30,137,31,137,30,30,31,7,31,77,31,16,31,252,31,253,31,196,31,196,30,111,31,18,31,166,31,166,30,166,29,183,31,229,31,134,31,67,31,5,31,16,31,157,31,192,31,192,30,246,31,243,31,243,30,123,31,153,31,167,31,156,31,143,31,143,30,109,31,109,30,225,31,123,31,95,31,23,31,102,31,225,31,225,30,16,31,16,30,16,29,208,31,100,31,88,31,186,31,186,30,205,31,96,31,107,31,39,31,30,31,16,31,187,31,44,31,247,31,247,30,247,29,167,31,82,31,49,31,49,30,10,31,89,31,83,31,204,31,204,30,70,31,128,31,87,31,116,31,142,31,92,31,111,31,241,31,114,31,223,31,223,30,88,31,97,31,97,30,97,29,224,31,4,31,125,31,125,30,248,31,242,31,75,31,139,31,139,30,139,29,197,31,197,30,177,31,125,31,135,31,166,31,27,31,27,30,27,29,22,31,148,31,148,30,52,31,133,31,62,31,151,31,151,30,95,31,95,30,55,31,67,31,175,31,77,31,115,31,115,30,115,29,145,31,239,31,239,30,142,31,25,31,126,31,28,31,28,30,90,31,24,31,178,31,43,31,202,31,246,31,27,31,157,31,157,30,231,31,231,30,180,31,88,31,88,30,106,31,44,31,18,31,85,31,57,31,127,31,72,31,24,31,24,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
