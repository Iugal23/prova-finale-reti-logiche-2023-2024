-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 976;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,27,0,104,0,241,0,169,0,70,0,101,0,0,0,97,0,246,0,0,0,161,0,217,0,88,0,20,0,40,0,127,0,187,0,0,0,86,0,0,0,157,0,139,0,59,0,88,0,78,0,1,0,144,0,95,0,0,0,192,0,111,0,42,0,224,0,79,0,206,0,234,0,146,0,150,0,41,0,0,0,0,0,0,0,38,0,0,0,0,0,194,0,179,0,0,0,0,0,242,0,248,0,0,0,156,0,128,0,17,0,196,0,0,0,160,0,251,0,149,0,83,0,16,0,156,0,0,0,143,0,0,0,26,0,248,0,110,0,129,0,250,0,213,0,75,0,58,0,94,0,246,0,143,0,243,0,136,0,228,0,178,0,49,0,64,0,153,0,27,0,172,0,41,0,212,0,17,0,87,0,163,0,252,0,204,0,0,0,220,0,239,0,0,0,0,0,194,0,0,0,244,0,41,0,241,0,77,0,206,0,251,0,0,0,132,0,17,0,223,0,127,0,0,0,20,0,156,0,0,0,61,0,215,0,203,0,38,0,88,0,123,0,0,0,135,0,27,0,184,0,168,0,0,0,181,0,255,0,171,0,237,0,106,0,111,0,176,0,96,0,24,0,129,0,16,0,0,0,209,0,156,0,62,0,0,0,242,0,139,0,86,0,137,0,184,0,197,0,0,0,169,0,0,0,0,0,0,0,37,0,228,0,0,0,34,0,197,0,113,0,118,0,147,0,47,0,233,0,0,0,131,0,0,0,105,0,219,0,0,0,137,0,32,0,86,0,126,0,0,0,113,0,199,0,248,0,147,0,168,0,81,0,84,0,72,0,132,0,145,0,67,0,230,0,21,0,198,0,77,0,124,0,133,0,0,0,0,0,113,0,192,0,152,0,159,0,187,0,11,0,134,0,171,0,94,0,89,0,1,0,133,0,60,0,0,0,97,0,97,0,224,0,0,0,56,0,31,0,171,0,109,0,185,0,0,0,0,0,123,0,0,0,241,0,147,0,0,0,167,0,20,0,73,0,59,0,60,0,0,0,207,0,0,0,67,0,0,0,169,0,72,0,55,0,22,0,236,0,103,0,111,0,242,0,33,0,149,0,197,0,0,0,0,0,41,0,0,0,148,0,120,0,204,0,236,0,91,0,136,0,245,0,62,0,0,0,0,0,98,0,122,0,0,0,120,0,92,0,60,0,210,0,180,0,8,0,182,0,0,0,0,0,40,0,79,0,0,0,92,0,30,0,182,0,22,0,0,0,96,0,243,0,56,0,243,0,215,0,100,0,238,0,141,0,231,0,199,0,153,0,61,0,29,0,168,0,6,0,1,0,178,0,132,0,38,0,63,0,47,0,0,0,75,0,0,0,79,0,21,0,105,0,57,0,0,0,66,0,251,0,34,0,0,0,34,0,156,0,252,0,242,0,0,0,7,0,58,0,214,0,35,0,35,0,42,0,0,0,0,0,0,0,117,0,68,0,98,0,152,0,210,0,61,0,181,0,0,0,227,0,195,0,243,0,0,0,0,0,40,0,0,0,219,0,23,0,25,0,123,0,0,0,177,0,21,0,33,0,9,0,46,0,92,0,246,0,181,0,38,0,0,0,164,0,171,0,185,0,206,0,189,0,0,0,187,0,162,0,189,0,5,0,180,0,48,0,180,0,126,0,0,0,38,0,201,0,0,0,182,0,1,0,0,0,252,0,18,0,0,0,149,0,0,0,66,0,243,0,41,0,233,0,89,0,208,0,110,0,0,0,0,0,176,0,0,0,230,0,74,0,71,0,120,0,0,0,172,0,44,0,160,0,212,0,0,0,0,0,176,0,116,0,209,0,154,0,26,0,60,0,64,0,248,0,188,0,228,0,218,0,106,0,127,0,0,0,164,0,194,0,190,0,16,0,128,0,185,0,0,0,73,0,56,0,0,0,9,0,130,0,221,0,37,0,111,0,175,0,7,0,85,0,8,0,132,0,176,0,0,0,158,0,212,0,80,0,28,0,0,0,253,0,0,0,104,0,207,0,144,0,137,0,127,0,48,0,205,0,98,0,0,0,50,0,57,0,124,0,226,0,29,0,229,0,83,0,0,0,0,0,111,0,255,0,134,0,143,0,0,0,67,0,77,0,96,0,167,0,186,0,158,0,160,0,164,0,49,0,0,0,0,0,0,0,58,0,98,0,125,0,0,0,219,0,0,0,47,0,247,0,94,0,242,0,170,0,0,0,0,0,105,0,202,0,0,0,7,0,145,0,249,0,0,0,14,0,25,0,173,0,199,0,231,0,143,0,9,0,0,0,0,0,190,0,54,0,196,0,0,0,66,0,233,0,93,0,197,0,52,0,169,0,11,0,217,0,106,0,197,0,84,0,143,0,0,0,204,0,0,0,98,0,0,0,0,0,220,0,148,0,0,0,76,0,133,0,235,0,205,0,71,0,46,0,88,0,73,0,158,0,97,0,202,0,0,0,52,0,185,0,2,0,90,0,0,0,38,0,232,0,38,0,0,0,59,0,44,0,131,0,250,0,97,0,118,0,0,0,177,0,33,0,232,0,119,0,215,0,34,0,5,0,142,0,103,0,0,0,7,0,48,0,11,0,210,0,29,0,23,0,60,0,91,0,15,0,89,0,1,0,106,0,132,0,149,0,83,0,190,0,242,0,156,0,204,0,44,0,211,0,40,0,211,0,102,0,214,0,56,0,240,0,89,0,13,0,59,0,19,0,0,0,204,0,25,0,136,0,229,0,47,0,0,0,0,0,0,0,126,0,76,0,210,0,149,0,197,0,0,0,148,0,0,0,0,0,0,0,252,0,13,0,72,0,160,0,227,0,127,0,130,0,255,0,98,0,230,0,159,0,163,0,22,0,143,0,133,0,65,0,174,0,7,0,180,0,0,0,0,0,0,0,0,0,120,0,0,0,17,0,27,0,62,0,62,0,92,0,21,0,91,0,194,0,97,0,58,0,48,0,42,0,243,0,124,0,145,0,242,0,147,0,44,0,83,0,186,0,102,0,229,0,64,0,41,0,0,0,220,0,25,0,154,0,173,0,71,0,174,0,239,0,252,0,47,0,213,0,81,0,237,0,170,0,0,0,99,0,0,0,103,0,0,0,70,0,215,0,236,0,161,0,0,0,15,0,34,0,246,0,20,0,139,0,128,0,63,0,77,0,69,0,183,0,120,0,113,0,232,0,181,0,0,0,228,0,30,0,43,0,236,0,138,0,179,0,215,0,34,0,0,0,33,0,123,0,59,0,0,0,111,0,123,0,190,0,60,0,97,0,155,0,167,0,50,0,215,0,30,0,100,0,143,0,186,0,14,0,0,0,100,0,186,0,229,0,42,0,0,0,0,0,181,0,126,0,205,0,246,0,62,0,9,0,147,0,126,0,134,0,141,0,0,0,0,0,25,0,171,0,0,0,0,0,6,0,49,0,1,0,205,0,38,0,208,0,208,0,192,0,96,0,90,0,86,0,74,0,167,0,0,0,22,0,54,0,108,0,0,0,50,0,190,0,243,0,88,0,0,0,218,0,54,0,125,0,156,0,181,0,142,0,0,0,0,0,159,0,3,0,0,0,127,0,156,0,235,0,41,0,2,0,31,0,185,0,23,0,249,0,0,0,0,0,152,0,135,0,0,0,247,0,0,0,38,0,0,0,119,0,108,0,0,0,184,0,30,0,0,0,109,0,182,0,194,0,176,0,132,0,118,0,195,0,0,0,69,0,42,0,0,0,0,0,108,0,196,0,235,0,18,0,165,0,54,0,1,0,114,0,47,0,251,0,0,0,238,0,191,0,91,0,225,0,212,0,161,0,234,0,242,0,28,0,132,0,250,0,0,0,143,0,0,0,5,0,0,0,179,0,208,0,0,0,61,0,29,0,0,0,186,0,155,0,0,0,198,0,108,0,162,0,214,0,118,0,0,0,35,0,48,0,254,0,15,0,167,0,153,0,0,0,0,0,90,0,215,0,33,0,230,0,169,0,172,0,205,0,0,0,224,0,239,0,209,0,160,0,144,0,0,0,0,0,0,0,64,0,0,0,0,0,176,0,0,0,0,0,76,0,232,0,25,0,50,0,154,0,116,0,172,0,88,0,176,0,175,0,99,0,171,0,0,0,0,0,0,0,196,0,190,0,82,0,92,0,248,0,136,0,152,0,204,0,43,0,0,0,58,0,29,0,37,0,0,0,132,0,112,0,16,0,203,0,251,0,31,0,26,0,18,0,18,0,0,0,24,0,63,0,81,0,0,0,64,0,0,0,168,0,56,0,25,0,170,0,203,0,119,0,108,0,226,0,3,0,115,0,91,0,195,0,199,0,67,0,244,0,0,0,0,0,69,0,226,0,213,0,0,0,187,0,0,0,90,0,0,0,240,0);
signal scenario_full  : scenario_type := (0,0,27,31,104,31,241,31,169,31,70,31,101,31,101,30,97,31,246,31,246,30,161,31,217,31,88,31,20,31,40,31,127,31,187,31,187,30,86,31,86,30,157,31,139,31,59,31,88,31,78,31,1,31,144,31,95,31,95,30,192,31,111,31,42,31,224,31,79,31,206,31,234,31,146,31,150,31,41,31,41,30,41,29,41,28,38,31,38,30,38,29,194,31,179,31,179,30,179,29,242,31,248,31,248,30,156,31,128,31,17,31,196,31,196,30,160,31,251,31,149,31,83,31,16,31,156,31,156,30,143,31,143,30,26,31,248,31,110,31,129,31,250,31,213,31,75,31,58,31,94,31,246,31,143,31,243,31,136,31,228,31,178,31,49,31,64,31,153,31,27,31,172,31,41,31,212,31,17,31,87,31,163,31,252,31,204,31,204,30,220,31,239,31,239,30,239,29,194,31,194,30,244,31,41,31,241,31,77,31,206,31,251,31,251,30,132,31,17,31,223,31,127,31,127,30,20,31,156,31,156,30,61,31,215,31,203,31,38,31,88,31,123,31,123,30,135,31,27,31,184,31,168,31,168,30,181,31,255,31,171,31,237,31,106,31,111,31,176,31,96,31,24,31,129,31,16,31,16,30,209,31,156,31,62,31,62,30,242,31,139,31,86,31,137,31,184,31,197,31,197,30,169,31,169,30,169,29,169,28,37,31,228,31,228,30,34,31,197,31,113,31,118,31,147,31,47,31,233,31,233,30,131,31,131,30,105,31,219,31,219,30,137,31,32,31,86,31,126,31,126,30,113,31,199,31,248,31,147,31,168,31,81,31,84,31,72,31,132,31,145,31,67,31,230,31,21,31,198,31,77,31,124,31,133,31,133,30,133,29,113,31,192,31,152,31,159,31,187,31,11,31,134,31,171,31,94,31,89,31,1,31,133,31,60,31,60,30,97,31,97,31,224,31,224,30,56,31,31,31,171,31,109,31,185,31,185,30,185,29,123,31,123,30,241,31,147,31,147,30,167,31,20,31,73,31,59,31,60,31,60,30,207,31,207,30,67,31,67,30,169,31,72,31,55,31,22,31,236,31,103,31,111,31,242,31,33,31,149,31,197,31,197,30,197,29,41,31,41,30,148,31,120,31,204,31,236,31,91,31,136,31,245,31,62,31,62,30,62,29,98,31,122,31,122,30,120,31,92,31,60,31,210,31,180,31,8,31,182,31,182,30,182,29,40,31,79,31,79,30,92,31,30,31,182,31,22,31,22,30,96,31,243,31,56,31,243,31,215,31,100,31,238,31,141,31,231,31,199,31,153,31,61,31,29,31,168,31,6,31,1,31,178,31,132,31,38,31,63,31,47,31,47,30,75,31,75,30,79,31,21,31,105,31,57,31,57,30,66,31,251,31,34,31,34,30,34,31,156,31,252,31,242,31,242,30,7,31,58,31,214,31,35,31,35,31,42,31,42,30,42,29,42,28,117,31,68,31,98,31,152,31,210,31,61,31,181,31,181,30,227,31,195,31,243,31,243,30,243,29,40,31,40,30,219,31,23,31,25,31,123,31,123,30,177,31,21,31,33,31,9,31,46,31,92,31,246,31,181,31,38,31,38,30,164,31,171,31,185,31,206,31,189,31,189,30,187,31,162,31,189,31,5,31,180,31,48,31,180,31,126,31,126,30,38,31,201,31,201,30,182,31,1,31,1,30,252,31,18,31,18,30,149,31,149,30,66,31,243,31,41,31,233,31,89,31,208,31,110,31,110,30,110,29,176,31,176,30,230,31,74,31,71,31,120,31,120,30,172,31,44,31,160,31,212,31,212,30,212,29,176,31,116,31,209,31,154,31,26,31,60,31,64,31,248,31,188,31,228,31,218,31,106,31,127,31,127,30,164,31,194,31,190,31,16,31,128,31,185,31,185,30,73,31,56,31,56,30,9,31,130,31,221,31,37,31,111,31,175,31,7,31,85,31,8,31,132,31,176,31,176,30,158,31,212,31,80,31,28,31,28,30,253,31,253,30,104,31,207,31,144,31,137,31,127,31,48,31,205,31,98,31,98,30,50,31,57,31,124,31,226,31,29,31,229,31,83,31,83,30,83,29,111,31,255,31,134,31,143,31,143,30,67,31,77,31,96,31,167,31,186,31,158,31,160,31,164,31,49,31,49,30,49,29,49,28,58,31,98,31,125,31,125,30,219,31,219,30,47,31,247,31,94,31,242,31,170,31,170,30,170,29,105,31,202,31,202,30,7,31,145,31,249,31,249,30,14,31,25,31,173,31,199,31,231,31,143,31,9,31,9,30,9,29,190,31,54,31,196,31,196,30,66,31,233,31,93,31,197,31,52,31,169,31,11,31,217,31,106,31,197,31,84,31,143,31,143,30,204,31,204,30,98,31,98,30,98,29,220,31,148,31,148,30,76,31,133,31,235,31,205,31,71,31,46,31,88,31,73,31,158,31,97,31,202,31,202,30,52,31,185,31,2,31,90,31,90,30,38,31,232,31,38,31,38,30,59,31,44,31,131,31,250,31,97,31,118,31,118,30,177,31,33,31,232,31,119,31,215,31,34,31,5,31,142,31,103,31,103,30,7,31,48,31,11,31,210,31,29,31,23,31,60,31,91,31,15,31,89,31,1,31,106,31,132,31,149,31,83,31,190,31,242,31,156,31,204,31,44,31,211,31,40,31,211,31,102,31,214,31,56,31,240,31,89,31,13,31,59,31,19,31,19,30,204,31,25,31,136,31,229,31,47,31,47,30,47,29,47,28,126,31,76,31,210,31,149,31,197,31,197,30,148,31,148,30,148,29,148,28,252,31,13,31,72,31,160,31,227,31,127,31,130,31,255,31,98,31,230,31,159,31,163,31,22,31,143,31,133,31,65,31,174,31,7,31,180,31,180,30,180,29,180,28,180,27,120,31,120,30,17,31,27,31,62,31,62,31,92,31,21,31,91,31,194,31,97,31,58,31,48,31,42,31,243,31,124,31,145,31,242,31,147,31,44,31,83,31,186,31,102,31,229,31,64,31,41,31,41,30,220,31,25,31,154,31,173,31,71,31,174,31,239,31,252,31,47,31,213,31,81,31,237,31,170,31,170,30,99,31,99,30,103,31,103,30,70,31,215,31,236,31,161,31,161,30,15,31,34,31,246,31,20,31,139,31,128,31,63,31,77,31,69,31,183,31,120,31,113,31,232,31,181,31,181,30,228,31,30,31,43,31,236,31,138,31,179,31,215,31,34,31,34,30,33,31,123,31,59,31,59,30,111,31,123,31,190,31,60,31,97,31,155,31,167,31,50,31,215,31,30,31,100,31,143,31,186,31,14,31,14,30,100,31,186,31,229,31,42,31,42,30,42,29,181,31,126,31,205,31,246,31,62,31,9,31,147,31,126,31,134,31,141,31,141,30,141,29,25,31,171,31,171,30,171,29,6,31,49,31,1,31,205,31,38,31,208,31,208,31,192,31,96,31,90,31,86,31,74,31,167,31,167,30,22,31,54,31,108,31,108,30,50,31,190,31,243,31,88,31,88,30,218,31,54,31,125,31,156,31,181,31,142,31,142,30,142,29,159,31,3,31,3,30,127,31,156,31,235,31,41,31,2,31,31,31,185,31,23,31,249,31,249,30,249,29,152,31,135,31,135,30,247,31,247,30,38,31,38,30,119,31,108,31,108,30,184,31,30,31,30,30,109,31,182,31,194,31,176,31,132,31,118,31,195,31,195,30,69,31,42,31,42,30,42,29,108,31,196,31,235,31,18,31,165,31,54,31,1,31,114,31,47,31,251,31,251,30,238,31,191,31,91,31,225,31,212,31,161,31,234,31,242,31,28,31,132,31,250,31,250,30,143,31,143,30,5,31,5,30,179,31,208,31,208,30,61,31,29,31,29,30,186,31,155,31,155,30,198,31,108,31,162,31,214,31,118,31,118,30,35,31,48,31,254,31,15,31,167,31,153,31,153,30,153,29,90,31,215,31,33,31,230,31,169,31,172,31,205,31,205,30,224,31,239,31,209,31,160,31,144,31,144,30,144,29,144,28,64,31,64,30,64,29,176,31,176,30,176,29,76,31,232,31,25,31,50,31,154,31,116,31,172,31,88,31,176,31,175,31,99,31,171,31,171,30,171,29,171,28,196,31,190,31,82,31,92,31,248,31,136,31,152,31,204,31,43,31,43,30,58,31,29,31,37,31,37,30,132,31,112,31,16,31,203,31,251,31,31,31,26,31,18,31,18,31,18,30,24,31,63,31,81,31,81,30,64,31,64,30,168,31,56,31,25,31,170,31,203,31,119,31,108,31,226,31,3,31,115,31,91,31,195,31,199,31,67,31,244,31,244,30,244,29,69,31,226,31,213,31,213,30,187,31,187,30,90,31,90,30,240,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
