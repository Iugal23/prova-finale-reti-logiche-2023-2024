-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 865;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (155,0,209,0,191,0,240,0,77,0,96,0,96,0,0,0,89,0,0,0,154,0,113,0,78,0,44,0,149,0,9,0,0,0,0,0,0,0,188,0,245,0,74,0,80,0,42,0,249,0,181,0,0,0,65,0,87,0,82,0,253,0,113,0,108,0,0,0,225,0,0,0,161,0,103,0,247,0,242,0,0,0,61,0,0,0,156,0,80,0,247,0,85,0,29,0,119,0,0,0,78,0,0,0,0,0,128,0,251,0,0,0,225,0,245,0,0,0,29,0,71,0,167,0,39,0,244,0,129,0,60,0,217,0,213,0,0,0,252,0,136,0,0,0,7,0,203,0,199,0,0,0,200,0,94,0,73,0,238,0,189,0,11,0,0,0,0,0,213,0,0,0,168,0,152,0,109,0,83,0,107,0,34,0,0,0,88,0,218,0,174,0,161,0,131,0,72,0,132,0,249,0,162,0,81,0,58,0,114,0,51,0,172,0,245,0,0,0,0,0,193,0,102,0,37,0,0,0,38,0,177,0,12,0,159,0,245,0,27,0,0,0,90,0,91,0,0,0,170,0,254,0,0,0,221,0,23,0,147,0,232,0,122,0,152,0,183,0,33,0,76,0,0,0,186,0,37,0,0,0,210,0,120,0,217,0,162,0,185,0,36,0,97,0,103,0,0,0,138,0,0,0,144,0,217,0,0,0,60,0,87,0,0,0,166,0,25,0,203,0,40,0,129,0,0,0,47,0,22,0,156,0,60,0,234,0,173,0,53,0,253,0,160,0,106,0,188,0,161,0,186,0,128,0,188,0,29,0,50,0,62,0,0,0,107,0,0,0,173,0,82,0,0,0,0,0,189,0,237,0,108,0,0,0,0,0,182,0,203,0,0,0,206,0,233,0,97,0,254,0,240,0,0,0,0,0,76,0,95,0,200,0,0,0,0,0,157,0,44,0,76,0,0,0,60,0,9,0,96,0,128,0,0,0,210,0,0,0,219,0,0,0,21,0,149,0,4,0,96,0,38,0,190,0,40,0,131,0,70,0,139,0,97,0,199,0,159,0,49,0,0,0,129,0,115,0,192,0,191,0,216,0,182,0,0,0,205,0,0,0,0,0,238,0,5,0,115,0,82,0,240,0,180,0,91,0,0,0,157,0,0,0,41,0,0,0,214,0,0,0,0,0,255,0,0,0,173,0,192,0,0,0,38,0,0,0,136,0,43,0,145,0,62,0,167,0,212,0,222,0,0,0,206,0,0,0,19,0,119,0,148,0,128,0,71,0,110,0,197,0,109,0,11,0,172,0,90,0,244,0,2,0,62,0,140,0,213,0,223,0,80,0,37,0,219,0,199,0,0,0,198,0,25,0,94,0,229,0,1,0,108,0,135,0,45,0,207,0,0,0,0,0,229,0,197,0,0,0,131,0,10,0,93,0,21,0,0,0,158,0,33,0,247,0,19,0,30,0,116,0,163,0,0,0,213,0,229,0,7,0,16,0,208,0,122,0,28,0,199,0,153,0,100,0,144,0,0,0,247,0,0,0,159,0,105,0,106,0,161,0,204,0,0,0,0,0,97,0,103,0,0,0,95,0,64,0,0,0,110,0,115,0,149,0,193,0,226,0,0,0,121,0,95,0,225,0,17,0,109,0,94,0,0,0,184,0,232,0,0,0,175,0,21,0,150,0,169,0,231,0,216,0,0,0,0,0,152,0,244,0,48,0,230,0,128,0,170,0,230,0,0,0,239,0,101,0,48,0,242,0,131,0,113,0,133,0,206,0,45,0,114,0,0,0,137,0,238,0,22,0,165,0,0,0,0,0,172,0,198,0,196,0,175,0,0,0,165,0,240,0,97,0,196,0,32,0,220,0,226,0,92,0,0,0,0,0,252,0,0,0,104,0,0,0,0,0,12,0,85,0,0,0,26,0,220,0,107,0,0,0,0,0,0,0,203,0,38,0,0,0,135,0,0,0,24,0,0,0,147,0,54,0,156,0,0,0,0,0,161,0,52,0,0,0,232,0,0,0,48,0,0,0,83,0,218,0,0,0,255,0,217,0,84,0,68,0,95,0,73,0,165,0,205,0,193,0,77,0,0,0,234,0,48,0,205,0,13,0,102,0,127,0,225,0,245,0,0,0,22,0,226,0,132,0,165,0,0,0,223,0,165,0,63,0,145,0,232,0,70,0,159,0,220,0,98,0,7,0,179,0,0,0,18,0,0,0,183,0,254,0,249,0,212,0,192,0,214,0,137,0,246,0,181,0,0,0,158,0,122,0,229,0,49,0,132,0,74,0,187,0,73,0,103,0,136,0,40,0,0,0,50,0,177,0,218,0,161,0,180,0,221,0,251,0,98,0,125,0,38,0,0,0,0,0,224,0,78,0,65,0,9,0,197,0,154,0,245,0,239,0,93,0,54,0,117,0,0,0,196,0,65,0,148,0,64,0,241,0,13,0,224,0,212,0,76,0,62,0,4,0,0,0,77,0,62,0,56,0,204,0,9,0,253,0,113,0,172,0,69,0,0,0,12,0,243,0,96,0,230,0,154,0,210,0,100,0,0,0,58,0,66,0,0,0,186,0,15,0,22,0,46,0,0,0,205,0,0,0,195,0,255,0,169,0,122,0,22,0,5,0,0,0,0,0,88,0,159,0,0,0,0,0,31,0,160,0,0,0,199,0,248,0,0,0,116,0,182,0,0,0,166,0,0,0,171,0,48,0,40,0,89,0,0,0,154,0,154,0,32,0,190,0,169,0,72,0,234,0,116,0,112,0,176,0,51,0,242,0,65,0,0,0,84,0,0,0,84,0,212,0,0,0,243,0,85,0,0,0,4,0,90,0,115,0,92,0,0,0,72,0,171,0,34,0,128,0,195,0,21,0,65,0,0,0,249,0,70,0,230,0,125,0,91,0,212,0,253,0,137,0,38,0,236,0,112,0,121,0,63,0,0,0,78,0,183,0,217,0,69,0,154,0,119,0,229,0,70,0,121,0,166,0,0,0,207,0,83,0,0,0,134,0,0,0,139,0,147,0,121,0,79,0,108,0,211,0,59,0,183,0,5,0,120,0,224,0,5,0,154,0,70,0,165,0,0,0,251,0,0,0,86,0,198,0,61,0,140,0,103,0,37,0,92,0,151,0,166,0,112,0,7,0,202,0,163,0,0,0,0,0,124,0,131,0,196,0,21,0,231,0,233,0,85,0,210,0,59,0,122,0,186,0,210,0,0,0,0,0,0,0,211,0,157,0,0,0,142,0,0,0,110,0,186,0,232,0,46,0,42,0,95,0,143,0,148,0,0,0,0,0,67,0,59,0,48,0,153,0,84,0,0,0,240,0,232,0,143,0,213,0,82,0,175,0,11,0,139,0,248,0,173,0,169,0,0,0,201,0,44,0,0,0,0,0,147,0,0,0,34,0,96,0,0,0,0,0,37,0,208,0,92,0,0,0,0,0,71,0,48,0,0,0,149,0,135,0,250,0,245,0,21,0,0,0,88,0,0,0,118,0,70,0,81,0,8,0,18,0,113,0,78,0,169,0,84,0,229,0,0,0,237,0,77,0,78,0,199,0,120,0,127,0,0,0,140,0,40,0,223,0,170,0,184,0,8,0,0,0,177,0,45,0,150,0,95,0,0,0,158,0,85,0,139,0,89,0,113,0,162,0,0,0,0,0,252,0,39,0,202,0,71,0,111,0,104,0,0,0,0,0,0,0,141,0,65,0,193,0,12,0,0,0,142,0,246,0,68,0,168,0,149,0,84,0,10,0,78,0,168,0,40,0,0,0,83,0,136,0,236,0,43,0,0,0,53,0,179,0,212,0,37,0,112,0,55,0,0,0,12,0,0,0,39,0,182,0,75,0,228,0,154,0,236,0,0,0,0,0,188,0);
signal scenario_full  : scenario_type := (155,31,209,31,191,31,240,31,77,31,96,31,96,31,96,30,89,31,89,30,154,31,113,31,78,31,44,31,149,31,9,31,9,30,9,29,9,28,188,31,245,31,74,31,80,31,42,31,249,31,181,31,181,30,65,31,87,31,82,31,253,31,113,31,108,31,108,30,225,31,225,30,161,31,103,31,247,31,242,31,242,30,61,31,61,30,156,31,80,31,247,31,85,31,29,31,119,31,119,30,78,31,78,30,78,29,128,31,251,31,251,30,225,31,245,31,245,30,29,31,71,31,167,31,39,31,244,31,129,31,60,31,217,31,213,31,213,30,252,31,136,31,136,30,7,31,203,31,199,31,199,30,200,31,94,31,73,31,238,31,189,31,11,31,11,30,11,29,213,31,213,30,168,31,152,31,109,31,83,31,107,31,34,31,34,30,88,31,218,31,174,31,161,31,131,31,72,31,132,31,249,31,162,31,81,31,58,31,114,31,51,31,172,31,245,31,245,30,245,29,193,31,102,31,37,31,37,30,38,31,177,31,12,31,159,31,245,31,27,31,27,30,90,31,91,31,91,30,170,31,254,31,254,30,221,31,23,31,147,31,232,31,122,31,152,31,183,31,33,31,76,31,76,30,186,31,37,31,37,30,210,31,120,31,217,31,162,31,185,31,36,31,97,31,103,31,103,30,138,31,138,30,144,31,217,31,217,30,60,31,87,31,87,30,166,31,25,31,203,31,40,31,129,31,129,30,47,31,22,31,156,31,60,31,234,31,173,31,53,31,253,31,160,31,106,31,188,31,161,31,186,31,128,31,188,31,29,31,50,31,62,31,62,30,107,31,107,30,173,31,82,31,82,30,82,29,189,31,237,31,108,31,108,30,108,29,182,31,203,31,203,30,206,31,233,31,97,31,254,31,240,31,240,30,240,29,76,31,95,31,200,31,200,30,200,29,157,31,44,31,76,31,76,30,60,31,9,31,96,31,128,31,128,30,210,31,210,30,219,31,219,30,21,31,149,31,4,31,96,31,38,31,190,31,40,31,131,31,70,31,139,31,97,31,199,31,159,31,49,31,49,30,129,31,115,31,192,31,191,31,216,31,182,31,182,30,205,31,205,30,205,29,238,31,5,31,115,31,82,31,240,31,180,31,91,31,91,30,157,31,157,30,41,31,41,30,214,31,214,30,214,29,255,31,255,30,173,31,192,31,192,30,38,31,38,30,136,31,43,31,145,31,62,31,167,31,212,31,222,31,222,30,206,31,206,30,19,31,119,31,148,31,128,31,71,31,110,31,197,31,109,31,11,31,172,31,90,31,244,31,2,31,62,31,140,31,213,31,223,31,80,31,37,31,219,31,199,31,199,30,198,31,25,31,94,31,229,31,1,31,108,31,135,31,45,31,207,31,207,30,207,29,229,31,197,31,197,30,131,31,10,31,93,31,21,31,21,30,158,31,33,31,247,31,19,31,30,31,116,31,163,31,163,30,213,31,229,31,7,31,16,31,208,31,122,31,28,31,199,31,153,31,100,31,144,31,144,30,247,31,247,30,159,31,105,31,106,31,161,31,204,31,204,30,204,29,97,31,103,31,103,30,95,31,64,31,64,30,110,31,115,31,149,31,193,31,226,31,226,30,121,31,95,31,225,31,17,31,109,31,94,31,94,30,184,31,232,31,232,30,175,31,21,31,150,31,169,31,231,31,216,31,216,30,216,29,152,31,244,31,48,31,230,31,128,31,170,31,230,31,230,30,239,31,101,31,48,31,242,31,131,31,113,31,133,31,206,31,45,31,114,31,114,30,137,31,238,31,22,31,165,31,165,30,165,29,172,31,198,31,196,31,175,31,175,30,165,31,240,31,97,31,196,31,32,31,220,31,226,31,92,31,92,30,92,29,252,31,252,30,104,31,104,30,104,29,12,31,85,31,85,30,26,31,220,31,107,31,107,30,107,29,107,28,203,31,38,31,38,30,135,31,135,30,24,31,24,30,147,31,54,31,156,31,156,30,156,29,161,31,52,31,52,30,232,31,232,30,48,31,48,30,83,31,218,31,218,30,255,31,217,31,84,31,68,31,95,31,73,31,165,31,205,31,193,31,77,31,77,30,234,31,48,31,205,31,13,31,102,31,127,31,225,31,245,31,245,30,22,31,226,31,132,31,165,31,165,30,223,31,165,31,63,31,145,31,232,31,70,31,159,31,220,31,98,31,7,31,179,31,179,30,18,31,18,30,183,31,254,31,249,31,212,31,192,31,214,31,137,31,246,31,181,31,181,30,158,31,122,31,229,31,49,31,132,31,74,31,187,31,73,31,103,31,136,31,40,31,40,30,50,31,177,31,218,31,161,31,180,31,221,31,251,31,98,31,125,31,38,31,38,30,38,29,224,31,78,31,65,31,9,31,197,31,154,31,245,31,239,31,93,31,54,31,117,31,117,30,196,31,65,31,148,31,64,31,241,31,13,31,224,31,212,31,76,31,62,31,4,31,4,30,77,31,62,31,56,31,204,31,9,31,253,31,113,31,172,31,69,31,69,30,12,31,243,31,96,31,230,31,154,31,210,31,100,31,100,30,58,31,66,31,66,30,186,31,15,31,22,31,46,31,46,30,205,31,205,30,195,31,255,31,169,31,122,31,22,31,5,31,5,30,5,29,88,31,159,31,159,30,159,29,31,31,160,31,160,30,199,31,248,31,248,30,116,31,182,31,182,30,166,31,166,30,171,31,48,31,40,31,89,31,89,30,154,31,154,31,32,31,190,31,169,31,72,31,234,31,116,31,112,31,176,31,51,31,242,31,65,31,65,30,84,31,84,30,84,31,212,31,212,30,243,31,85,31,85,30,4,31,90,31,115,31,92,31,92,30,72,31,171,31,34,31,128,31,195,31,21,31,65,31,65,30,249,31,70,31,230,31,125,31,91,31,212,31,253,31,137,31,38,31,236,31,112,31,121,31,63,31,63,30,78,31,183,31,217,31,69,31,154,31,119,31,229,31,70,31,121,31,166,31,166,30,207,31,83,31,83,30,134,31,134,30,139,31,147,31,121,31,79,31,108,31,211,31,59,31,183,31,5,31,120,31,224,31,5,31,154,31,70,31,165,31,165,30,251,31,251,30,86,31,198,31,61,31,140,31,103,31,37,31,92,31,151,31,166,31,112,31,7,31,202,31,163,31,163,30,163,29,124,31,131,31,196,31,21,31,231,31,233,31,85,31,210,31,59,31,122,31,186,31,210,31,210,30,210,29,210,28,211,31,157,31,157,30,142,31,142,30,110,31,186,31,232,31,46,31,42,31,95,31,143,31,148,31,148,30,148,29,67,31,59,31,48,31,153,31,84,31,84,30,240,31,232,31,143,31,213,31,82,31,175,31,11,31,139,31,248,31,173,31,169,31,169,30,201,31,44,31,44,30,44,29,147,31,147,30,34,31,96,31,96,30,96,29,37,31,208,31,92,31,92,30,92,29,71,31,48,31,48,30,149,31,135,31,250,31,245,31,21,31,21,30,88,31,88,30,118,31,70,31,81,31,8,31,18,31,113,31,78,31,169,31,84,31,229,31,229,30,237,31,77,31,78,31,199,31,120,31,127,31,127,30,140,31,40,31,223,31,170,31,184,31,8,31,8,30,177,31,45,31,150,31,95,31,95,30,158,31,85,31,139,31,89,31,113,31,162,31,162,30,162,29,252,31,39,31,202,31,71,31,111,31,104,31,104,30,104,29,104,28,141,31,65,31,193,31,12,31,12,30,142,31,246,31,68,31,168,31,149,31,84,31,10,31,78,31,168,31,40,31,40,30,83,31,136,31,236,31,43,31,43,30,53,31,179,31,212,31,37,31,112,31,55,31,55,30,12,31,12,30,39,31,182,31,75,31,228,31,154,31,236,31,236,30,236,29,188,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
