-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 867;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,173,0,56,0,67,0,100,0,247,0,72,0,212,0,120,0,243,0,10,0,195,0,4,0,59,0,200,0,0,0,124,0,0,0,98,0,0,0,249,0,64,0,176,0,214,0,83,0,40,0,137,0,10,0,38,0,153,0,2,0,0,0,3,0,73,0,101,0,154,0,5,0,52,0,213,0,0,0,222,0,240,0,207,0,54,0,190,0,0,0,208,0,207,0,65,0,234,0,0,0,198,0,73,0,25,0,68,0,89,0,135,0,254,0,42,0,189,0,0,0,39,0,0,0,251,0,55,0,255,0,45,0,0,0,107,0,189,0,154,0,78,0,154,0,194,0,230,0,157,0,242,0,29,0,101,0,0,0,139,0,170,0,170,0,149,0,139,0,129,0,197,0,93,0,0,0,0,0,19,0,240,0,0,0,208,0,247,0,0,0,66,0,137,0,75,0,167,0,145,0,199,0,192,0,187,0,0,0,123,0,230,0,0,0,199,0,214,0,189,0,49,0,114,0,142,0,96,0,59,0,34,0,62,0,138,0,136,0,234,0,27,0,42,0,159,0,85,0,207,0,9,0,149,0,236,0,167,0,33,0,28,0,173,0,131,0,43,0,243,0,48,0,0,0,0,0,243,0,0,0,200,0,54,0,93,0,153,0,10,0,146,0,0,0,0,0,28,0,220,0,243,0,0,0,0,0,208,0,201,0,201,0,141,0,0,0,143,0,0,0,91,0,0,0,104,0,69,0,71,0,39,0,0,0,200,0,16,0,56,0,56,0,221,0,62,0,226,0,74,0,0,0,97,0,197,0,75,0,250,0,31,0,162,0,0,0,149,0,127,0,78,0,116,0,176,0,201,0,174,0,8,0,78,0,48,0,13,0,139,0,252,0,0,0,69,0,93,0,0,0,0,0,43,0,62,0,164,0,114,0,113,0,68,0,107,0,160,0,0,0,18,0,0,0,88,0,0,0,138,0,0,0,117,0,117,0,5,0,237,0,254,0,37,0,137,0,44,0,0,0,0,0,233,0,18,0,59,0,151,0,92,0,251,0,183,0,28,0,170,0,18,0,137,0,0,0,196,0,208,0,51,0,59,0,218,0,120,0,113,0,13,0,146,0,71,0,247,0,42,0,0,0,0,0,159,0,95,0,99,0,228,0,20,0,0,0,166,0,78,0,111,0,242,0,5,0,42,0,127,0,183,0,92,0,231,0,0,0,0,0,179,0,61,0,0,0,0,0,160,0,136,0,13,0,248,0,0,0,67,0,126,0,0,0,104,0,0,0,104,0,0,0,45,0,166,0,0,0,0,0,226,0,152,0,131,0,0,0,107,0,40,0,135,0,202,0,208,0,249,0,0,0,240,0,0,0,166,0,125,0,0,0,0,0,252,0,173,0,172,0,192,0,210,0,110,0,122,0,34,0,110,0,134,0,0,0,68,0,0,0,188,0,216,0,104,0,236,0,0,0,247,0,0,0,47,0,185,0,0,0,68,0,0,0,205,0,195,0,84,0,124,0,66,0,107,0,150,0,159,0,42,0,0,0,90,0,243,0,141,0,228,0,225,0,0,0,211,0,0,0,0,0,0,0,0,0,15,0,193,0,0,0,184,0,38,0,212,0,56,0,230,0,194,0,117,0,0,0,185,0,0,0,32,0,12,0,251,0,0,0,199,0,0,0,78,0,0,0,25,0,0,0,224,0,207,0,29,0,0,0,71,0,0,0,83,0,165,0,144,0,219,0,0,0,131,0,76,0,0,0,97,0,213,0,211,0,0,0,62,0,16,0,219,0,0,0,251,0,94,0,89,0,130,0,33,0,212,0,215,0,219,0,89,0,93,0,214,0,0,0,128,0,136,0,8,0,18,0,72,0,57,0,147,0,207,0,73,0,178,0,234,0,42,0,0,0,64,0,37,0,132,0,0,0,130,0,134,0,194,0,24,0,0,0,154,0,94,0,182,0,108,0,175,0,0,0,48,0,53,0,126,0,85,0,81,0,50,0,28,0,0,0,73,0,204,0,0,0,60,0,28,0,87,0,107,0,36,0,0,0,16,0,169,0,237,0,252,0,0,0,118,0,0,0,0,0,73,0,34,0,195,0,164,0,94,0,75,0,6,0,180,0,0,0,177,0,0,0,54,0,200,0,0,0,195,0,213,0,101,0,0,0,87,0,64,0,248,0,112,0,254,0,0,0,0,0,66,0,159,0,228,0,220,0,94,0,194,0,25,0,14,0,251,0,108,0,5,0,0,0,120,0,100,0,245,0,0,0,58,0,92,0,0,0,0,0,242,0,121,0,168,0,118,0,249,0,50,0,0,0,3,0,112,0,99,0,0,0,0,0,55,0,1,0,0,0,248,0,83,0,237,0,151,0,70,0,8,0,140,0,186,0,119,0,11,0,129,0,223,0,162,0,59,0,106,0,73,0,0,0,116,0,150,0,235,0,0,0,206,0,0,0,128,0,236,0,194,0,136,0,122,0,2,0,113,0,0,0,0,0,98,0,169,0,0,0,19,0,30,0,68,0,60,0,0,0,136,0,145,0,52,0,67,0,65,0,170,0,0,0,166,0,93,0,200,0,211,0,0,0,27,0,7,0,110,0,224,0,28,0,22,0,186,0,161,0,14,0,78,0,0,0,137,0,8,0,0,0,255,0,224,0,0,0,131,0,120,0,75,0,102,0,159,0,90,0,114,0,98,0,0,0,0,0,80,0,245,0,0,0,174,0,207,0,0,0,86,0,22,0,59,0,119,0,122,0,216,0,109,0,24,0,242,0,105,0,180,0,255,0,122,0,106,0,39,0,121,0,195,0,3,0,223,0,142,0,91,0,0,0,0,0,0,0,36,0,162,0,242,0,234,0,23,0,119,0,205,0,0,0,0,0,109,0,226,0,4,0,202,0,0,0,166,0,224,0,0,0,0,0,132,0,65,0,13,0,188,0,240,0,0,0,236,0,23,0,192,0,0,0,138,0,0,0,106,0,226,0,224,0,118,0,94,0,255,0,0,0,93,0,178,0,246,0,119,0,190,0,218,0,108,0,33,0,0,0,141,0,181,0,67,0,195,0,162,0,249,0,236,0,0,0,50,0,75,0,109,0,0,0,189,0,188,0,144,0,0,0,66,0,200,0,254,0,55,0,0,0,116,0,160,0,226,0,61,0,181,0,51,0,30,0,0,0,94,0,41,0,229,0,226,0,0,0,0,0,129,0,14,0,209,0,0,0,0,0,24,0,0,0,0,0,214,0,0,0,131,0,82,0,151,0,112,0,20,0,219,0,90,0,0,0,140,0,173,0,117,0,243,0,62,0,144,0,42,0,0,0,90,0,0,0,122,0,223,0,0,0,48,0,142,0,58,0,240,0,79,0,235,0,0,0,138,0,228,0,130,0,247,0,156,0,129,0,97,0,89,0,21,0,90,0,29,0,137,0,0,0,204,0,69,0,234,0,208,0,240,0,238,0,43,0,0,0,86,0,149,0,57,0,196,0,223,0,99,0,171,0,132,0,0,0,52,0,79,0,197,0,76,0,0,0,0,0,25,0,0,0,240,0,0,0,0,0,112,0,14,0,196,0,0,0,61,0,0,0,222,0,86,0,181,0,156,0,119,0,100,0,91,0,17,0,38,0,55,0,168,0,130,0,169,0,206,0,2,0,0,0,0,0,39,0,0,0,0,0,10,0,35,0,0,0,136,0,85,0,8,0,95,0,106,0,120,0,195,0,140,0,181,0,128,0,239,0,239,0,87,0,0,0,92,0,251,0,0,0,196,0,24,0,0,0,229,0,0,0,139,0,141,0,214,0,158,0,110,0,155,0,87,0,116,0,47,0,187,0,0,0,0,0,41,0,124,0,219,0,135,0,155,0,195,0,68,0,0,0,216,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,173,31,56,31,67,31,100,31,247,31,72,31,212,31,120,31,243,31,10,31,195,31,4,31,59,31,200,31,200,30,124,31,124,30,98,31,98,30,249,31,64,31,176,31,214,31,83,31,40,31,137,31,10,31,38,31,153,31,2,31,2,30,3,31,73,31,101,31,154,31,5,31,52,31,213,31,213,30,222,31,240,31,207,31,54,31,190,31,190,30,208,31,207,31,65,31,234,31,234,30,198,31,73,31,25,31,68,31,89,31,135,31,254,31,42,31,189,31,189,30,39,31,39,30,251,31,55,31,255,31,45,31,45,30,107,31,189,31,154,31,78,31,154,31,194,31,230,31,157,31,242,31,29,31,101,31,101,30,139,31,170,31,170,31,149,31,139,31,129,31,197,31,93,31,93,30,93,29,19,31,240,31,240,30,208,31,247,31,247,30,66,31,137,31,75,31,167,31,145,31,199,31,192,31,187,31,187,30,123,31,230,31,230,30,199,31,214,31,189,31,49,31,114,31,142,31,96,31,59,31,34,31,62,31,138,31,136,31,234,31,27,31,42,31,159,31,85,31,207,31,9,31,149,31,236,31,167,31,33,31,28,31,173,31,131,31,43,31,243,31,48,31,48,30,48,29,243,31,243,30,200,31,54,31,93,31,153,31,10,31,146,31,146,30,146,29,28,31,220,31,243,31,243,30,243,29,208,31,201,31,201,31,141,31,141,30,143,31,143,30,91,31,91,30,104,31,69,31,71,31,39,31,39,30,200,31,16,31,56,31,56,31,221,31,62,31,226,31,74,31,74,30,97,31,197,31,75,31,250,31,31,31,162,31,162,30,149,31,127,31,78,31,116,31,176,31,201,31,174,31,8,31,78,31,48,31,13,31,139,31,252,31,252,30,69,31,93,31,93,30,93,29,43,31,62,31,164,31,114,31,113,31,68,31,107,31,160,31,160,30,18,31,18,30,88,31,88,30,138,31,138,30,117,31,117,31,5,31,237,31,254,31,37,31,137,31,44,31,44,30,44,29,233,31,18,31,59,31,151,31,92,31,251,31,183,31,28,31,170,31,18,31,137,31,137,30,196,31,208,31,51,31,59,31,218,31,120,31,113,31,13,31,146,31,71,31,247,31,42,31,42,30,42,29,159,31,95,31,99,31,228,31,20,31,20,30,166,31,78,31,111,31,242,31,5,31,42,31,127,31,183,31,92,31,231,31,231,30,231,29,179,31,61,31,61,30,61,29,160,31,136,31,13,31,248,31,248,30,67,31,126,31,126,30,104,31,104,30,104,31,104,30,45,31,166,31,166,30,166,29,226,31,152,31,131,31,131,30,107,31,40,31,135,31,202,31,208,31,249,31,249,30,240,31,240,30,166,31,125,31,125,30,125,29,252,31,173,31,172,31,192,31,210,31,110,31,122,31,34,31,110,31,134,31,134,30,68,31,68,30,188,31,216,31,104,31,236,31,236,30,247,31,247,30,47,31,185,31,185,30,68,31,68,30,205,31,195,31,84,31,124,31,66,31,107,31,150,31,159,31,42,31,42,30,90,31,243,31,141,31,228,31,225,31,225,30,211,31,211,30,211,29,211,28,211,27,15,31,193,31,193,30,184,31,38,31,212,31,56,31,230,31,194,31,117,31,117,30,185,31,185,30,32,31,12,31,251,31,251,30,199,31,199,30,78,31,78,30,25,31,25,30,224,31,207,31,29,31,29,30,71,31,71,30,83,31,165,31,144,31,219,31,219,30,131,31,76,31,76,30,97,31,213,31,211,31,211,30,62,31,16,31,219,31,219,30,251,31,94,31,89,31,130,31,33,31,212,31,215,31,219,31,89,31,93,31,214,31,214,30,128,31,136,31,8,31,18,31,72,31,57,31,147,31,207,31,73,31,178,31,234,31,42,31,42,30,64,31,37,31,132,31,132,30,130,31,134,31,194,31,24,31,24,30,154,31,94,31,182,31,108,31,175,31,175,30,48,31,53,31,126,31,85,31,81,31,50,31,28,31,28,30,73,31,204,31,204,30,60,31,28,31,87,31,107,31,36,31,36,30,16,31,169,31,237,31,252,31,252,30,118,31,118,30,118,29,73,31,34,31,195,31,164,31,94,31,75,31,6,31,180,31,180,30,177,31,177,30,54,31,200,31,200,30,195,31,213,31,101,31,101,30,87,31,64,31,248,31,112,31,254,31,254,30,254,29,66,31,159,31,228,31,220,31,94,31,194,31,25,31,14,31,251,31,108,31,5,31,5,30,120,31,100,31,245,31,245,30,58,31,92,31,92,30,92,29,242,31,121,31,168,31,118,31,249,31,50,31,50,30,3,31,112,31,99,31,99,30,99,29,55,31,1,31,1,30,248,31,83,31,237,31,151,31,70,31,8,31,140,31,186,31,119,31,11,31,129,31,223,31,162,31,59,31,106,31,73,31,73,30,116,31,150,31,235,31,235,30,206,31,206,30,128,31,236,31,194,31,136,31,122,31,2,31,113,31,113,30,113,29,98,31,169,31,169,30,19,31,30,31,68,31,60,31,60,30,136,31,145,31,52,31,67,31,65,31,170,31,170,30,166,31,93,31,200,31,211,31,211,30,27,31,7,31,110,31,224,31,28,31,22,31,186,31,161,31,14,31,78,31,78,30,137,31,8,31,8,30,255,31,224,31,224,30,131,31,120,31,75,31,102,31,159,31,90,31,114,31,98,31,98,30,98,29,80,31,245,31,245,30,174,31,207,31,207,30,86,31,22,31,59,31,119,31,122,31,216,31,109,31,24,31,242,31,105,31,180,31,255,31,122,31,106,31,39,31,121,31,195,31,3,31,223,31,142,31,91,31,91,30,91,29,91,28,36,31,162,31,242,31,234,31,23,31,119,31,205,31,205,30,205,29,109,31,226,31,4,31,202,31,202,30,166,31,224,31,224,30,224,29,132,31,65,31,13,31,188,31,240,31,240,30,236,31,23,31,192,31,192,30,138,31,138,30,106,31,226,31,224,31,118,31,94,31,255,31,255,30,93,31,178,31,246,31,119,31,190,31,218,31,108,31,33,31,33,30,141,31,181,31,67,31,195,31,162,31,249,31,236,31,236,30,50,31,75,31,109,31,109,30,189,31,188,31,144,31,144,30,66,31,200,31,254,31,55,31,55,30,116,31,160,31,226,31,61,31,181,31,51,31,30,31,30,30,94,31,41,31,229,31,226,31,226,30,226,29,129,31,14,31,209,31,209,30,209,29,24,31,24,30,24,29,214,31,214,30,131,31,82,31,151,31,112,31,20,31,219,31,90,31,90,30,140,31,173,31,117,31,243,31,62,31,144,31,42,31,42,30,90,31,90,30,122,31,223,31,223,30,48,31,142,31,58,31,240,31,79,31,235,31,235,30,138,31,228,31,130,31,247,31,156,31,129,31,97,31,89,31,21,31,90,31,29,31,137,31,137,30,204,31,69,31,234,31,208,31,240,31,238,31,43,31,43,30,86,31,149,31,57,31,196,31,223,31,99,31,171,31,132,31,132,30,52,31,79,31,197,31,76,31,76,30,76,29,25,31,25,30,240,31,240,30,240,29,112,31,14,31,196,31,196,30,61,31,61,30,222,31,86,31,181,31,156,31,119,31,100,31,91,31,17,31,38,31,55,31,168,31,130,31,169,31,206,31,2,31,2,30,2,29,39,31,39,30,39,29,10,31,35,31,35,30,136,31,85,31,8,31,95,31,106,31,120,31,195,31,140,31,181,31,128,31,239,31,239,31,87,31,87,30,92,31,251,31,251,30,196,31,24,31,24,30,229,31,229,30,139,31,141,31,214,31,158,31,110,31,155,31,87,31,116,31,47,31,187,31,187,30,187,29,41,31,124,31,219,31,135,31,155,31,195,31,68,31,68,30,216,31,216,30,216,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
