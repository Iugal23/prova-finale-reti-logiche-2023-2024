-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_867 is
end project_tb_867;

architecture project_tb_arch_867 of project_tb_867 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 820;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,221,0,7,0,18,0,105,0,226,0,43,0,211,0,84,0,128,0,0,0,28,0,194,0,131,0,85,0,124,0,159,0,111,0,206,0,243,0,80,0,24,0,195,0,0,0,218,0,0,0,226,0,71,0,0,0,240,0,0,0,245,0,232,0,137,0,205,0,246,0,220,0,116,0,0,0,232,0,50,0,121,0,228,0,119,0,3,0,49,0,0,0,150,0,131,0,234,0,108,0,245,0,218,0,0,0,21,0,164,0,105,0,235,0,100,0,152,0,0,0,0,0,177,0,75,0,205,0,0,0,168,0,205,0,212,0,208,0,238,0,0,0,200,0,31,0,131,0,79,0,0,0,102,0,72,0,63,0,0,0,0,0,27,0,254,0,106,0,19,0,127,0,195,0,0,0,0,0,0,0,119,0,252,0,69,0,0,0,170,0,144,0,0,0,0,0,90,0,0,0,0,0,7,0,248,0,191,0,0,0,228,0,177,0,92,0,217,0,7,0,202,0,104,0,0,0,0,0,157,0,0,0,88,0,131,0,0,0,31,0,217,0,10,0,224,0,43,0,116,0,0,0,28,0,11,0,72,0,170,0,0,0,0,0,77,0,105,0,86,0,216,0,185,0,207,0,0,0,178,0,7,0,60,0,0,0,124,0,0,0,79,0,241,0,255,0,12,0,0,0,0,0,30,0,0,0,225,0,209,0,166,0,191,0,79,0,0,0,28,0,152,0,45,0,26,0,141,0,120,0,0,0,8,0,230,0,53,0,198,0,167,0,0,0,97,0,81,0,134,0,0,0,48,0,246,0,163,0,203,0,112,0,137,0,62,0,53,0,0,0,58,0,153,0,147,0,137,0,214,0,229,0,241,0,226,0,205,0,79,0,0,0,104,0,196,0,31,0,36,0,220,0,181,0,28,0,129,0,0,0,183,0,64,0,4,0,218,0,0,0,0,0,0,0,77,0,195,0,115,0,28,0,185,0,58,0,176,0,141,0,65,0,141,0,5,0,0,0,92,0,45,0,146,0,0,0,76,0,238,0,157,0,121,0,126,0,153,0,0,0,82,0,13,0,172,0,34,0,20,0,79,0,18,0,42,0,94,0,112,0,184,0,0,0,153,0,0,0,0,0,198,0,121,0,23,0,209,0,93,0,138,0,24,0,184,0,179,0,77,0,122,0,0,0,225,0,125,0,226,0,33,0,214,0,81,0,73,0,0,0,0,0,65,0,165,0,0,0,78,0,1,0,141,0,130,0,109,0,201,0,227,0,9,0,58,0,82,0,218,0,195,0,154,0,189,0,126,0,110,0,62,0,119,0,0,0,206,0,0,0,28,0,28,0,0,0,0,0,199,0,28,0,86,0,115,0,4,0,119,0,0,0,0,0,63,0,31,0,0,0,0,0,175,0,0,0,67,0,144,0,0,0,172,0,222,0,8,0,148,0,0,0,221,0,146,0,120,0,88,0,94,0,80,0,127,0,144,0,239,0,118,0,89,0,198,0,172,0,46,0,123,0,55,0,7,0,149,0,62,0,24,0,0,0,43,0,33,0,0,0,115,0,217,0,206,0,186,0,14,0,254,0,147,0,154,0,141,0,134,0,24,0,187,0,0,0,55,0,155,0,186,0,107,0,123,0,61,0,207,0,7,0,130,0,10,0,114,0,138,0,0,0,16,0,104,0,1,0,153,0,182,0,0,0,0,0,66,0,243,0,0,0,151,0,118,0,143,0,176,0,93,0,169,0,154,0,113,0,161,0,2,0,134,0,194,0,218,0,0,0,0,0,227,0,0,0,215,0,0,0,0,0,49,0,96,0,12,0,219,0,0,0,226,0,93,0,216,0,240,0,0,0,142,0,195,0,173,0,108,0,48,0,20,0,167,0,0,0,154,0,63,0,132,0,123,0,248,0,19,0,0,0,153,0,154,0,61,0,106,0,0,0,212,0,68,0,200,0,56,0,233,0,185,0,177,0,187,0,0,0,16,0,140,0,164,0,3,0,70,0,82,0,0,0,221,0,52,0,208,0,114,0,201,0,203,0,191,0,225,0,75,0,69,0,128,0,0,0,0,0,189,0,0,0,247,0,68,0,75,0,180,0,0,0,154,0,221,0,26,0,16,0,8,0,228,0,243,0,0,0,200,0,71,0,152,0,115,0,175,0,238,0,224,0,136,0,60,0,146,0,231,0,32,0,0,0,10,0,219,0,233,0,0,0,126,0,0,0,194,0,125,0,170,0,118,0,0,0,7,0,1,0,0,0,94,0,255,0,39,0,182,0,0,0,0,0,28,0,0,0,196,0,124,0,147,0,191,0,0,0,224,0,185,0,0,0,61,0,187,0,0,0,17,0,19,0,221,0,144,0,62,0,226,0,0,0,117,0,78,0,0,0,239,0,248,0,112,0,21,0,80,0,186,0,21,0,212,0,176,0,228,0,246,0,93,0,78,0,238,0,214,0,68,0,0,0,82,0,108,0,0,0,0,0,125,0,47,0,0,0,82,0,0,0,207,0,60,0,42,0,0,0,83,0,0,0,0,0,0,0,100,0,151,0,165,0,0,0,167,0,56,0,0,0,193,0,0,0,91,0,36,0,0,0,242,0,30,0,10,0,202,0,171,0,102,0,0,0,31,0,0,0,162,0,235,0,223,0,243,0,193,0,0,0,199,0,1,0,16,0,27,0,0,0,0,0,233,0,85,0,145,0,71,0,68,0,245,0,79,0,184,0,236,0,43,0,60,0,228,0,0,0,190,0,230,0,181,0,175,0,89,0,100,0,25,0,101,0,164,0,0,0,124,0,224,0,8,0,245,0,105,0,125,0,109,0,0,0,170,0,84,0,153,0,47,0,194,0,99,0,175,0,95,0,221,0,133,0,151,0,110,0,125,0,250,0,61,0,178,0,121,0,40,0,0,0,28,0,231,0,77,0,98,0,120,0,76,0,97,0,9,0,203,0,157,0,211,0,202,0,0,0,100,0,57,0,137,0,117,0,32,0,0,0,125,0,158,0,222,0,69,0,156,0,202,0,236,0,74,0,0,0,53,0,122,0,120,0,66,0,10,0,251,0,172,0,63,0,181,0,0,0,47,0,41,0,175,0,14,0,97,0,104,0,147,0,36,0,91,0,202,0,148,0,63,0,205,0,0,0,241,0,122,0,224,0,0,0,0,0,73,0,170,0,202,0,172,0,0,0,27,0,139,0,210,0,98,0,144,0,23,0,55,0,159,0,43,0,244,0,0,0,0,0,159,0,0,0,163,0,180,0,188,0,185,0,98,0,0,0,0,0,0,0,245,0,250,0,133,0,0,0,111,0,214,0,171,0,47,0,86,0,71,0,87,0,0,0,247,0,54,0,96,0,52,0,0,0,177,0,0,0,118,0,0,0,167,0,122,0,142,0,29,0,200,0,0,0,245,0,189,0,39,0,115,0,145,0,136,0,184,0,208,0,232,0,0,0,24,0,123,0,70,0,181,0,215,0,150,0,175,0,16,0,247,0,78,0,44,0,66,0,147,0,178,0,248,0,82,0,59,0,89,0,64,0,59,0,163,0,80,0,88,0,0,0,152,0,0,0,27,0,0,0,176,0,87,0,173,0,0,0,52,0,236,0,49,0,0,0,7,0,0,0,0,0,112,0,0,0,0,0,0,0,48,0,7,0,65,0,82,0,1,0,0,0,241,0);
signal scenario_full  : scenario_type := (0,0,221,31,7,31,18,31,105,31,226,31,43,31,211,31,84,31,128,31,128,30,28,31,194,31,131,31,85,31,124,31,159,31,111,31,206,31,243,31,80,31,24,31,195,31,195,30,218,31,218,30,226,31,71,31,71,30,240,31,240,30,245,31,232,31,137,31,205,31,246,31,220,31,116,31,116,30,232,31,50,31,121,31,228,31,119,31,3,31,49,31,49,30,150,31,131,31,234,31,108,31,245,31,218,31,218,30,21,31,164,31,105,31,235,31,100,31,152,31,152,30,152,29,177,31,75,31,205,31,205,30,168,31,205,31,212,31,208,31,238,31,238,30,200,31,31,31,131,31,79,31,79,30,102,31,72,31,63,31,63,30,63,29,27,31,254,31,106,31,19,31,127,31,195,31,195,30,195,29,195,28,119,31,252,31,69,31,69,30,170,31,144,31,144,30,144,29,90,31,90,30,90,29,7,31,248,31,191,31,191,30,228,31,177,31,92,31,217,31,7,31,202,31,104,31,104,30,104,29,157,31,157,30,88,31,131,31,131,30,31,31,217,31,10,31,224,31,43,31,116,31,116,30,28,31,11,31,72,31,170,31,170,30,170,29,77,31,105,31,86,31,216,31,185,31,207,31,207,30,178,31,7,31,60,31,60,30,124,31,124,30,79,31,241,31,255,31,12,31,12,30,12,29,30,31,30,30,225,31,209,31,166,31,191,31,79,31,79,30,28,31,152,31,45,31,26,31,141,31,120,31,120,30,8,31,230,31,53,31,198,31,167,31,167,30,97,31,81,31,134,31,134,30,48,31,246,31,163,31,203,31,112,31,137,31,62,31,53,31,53,30,58,31,153,31,147,31,137,31,214,31,229,31,241,31,226,31,205,31,79,31,79,30,104,31,196,31,31,31,36,31,220,31,181,31,28,31,129,31,129,30,183,31,64,31,4,31,218,31,218,30,218,29,218,28,77,31,195,31,115,31,28,31,185,31,58,31,176,31,141,31,65,31,141,31,5,31,5,30,92,31,45,31,146,31,146,30,76,31,238,31,157,31,121,31,126,31,153,31,153,30,82,31,13,31,172,31,34,31,20,31,79,31,18,31,42,31,94,31,112,31,184,31,184,30,153,31,153,30,153,29,198,31,121,31,23,31,209,31,93,31,138,31,24,31,184,31,179,31,77,31,122,31,122,30,225,31,125,31,226,31,33,31,214,31,81,31,73,31,73,30,73,29,65,31,165,31,165,30,78,31,1,31,141,31,130,31,109,31,201,31,227,31,9,31,58,31,82,31,218,31,195,31,154,31,189,31,126,31,110,31,62,31,119,31,119,30,206,31,206,30,28,31,28,31,28,30,28,29,199,31,28,31,86,31,115,31,4,31,119,31,119,30,119,29,63,31,31,31,31,30,31,29,175,31,175,30,67,31,144,31,144,30,172,31,222,31,8,31,148,31,148,30,221,31,146,31,120,31,88,31,94,31,80,31,127,31,144,31,239,31,118,31,89,31,198,31,172,31,46,31,123,31,55,31,7,31,149,31,62,31,24,31,24,30,43,31,33,31,33,30,115,31,217,31,206,31,186,31,14,31,254,31,147,31,154,31,141,31,134,31,24,31,187,31,187,30,55,31,155,31,186,31,107,31,123,31,61,31,207,31,7,31,130,31,10,31,114,31,138,31,138,30,16,31,104,31,1,31,153,31,182,31,182,30,182,29,66,31,243,31,243,30,151,31,118,31,143,31,176,31,93,31,169,31,154,31,113,31,161,31,2,31,134,31,194,31,218,31,218,30,218,29,227,31,227,30,215,31,215,30,215,29,49,31,96,31,12,31,219,31,219,30,226,31,93,31,216,31,240,31,240,30,142,31,195,31,173,31,108,31,48,31,20,31,167,31,167,30,154,31,63,31,132,31,123,31,248,31,19,31,19,30,153,31,154,31,61,31,106,31,106,30,212,31,68,31,200,31,56,31,233,31,185,31,177,31,187,31,187,30,16,31,140,31,164,31,3,31,70,31,82,31,82,30,221,31,52,31,208,31,114,31,201,31,203,31,191,31,225,31,75,31,69,31,128,31,128,30,128,29,189,31,189,30,247,31,68,31,75,31,180,31,180,30,154,31,221,31,26,31,16,31,8,31,228,31,243,31,243,30,200,31,71,31,152,31,115,31,175,31,238,31,224,31,136,31,60,31,146,31,231,31,32,31,32,30,10,31,219,31,233,31,233,30,126,31,126,30,194,31,125,31,170,31,118,31,118,30,7,31,1,31,1,30,94,31,255,31,39,31,182,31,182,30,182,29,28,31,28,30,196,31,124,31,147,31,191,31,191,30,224,31,185,31,185,30,61,31,187,31,187,30,17,31,19,31,221,31,144,31,62,31,226,31,226,30,117,31,78,31,78,30,239,31,248,31,112,31,21,31,80,31,186,31,21,31,212,31,176,31,228,31,246,31,93,31,78,31,238,31,214,31,68,31,68,30,82,31,108,31,108,30,108,29,125,31,47,31,47,30,82,31,82,30,207,31,60,31,42,31,42,30,83,31,83,30,83,29,83,28,100,31,151,31,165,31,165,30,167,31,56,31,56,30,193,31,193,30,91,31,36,31,36,30,242,31,30,31,10,31,202,31,171,31,102,31,102,30,31,31,31,30,162,31,235,31,223,31,243,31,193,31,193,30,199,31,1,31,16,31,27,31,27,30,27,29,233,31,85,31,145,31,71,31,68,31,245,31,79,31,184,31,236,31,43,31,60,31,228,31,228,30,190,31,230,31,181,31,175,31,89,31,100,31,25,31,101,31,164,31,164,30,124,31,224,31,8,31,245,31,105,31,125,31,109,31,109,30,170,31,84,31,153,31,47,31,194,31,99,31,175,31,95,31,221,31,133,31,151,31,110,31,125,31,250,31,61,31,178,31,121,31,40,31,40,30,28,31,231,31,77,31,98,31,120,31,76,31,97,31,9,31,203,31,157,31,211,31,202,31,202,30,100,31,57,31,137,31,117,31,32,31,32,30,125,31,158,31,222,31,69,31,156,31,202,31,236,31,74,31,74,30,53,31,122,31,120,31,66,31,10,31,251,31,172,31,63,31,181,31,181,30,47,31,41,31,175,31,14,31,97,31,104,31,147,31,36,31,91,31,202,31,148,31,63,31,205,31,205,30,241,31,122,31,224,31,224,30,224,29,73,31,170,31,202,31,172,31,172,30,27,31,139,31,210,31,98,31,144,31,23,31,55,31,159,31,43,31,244,31,244,30,244,29,159,31,159,30,163,31,180,31,188,31,185,31,98,31,98,30,98,29,98,28,245,31,250,31,133,31,133,30,111,31,214,31,171,31,47,31,86,31,71,31,87,31,87,30,247,31,54,31,96,31,52,31,52,30,177,31,177,30,118,31,118,30,167,31,122,31,142,31,29,31,200,31,200,30,245,31,189,31,39,31,115,31,145,31,136,31,184,31,208,31,232,31,232,30,24,31,123,31,70,31,181,31,215,31,150,31,175,31,16,31,247,31,78,31,44,31,66,31,147,31,178,31,248,31,82,31,59,31,89,31,64,31,59,31,163,31,80,31,88,31,88,30,152,31,152,30,27,31,27,30,176,31,87,31,173,31,173,30,52,31,236,31,49,31,49,30,7,31,7,30,7,29,112,31,112,30,112,29,112,28,48,31,7,31,65,31,82,31,1,31,1,30,241,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
