-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_926 is
end project_tb_926;

architecture project_tb_arch_926 of project_tb_926 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 987;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (235,0,230,0,107,0,206,0,0,0,199,0,229,0,0,0,185,0,58,0,125,0,53,0,128,0,0,0,169,0,230,0,21,0,216,0,92,0,0,0,83,0,67,0,142,0,227,0,123,0,19,0,173,0,121,0,108,0,243,0,125,0,214,0,141,0,21,0,68,0,113,0,12,0,142,0,215,0,0,0,180,0,41,0,196,0,0,0,83,0,44,0,189,0,249,0,225,0,110,0,159,0,159,0,0,0,168,0,252,0,50,0,252,0,137,0,207,0,1,0,61,0,88,0,90,0,0,0,0,0,35,0,0,0,0,0,131,0,126,0,27,0,77,0,177,0,152,0,97,0,226,0,0,0,0,0,159,0,0,0,83,0,107,0,157,0,172,0,36,0,0,0,32,0,62,0,136,0,0,0,243,0,145,0,56,0,50,0,250,0,0,0,135,0,118,0,0,0,7,0,4,0,216,0,83,0,23,0,144,0,123,0,64,0,242,0,98,0,162,0,253,0,75,0,25,0,102,0,142,0,35,0,149,0,180,0,238,0,0,0,0,0,0,0,114,0,233,0,240,0,2,0,191,0,14,0,0,0,248,0,0,0,70,0,138,0,169,0,1,0,208,0,228,0,143,0,49,0,0,0,249,0,57,0,132,0,130,0,104,0,243,0,87,0,0,0,119,0,0,0,153,0,71,0,48,0,173,0,0,0,133,0,141,0,0,0,0,0,143,0,181,0,0,0,243,0,10,0,117,0,167,0,156,0,106,0,207,0,172,0,192,0,102,0,135,0,81,0,152,0,0,0,136,0,0,0,0,0,0,0,0,0,202,0,0,0,53,0,159,0,185,0,0,0,160,0,95,0,27,0,82,0,0,0,175,0,243,0,0,0,194,0,0,0,231,0,147,0,204,0,16,0,0,0,150,0,31,0,231,0,0,0,2,0,130,0,9,0,52,0,231,0,247,0,53,0,0,0,208,0,8,0,74,0,173,0,17,0,45,0,0,0,0,0,107,0,169,0,0,0,0,0,76,0,45,0,102,0,156,0,80,0,193,0,43,0,0,0,190,0,0,0,212,0,204,0,163,0,136,0,0,0,50,0,0,0,18,0,102,0,21,0,10,0,120,0,168,0,73,0,0,0,163,0,234,0,0,0,55,0,188,0,31,0,0,0,165,0,243,0,168,0,130,0,16,0,63,0,167,0,42,0,0,0,88,0,0,0,216,0,55,0,185,0,92,0,0,0,235,0,112,0,100,0,104,0,181,0,242,0,79,0,95,0,58,0,47,0,230,0,146,0,32,0,0,0,231,0,11,0,244,0,250,0,143,0,0,0,0,0,0,0,46,0,102,0,242,0,238,0,249,0,0,0,222,0,0,0,178,0,175,0,222,0,0,0,0,0,175,0,0,0,217,0,0,0,65,0,153,0,213,0,6,0,214,0,142,0,62,0,250,0,187,0,27,0,0,0,45,0,24,0,124,0,178,0,0,0,174,0,246,0,97,0,34,0,203,0,227,0,49,0,249,0,85,0,0,0,235,0,102,0,0,0,0,0,0,0,226,0,87,0,172,0,148,0,86,0,6,0,154,0,204,0,202,0,229,0,0,0,0,0,0,0,0,0,0,0,164,0,0,0,152,0,186,0,0,0,39,0,0,0,109,0,223,0,44,0,48,0,43,0,41,0,252,0,119,0,148,0,85,0,12,0,135,0,180,0,0,0,181,0,203,0,165,0,0,0,229,0,0,0,190,0,188,0,0,0,140,0,41,0,101,0,0,0,0,0,2,0,0,0,0,0,0,0,152,0,148,0,178,0,74,0,192,0,99,0,115,0,206,0,0,0,171,0,0,0,147,0,4,0,43,0,0,0,19,0,12,0,108,0,230,0,0,0,5,0,0,0,163,0,0,0,228,0,2,0,76,0,30,0,0,0,94,0,0,0,119,0,58,0,131,0,0,0,48,0,236,0,136,0,197,0,176,0,74,0,180,0,231,0,42,0,25,0,45,0,35,0,162,0,240,0,45,0,253,0,183,0,48,0,210,0,181,0,0,0,0,0,166,0,0,0,18,0,10,0,125,0,0,0,165,0,250,0,185,0,212,0,81,0,61,0,220,0,180,0,210,0,196,0,186,0,237,0,0,0,58,0,0,0,0,0,9,0,138,0,153,0,15,0,0,0,0,0,64,0,82,0,99,0,185,0,16,0,37,0,233,0,177,0,244,0,0,0,62,0,86,0,50,0,141,0,125,0,38,0,253,0,4,0,168,0,162,0,180,0,0,0,22,0,0,0,19,0,33,0,95,0,125,0,95,0,185,0,110,0,152,0,140,0,55,0,61,0,160,0,70,0,237,0,212,0,90,0,0,0,177,0,125,0,0,0,0,0,255,0,64,0,121,0,155,0,0,0,225,0,19,0,218,0,248,0,34,0,0,0,14,0,146,0,194,0,224,0,78,0,0,0,0,0,66,0,238,0,39,0,100,0,188,0,0,0,139,0,186,0,0,0,211,0,225,0,94,0,85,0,1,0,171,0,0,0,166,0,34,0,105,0,0,0,50,0,128,0,221,0,251,0,195,0,9,0,135,0,70,0,25,0,172,0,161,0,74,0,50,0,241,0,74,0,218,0,0,0,241,0,20,0,149,0,0,0,0,0,185,0,51,0,193,0,0,0,191,0,103,0,146,0,244,0,2,0,28,0,13,0,55,0,0,0,0,0,238,0,0,0,0,0,216,0,0,0,124,0,114,0,72,0,11,0,211,0,86,0,250,0,15,0,216,0,119,0,0,0,239,0,100,0,85,0,104,0,174,0,59,0,255,0,0,0,167,0,197,0,38,0,225,0,249,0,117,0,9,0,67,0,0,0,81,0,250,0,206,0,0,0,215,0,11,0,205,0,120,0,233,0,17,0,82,0,97,0,141,0,47,0,29,0,112,0,170,0,98,0,0,0,33,0,27,0,0,0,15,0,91,0,20,0,17,0,196,0,51,0,117,0,237,0,1,0,61,0,177,0,252,0,113,0,160,0,78,0,69,0,197,0,102,0,118,0,0,0,0,0,191,0,234,0,255,0,9,0,201,0,0,0,161,0,95,0,0,0,133,0,98,0,94,0,68,0,253,0,202,0,5,0,153,0,0,0,67,0,0,0,245,0,152,0,201,0,190,0,185,0,38,0,212,0,110,0,0,0,0,0,177,0,141,0,144,0,12,0,77,0,61,0,0,0,167,0,0,0,87,0,102,0,104,0,192,0,146,0,0,0,171,0,85,0,11,0,0,0,0,0,0,0,87,0,0,0,81,0,236,0,0,0,73,0,184,0,219,0,174,0,85,0,116,0,83,0,182,0,94,0,0,0,0,0,139,0,119,0,151,0,73,0,242,0,194,0,40,0,139,0,134,0,152,0,42,0,45,0,0,0,175,0,18,0,5,0,4,0,231,0,202,0,122,0,0,0,0,0,0,0,246,0,228,0,0,0,0,0,57,0,18,0,137,0,163,0,234,0,194,0,50,0,0,0,41,0,0,0,0,0,140,0,0,0,0,0,248,0,0,0,241,0,107,0,1,0,82,0,212,0,0,0,107,0,111,0,0,0,0,0,210,0,0,0,36,0,75,0,0,0,65,0,37,0,178,0,0,0,237,0,134,0,54,0,135,0,0,0,252,0,202,0,24,0,187,0,92,0,45,0,161,0,165,0,0,0,26,0,47,0,3,0,250,0,39,0,192,0,25,0,214,0,176,0,139,0,0,0,144,0,218,0,245,0,133,0,0,0,7,0,34,0,69,0,0,0,0,0,0,0,131,0,198,0,239,0,128,0,182,0,214,0,172,0,0,0,95,0,152,0,6,0,0,0,189,0,51,0,0,0,160,0,147,0,0,0,123,0,162,0,0,0,254,0,165,0,196,0,19,0,139,0,29,0,0,0,50,0,133,0,94,0,19,0,0,0,0,0,79,0,250,0,236,0,53,0,106,0,199,0,222,0,127,0,205,0,46,0,26,0,0,0,73,0,225,0,53,0,202,0,188,0,221,0,0,0,42,0,231,0,204,0,73,0,96,0,206,0,20,0,101,0,184,0,140,0,0,0,0,0,35,0,166,0,38,0,229,0,0,0,0,0,158,0,158,0,170,0,211,0,59,0,250,0,245,0,36,0,0,0,78,0,0,0,18,0,6,0,117,0,210,0,0,0,58,0,3,0,36,0,8,0,0,0,129,0,158,0,0,0,238,0,113,0,0,0,251,0,169,0,188,0,78,0,0,0,0,0,248,0,19,0,36,0,179,0,0,0,0,0,219,0,19,0,246,0,45,0,237,0,0,0,145,0,0,0,19,0,146,0,0,0,239,0,254,0,178,0,0,0,139,0,48,0,186,0,0,0,43,0,32,0,213,0,239,0,209,0,103,0,158,0,249,0,254,0,0,0,158,0,160,0,169,0,102,0,130,0);
signal scenario_full  : scenario_type := (235,31,230,31,107,31,206,31,206,30,199,31,229,31,229,30,185,31,58,31,125,31,53,31,128,31,128,30,169,31,230,31,21,31,216,31,92,31,92,30,83,31,67,31,142,31,227,31,123,31,19,31,173,31,121,31,108,31,243,31,125,31,214,31,141,31,21,31,68,31,113,31,12,31,142,31,215,31,215,30,180,31,41,31,196,31,196,30,83,31,44,31,189,31,249,31,225,31,110,31,159,31,159,31,159,30,168,31,252,31,50,31,252,31,137,31,207,31,1,31,61,31,88,31,90,31,90,30,90,29,35,31,35,30,35,29,131,31,126,31,27,31,77,31,177,31,152,31,97,31,226,31,226,30,226,29,159,31,159,30,83,31,107,31,157,31,172,31,36,31,36,30,32,31,62,31,136,31,136,30,243,31,145,31,56,31,50,31,250,31,250,30,135,31,118,31,118,30,7,31,4,31,216,31,83,31,23,31,144,31,123,31,64,31,242,31,98,31,162,31,253,31,75,31,25,31,102,31,142,31,35,31,149,31,180,31,238,31,238,30,238,29,238,28,114,31,233,31,240,31,2,31,191,31,14,31,14,30,248,31,248,30,70,31,138,31,169,31,1,31,208,31,228,31,143,31,49,31,49,30,249,31,57,31,132,31,130,31,104,31,243,31,87,31,87,30,119,31,119,30,153,31,71,31,48,31,173,31,173,30,133,31,141,31,141,30,141,29,143,31,181,31,181,30,243,31,10,31,117,31,167,31,156,31,106,31,207,31,172,31,192,31,102,31,135,31,81,31,152,31,152,30,136,31,136,30,136,29,136,28,136,27,202,31,202,30,53,31,159,31,185,31,185,30,160,31,95,31,27,31,82,31,82,30,175,31,243,31,243,30,194,31,194,30,231,31,147,31,204,31,16,31,16,30,150,31,31,31,231,31,231,30,2,31,130,31,9,31,52,31,231,31,247,31,53,31,53,30,208,31,8,31,74,31,173,31,17,31,45,31,45,30,45,29,107,31,169,31,169,30,169,29,76,31,45,31,102,31,156,31,80,31,193,31,43,31,43,30,190,31,190,30,212,31,204,31,163,31,136,31,136,30,50,31,50,30,18,31,102,31,21,31,10,31,120,31,168,31,73,31,73,30,163,31,234,31,234,30,55,31,188,31,31,31,31,30,165,31,243,31,168,31,130,31,16,31,63,31,167,31,42,31,42,30,88,31,88,30,216,31,55,31,185,31,92,31,92,30,235,31,112,31,100,31,104,31,181,31,242,31,79,31,95,31,58,31,47,31,230,31,146,31,32,31,32,30,231,31,11,31,244,31,250,31,143,31,143,30,143,29,143,28,46,31,102,31,242,31,238,31,249,31,249,30,222,31,222,30,178,31,175,31,222,31,222,30,222,29,175,31,175,30,217,31,217,30,65,31,153,31,213,31,6,31,214,31,142,31,62,31,250,31,187,31,27,31,27,30,45,31,24,31,124,31,178,31,178,30,174,31,246,31,97,31,34,31,203,31,227,31,49,31,249,31,85,31,85,30,235,31,102,31,102,30,102,29,102,28,226,31,87,31,172,31,148,31,86,31,6,31,154,31,204,31,202,31,229,31,229,30,229,29,229,28,229,27,229,26,164,31,164,30,152,31,186,31,186,30,39,31,39,30,109,31,223,31,44,31,48,31,43,31,41,31,252,31,119,31,148,31,85,31,12,31,135,31,180,31,180,30,181,31,203,31,165,31,165,30,229,31,229,30,190,31,188,31,188,30,140,31,41,31,101,31,101,30,101,29,2,31,2,30,2,29,2,28,152,31,148,31,178,31,74,31,192,31,99,31,115,31,206,31,206,30,171,31,171,30,147,31,4,31,43,31,43,30,19,31,12,31,108,31,230,31,230,30,5,31,5,30,163,31,163,30,228,31,2,31,76,31,30,31,30,30,94,31,94,30,119,31,58,31,131,31,131,30,48,31,236,31,136,31,197,31,176,31,74,31,180,31,231,31,42,31,25,31,45,31,35,31,162,31,240,31,45,31,253,31,183,31,48,31,210,31,181,31,181,30,181,29,166,31,166,30,18,31,10,31,125,31,125,30,165,31,250,31,185,31,212,31,81,31,61,31,220,31,180,31,210,31,196,31,186,31,237,31,237,30,58,31,58,30,58,29,9,31,138,31,153,31,15,31,15,30,15,29,64,31,82,31,99,31,185,31,16,31,37,31,233,31,177,31,244,31,244,30,62,31,86,31,50,31,141,31,125,31,38,31,253,31,4,31,168,31,162,31,180,31,180,30,22,31,22,30,19,31,33,31,95,31,125,31,95,31,185,31,110,31,152,31,140,31,55,31,61,31,160,31,70,31,237,31,212,31,90,31,90,30,177,31,125,31,125,30,125,29,255,31,64,31,121,31,155,31,155,30,225,31,19,31,218,31,248,31,34,31,34,30,14,31,146,31,194,31,224,31,78,31,78,30,78,29,66,31,238,31,39,31,100,31,188,31,188,30,139,31,186,31,186,30,211,31,225,31,94,31,85,31,1,31,171,31,171,30,166,31,34,31,105,31,105,30,50,31,128,31,221,31,251,31,195,31,9,31,135,31,70,31,25,31,172,31,161,31,74,31,50,31,241,31,74,31,218,31,218,30,241,31,20,31,149,31,149,30,149,29,185,31,51,31,193,31,193,30,191,31,103,31,146,31,244,31,2,31,28,31,13,31,55,31,55,30,55,29,238,31,238,30,238,29,216,31,216,30,124,31,114,31,72,31,11,31,211,31,86,31,250,31,15,31,216,31,119,31,119,30,239,31,100,31,85,31,104,31,174,31,59,31,255,31,255,30,167,31,197,31,38,31,225,31,249,31,117,31,9,31,67,31,67,30,81,31,250,31,206,31,206,30,215,31,11,31,205,31,120,31,233,31,17,31,82,31,97,31,141,31,47,31,29,31,112,31,170,31,98,31,98,30,33,31,27,31,27,30,15,31,91,31,20,31,17,31,196,31,51,31,117,31,237,31,1,31,61,31,177,31,252,31,113,31,160,31,78,31,69,31,197,31,102,31,118,31,118,30,118,29,191,31,234,31,255,31,9,31,201,31,201,30,161,31,95,31,95,30,133,31,98,31,94,31,68,31,253,31,202,31,5,31,153,31,153,30,67,31,67,30,245,31,152,31,201,31,190,31,185,31,38,31,212,31,110,31,110,30,110,29,177,31,141,31,144,31,12,31,77,31,61,31,61,30,167,31,167,30,87,31,102,31,104,31,192,31,146,31,146,30,171,31,85,31,11,31,11,30,11,29,11,28,87,31,87,30,81,31,236,31,236,30,73,31,184,31,219,31,174,31,85,31,116,31,83,31,182,31,94,31,94,30,94,29,139,31,119,31,151,31,73,31,242,31,194,31,40,31,139,31,134,31,152,31,42,31,45,31,45,30,175,31,18,31,5,31,4,31,231,31,202,31,122,31,122,30,122,29,122,28,246,31,228,31,228,30,228,29,57,31,18,31,137,31,163,31,234,31,194,31,50,31,50,30,41,31,41,30,41,29,140,31,140,30,140,29,248,31,248,30,241,31,107,31,1,31,82,31,212,31,212,30,107,31,111,31,111,30,111,29,210,31,210,30,36,31,75,31,75,30,65,31,37,31,178,31,178,30,237,31,134,31,54,31,135,31,135,30,252,31,202,31,24,31,187,31,92,31,45,31,161,31,165,31,165,30,26,31,47,31,3,31,250,31,39,31,192,31,25,31,214,31,176,31,139,31,139,30,144,31,218,31,245,31,133,31,133,30,7,31,34,31,69,31,69,30,69,29,69,28,131,31,198,31,239,31,128,31,182,31,214,31,172,31,172,30,95,31,152,31,6,31,6,30,189,31,51,31,51,30,160,31,147,31,147,30,123,31,162,31,162,30,254,31,165,31,196,31,19,31,139,31,29,31,29,30,50,31,133,31,94,31,19,31,19,30,19,29,79,31,250,31,236,31,53,31,106,31,199,31,222,31,127,31,205,31,46,31,26,31,26,30,73,31,225,31,53,31,202,31,188,31,221,31,221,30,42,31,231,31,204,31,73,31,96,31,206,31,20,31,101,31,184,31,140,31,140,30,140,29,35,31,166,31,38,31,229,31,229,30,229,29,158,31,158,31,170,31,211,31,59,31,250,31,245,31,36,31,36,30,78,31,78,30,18,31,6,31,117,31,210,31,210,30,58,31,3,31,36,31,8,31,8,30,129,31,158,31,158,30,238,31,113,31,113,30,251,31,169,31,188,31,78,31,78,30,78,29,248,31,19,31,36,31,179,31,179,30,179,29,219,31,19,31,246,31,45,31,237,31,237,30,145,31,145,30,19,31,146,31,146,30,239,31,254,31,178,31,178,30,139,31,48,31,186,31,186,30,43,31,32,31,213,31,239,31,209,31,103,31,158,31,249,31,254,31,254,30,158,31,160,31,169,31,102,31,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
