-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 792;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (33,0,84,0,0,0,129,0,152,0,155,0,61,0,180,0,244,0,9,0,20,0,201,0,119,0,148,0,0,0,20,0,171,0,146,0,0,0,150,0,64,0,81,0,77,0,118,0,176,0,99,0,22,0,85,0,73,0,208,0,60,0,121,0,190,0,132,0,181,0,140,0,41,0,159,0,0,0,47,0,204,0,179,0,0,0,30,0,168,0,125,0,34,0,118,0,34,0,155,0,123,0,0,0,61,0,3,0,50,0,0,0,0,0,62,0,16,0,162,0,153,0,86,0,39,0,0,0,188,0,194,0,0,0,118,0,155,0,142,0,38,0,95,0,144,0,0,0,8,0,157,0,153,0,92,0,6,0,176,0,252,0,36,0,0,0,28,0,104,0,113,0,0,0,201,0,95,0,12,0,251,0,77,0,182,0,0,0,103,0,32,0,63,0,0,0,136,0,79,0,8,0,50,0,0,0,92,0,40,0,0,0,54,0,0,0,0,0,101,0,139,0,0,0,0,0,12,0,124,0,96,0,137,0,101,0,223,0,93,0,148,0,80,0,85,0,105,0,0,0,86,0,0,0,115,0,218,0,52,0,51,0,21,0,104,0,54,0,0,0,34,0,228,0,48,0,34,0,2,0,95,0,250,0,0,0,25,0,76,0,1,0,190,0,93,0,0,0,0,0,138,0,79,0,195,0,0,0,234,0,87,0,118,0,0,0,211,0,0,0,208,0,91,0,17,0,95,0,177,0,40,0,0,0,107,0,156,0,80,0,131,0,236,0,121,0,46,0,0,0,0,0,165,0,249,0,99,0,62,0,57,0,0,0,190,0,101,0,0,0,136,0,159,0,0,0,78,0,198,0,194,0,161,0,133,0,236,0,0,0,220,0,241,0,192,0,71,0,79,0,7,0,0,0,80,0,184,0,252,0,188,0,0,0,100,0,48,0,156,0,188,0,0,0,0,0,193,0,4,0,8,0,40,0,183,0,133,0,153,0,148,0,0,0,91,0,90,0,13,0,97,0,157,0,64,0,75,0,245,0,0,0,157,0,51,0,76,0,0,0,127,0,90,0,184,0,61,0,77,0,0,0,76,0,84,0,0,0,56,0,0,0,156,0,0,0,37,0,72,0,116,0,108,0,226,0,247,0,38,0,163,0,131,0,0,0,195,0,51,0,99,0,161,0,215,0,231,0,2,0,118,0,161,0,137,0,60,0,26,0,198,0,0,0,147,0,255,0,82,0,225,0,92,0,34,0,201,0,203,0,0,0,78,0,92,0,100,0,135,0,55,0,170,0,0,0,94,0,182,0,79,0,49,0,232,0,167,0,18,0,48,0,26,0,88,0,55,0,22,0,216,0,0,0,41,0,40,0,251,0,91,0,124,0,100,0,161,0,73,0,110,0,0,0,253,0,0,0,22,0,84,0,78,0,0,0,166,0,0,0,161,0,144,0,195,0,151,0,83,0,130,0,167,0,24,0,176,0,102,0,0,0,114,0,156,0,0,0,18,0,0,0,0,0,189,0,107,0,51,0,250,0,229,0,0,0,0,0,10,0,119,0,80,0,0,0,0,0,140,0,143,0,0,0,228,0,180,0,155,0,134,0,0,0,76,0,26,0,151,0,190,0,186,0,198,0,0,0,222,0,252,0,0,0,95,0,253,0,109,0,0,0,0,0,86,0,156,0,0,0,36,0,141,0,126,0,0,0,130,0,168,0,34,0,17,0,153,0,0,0,227,0,120,0,0,0,146,0,0,0,110,0,249,0,78,0,1,0,127,0,218,0,152,0,0,0,229,0,142,0,5,0,0,0,73,0,200,0,0,0,51,0,166,0,0,0,0,0,173,0,65,0,0,0,54,0,66,0,0,0,180,0,160,0,0,0,0,0,174,0,0,0,5,0,223,0,245,0,66,0,206,0,79,0,118,0,34,0,234,0,170,0,31,0,246,0,138,0,240,0,145,0,104,0,0,0,231,0,25,0,192,0,64,0,0,0,109,0,232,0,177,0,165,0,188,0,200,0,243,0,33,0,246,0,0,0,93,0,70,0,232,0,195,0,6,0,230,0,135,0,0,0,133,0,91,0,159,0,187,0,134,0,255,0,222,0,74,0,99,0,150,0,130,0,137,0,185,0,0,0,140,0,150,0,227,0,0,0,166,0,81,0,219,0,237,0,200,0,30,0,243,0,0,0,57,0,0,0,76,0,167,0,204,0,63,0,192,0,191,0,85,0,173,0,244,0,114,0,51,0,181,0,90,0,249,0,67,0,157,0,0,0,87,0,118,0,36,0,32,0,38,0,246,0,0,0,0,0,105,0,23,0,132,0,0,0,0,0,6,0,113,0,192,0,0,0,134,0,249,0,231,0,183,0,14,0,171,0,49,0,178,0,0,0,174,0,54,0,30,0,228,0,127,0,172,0,191,0,79,0,0,0,214,0,51,0,0,0,187,0,47,0,109,0,0,0,61,0,248,0,109,0,61,0,49,0,243,0,39,0,225,0,105,0,222,0,191,0,192,0,0,0,128,0,130,0,217,0,193,0,0,0,176,0,49,0,96,0,1,0,0,0,13,0,0,0,222,0,161,0,160,0,1,0,0,0,118,0,115,0,114,0,170,0,164,0,236,0,219,0,179,0,80,0,117,0,90,0,0,0,234,0,122,0,0,0,0,0,86,0,79,0,28,0,245,0,177,0,117,0,110,0,0,0,197,0,45,0,0,0,137,0,38,0,59,0,40,0,156,0,90,0,208,0,157,0,25,0,172,0,190,0,215,0,219,0,0,0,127,0,36,0,186,0,43,0,0,0,64,0,161,0,70,0,80,0,146,0,0,0,175,0,26,0,84,0,253,0,0,0,0,0,100,0,42,0,70,0,0,0,118,0,14,0,45,0,0,0,181,0,44,0,34,0,68,0,187,0,120,0,0,0,133,0,66,0,214,0,83,0,218,0,212,0,238,0,0,0,56,0,28,0,57,0,15,0,60,0,0,0,89,0,75,0,146,0,62,0,79,0,149,0,174,0,140,0,105,0,225,0,71,0,0,0,154,0,0,0,0,0,197,0,0,0,205,0,102,0,251,0,20,0,123,0,78,0,85,0,193,0,203,0,118,0,235,0,83,0,0,0,156,0,237,0,20,0,28,0,0,0,214,0,0,0,183,0,0,0,190,0,0,0,154,0,80,0,252,0,26,0,0,0,0,0,169,0,115,0,159,0,135,0,137,0,131,0,0,0,203,0,190,0,0,0,0,0,88,0,157,0,0,0,0,0,0,0,138,0,0,0,223,0,191,0,32,0,182,0,133,0,133,0,136,0,191,0,194,0,134,0,0,0,28,0,165,0,218,0,113,0,125,0,149,0,181,0,90,0,191,0,0,0,204,0,54,0,238,0,183,0,220,0,18,0,65,0,72,0,84,0,0,0,141,0,0,0,0,0,73,0,23,0,254,0,226,0,174,0,168,0,124,0,0,0,158,0,0,0,92,0,240,0,34,0,165,0,39,0,0,0,0,0,95,0,213,0,220,0,236,0,0,0,190,0,110,0,140,0,186,0,151,0,0,0);
signal scenario_full  : scenario_type := (33,31,84,31,84,30,129,31,152,31,155,31,61,31,180,31,244,31,9,31,20,31,201,31,119,31,148,31,148,30,20,31,171,31,146,31,146,30,150,31,64,31,81,31,77,31,118,31,176,31,99,31,22,31,85,31,73,31,208,31,60,31,121,31,190,31,132,31,181,31,140,31,41,31,159,31,159,30,47,31,204,31,179,31,179,30,30,31,168,31,125,31,34,31,118,31,34,31,155,31,123,31,123,30,61,31,3,31,50,31,50,30,50,29,62,31,16,31,162,31,153,31,86,31,39,31,39,30,188,31,194,31,194,30,118,31,155,31,142,31,38,31,95,31,144,31,144,30,8,31,157,31,153,31,92,31,6,31,176,31,252,31,36,31,36,30,28,31,104,31,113,31,113,30,201,31,95,31,12,31,251,31,77,31,182,31,182,30,103,31,32,31,63,31,63,30,136,31,79,31,8,31,50,31,50,30,92,31,40,31,40,30,54,31,54,30,54,29,101,31,139,31,139,30,139,29,12,31,124,31,96,31,137,31,101,31,223,31,93,31,148,31,80,31,85,31,105,31,105,30,86,31,86,30,115,31,218,31,52,31,51,31,21,31,104,31,54,31,54,30,34,31,228,31,48,31,34,31,2,31,95,31,250,31,250,30,25,31,76,31,1,31,190,31,93,31,93,30,93,29,138,31,79,31,195,31,195,30,234,31,87,31,118,31,118,30,211,31,211,30,208,31,91,31,17,31,95,31,177,31,40,31,40,30,107,31,156,31,80,31,131,31,236,31,121,31,46,31,46,30,46,29,165,31,249,31,99,31,62,31,57,31,57,30,190,31,101,31,101,30,136,31,159,31,159,30,78,31,198,31,194,31,161,31,133,31,236,31,236,30,220,31,241,31,192,31,71,31,79,31,7,31,7,30,80,31,184,31,252,31,188,31,188,30,100,31,48,31,156,31,188,31,188,30,188,29,193,31,4,31,8,31,40,31,183,31,133,31,153,31,148,31,148,30,91,31,90,31,13,31,97,31,157,31,64,31,75,31,245,31,245,30,157,31,51,31,76,31,76,30,127,31,90,31,184,31,61,31,77,31,77,30,76,31,84,31,84,30,56,31,56,30,156,31,156,30,37,31,72,31,116,31,108,31,226,31,247,31,38,31,163,31,131,31,131,30,195,31,51,31,99,31,161,31,215,31,231,31,2,31,118,31,161,31,137,31,60,31,26,31,198,31,198,30,147,31,255,31,82,31,225,31,92,31,34,31,201,31,203,31,203,30,78,31,92,31,100,31,135,31,55,31,170,31,170,30,94,31,182,31,79,31,49,31,232,31,167,31,18,31,48,31,26,31,88,31,55,31,22,31,216,31,216,30,41,31,40,31,251,31,91,31,124,31,100,31,161,31,73,31,110,31,110,30,253,31,253,30,22,31,84,31,78,31,78,30,166,31,166,30,161,31,144,31,195,31,151,31,83,31,130,31,167,31,24,31,176,31,102,31,102,30,114,31,156,31,156,30,18,31,18,30,18,29,189,31,107,31,51,31,250,31,229,31,229,30,229,29,10,31,119,31,80,31,80,30,80,29,140,31,143,31,143,30,228,31,180,31,155,31,134,31,134,30,76,31,26,31,151,31,190,31,186,31,198,31,198,30,222,31,252,31,252,30,95,31,253,31,109,31,109,30,109,29,86,31,156,31,156,30,36,31,141,31,126,31,126,30,130,31,168,31,34,31,17,31,153,31,153,30,227,31,120,31,120,30,146,31,146,30,110,31,249,31,78,31,1,31,127,31,218,31,152,31,152,30,229,31,142,31,5,31,5,30,73,31,200,31,200,30,51,31,166,31,166,30,166,29,173,31,65,31,65,30,54,31,66,31,66,30,180,31,160,31,160,30,160,29,174,31,174,30,5,31,223,31,245,31,66,31,206,31,79,31,118,31,34,31,234,31,170,31,31,31,246,31,138,31,240,31,145,31,104,31,104,30,231,31,25,31,192,31,64,31,64,30,109,31,232,31,177,31,165,31,188,31,200,31,243,31,33,31,246,31,246,30,93,31,70,31,232,31,195,31,6,31,230,31,135,31,135,30,133,31,91,31,159,31,187,31,134,31,255,31,222,31,74,31,99,31,150,31,130,31,137,31,185,31,185,30,140,31,150,31,227,31,227,30,166,31,81,31,219,31,237,31,200,31,30,31,243,31,243,30,57,31,57,30,76,31,167,31,204,31,63,31,192,31,191,31,85,31,173,31,244,31,114,31,51,31,181,31,90,31,249,31,67,31,157,31,157,30,87,31,118,31,36,31,32,31,38,31,246,31,246,30,246,29,105,31,23,31,132,31,132,30,132,29,6,31,113,31,192,31,192,30,134,31,249,31,231,31,183,31,14,31,171,31,49,31,178,31,178,30,174,31,54,31,30,31,228,31,127,31,172,31,191,31,79,31,79,30,214,31,51,31,51,30,187,31,47,31,109,31,109,30,61,31,248,31,109,31,61,31,49,31,243,31,39,31,225,31,105,31,222,31,191,31,192,31,192,30,128,31,130,31,217,31,193,31,193,30,176,31,49,31,96,31,1,31,1,30,13,31,13,30,222,31,161,31,160,31,1,31,1,30,118,31,115,31,114,31,170,31,164,31,236,31,219,31,179,31,80,31,117,31,90,31,90,30,234,31,122,31,122,30,122,29,86,31,79,31,28,31,245,31,177,31,117,31,110,31,110,30,197,31,45,31,45,30,137,31,38,31,59,31,40,31,156,31,90,31,208,31,157,31,25,31,172,31,190,31,215,31,219,31,219,30,127,31,36,31,186,31,43,31,43,30,64,31,161,31,70,31,80,31,146,31,146,30,175,31,26,31,84,31,253,31,253,30,253,29,100,31,42,31,70,31,70,30,118,31,14,31,45,31,45,30,181,31,44,31,34,31,68,31,187,31,120,31,120,30,133,31,66,31,214,31,83,31,218,31,212,31,238,31,238,30,56,31,28,31,57,31,15,31,60,31,60,30,89,31,75,31,146,31,62,31,79,31,149,31,174,31,140,31,105,31,225,31,71,31,71,30,154,31,154,30,154,29,197,31,197,30,205,31,102,31,251,31,20,31,123,31,78,31,85,31,193,31,203,31,118,31,235,31,83,31,83,30,156,31,237,31,20,31,28,31,28,30,214,31,214,30,183,31,183,30,190,31,190,30,154,31,80,31,252,31,26,31,26,30,26,29,169,31,115,31,159,31,135,31,137,31,131,31,131,30,203,31,190,31,190,30,190,29,88,31,157,31,157,30,157,29,157,28,138,31,138,30,223,31,191,31,32,31,182,31,133,31,133,31,136,31,191,31,194,31,134,31,134,30,28,31,165,31,218,31,113,31,125,31,149,31,181,31,90,31,191,31,191,30,204,31,54,31,238,31,183,31,220,31,18,31,65,31,72,31,84,31,84,30,141,31,141,30,141,29,73,31,23,31,254,31,226,31,174,31,168,31,124,31,124,30,158,31,158,30,92,31,240,31,34,31,165,31,39,31,39,30,39,29,95,31,213,31,220,31,236,31,236,30,190,31,110,31,140,31,186,31,151,31,151,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
