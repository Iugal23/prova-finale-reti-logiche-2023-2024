-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_373 is
end project_tb_373;

architecture project_tb_arch_373 of project_tb_373 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 504;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (141,0,184,0,148,0,46,0,237,0,25,0,209,0,249,0,224,0,0,0,154,0,27,0,0,0,202,0,84,0,94,0,46,0,57,0,95,0,155,0,216,0,0,0,102,0,221,0,0,0,244,0,86,0,116,0,0,0,36,0,101,0,40,0,106,0,32,0,83,0,182,0,26,0,127,0,92,0,0,0,105,0,119,0,194,0,0,0,145,0,24,0,18,0,250,0,118,0,152,0,0,0,157,0,0,0,0,0,44,0,131,0,0,0,206,0,112,0,0,0,128,0,28,0,55,0,125,0,51,0,0,0,64,0,0,0,237,0,138,0,0,0,197,0,0,0,0,0,202,0,113,0,24,0,164,0,128,0,67,0,0,0,0,0,145,0,193,0,0,0,133,0,113,0,205,0,255,0,7,0,161,0,245,0,254,0,0,0,80,0,129,0,128,0,42,0,234,0,76,0,254,0,105,0,73,0,110,0,0,0,143,0,0,0,137,0,126,0,36,0,9,0,0,0,232,0,214,0,137,0,202,0,117,0,0,0,243,0,248,0,194,0,125,0,0,0,0,0,16,0,0,0,255,0,26,0,117,0,46,0,0,0,128,0,0,0,141,0,205,0,0,0,241,0,22,0,0,0,176,0,246,0,0,0,18,0,233,0,101,0,8,0,102,0,138,0,119,0,61,0,64,0,32,0,77,0,28,0,70,0,26,0,109,0,0,0,119,0,33,0,111,0,234,0,166,0,166,0,39,0,0,0,166,0,114,0,130,0,74,0,32,0,0,0,150,0,109,0,135,0,176,0,254,0,204,0,249,0,198,0,100,0,0,0,156,0,236,0,88,0,214,0,26,0,0,0,83,0,219,0,253,0,101,0,0,0,136,0,118,0,57,0,106,0,155,0,2,0,176,0,0,0,90,0,134,0,0,0,110,0,0,0,126,0,67,0,0,0,179,0,23,0,220,0,157,0,69,0,17,0,12,0,139,0,92,0,209,0,78,0,0,0,0,0,84,0,5,0,163,0,0,0,0,0,131,0,143,0,104,0,37,0,197,0,0,0,0,0,54,0,0,0,51,0,30,0,0,0,100,0,22,0,0,0,85,0,6,0,117,0,135,0,112,0,0,0,27,0,52,0,0,0,253,0,81,0,188,0,15,0,242,0,185,0,147,0,199,0,252,0,55,0,12,0,18,0,251,0,90,0,221,0,0,0,0,0,10,0,106,0,211,0,181,0,0,0,47,0,52,0,2,0,57,0,34,0,23,0,160,0,78,0,23,0,108,0,0,0,130,0,73,0,28,0,131,0,145,0,48,0,40,0,244,0,198,0,211,0,164,0,60,0,144,0,172,0,50,0,208,0,1,0,211,0,0,0,0,0,0,0,177,0,202,0,141,0,166,0,0,0,187,0,33,0,193,0,122,0,248,0,22,0,199,0,0,0,231,0,100,0,106,0,178,0,0,0,0,0,69,0,196,0,81,0,0,0,88,0,161,0,15,0,194,0,0,0,9,0,0,0,54,0,185,0,89,0,36,0,219,0,79,0,0,0,153,0,90,0,0,0,220,0,111,0,203,0,218,0,187,0,19,0,0,0,195,0,22,0,0,0,0,0,104,0,151,0,77,0,183,0,41,0,69,0,166,0,121,0,228,0,218,0,200,0,217,0,153,0,239,0,20,0,57,0,112,0,49,0,159,0,170,0,144,0,0,0,3,0,124,0,102,0,0,0,168,0,192,0,0,0,12,0,0,0,226,0,0,0,21,0,0,0,167,0,62,0,240,0,7,0,134,0,126,0,193,0,0,0,205,0,50,0,224,0,44,0,102,0,13,0,144,0,39,0,211,0,219,0,148,0,153,0,0,0,189,0,43,0,0,0,0,0,58,0,34,0,159,0,0,0,54,0,0,0,82,0,40,0,0,0,194,0,21,0,13,0,0,0,213,0,154,0,155,0,187,0,23,0,4,0,79,0,72,0,93,0,204,0,0,0,166,0,104,0,11,0,116,0,0,0,184,0,0,0,216,0,164,0,85,0,254,0,229,0,239,0,60,0,49,0,0,0,33,0,0,0,0,0,134,0,0,0,46,0,65,0,151,0,0,0,168,0,108,0,147,0,238,0,180,0,187,0,220,0,0,0,18,0,234,0,222,0,55,0,120,0,121,0,0,0,191,0,0,0,19,0,184,0,19,0,0,0,105,0,154,0,237,0,196,0,195,0,14,0,34,0,37,0,221,0,89,0,8,0,8,0,235,0,235,0,179,0,34,0,186,0,43,0);
signal scenario_full  : scenario_type := (141,31,184,31,148,31,46,31,237,31,25,31,209,31,249,31,224,31,224,30,154,31,27,31,27,30,202,31,84,31,94,31,46,31,57,31,95,31,155,31,216,31,216,30,102,31,221,31,221,30,244,31,86,31,116,31,116,30,36,31,101,31,40,31,106,31,32,31,83,31,182,31,26,31,127,31,92,31,92,30,105,31,119,31,194,31,194,30,145,31,24,31,18,31,250,31,118,31,152,31,152,30,157,31,157,30,157,29,44,31,131,31,131,30,206,31,112,31,112,30,128,31,28,31,55,31,125,31,51,31,51,30,64,31,64,30,237,31,138,31,138,30,197,31,197,30,197,29,202,31,113,31,24,31,164,31,128,31,67,31,67,30,67,29,145,31,193,31,193,30,133,31,113,31,205,31,255,31,7,31,161,31,245,31,254,31,254,30,80,31,129,31,128,31,42,31,234,31,76,31,254,31,105,31,73,31,110,31,110,30,143,31,143,30,137,31,126,31,36,31,9,31,9,30,232,31,214,31,137,31,202,31,117,31,117,30,243,31,248,31,194,31,125,31,125,30,125,29,16,31,16,30,255,31,26,31,117,31,46,31,46,30,128,31,128,30,141,31,205,31,205,30,241,31,22,31,22,30,176,31,246,31,246,30,18,31,233,31,101,31,8,31,102,31,138,31,119,31,61,31,64,31,32,31,77,31,28,31,70,31,26,31,109,31,109,30,119,31,33,31,111,31,234,31,166,31,166,31,39,31,39,30,166,31,114,31,130,31,74,31,32,31,32,30,150,31,109,31,135,31,176,31,254,31,204,31,249,31,198,31,100,31,100,30,156,31,236,31,88,31,214,31,26,31,26,30,83,31,219,31,253,31,101,31,101,30,136,31,118,31,57,31,106,31,155,31,2,31,176,31,176,30,90,31,134,31,134,30,110,31,110,30,126,31,67,31,67,30,179,31,23,31,220,31,157,31,69,31,17,31,12,31,139,31,92,31,209,31,78,31,78,30,78,29,84,31,5,31,163,31,163,30,163,29,131,31,143,31,104,31,37,31,197,31,197,30,197,29,54,31,54,30,51,31,30,31,30,30,100,31,22,31,22,30,85,31,6,31,117,31,135,31,112,31,112,30,27,31,52,31,52,30,253,31,81,31,188,31,15,31,242,31,185,31,147,31,199,31,252,31,55,31,12,31,18,31,251,31,90,31,221,31,221,30,221,29,10,31,106,31,211,31,181,31,181,30,47,31,52,31,2,31,57,31,34,31,23,31,160,31,78,31,23,31,108,31,108,30,130,31,73,31,28,31,131,31,145,31,48,31,40,31,244,31,198,31,211,31,164,31,60,31,144,31,172,31,50,31,208,31,1,31,211,31,211,30,211,29,211,28,177,31,202,31,141,31,166,31,166,30,187,31,33,31,193,31,122,31,248,31,22,31,199,31,199,30,231,31,100,31,106,31,178,31,178,30,178,29,69,31,196,31,81,31,81,30,88,31,161,31,15,31,194,31,194,30,9,31,9,30,54,31,185,31,89,31,36,31,219,31,79,31,79,30,153,31,90,31,90,30,220,31,111,31,203,31,218,31,187,31,19,31,19,30,195,31,22,31,22,30,22,29,104,31,151,31,77,31,183,31,41,31,69,31,166,31,121,31,228,31,218,31,200,31,217,31,153,31,239,31,20,31,57,31,112,31,49,31,159,31,170,31,144,31,144,30,3,31,124,31,102,31,102,30,168,31,192,31,192,30,12,31,12,30,226,31,226,30,21,31,21,30,167,31,62,31,240,31,7,31,134,31,126,31,193,31,193,30,205,31,50,31,224,31,44,31,102,31,13,31,144,31,39,31,211,31,219,31,148,31,153,31,153,30,189,31,43,31,43,30,43,29,58,31,34,31,159,31,159,30,54,31,54,30,82,31,40,31,40,30,194,31,21,31,13,31,13,30,213,31,154,31,155,31,187,31,23,31,4,31,79,31,72,31,93,31,204,31,204,30,166,31,104,31,11,31,116,31,116,30,184,31,184,30,216,31,164,31,85,31,254,31,229,31,239,31,60,31,49,31,49,30,33,31,33,30,33,29,134,31,134,30,46,31,65,31,151,31,151,30,168,31,108,31,147,31,238,31,180,31,187,31,220,31,220,30,18,31,234,31,222,31,55,31,120,31,121,31,121,30,191,31,191,30,19,31,184,31,19,31,19,30,105,31,154,31,237,31,196,31,195,31,14,31,34,31,37,31,221,31,89,31,8,31,8,31,235,31,235,31,179,31,34,31,186,31,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
