-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_154 is
end project_tb_154;

architecture project_tb_arch_154 of project_tb_154 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 266;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,31,0,13,0,65,0,35,0,250,0,0,0,74,0,113,0,175,0,60,0,0,0,86,0,164,0,117,0,0,0,0,0,0,0,211,0,145,0,0,0,28,0,207,0,18,0,238,0,0,0,45,0,11,0,33,0,177,0,0,0,28,0,78,0,102,0,254,0,226,0,71,0,44,0,0,0,210,0,173,0,2,0,24,0,0,0,4,0,75,0,183,0,93,0,18,0,185,0,2,0,225,0,187,0,237,0,138,0,253,0,47,0,238,0,35,0,0,0,65,0,72,0,217,0,0,0,188,0,7,0,233,0,109,0,238,0,115,0,49,0,30,0,73,0,131,0,143,0,47,0,189,0,33,0,1,0,108,0,98,0,238,0,0,0,110,0,0,0,198,0,60,0,96,0,107,0,0,0,211,0,0,0,0,0,215,0,4,0,64,0,124,0,112,0,206,0,100,0,7,0,114,0,199,0,83,0,223,0,108,0,148,0,0,0,48,0,88,0,214,0,40,0,0,0,175,0,60,0,54,0,0,0,158,0,0,0,64,0,237,0,244,0,202,0,179,0,251,0,30,0,55,0,0,0,0,0,52,0,241,0,80,0,164,0,195,0,0,0,206,0,193,0,0,0,0,0,71,0,14,0,179,0,0,0,113,0,232,0,0,0,188,0,193,0,220,0,158,0,8,0,12,0,108,0,142,0,128,0,198,0,0,0,220,0,221,0,0,0,91,0,202,0,27,0,134,0,1,0,99,0,240,0,234,0,0,0,204,0,67,0,0,0,205,0,0,0,0,0,237,0,69,0,0,0,80,0,0,0,0,0,238,0,232,0,54,0,55,0,245,0,44,0,64,0,0,0,80,0,110,0,3,0,0,0,90,0,62,0,0,0,205,0,146,0,158,0,138,0,140,0,176,0,253,0,93,0,76,0,246,0,95,0,5,0,55,0,116,0,164,0,17,0,93,0,110,0,158,0,0,0,105,0,202,0,0,0,180,0,25,0,0,0,14,0,0,0,176,0,225,0,0,0,239,0,148,0,164,0,171,0,171,0,98,0,115,0,15,0,54,0,220,0,0,0,64,0,0,0,0,0,0,0,0,0,34,0,0,0,167,0,252,0,111,0,64,0,213,0,62,0,127,0,43,0,82,0,171,0,0,0,140,0,179,0,212,0,250,0,56,0,139,0,188,0,160,0,29,0,0,0);
signal scenario_full  : scenario_type := (0,0,31,31,13,31,65,31,35,31,250,31,250,30,74,31,113,31,175,31,60,31,60,30,86,31,164,31,117,31,117,30,117,29,117,28,211,31,145,31,145,30,28,31,207,31,18,31,238,31,238,30,45,31,11,31,33,31,177,31,177,30,28,31,78,31,102,31,254,31,226,31,71,31,44,31,44,30,210,31,173,31,2,31,24,31,24,30,4,31,75,31,183,31,93,31,18,31,185,31,2,31,225,31,187,31,237,31,138,31,253,31,47,31,238,31,35,31,35,30,65,31,72,31,217,31,217,30,188,31,7,31,233,31,109,31,238,31,115,31,49,31,30,31,73,31,131,31,143,31,47,31,189,31,33,31,1,31,108,31,98,31,238,31,238,30,110,31,110,30,198,31,60,31,96,31,107,31,107,30,211,31,211,30,211,29,215,31,4,31,64,31,124,31,112,31,206,31,100,31,7,31,114,31,199,31,83,31,223,31,108,31,148,31,148,30,48,31,88,31,214,31,40,31,40,30,175,31,60,31,54,31,54,30,158,31,158,30,64,31,237,31,244,31,202,31,179,31,251,31,30,31,55,31,55,30,55,29,52,31,241,31,80,31,164,31,195,31,195,30,206,31,193,31,193,30,193,29,71,31,14,31,179,31,179,30,113,31,232,31,232,30,188,31,193,31,220,31,158,31,8,31,12,31,108,31,142,31,128,31,198,31,198,30,220,31,221,31,221,30,91,31,202,31,27,31,134,31,1,31,99,31,240,31,234,31,234,30,204,31,67,31,67,30,205,31,205,30,205,29,237,31,69,31,69,30,80,31,80,30,80,29,238,31,232,31,54,31,55,31,245,31,44,31,64,31,64,30,80,31,110,31,3,31,3,30,90,31,62,31,62,30,205,31,146,31,158,31,138,31,140,31,176,31,253,31,93,31,76,31,246,31,95,31,5,31,55,31,116,31,164,31,17,31,93,31,110,31,158,31,158,30,105,31,202,31,202,30,180,31,25,31,25,30,14,31,14,30,176,31,225,31,225,30,239,31,148,31,164,31,171,31,171,31,98,31,115,31,15,31,54,31,220,31,220,30,64,31,64,30,64,29,64,28,64,27,34,31,34,30,167,31,252,31,111,31,64,31,213,31,62,31,127,31,43,31,82,31,171,31,171,30,140,31,179,31,212,31,250,31,56,31,139,31,188,31,160,31,29,31,29,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
