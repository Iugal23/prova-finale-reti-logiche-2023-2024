-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 518;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (61,0,158,0,253,0,111,0,0,0,178,0,52,0,174,0,19,0,0,0,0,0,0,0,54,0,20,0,110,0,40,0,250,0,130,0,68,0,39,0,185,0,229,0,197,0,105,0,0,0,197,0,239,0,185,0,132,0,117,0,182,0,0,0,216,0,153,0,153,0,0,0,250,0,34,0,0,0,113,0,106,0,121,0,161,0,98,0,54,0,0,0,130,0,57,0,174,0,64,0,179,0,179,0,64,0,87,0,196,0,78,0,217,0,33,0,52,0,0,0,106,0,240,0,156,0,37,0,174,0,224,0,139,0,0,0,0,0,129,0,30,0,167,0,0,0,42,0,204,0,0,0,22,0,20,0,100,0,17,0,54,0,35,0,0,0,20,0,68,0,139,0,230,0,101,0,97,0,196,0,0,0,229,0,129,0,0,0,166,0,134,0,22,0,250,0,33,0,0,0,238,0,116,0,42,0,11,0,31,0,167,0,118,0,86,0,119,0,169,0,44,0,2,0,0,0,200,0,174,0,177,0,222,0,105,0,0,0,15,0,0,0,29,0,10,0,156,0,23,0,226,0,147,0,26,0,107,0,220,0,4,0,64,0,147,0,202,0,183,0,137,0,57,0,82,0,137,0,179,0,139,0,239,0,0,0,0,0,104,0,188,0,215,0,90,0,196,0,254,0,178,0,59,0,85,0,0,0,166,0,0,0,16,0,73,0,148,0,10,0,244,0,235,0,0,0,15,0,0,0,151,0,0,0,212,0,0,0,163,0,173,0,3,0,74,0,0,0,137,0,54,0,70,0,237,0,216,0,50,0,237,0,0,0,67,0,120,0,83,0,0,0,157,0,30,0,94,0,138,0,0,0,158,0,114,0,214,0,16,0,213,0,0,0,151,0,102,0,28,0,98,0,247,0,106,0,61,0,0,0,108,0,103,0,0,0,14,0,138,0,43,0,191,0,16,0,153,0,20,0,23,0,9,0,11,0,199,0,233,0,129,0,205,0,131,0,204,0,84,0,24,0,249,0,41,0,230,0,36,0,0,0,65,0,125,0,226,0,157,0,0,0,64,0,0,0,136,0,0,0,194,0,4,0,114,0,95,0,23,0,194,0,195,0,176,0,0,0,23,0,224,0,242,0,0,0,31,0,200,0,0,0,136,0,147,0,89,0,17,0,40,0,206,0,27,0,0,0,0,0,127,0,0,0,227,0,51,0,249,0,0,0,171,0,0,0,190,0,180,0,76,0,80,0,59,0,102,0,0,0,204,0,0,0,95,0,95,0,0,0,153,0,195,0,1,0,0,0,70,0,248,0,0,0,0,0,90,0,229,0,27,0,51,0,26,0,0,0,57,0,171,0,84,0,197,0,166,0,159,0,197,0,222,0,0,0,233,0,52,0,112,0,181,0,8,0,142,0,121,0,20,0,108,0,14,0,0,0,0,0,171,0,0,0,0,0,97,0,131,0,60,0,136,0,60,0,174,0,195,0,3,0,0,0,145,0,35,0,218,0,40,0,44,0,239,0,233,0,0,0,229,0,93,0,52,0,182,0,82,0,63,0,5,0,181,0,36,0,23,0,49,0,205,0,0,0,0,0,228,0,197,0,84,0,134,0,55,0,64,0,200,0,0,0,65,0,44,0,81,0,229,0,114,0,183,0,49,0,0,0,8,0,55,0,181,0,128,0,82,0,228,0,51,0,42,0,101,0,246,0,0,0,113,0,55,0,40,0,101,0,117,0,0,0,150,0,245,0,89,0,182,0,148,0,0,0,224,0,18,0,7,0,0,0,25,0,79,0,241,0,63,0,141,0,132,0,173,0,241,0,0,0,155,0,204,0,0,0,195,0,66,0,183,0,79,0,76,0,246,0,58,0,114,0,43,0,151,0,75,0,117,0,23,0,0,0,10,0,179,0,46,0,138,0,0,0,235,0,194,0,252,0,178,0,25,0,147,0,0,0,202,0,55,0,21,0,161,0,0,0,45,0,114,0,185,0,60,0,227,0,53,0,224,0,0,0,12,0,0,0,39,0,49,0,0,0,31,0,71,0,66,0,192,0,124,0,114,0,251,0,30,0,169,0,117,0,0,0,10,0,9,0,66,0,255,0,100,0,149,0,233,0,18,0,32,0,145,0,0,0,105,0,175,0,37,0,250,0,58,0,140,0,0,0,0,0,54,0,190,0,169,0,197,0,102,0,141,0,25,0,0,0,74,0,243,0,0,0,133,0,0,0,38,0,103,0,0,0,156,0,0,0,192,0,94,0,221,0,44,0,117,0,65,0,0,0,133,0,33,0,222,0,157,0,2,0,76,0,251,0,155,0,10,0,206,0);
signal scenario_full  : scenario_type := (61,31,158,31,253,31,111,31,111,30,178,31,52,31,174,31,19,31,19,30,19,29,19,28,54,31,20,31,110,31,40,31,250,31,130,31,68,31,39,31,185,31,229,31,197,31,105,31,105,30,197,31,239,31,185,31,132,31,117,31,182,31,182,30,216,31,153,31,153,31,153,30,250,31,34,31,34,30,113,31,106,31,121,31,161,31,98,31,54,31,54,30,130,31,57,31,174,31,64,31,179,31,179,31,64,31,87,31,196,31,78,31,217,31,33,31,52,31,52,30,106,31,240,31,156,31,37,31,174,31,224,31,139,31,139,30,139,29,129,31,30,31,167,31,167,30,42,31,204,31,204,30,22,31,20,31,100,31,17,31,54,31,35,31,35,30,20,31,68,31,139,31,230,31,101,31,97,31,196,31,196,30,229,31,129,31,129,30,166,31,134,31,22,31,250,31,33,31,33,30,238,31,116,31,42,31,11,31,31,31,167,31,118,31,86,31,119,31,169,31,44,31,2,31,2,30,200,31,174,31,177,31,222,31,105,31,105,30,15,31,15,30,29,31,10,31,156,31,23,31,226,31,147,31,26,31,107,31,220,31,4,31,64,31,147,31,202,31,183,31,137,31,57,31,82,31,137,31,179,31,139,31,239,31,239,30,239,29,104,31,188,31,215,31,90,31,196,31,254,31,178,31,59,31,85,31,85,30,166,31,166,30,16,31,73,31,148,31,10,31,244,31,235,31,235,30,15,31,15,30,151,31,151,30,212,31,212,30,163,31,173,31,3,31,74,31,74,30,137,31,54,31,70,31,237,31,216,31,50,31,237,31,237,30,67,31,120,31,83,31,83,30,157,31,30,31,94,31,138,31,138,30,158,31,114,31,214,31,16,31,213,31,213,30,151,31,102,31,28,31,98,31,247,31,106,31,61,31,61,30,108,31,103,31,103,30,14,31,138,31,43,31,191,31,16,31,153,31,20,31,23,31,9,31,11,31,199,31,233,31,129,31,205,31,131,31,204,31,84,31,24,31,249,31,41,31,230,31,36,31,36,30,65,31,125,31,226,31,157,31,157,30,64,31,64,30,136,31,136,30,194,31,4,31,114,31,95,31,23,31,194,31,195,31,176,31,176,30,23,31,224,31,242,31,242,30,31,31,200,31,200,30,136,31,147,31,89,31,17,31,40,31,206,31,27,31,27,30,27,29,127,31,127,30,227,31,51,31,249,31,249,30,171,31,171,30,190,31,180,31,76,31,80,31,59,31,102,31,102,30,204,31,204,30,95,31,95,31,95,30,153,31,195,31,1,31,1,30,70,31,248,31,248,30,248,29,90,31,229,31,27,31,51,31,26,31,26,30,57,31,171,31,84,31,197,31,166,31,159,31,197,31,222,31,222,30,233,31,52,31,112,31,181,31,8,31,142,31,121,31,20,31,108,31,14,31,14,30,14,29,171,31,171,30,171,29,97,31,131,31,60,31,136,31,60,31,174,31,195,31,3,31,3,30,145,31,35,31,218,31,40,31,44,31,239,31,233,31,233,30,229,31,93,31,52,31,182,31,82,31,63,31,5,31,181,31,36,31,23,31,49,31,205,31,205,30,205,29,228,31,197,31,84,31,134,31,55,31,64,31,200,31,200,30,65,31,44,31,81,31,229,31,114,31,183,31,49,31,49,30,8,31,55,31,181,31,128,31,82,31,228,31,51,31,42,31,101,31,246,31,246,30,113,31,55,31,40,31,101,31,117,31,117,30,150,31,245,31,89,31,182,31,148,31,148,30,224,31,18,31,7,31,7,30,25,31,79,31,241,31,63,31,141,31,132,31,173,31,241,31,241,30,155,31,204,31,204,30,195,31,66,31,183,31,79,31,76,31,246,31,58,31,114,31,43,31,151,31,75,31,117,31,23,31,23,30,10,31,179,31,46,31,138,31,138,30,235,31,194,31,252,31,178,31,25,31,147,31,147,30,202,31,55,31,21,31,161,31,161,30,45,31,114,31,185,31,60,31,227,31,53,31,224,31,224,30,12,31,12,30,39,31,49,31,49,30,31,31,71,31,66,31,192,31,124,31,114,31,251,31,30,31,169,31,117,31,117,30,10,31,9,31,66,31,255,31,100,31,149,31,233,31,18,31,32,31,145,31,145,30,105,31,175,31,37,31,250,31,58,31,140,31,140,30,140,29,54,31,190,31,169,31,197,31,102,31,141,31,25,31,25,30,74,31,243,31,243,30,133,31,133,30,38,31,103,31,103,30,156,31,156,30,192,31,94,31,221,31,44,31,117,31,65,31,65,30,133,31,33,31,222,31,157,31,2,31,76,31,251,31,155,31,10,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
