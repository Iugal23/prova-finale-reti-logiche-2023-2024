-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_88 is
end project_tb_88;

architecture project_tb_arch_88 of project_tb_88 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 241;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (198,0,128,0,8,0,204,0,180,0,229,0,197,0,246,0,22,0,90,0,2,0,0,0,0,0,235,0,17,0,27,0,0,0,118,0,113,0,216,0,8,0,75,0,5,0,0,0,0,0,156,0,54,0,43,0,21,0,251,0,151,0,195,0,0,0,52,0,217,0,0,0,51,0,196,0,0,0,180,0,158,0,254,0,246,0,8,0,118,0,0,0,251,0,200,0,179,0,0,0,130,0,185,0,22,0,0,0,74,0,0,0,218,0,33,0,0,0,0,0,0,0,247,0,111,0,204,0,199,0,191,0,123,0,4,0,73,0,0,0,140,0,16,0,83,0,178,0,0,0,168,0,0,0,162,0,6,0,0,0,56,0,6,0,251,0,0,0,133,0,84,0,36,0,116,0,18,0,247,0,146,0,0,0,104,0,112,0,0,0,232,0,226,0,83,0,90,0,0,0,97,0,126,0,0,0,0,0,0,0,146,0,30,0,172,0,0,0,0,0,62,0,0,0,0,0,0,0,191,0,192,0,99,0,18,0,66,0,150,0,117,0,214,0,144,0,105,0,77,0,158,0,228,0,250,0,2,0,0,0,249,0,33,0,0,0,1,0,160,0,0,0,146,0,0,0,0,0,171,0,206,0,7,0,166,0,15,0,235,0,81,0,180,0,101,0,94,0,0,0,231,0,10,0,8,0,36,0,0,0,63,0,67,0,71,0,14,0,0,0,76,0,12,0,0,0,143,0,139,0,246,0,0,0,52,0,94,0,227,0,44,0,235,0,0,0,122,0,0,0,137,0,14,0,129,0,0,0,16,0,165,0,99,0,1,0,0,0,130,0,0,0,32,0,237,0,206,0,37,0,0,0,92,0,2,0,59,0,179,0,138,0,62,0,0,0,228,0,68,0,0,0,42,0,61,0,11,0,0,0,0,0,228,0,39,0,0,0,0,0,0,0,0,0,130,0,84,0,69,0,0,0,28,0,177,0,119,0,75,0,0,0,155,0,242,0,36,0,0,0,0,0,0,0,73,0,53,0,94,0,233,0,201,0,186,0,246,0,103,0,206,0,245,0,156,0,136,0,166,0,116,0);
signal scenario_full  : scenario_type := (198,31,128,31,8,31,204,31,180,31,229,31,197,31,246,31,22,31,90,31,2,31,2,30,2,29,235,31,17,31,27,31,27,30,118,31,113,31,216,31,8,31,75,31,5,31,5,30,5,29,156,31,54,31,43,31,21,31,251,31,151,31,195,31,195,30,52,31,217,31,217,30,51,31,196,31,196,30,180,31,158,31,254,31,246,31,8,31,118,31,118,30,251,31,200,31,179,31,179,30,130,31,185,31,22,31,22,30,74,31,74,30,218,31,33,31,33,30,33,29,33,28,247,31,111,31,204,31,199,31,191,31,123,31,4,31,73,31,73,30,140,31,16,31,83,31,178,31,178,30,168,31,168,30,162,31,6,31,6,30,56,31,6,31,251,31,251,30,133,31,84,31,36,31,116,31,18,31,247,31,146,31,146,30,104,31,112,31,112,30,232,31,226,31,83,31,90,31,90,30,97,31,126,31,126,30,126,29,126,28,146,31,30,31,172,31,172,30,172,29,62,31,62,30,62,29,62,28,191,31,192,31,99,31,18,31,66,31,150,31,117,31,214,31,144,31,105,31,77,31,158,31,228,31,250,31,2,31,2,30,249,31,33,31,33,30,1,31,160,31,160,30,146,31,146,30,146,29,171,31,206,31,7,31,166,31,15,31,235,31,81,31,180,31,101,31,94,31,94,30,231,31,10,31,8,31,36,31,36,30,63,31,67,31,71,31,14,31,14,30,76,31,12,31,12,30,143,31,139,31,246,31,246,30,52,31,94,31,227,31,44,31,235,31,235,30,122,31,122,30,137,31,14,31,129,31,129,30,16,31,165,31,99,31,1,31,1,30,130,31,130,30,32,31,237,31,206,31,37,31,37,30,92,31,2,31,59,31,179,31,138,31,62,31,62,30,228,31,68,31,68,30,42,31,61,31,11,31,11,30,11,29,228,31,39,31,39,30,39,29,39,28,39,27,130,31,84,31,69,31,69,30,28,31,177,31,119,31,75,31,75,30,155,31,242,31,36,31,36,30,36,29,36,28,73,31,53,31,94,31,233,31,201,31,186,31,246,31,103,31,206,31,245,31,156,31,136,31,166,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
