-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 819;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,0,0,171,0,171,0,0,0,220,0,158,0,196,0,91,0,0,0,155,0,0,0,0,0,0,0,27,0,124,0,43,0,136,0,67,0,129,0,128,0,0,0,151,0,203,0,69,0,75,0,70,0,0,0,47,0,212,0,0,0,198,0,0,0,168,0,83,0,169,0,0,0,216,0,172,0,160,0,159,0,108,0,77,0,32,0,53,0,85,0,0,0,158,0,185,0,117,0,0,0,0,0,0,0,0,0,222,0,253,0,161,0,177,0,178,0,187,0,139,0,6,0,221,0,129,0,0,0,122,0,94,0,239,0,0,0,155,0,138,0,90,0,204,0,10,0,237,0,0,0,46,0,84,0,26,0,0,0,121,0,0,0,243,0,0,0,0,0,169,0,116,0,148,0,230,0,0,0,146,0,189,0,85,0,197,0,62,0,35,0,127,0,0,0,142,0,32,0,0,0,40,0,131,0,176,0,110,0,91,0,0,0,238,0,0,0,67,0,169,0,28,0,65,0,187,0,147,0,100,0,0,0,150,0,0,0,239,0,254,0,20,0,186,0,24,0,96,0,0,0,215,0,64,0,0,0,76,0,83,0,181,0,0,0,101,0,155,0,227,0,158,0,0,0,235,0,102,0,214,0,0,0,42,0,0,0,44,0,137,0,101,0,114,0,114,0,67,0,240,0,0,0,127,0,176,0,0,0,0,0,33,0,0,0,51,0,0,0,116,0,80,0,40,0,105,0,178,0,121,0,68,0,84,0,25,0,43,0,0,0,236,0,227,0,228,0,150,0,220,0,0,0,206,0,103,0,57,0,0,0,148,0,162,0,0,0,0,0,74,0,34,0,117,0,198,0,228,0,111,0,149,0,5,0,95,0,0,0,189,0,6,0,184,0,118,0,163,0,203,0,156,0,103,0,125,0,202,0,0,0,40,0,198,0,220,0,198,0,0,0,0,0,0,0,111,0,215,0,40,0,0,0,81,0,9,0,171,0,201,0,36,0,81,0,147,0,236,0,9,0,253,0,240,0,61,0,130,0,207,0,0,0,148,0,226,0,173,0,108,0,222,0,245,0,18,0,224,0,193,0,37,0,0,0,18,0,108,0,249,0,149,0,201,0,118,0,180,0,174,0,15,0,224,0,33,0,213,0,229,0,213,0,244,0,53,0,0,0,214,0,54,0,118,0,84,0,0,0,155,0,100,0,179,0,75,0,65,0,0,0,117,0,0,0,191,0,0,0,151,0,176,0,249,0,170,0,25,0,51,0,209,0,36,0,149,0,46,0,33,0,20,0,196,0,229,0,109,0,7,0,208,0,0,0,45,0,45,0,0,0,183,0,128,0,156,0,114,0,87,0,172,0,8,0,30,0,177,0,203,0,168,0,0,0,55,0,199,0,187,0,135,0,37,0,97,0,198,0,138,0,141,0,152,0,0,0,153,0,85,0,237,0,215,0,5,0,91,0,92,0,136,0,153,0,0,0,221,0,77,0,15,0,0,0,0,0,101,0,145,0,133,0,229,0,37,0,225,0,0,0,140,0,23,0,210,0,199,0,0,0,0,0,93,0,37,0,61,0,21,0,0,0,0,0,74,0,108,0,81,0,103,0,61,0,113,0,0,0,1,0,253,0,254,0,175,0,185,0,144,0,90,0,72,0,223,0,83,0,253,0,0,0,77,0,200,0,72,0,13,0,76,0,176,0,0,0,243,0,65,0,172,0,0,0,128,0,139,0,17,0,0,0,0,0,245,0,52,0,250,0,208,0,162,0,157,0,115,0,0,0,175,0,200,0,0,0,194,0,145,0,27,0,0,0,162,0,92,0,218,0,91,0,0,0,0,0,251,0,0,0,134,0,77,0,138,0,171,0,50,0,0,0,18,0,215,0,103,0,14,0,25,0,33,0,148,0,136,0,45,0,0,0,0,0,0,0,0,0,105,0,0,0,118,0,29,0,62,0,221,0,251,0,198,0,207,0,164,0,28,0,5,0,120,0,195,0,166,0,0,0,0,0,0,0,69,0,0,0,0,0,126,0,118,0,63,0,204,0,202,0,0,0,0,0,0,0,147,0,96,0,149,0,201,0,0,0,31,0,153,0,3,0,4,0,176,0,96,0,0,0,0,0,240,0,88,0,167,0,45,0,52,0,251,0,12,0,230,0,4,0,0,0,3,0,0,0,137,0,121,0,53,0,0,0,141,0,101,0,183,0,238,0,254,0,161,0,86,0,201,0,156,0,107,0,38,0,148,0,230,0,21,0,187,0,0,0,82,0,58,0,0,0,40,0,0,0,38,0,127,0,73,0,169,0,0,0,163,0,77,0,164,0,214,0,123,0,84,0,61,0,0,0,0,0,4,0,30,0,155,0,242,0,238,0,237,0,212,0,134,0,0,0,213,0,109,0,143,0,111,0,0,0,78,0,231,0,198,0,239,0,202,0,0,0,84,0,17,0,129,0,20,0,0,0,0,0,0,0,0,0,117,0,89,0,182,0,20,0,101,0,206,0,243,0,25,0,26,0,243,0,197,0,0,0,183,0,139,0,48,0,48,0,2,0,137,0,188,0,197,0,0,0,11,0,231,0,252,0,94,0,59,0,139,0,0,0,77,0,58,0,107,0,169,0,139,0,0,0,0,0,50,0,0,0,0,0,204,0,48,0,0,0,116,0,0,0,40,0,93,0,80,0,0,0,128,0,140,0,96,0,61,0,248,0,8,0,0,0,90,0,0,0,205,0,153,0,108,0,225,0,72,0,0,0,144,0,145,0,106,0,0,0,169,0,0,0,86,0,250,0,0,0,248,0,12,0,0,0,26,0,17,0,216,0,255,0,151,0,76,0,162,0,0,0,36,0,0,0,161,0,32,0,17,0,234,0,166,0,111,0,33,0,235,0,210,0,75,0,185,0,210,0,206,0,93,0,58,0,171,0,159,0,134,0,0,0,90,0,114,0,0,0,16,0,82,0,122,0,138,0,26,0,31,0,159,0,191,0,0,0,227,0,138,0,3,0,184,0,131,0,31,0,100,0,73,0,94,0,0,0,6,0,194,0,94,0,123,0,112,0,197,0,80,0,0,0,23,0,101,0,131,0,97,0,237,0,0,0,0,0,98,0,235,0,144,0,137,0,99,0,45,0,0,0,93,0,246,0,122,0,69,0,27,0,212,0,36,0,152,0,139,0,120,0,227,0,120,0,35,0,41,0,208,0,136,0,4,0,66,0,249,0,0,0,170,0,52,0,189,0,69,0,92,0,90,0,79,0,154,0,165,0,131,0,209,0,186,0,0,0,65,0,0,0,223,0,37,0,149,0,197,0,231,0,174,0,64,0,248,0,28,0,26,0,104,0,36,0,9,0,0,0,0,0,148,0,219,0,87,0,60,0,175,0,0,0,116,0,21,0,156,0,190,0,219,0,0,0,0,0,129,0,212,0,222,0,113,0,113,0,125,0,220,0,139,0,55,0,201,0,0,0,151,0,117,0,0,0,172,0,0,0,85,0,0,0,0,0,84,0,92,0,10,0,190,0,17,0,92,0,174,0,200,0,160,0,130,0,6,0,18,0,0,0,96,0,144,0,0,0,10,0,40,0,18,0,194,0,0,0,93,0,209,0,31,0,15,0,0,0,187,0,176,0,83,0,0,0,123,0,224,0,140,0,107,0,191,0,111,0,145,0,151,0,141,0);
signal scenario_full  : scenario_type := (250,31,250,30,171,31,171,31,171,30,220,31,158,31,196,31,91,31,91,30,155,31,155,30,155,29,155,28,27,31,124,31,43,31,136,31,67,31,129,31,128,31,128,30,151,31,203,31,69,31,75,31,70,31,70,30,47,31,212,31,212,30,198,31,198,30,168,31,83,31,169,31,169,30,216,31,172,31,160,31,159,31,108,31,77,31,32,31,53,31,85,31,85,30,158,31,185,31,117,31,117,30,117,29,117,28,117,27,222,31,253,31,161,31,177,31,178,31,187,31,139,31,6,31,221,31,129,31,129,30,122,31,94,31,239,31,239,30,155,31,138,31,90,31,204,31,10,31,237,31,237,30,46,31,84,31,26,31,26,30,121,31,121,30,243,31,243,30,243,29,169,31,116,31,148,31,230,31,230,30,146,31,189,31,85,31,197,31,62,31,35,31,127,31,127,30,142,31,32,31,32,30,40,31,131,31,176,31,110,31,91,31,91,30,238,31,238,30,67,31,169,31,28,31,65,31,187,31,147,31,100,31,100,30,150,31,150,30,239,31,254,31,20,31,186,31,24,31,96,31,96,30,215,31,64,31,64,30,76,31,83,31,181,31,181,30,101,31,155,31,227,31,158,31,158,30,235,31,102,31,214,31,214,30,42,31,42,30,44,31,137,31,101,31,114,31,114,31,67,31,240,31,240,30,127,31,176,31,176,30,176,29,33,31,33,30,51,31,51,30,116,31,80,31,40,31,105,31,178,31,121,31,68,31,84,31,25,31,43,31,43,30,236,31,227,31,228,31,150,31,220,31,220,30,206,31,103,31,57,31,57,30,148,31,162,31,162,30,162,29,74,31,34,31,117,31,198,31,228,31,111,31,149,31,5,31,95,31,95,30,189,31,6,31,184,31,118,31,163,31,203,31,156,31,103,31,125,31,202,31,202,30,40,31,198,31,220,31,198,31,198,30,198,29,198,28,111,31,215,31,40,31,40,30,81,31,9,31,171,31,201,31,36,31,81,31,147,31,236,31,9,31,253,31,240,31,61,31,130,31,207,31,207,30,148,31,226,31,173,31,108,31,222,31,245,31,18,31,224,31,193,31,37,31,37,30,18,31,108,31,249,31,149,31,201,31,118,31,180,31,174,31,15,31,224,31,33,31,213,31,229,31,213,31,244,31,53,31,53,30,214,31,54,31,118,31,84,31,84,30,155,31,100,31,179,31,75,31,65,31,65,30,117,31,117,30,191,31,191,30,151,31,176,31,249,31,170,31,25,31,51,31,209,31,36,31,149,31,46,31,33,31,20,31,196,31,229,31,109,31,7,31,208,31,208,30,45,31,45,31,45,30,183,31,128,31,156,31,114,31,87,31,172,31,8,31,30,31,177,31,203,31,168,31,168,30,55,31,199,31,187,31,135,31,37,31,97,31,198,31,138,31,141,31,152,31,152,30,153,31,85,31,237,31,215,31,5,31,91,31,92,31,136,31,153,31,153,30,221,31,77,31,15,31,15,30,15,29,101,31,145,31,133,31,229,31,37,31,225,31,225,30,140,31,23,31,210,31,199,31,199,30,199,29,93,31,37,31,61,31,21,31,21,30,21,29,74,31,108,31,81,31,103,31,61,31,113,31,113,30,1,31,253,31,254,31,175,31,185,31,144,31,90,31,72,31,223,31,83,31,253,31,253,30,77,31,200,31,72,31,13,31,76,31,176,31,176,30,243,31,65,31,172,31,172,30,128,31,139,31,17,31,17,30,17,29,245,31,52,31,250,31,208,31,162,31,157,31,115,31,115,30,175,31,200,31,200,30,194,31,145,31,27,31,27,30,162,31,92,31,218,31,91,31,91,30,91,29,251,31,251,30,134,31,77,31,138,31,171,31,50,31,50,30,18,31,215,31,103,31,14,31,25,31,33,31,148,31,136,31,45,31,45,30,45,29,45,28,45,27,105,31,105,30,118,31,29,31,62,31,221,31,251,31,198,31,207,31,164,31,28,31,5,31,120,31,195,31,166,31,166,30,166,29,166,28,69,31,69,30,69,29,126,31,118,31,63,31,204,31,202,31,202,30,202,29,202,28,147,31,96,31,149,31,201,31,201,30,31,31,153,31,3,31,4,31,176,31,96,31,96,30,96,29,240,31,88,31,167,31,45,31,52,31,251,31,12,31,230,31,4,31,4,30,3,31,3,30,137,31,121,31,53,31,53,30,141,31,101,31,183,31,238,31,254,31,161,31,86,31,201,31,156,31,107,31,38,31,148,31,230,31,21,31,187,31,187,30,82,31,58,31,58,30,40,31,40,30,38,31,127,31,73,31,169,31,169,30,163,31,77,31,164,31,214,31,123,31,84,31,61,31,61,30,61,29,4,31,30,31,155,31,242,31,238,31,237,31,212,31,134,31,134,30,213,31,109,31,143,31,111,31,111,30,78,31,231,31,198,31,239,31,202,31,202,30,84,31,17,31,129,31,20,31,20,30,20,29,20,28,20,27,117,31,89,31,182,31,20,31,101,31,206,31,243,31,25,31,26,31,243,31,197,31,197,30,183,31,139,31,48,31,48,31,2,31,137,31,188,31,197,31,197,30,11,31,231,31,252,31,94,31,59,31,139,31,139,30,77,31,58,31,107,31,169,31,139,31,139,30,139,29,50,31,50,30,50,29,204,31,48,31,48,30,116,31,116,30,40,31,93,31,80,31,80,30,128,31,140,31,96,31,61,31,248,31,8,31,8,30,90,31,90,30,205,31,153,31,108,31,225,31,72,31,72,30,144,31,145,31,106,31,106,30,169,31,169,30,86,31,250,31,250,30,248,31,12,31,12,30,26,31,17,31,216,31,255,31,151,31,76,31,162,31,162,30,36,31,36,30,161,31,32,31,17,31,234,31,166,31,111,31,33,31,235,31,210,31,75,31,185,31,210,31,206,31,93,31,58,31,171,31,159,31,134,31,134,30,90,31,114,31,114,30,16,31,82,31,122,31,138,31,26,31,31,31,159,31,191,31,191,30,227,31,138,31,3,31,184,31,131,31,31,31,100,31,73,31,94,31,94,30,6,31,194,31,94,31,123,31,112,31,197,31,80,31,80,30,23,31,101,31,131,31,97,31,237,31,237,30,237,29,98,31,235,31,144,31,137,31,99,31,45,31,45,30,93,31,246,31,122,31,69,31,27,31,212,31,36,31,152,31,139,31,120,31,227,31,120,31,35,31,41,31,208,31,136,31,4,31,66,31,249,31,249,30,170,31,52,31,189,31,69,31,92,31,90,31,79,31,154,31,165,31,131,31,209,31,186,31,186,30,65,31,65,30,223,31,37,31,149,31,197,31,231,31,174,31,64,31,248,31,28,31,26,31,104,31,36,31,9,31,9,30,9,29,148,31,219,31,87,31,60,31,175,31,175,30,116,31,21,31,156,31,190,31,219,31,219,30,219,29,129,31,212,31,222,31,113,31,113,31,125,31,220,31,139,31,55,31,201,31,201,30,151,31,117,31,117,30,172,31,172,30,85,31,85,30,85,29,84,31,92,31,10,31,190,31,17,31,92,31,174,31,200,31,160,31,130,31,6,31,18,31,18,30,96,31,144,31,144,30,10,31,40,31,18,31,194,31,194,30,93,31,209,31,31,31,15,31,15,30,187,31,176,31,83,31,83,30,123,31,224,31,140,31,107,31,191,31,111,31,145,31,151,31,141,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
