-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 301;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,241,0,220,0,0,0,203,0,0,0,41,0,30,0,186,0,61,0,42,0,78,0,70,0,215,0,108,0,226,0,224,0,153,0,61,0,205,0,225,0,145,0,0,0,1,0,98,0,75,0,28,0,220,0,0,0,53,0,248,0,139,0,164,0,192,0,196,0,115,0,199,0,96,0,202,0,139,0,158,0,38,0,0,0,149,0,123,0,162,0,61,0,9,0,0,0,203,0,188,0,12,0,29,0,0,0,211,0,171,0,41,0,106,0,0,0,105,0,41,0,11,0,17,0,186,0,0,0,151,0,102,0,221,0,121,0,58,0,0,0,214,0,31,0,61,0,216,0,15,0,52,0,147,0,123,0,54,0,137,0,158,0,149,0,41,0,182,0,0,0,0,0,155,0,0,0,11,0,220,0,0,0,185,0,238,0,1,0,215,0,0,0,229,0,27,0,105,0,0,0,93,0,183,0,165,0,206,0,30,0,223,0,0,0,80,0,163,0,126,0,13,0,58,0,0,0,0,0,233,0,191,0,224,0,0,0,36,0,64,0,196,0,208,0,67,0,134,0,103,0,12,0,198,0,60,0,218,0,180,0,191,0,163,0,0,0,0,0,0,0,14,0,244,0,241,0,18,0,66,0,57,0,209,0,164,0,169,0,202,0,236,0,129,0,0,0,37,0,132,0,228,0,140,0,209,0,202,0,0,0,74,0,179,0,157,0,6,0,184,0,97,0,0,0,0,0,64,0,8,0,58,0,108,0,0,0,142,0,141,0,189,0,233,0,169,0,0,0,182,0,67,0,50,0,214,0,199,0,232,0,245,0,62,0,30,0,137,0,42,0,44,0,37,0,236,0,130,0,206,0,0,0,110,0,179,0,97,0,232,0,158,0,237,0,0,0,0,0,79,0,0,0,168,0,245,0,248,0,26,0,191,0,30,0,25,0,0,0,202,0,164,0,250,0,0,0,74,0,37,0,174,0,49,0,228,0,188,0,0,0,0,0,248,0,5,0,0,0,94,0,242,0,44,0,154,0,160,0,137,0,0,0,226,0,234,0,26,0,0,0,133,0,135,0,175,0,229,0,54,0,64,0,0,0,184,0,106,0,194,0,130,0,0,0,79,0,247,0,0,0,63,0,40,0,243,0,0,0,0,0,44,0,0,0,242,0,156,0,94,0,168,0,234,0,65,0,94,0,93,0,128,0,240,0,198,0,237,0,28,0,74,0,20,0,232,0,139,0,46,0,121,0,41,0,0,0,125,0,145,0,126,0,18,0,162,0,41,0,26,0,209,0,105,0,186,0,118,0,0,0,179,0,51,0,195,0,53,0,23,0,124,0,129,0,65,0,3,0,0,0);
signal scenario_full  : scenario_type := (0,0,241,31,220,31,220,30,203,31,203,30,41,31,30,31,186,31,61,31,42,31,78,31,70,31,215,31,108,31,226,31,224,31,153,31,61,31,205,31,225,31,145,31,145,30,1,31,98,31,75,31,28,31,220,31,220,30,53,31,248,31,139,31,164,31,192,31,196,31,115,31,199,31,96,31,202,31,139,31,158,31,38,31,38,30,149,31,123,31,162,31,61,31,9,31,9,30,203,31,188,31,12,31,29,31,29,30,211,31,171,31,41,31,106,31,106,30,105,31,41,31,11,31,17,31,186,31,186,30,151,31,102,31,221,31,121,31,58,31,58,30,214,31,31,31,61,31,216,31,15,31,52,31,147,31,123,31,54,31,137,31,158,31,149,31,41,31,182,31,182,30,182,29,155,31,155,30,11,31,220,31,220,30,185,31,238,31,1,31,215,31,215,30,229,31,27,31,105,31,105,30,93,31,183,31,165,31,206,31,30,31,223,31,223,30,80,31,163,31,126,31,13,31,58,31,58,30,58,29,233,31,191,31,224,31,224,30,36,31,64,31,196,31,208,31,67,31,134,31,103,31,12,31,198,31,60,31,218,31,180,31,191,31,163,31,163,30,163,29,163,28,14,31,244,31,241,31,18,31,66,31,57,31,209,31,164,31,169,31,202,31,236,31,129,31,129,30,37,31,132,31,228,31,140,31,209,31,202,31,202,30,74,31,179,31,157,31,6,31,184,31,97,31,97,30,97,29,64,31,8,31,58,31,108,31,108,30,142,31,141,31,189,31,233,31,169,31,169,30,182,31,67,31,50,31,214,31,199,31,232,31,245,31,62,31,30,31,137,31,42,31,44,31,37,31,236,31,130,31,206,31,206,30,110,31,179,31,97,31,232,31,158,31,237,31,237,30,237,29,79,31,79,30,168,31,245,31,248,31,26,31,191,31,30,31,25,31,25,30,202,31,164,31,250,31,250,30,74,31,37,31,174,31,49,31,228,31,188,31,188,30,188,29,248,31,5,31,5,30,94,31,242,31,44,31,154,31,160,31,137,31,137,30,226,31,234,31,26,31,26,30,133,31,135,31,175,31,229,31,54,31,64,31,64,30,184,31,106,31,194,31,130,31,130,30,79,31,247,31,247,30,63,31,40,31,243,31,243,30,243,29,44,31,44,30,242,31,156,31,94,31,168,31,234,31,65,31,94,31,93,31,128,31,240,31,198,31,237,31,28,31,74,31,20,31,232,31,139,31,46,31,121,31,41,31,41,30,125,31,145,31,126,31,18,31,162,31,41,31,26,31,209,31,105,31,186,31,118,31,118,30,179,31,51,31,195,31,53,31,23,31,124,31,129,31,65,31,3,31,3,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
