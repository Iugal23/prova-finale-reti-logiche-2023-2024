-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 364;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,0,0,0,0,66,0,251,0,215,0,0,0,0,0,79,0,239,0,0,0,103,0,205,0,0,0,0,0,162,0,3,0,24,0,167,0,0,0,54,0,251,0,107,0,92,0,0,0,0,0,151,0,29,0,182,0,70,0,111,0,123,0,62,0,204,0,60,0,169,0,36,0,0,0,77,0,0,0,0,0,0,0,0,0,133,0,191,0,0,0,99,0,0,0,165,0,0,0,238,0,0,0,200,0,36,0,4,0,187,0,251,0,5,0,89,0,0,0,242,0,0,0,73,0,238,0,2,0,221,0,239,0,249,0,0,0,159,0,26,0,176,0,75,0,0,0,19,0,190,0,20,0,0,0,73,0,107,0,0,0,235,0,116,0,43,0,173,0,78,0,255,0,0,0,236,0,93,0,66,0,20,0,238,0,125,0,192,0,0,0,143,0,97,0,196,0,92,0,170,0,0,0,217,0,0,0,162,0,210,0,19,0,118,0,42,0,76,0,176,0,45,0,39,0,191,0,182,0,162,0,127,0,47,0,0,0,51,0,245,0,96,0,4,0,183,0,101,0,125,0,227,0,221,0,240,0,0,0,18,0,19,0,216,0,52,0,92,0,0,0,0,0,248,0,190,0,162,0,25,0,112,0,228,0,16,0,0,0,22,0,138,0,0,0,75,0,180,0,0,0,181,0,118,0,167,0,0,0,0,0,125,0,155,0,201,0,147,0,169,0,151,0,46,0,53,0,23,0,162,0,29,0,233,0,73,0,122,0,123,0,2,0,218,0,230,0,105,0,19,0,127,0,134,0,39,0,14,0,235,0,0,0,181,0,172,0,0,0,210,0,121,0,0,0,198,0,138,0,178,0,30,0,19,0,0,0,0,0,86,0,198,0,166,0,45,0,111,0,86,0,0,0,6,0,163,0,183,0,4,0,157,0,0,0,205,0,14,0,51,0,32,0,16,0,243,0,167,0,10,0,197,0,0,0,0,0,0,0,0,0,0,0,181,0,80,0,0,0,87,0,250,0,42,0,220,0,230,0,0,0,66,0,0,0,25,0,99,0,172,0,41,0,37,0,185,0,233,0,189,0,200,0,75,0,211,0,249,0,164,0,218,0,39,0,213,0,192,0,30,0,193,0,135,0,53,0,21,0,52,0,0,0,158,0,251,0,0,0,238,0,140,0,180,0,0,0,0,0,6,0,135,0,2,0,118,0,0,0,223,0,103,0,211,0,0,0,64,0,199,0,110,0,0,0,0,0,192,0,0,0,43,0,242,0,78,0,0,0,125,0,119,0,123,0,29,0,211,0,0,0,0,0,114,0,123,0,0,0,136,0,142,0,179,0,181,0,60,0,228,0,133,0,0,0,110,0,22,0,183,0,0,0,0,0,81,0,135,0,222,0,16,0,0,0,66,0,7,0,143,0,88,0,189,0,211,0,10,0,111,0,100,0,16,0,182,0,0,0,88,0,24,0,105,0,0,0,0,0,0,0,0,0,84,0,0,0,227,0,0,0,229,0,51,0,232,0,117,0,145,0,0,0,0,0,0,0,27,0,39,0,0,0,116,0,188,0,42,0,16,0,87,0,152,0,14,0,0,0,31,0,50,0,77,0,227,0,110,0,228,0,157,0,242,0,143,0);
signal scenario_full  : scenario_type := (69,31,69,30,69,29,66,31,251,31,215,31,215,30,215,29,79,31,239,31,239,30,103,31,205,31,205,30,205,29,162,31,3,31,24,31,167,31,167,30,54,31,251,31,107,31,92,31,92,30,92,29,151,31,29,31,182,31,70,31,111,31,123,31,62,31,204,31,60,31,169,31,36,31,36,30,77,31,77,30,77,29,77,28,77,27,133,31,191,31,191,30,99,31,99,30,165,31,165,30,238,31,238,30,200,31,36,31,4,31,187,31,251,31,5,31,89,31,89,30,242,31,242,30,73,31,238,31,2,31,221,31,239,31,249,31,249,30,159,31,26,31,176,31,75,31,75,30,19,31,190,31,20,31,20,30,73,31,107,31,107,30,235,31,116,31,43,31,173,31,78,31,255,31,255,30,236,31,93,31,66,31,20,31,238,31,125,31,192,31,192,30,143,31,97,31,196,31,92,31,170,31,170,30,217,31,217,30,162,31,210,31,19,31,118,31,42,31,76,31,176,31,45,31,39,31,191,31,182,31,162,31,127,31,47,31,47,30,51,31,245,31,96,31,4,31,183,31,101,31,125,31,227,31,221,31,240,31,240,30,18,31,19,31,216,31,52,31,92,31,92,30,92,29,248,31,190,31,162,31,25,31,112,31,228,31,16,31,16,30,22,31,138,31,138,30,75,31,180,31,180,30,181,31,118,31,167,31,167,30,167,29,125,31,155,31,201,31,147,31,169,31,151,31,46,31,53,31,23,31,162,31,29,31,233,31,73,31,122,31,123,31,2,31,218,31,230,31,105,31,19,31,127,31,134,31,39,31,14,31,235,31,235,30,181,31,172,31,172,30,210,31,121,31,121,30,198,31,138,31,178,31,30,31,19,31,19,30,19,29,86,31,198,31,166,31,45,31,111,31,86,31,86,30,6,31,163,31,183,31,4,31,157,31,157,30,205,31,14,31,51,31,32,31,16,31,243,31,167,31,10,31,197,31,197,30,197,29,197,28,197,27,197,26,181,31,80,31,80,30,87,31,250,31,42,31,220,31,230,31,230,30,66,31,66,30,25,31,99,31,172,31,41,31,37,31,185,31,233,31,189,31,200,31,75,31,211,31,249,31,164,31,218,31,39,31,213,31,192,31,30,31,193,31,135,31,53,31,21,31,52,31,52,30,158,31,251,31,251,30,238,31,140,31,180,31,180,30,180,29,6,31,135,31,2,31,118,31,118,30,223,31,103,31,211,31,211,30,64,31,199,31,110,31,110,30,110,29,192,31,192,30,43,31,242,31,78,31,78,30,125,31,119,31,123,31,29,31,211,31,211,30,211,29,114,31,123,31,123,30,136,31,142,31,179,31,181,31,60,31,228,31,133,31,133,30,110,31,22,31,183,31,183,30,183,29,81,31,135,31,222,31,16,31,16,30,66,31,7,31,143,31,88,31,189,31,211,31,10,31,111,31,100,31,16,31,182,31,182,30,88,31,24,31,105,31,105,30,105,29,105,28,105,27,84,31,84,30,227,31,227,30,229,31,51,31,232,31,117,31,145,31,145,30,145,29,145,28,27,31,39,31,39,30,116,31,188,31,42,31,16,31,87,31,152,31,14,31,14,30,31,31,50,31,77,31,227,31,110,31,228,31,157,31,242,31,143,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
