-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_49 is
end project_tb_49;

architecture project_tb_arch_49 of project_tb_49 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 225;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (146,0,150,0,59,0,19,0,236,0,5,0,0,0,49,0,0,0,132,0,32,0,0,0,199,0,247,0,142,0,163,0,241,0,168,0,200,0,178,0,156,0,104,0,218,0,229,0,104,0,216,0,197,0,219,0,0,0,2,0,168,0,68,0,230,0,69,0,193,0,0,0,0,0,113,0,224,0,81,0,0,0,2,0,156,0,9,0,133,0,0,0,234,0,186,0,0,0,84,0,202,0,188,0,102,0,46,0,98,0,0,0,74,0,67,0,101,0,176,0,198,0,90,0,163,0,165,0,217,0,97,0,0,0,233,0,168,0,0,0,192,0,145,0,119,0,10,0,66,0,143,0,204,0,42,0,136,0,202,0,14,0,129,0,41,0,138,0,50,0,0,0,0,0,249,0,221,0,153,0,0,0,161,0,22,0,169,0,120,0,0,0,46,0,0,0,100,0,255,0,89,0,204,0,65,0,80,0,0,0,131,0,0,0,158,0,0,0,0,0,137,0,25,0,133,0,89,0,151,0,133,0,54,0,0,0,200,0,72,0,174,0,162,0,248,0,31,0,148,0,78,0,82,0,96,0,0,0,155,0,246,0,242,0,45,0,255,0,241,0,126,0,74,0,191,0,112,0,0,0,241,0,213,0,153,0,129,0,0,0,203,0,177,0,0,0,156,0,0,0,103,0,22,0,47,0,217,0,132,0,40,0,192,0,35,0,134,0,93,0,54,0,238,0,0,0,0,0,73,0,36,0,74,0,0,0,82,0,0,0,220,0,147,0,102,0,11,0,19,0,247,0,117,0,178,0,109,0,0,0,56,0,57,0,54,0,70,0,85,0,151,0,249,0,156,0,0,0,188,0,221,0,103,0,0,0,64,0,125,0,77,0,72,0,243,0,70,0,30,0,240,0,125,0,0,0,234,0,110,0,157,0,210,0,112,0,244,0,0,0,236,0,97,0,79,0,147,0,0,0,67,0,74,0,121,0,164,0,183,0,77,0,194,0,14,0,0,0,9,0);
signal scenario_full  : scenario_type := (146,31,150,31,59,31,19,31,236,31,5,31,5,30,49,31,49,30,132,31,32,31,32,30,199,31,247,31,142,31,163,31,241,31,168,31,200,31,178,31,156,31,104,31,218,31,229,31,104,31,216,31,197,31,219,31,219,30,2,31,168,31,68,31,230,31,69,31,193,31,193,30,193,29,113,31,224,31,81,31,81,30,2,31,156,31,9,31,133,31,133,30,234,31,186,31,186,30,84,31,202,31,188,31,102,31,46,31,98,31,98,30,74,31,67,31,101,31,176,31,198,31,90,31,163,31,165,31,217,31,97,31,97,30,233,31,168,31,168,30,192,31,145,31,119,31,10,31,66,31,143,31,204,31,42,31,136,31,202,31,14,31,129,31,41,31,138,31,50,31,50,30,50,29,249,31,221,31,153,31,153,30,161,31,22,31,169,31,120,31,120,30,46,31,46,30,100,31,255,31,89,31,204,31,65,31,80,31,80,30,131,31,131,30,158,31,158,30,158,29,137,31,25,31,133,31,89,31,151,31,133,31,54,31,54,30,200,31,72,31,174,31,162,31,248,31,31,31,148,31,78,31,82,31,96,31,96,30,155,31,246,31,242,31,45,31,255,31,241,31,126,31,74,31,191,31,112,31,112,30,241,31,213,31,153,31,129,31,129,30,203,31,177,31,177,30,156,31,156,30,103,31,22,31,47,31,217,31,132,31,40,31,192,31,35,31,134,31,93,31,54,31,238,31,238,30,238,29,73,31,36,31,74,31,74,30,82,31,82,30,220,31,147,31,102,31,11,31,19,31,247,31,117,31,178,31,109,31,109,30,56,31,57,31,54,31,70,31,85,31,151,31,249,31,156,31,156,30,188,31,221,31,103,31,103,30,64,31,125,31,77,31,72,31,243,31,70,31,30,31,240,31,125,31,125,30,234,31,110,31,157,31,210,31,112,31,244,31,244,30,236,31,97,31,79,31,147,31,147,30,67,31,74,31,121,31,164,31,183,31,77,31,194,31,14,31,14,30,9,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
