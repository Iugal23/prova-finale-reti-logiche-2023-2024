-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_985 is
end project_tb_985;

architecture project_tb_arch_985 of project_tb_985 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 902;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (200,0,32,0,197,0,106,0,172,0,245,0,7,0,13,0,217,0,156,0,68,0,175,0,57,0,89,0,188,0,176,0,121,0,0,0,22,0,0,0,224,0,157,0,176,0,62,0,104,0,98,0,249,0,249,0,0,0,148,0,97,0,255,0,87,0,117,0,2,0,31,0,91,0,186,0,50,0,42,0,118,0,0,0,0,0,76,0,246,0,251,0,23,0,105,0,135,0,0,0,0,0,136,0,30,0,8,0,0,0,147,0,222,0,100,0,177,0,255,0,0,0,127,0,88,0,235,0,230,0,0,0,136,0,178,0,218,0,91,0,0,0,0,0,0,0,122,0,214,0,95,0,0,0,42,0,253,0,225,0,186,0,0,0,0,0,87,0,9,0,61,0,145,0,43,0,89,0,71,0,0,0,0,0,94,0,211,0,56,0,0,0,170,0,252,0,42,0,56,0,100,0,217,0,143,0,243,0,0,0,171,0,0,0,87,0,151,0,252,0,247,0,178,0,0,0,255,0,162,0,222,0,148,0,89,0,184,0,0,0,18,0,92,0,108,0,68,0,59,0,101,0,13,0,78,0,138,0,227,0,0,0,0,0,197,0,129,0,125,0,0,0,244,0,248,0,0,0,115,0,18,0,84,0,0,0,100,0,141,0,66,0,233,0,88,0,122,0,0,0,193,0,55,0,206,0,0,0,241,0,46,0,0,0,0,0,209,0,150,0,26,0,86,0,0,0,18,0,77,0,134,0,0,0,153,0,39,0,110,0,0,0,160,0,0,0,43,0,0,0,46,0,213,0,150,0,56,0,55,0,167,0,236,0,239,0,59,0,244,0,233,0,0,0,0,0,133,0,74,0,203,0,113,0,142,0,0,0,52,0,135,0,0,0,195,0,237,0,0,0,94,0,19,0,0,0,175,0,0,0,28,0,0,0,138,0,62,0,73,0,196,0,0,0,219,0,169,0,86,0,0,0,50,0,208,0,85,0,0,0,0,0,217,0,196,0,173,0,168,0,0,0,0,0,13,0,0,0,0,0,62,0,203,0,179,0,206,0,184,0,0,0,5,0,77,0,6,0,153,0,7,0,32,0,206,0,106,0,5,0,0,0,0,0,78,0,92,0,210,0,83,0,32,0,0,0,186,0,90,0,168,0,235,0,111,0,162,0,33,0,119,0,116,0,89,0,204,0,0,0,217,0,44,0,70,0,244,0,192,0,176,0,0,0,153,0,0,0,166,0,0,0,182,0,63,0,235,0,50,0,250,0,0,0,234,0,98,0,143,0,122,0,97,0,197,0,0,0,0,0,84,0,0,0,82,0,77,0,255,0,0,0,138,0,12,0,143,0,63,0,52,0,237,0,121,0,0,0,0,0,132,0,28,0,54,0,136,0,127,0,222,0,241,0,0,0,135,0,0,0,0,0,170,0,242,0,248,0,180,0,201,0,239,0,128,0,0,0,203,0,179,0,15,0,15,0,197,0,0,0,128,0,97,0,107,0,108,0,39,0,0,0,195,0,204,0,162,0,0,0,189,0,98,0,90,0,198,0,0,0,0,0,235,0,212,0,0,0,95,0,56,0,19,0,178,0,120,0,82,0,110,0,149,0,101,0,235,0,179,0,73,0,182,0,0,0,0,0,0,0,153,0,38,0,125,0,209,0,147,0,152,0,235,0,0,0,61,0,158,0,134,0,184,0,191,0,159,0,166,0,36,0,149,0,126,0,160,0,213,0,70,0,26,0,250,0,121,0,0,0,0,0,178,0,43,0,18,0,69,0,99,0,175,0,120,0,244,0,170,0,111,0,1,0,130,0,160,0,197,0,138,0,0,0,18,0,170,0,67,0,239,0,198,0,40,0,101,0,0,0,180,0,157,0,178,0,103,0,64,0,36,0,100,0,109,0,250,0,180,0,124,0,168,0,75,0,206,0,179,0,149,0,200,0,38,0,141,0,126,0,9,0,225,0,0,0,0,0,92,0,130,0,32,0,0,0,147,0,0,0,101,0,0,0,226,0,138,0,194,0,226,0,176,0,17,0,222,0,98,0,249,0,38,0,120,0,155,0,80,0,0,0,22,0,156,0,102,0,212,0,116,0,229,0,40,0,76,0,179,0,109,0,0,0,0,0,101,0,91,0,161,0,44,0,202,0,212,0,78,0,220,0,0,0,237,0,240,0,99,0,0,0,128,0,91,0,135,0,58,0,5,0,0,0,0,0,105,0,229,0,236,0,255,0,0,0,105,0,137,0,0,0,24,0,24,0,0,0,0,0,0,0,214,0,62,0,248,0,218,0,206,0,37,0,0,0,149,0,0,0,0,0,205,0,45,0,56,0,176,0,151,0,7,0,0,0,77,0,0,0,145,0,249,0,254,0,120,0,188,0,86,0,95,0,148,0,16,0,161,0,33,0,46,0,217,0,0,0,246,0,38,0,14,0,98,0,253,0,236,0,191,0,0,0,8,0,178,0,27,0,49,0,94,0,98,0,13,0,218,0,14,0,24,0,162,0,211,0,137,0,0,0,213,0,62,0,11,0,251,0,44,0,10,0,6,0,229,0,172,0,189,0,105,0,249,0,115,0,0,0,213,0,235,0,159,0,65,0,0,0,45,0,0,0,11,0,235,0,115,0,32,0,101,0,0,0,130,0,182,0,192,0,48,0,137,0,188,0,145,0,191,0,116,0,223,0,64,0,149,0,0,0,176,0,212,0,172,0,218,0,170,0,91,0,202,0,0,0,229,0,153,0,139,0,163,0,101,0,0,0,0,0,196,0,0,0,164,0,198,0,162,0,75,0,174,0,176,0,0,0,99,0,32,0,0,0,237,0,206,0,227,0,111,0,26,0,73,0,0,0,224,0,56,0,151,0,123,0,31,0,138,0,115,0,118,0,133,0,201,0,61,0,0,0,0,0,0,0,32,0,27,0,0,0,240,0,19,0,249,0,110,0,124,0,46,0,81,0,79,0,119,0,59,0,65,0,149,0,113,0,0,0,148,0,41,0,0,0,0,0,203,0,34,0,42,0,0,0,116,0,144,0,0,0,0,0,252,0,0,0,0,0,126,0,192,0,1,0,85,0,76,0,175,0,125,0,0,0,252,0,231,0,18,0,164,0,86,0,158,0,0,0,247,0,0,0,216,0,128,0,79,0,0,0,201,0,186,0,87,0,117,0,172,0,180,0,218,0,49,0,183,0,186,0,114,0,121,0,34,0,104,0,35,0,110,0,36,0,231,0,137,0,186,0,41,0,21,0,228,0,113,0,187,0,189,0,0,0,0,0,116,0,140,0,206,0,62,0,0,0,67,0,193,0,0,0,133,0,0,0,116,0,105,0,254,0,17,0,252,0,62,0,31,0,124,0,42,0,141,0,3,0,0,0,0,0,187,0,99,0,201,0,245,0,133,0,66,0,116,0,75,0,244,0,79,0,24,0,32,0,0,0,0,0,198,0,0,0,116,0,180,0,27,0,0,0,0,0,59,0,0,0,208,0,219,0,139,0,24,0,104,0,114,0,226,0,0,0,0,0,218,0,230,0,191,0,0,0,196,0,65,0,0,0,164,0,38,0,232,0,51,0,158,0,249,0,96,0,12,0,236,0,0,0,0,0,133,0,69,0,0,0,0,0,108,0,3,0,13,0,72,0,118,0,145,0,169,0,0,0,188,0,109,0,0,0,0,0,0,0,37,0,0,0,69,0,0,0,149,0,8,0,0,0,212,0,0,0,55,0,37,0,111,0,143,0,120,0,0,0,43,0,38,0,0,0,162,0,0,0,168,0,56,0,251,0,0,0,208,0,0,0,32,0,0,0,204,0,106,0,109,0,60,0,62,0,0,0,0,0,180,0,71,0,186,0,28,0,158,0,226,0,0,0,17,0,59,0,32,0,132,0,138,0,175,0,2,0,0,0,0,0,25,0,0,0,10,0,28,0,19,0,152,0,151,0,144,0,0,0,66,0,38,0,70,0,0,0,91,0,82,0,10,0,10,0,109,0,0,0,69,0,15,0,155,0,70,0,71,0,0,0,241,0,34,0,0,0,193,0,124,0,243,0);
signal scenario_full  : scenario_type := (200,31,32,31,197,31,106,31,172,31,245,31,7,31,13,31,217,31,156,31,68,31,175,31,57,31,89,31,188,31,176,31,121,31,121,30,22,31,22,30,224,31,157,31,176,31,62,31,104,31,98,31,249,31,249,31,249,30,148,31,97,31,255,31,87,31,117,31,2,31,31,31,91,31,186,31,50,31,42,31,118,31,118,30,118,29,76,31,246,31,251,31,23,31,105,31,135,31,135,30,135,29,136,31,30,31,8,31,8,30,147,31,222,31,100,31,177,31,255,31,255,30,127,31,88,31,235,31,230,31,230,30,136,31,178,31,218,31,91,31,91,30,91,29,91,28,122,31,214,31,95,31,95,30,42,31,253,31,225,31,186,31,186,30,186,29,87,31,9,31,61,31,145,31,43,31,89,31,71,31,71,30,71,29,94,31,211,31,56,31,56,30,170,31,252,31,42,31,56,31,100,31,217,31,143,31,243,31,243,30,171,31,171,30,87,31,151,31,252,31,247,31,178,31,178,30,255,31,162,31,222,31,148,31,89,31,184,31,184,30,18,31,92,31,108,31,68,31,59,31,101,31,13,31,78,31,138,31,227,31,227,30,227,29,197,31,129,31,125,31,125,30,244,31,248,31,248,30,115,31,18,31,84,31,84,30,100,31,141,31,66,31,233,31,88,31,122,31,122,30,193,31,55,31,206,31,206,30,241,31,46,31,46,30,46,29,209,31,150,31,26,31,86,31,86,30,18,31,77,31,134,31,134,30,153,31,39,31,110,31,110,30,160,31,160,30,43,31,43,30,46,31,213,31,150,31,56,31,55,31,167,31,236,31,239,31,59,31,244,31,233,31,233,30,233,29,133,31,74,31,203,31,113,31,142,31,142,30,52,31,135,31,135,30,195,31,237,31,237,30,94,31,19,31,19,30,175,31,175,30,28,31,28,30,138,31,62,31,73,31,196,31,196,30,219,31,169,31,86,31,86,30,50,31,208,31,85,31,85,30,85,29,217,31,196,31,173,31,168,31,168,30,168,29,13,31,13,30,13,29,62,31,203,31,179,31,206,31,184,31,184,30,5,31,77,31,6,31,153,31,7,31,32,31,206,31,106,31,5,31,5,30,5,29,78,31,92,31,210,31,83,31,32,31,32,30,186,31,90,31,168,31,235,31,111,31,162,31,33,31,119,31,116,31,89,31,204,31,204,30,217,31,44,31,70,31,244,31,192,31,176,31,176,30,153,31,153,30,166,31,166,30,182,31,63,31,235,31,50,31,250,31,250,30,234,31,98,31,143,31,122,31,97,31,197,31,197,30,197,29,84,31,84,30,82,31,77,31,255,31,255,30,138,31,12,31,143,31,63,31,52,31,237,31,121,31,121,30,121,29,132,31,28,31,54,31,136,31,127,31,222,31,241,31,241,30,135,31,135,30,135,29,170,31,242,31,248,31,180,31,201,31,239,31,128,31,128,30,203,31,179,31,15,31,15,31,197,31,197,30,128,31,97,31,107,31,108,31,39,31,39,30,195,31,204,31,162,31,162,30,189,31,98,31,90,31,198,31,198,30,198,29,235,31,212,31,212,30,95,31,56,31,19,31,178,31,120,31,82,31,110,31,149,31,101,31,235,31,179,31,73,31,182,31,182,30,182,29,182,28,153,31,38,31,125,31,209,31,147,31,152,31,235,31,235,30,61,31,158,31,134,31,184,31,191,31,159,31,166,31,36,31,149,31,126,31,160,31,213,31,70,31,26,31,250,31,121,31,121,30,121,29,178,31,43,31,18,31,69,31,99,31,175,31,120,31,244,31,170,31,111,31,1,31,130,31,160,31,197,31,138,31,138,30,18,31,170,31,67,31,239,31,198,31,40,31,101,31,101,30,180,31,157,31,178,31,103,31,64,31,36,31,100,31,109,31,250,31,180,31,124,31,168,31,75,31,206,31,179,31,149,31,200,31,38,31,141,31,126,31,9,31,225,31,225,30,225,29,92,31,130,31,32,31,32,30,147,31,147,30,101,31,101,30,226,31,138,31,194,31,226,31,176,31,17,31,222,31,98,31,249,31,38,31,120,31,155,31,80,31,80,30,22,31,156,31,102,31,212,31,116,31,229,31,40,31,76,31,179,31,109,31,109,30,109,29,101,31,91,31,161,31,44,31,202,31,212,31,78,31,220,31,220,30,237,31,240,31,99,31,99,30,128,31,91,31,135,31,58,31,5,31,5,30,5,29,105,31,229,31,236,31,255,31,255,30,105,31,137,31,137,30,24,31,24,31,24,30,24,29,24,28,214,31,62,31,248,31,218,31,206,31,37,31,37,30,149,31,149,30,149,29,205,31,45,31,56,31,176,31,151,31,7,31,7,30,77,31,77,30,145,31,249,31,254,31,120,31,188,31,86,31,95,31,148,31,16,31,161,31,33,31,46,31,217,31,217,30,246,31,38,31,14,31,98,31,253,31,236,31,191,31,191,30,8,31,178,31,27,31,49,31,94,31,98,31,13,31,218,31,14,31,24,31,162,31,211,31,137,31,137,30,213,31,62,31,11,31,251,31,44,31,10,31,6,31,229,31,172,31,189,31,105,31,249,31,115,31,115,30,213,31,235,31,159,31,65,31,65,30,45,31,45,30,11,31,235,31,115,31,32,31,101,31,101,30,130,31,182,31,192,31,48,31,137,31,188,31,145,31,191,31,116,31,223,31,64,31,149,31,149,30,176,31,212,31,172,31,218,31,170,31,91,31,202,31,202,30,229,31,153,31,139,31,163,31,101,31,101,30,101,29,196,31,196,30,164,31,198,31,162,31,75,31,174,31,176,31,176,30,99,31,32,31,32,30,237,31,206,31,227,31,111,31,26,31,73,31,73,30,224,31,56,31,151,31,123,31,31,31,138,31,115,31,118,31,133,31,201,31,61,31,61,30,61,29,61,28,32,31,27,31,27,30,240,31,19,31,249,31,110,31,124,31,46,31,81,31,79,31,119,31,59,31,65,31,149,31,113,31,113,30,148,31,41,31,41,30,41,29,203,31,34,31,42,31,42,30,116,31,144,31,144,30,144,29,252,31,252,30,252,29,126,31,192,31,1,31,85,31,76,31,175,31,125,31,125,30,252,31,231,31,18,31,164,31,86,31,158,31,158,30,247,31,247,30,216,31,128,31,79,31,79,30,201,31,186,31,87,31,117,31,172,31,180,31,218,31,49,31,183,31,186,31,114,31,121,31,34,31,104,31,35,31,110,31,36,31,231,31,137,31,186,31,41,31,21,31,228,31,113,31,187,31,189,31,189,30,189,29,116,31,140,31,206,31,62,31,62,30,67,31,193,31,193,30,133,31,133,30,116,31,105,31,254,31,17,31,252,31,62,31,31,31,124,31,42,31,141,31,3,31,3,30,3,29,187,31,99,31,201,31,245,31,133,31,66,31,116,31,75,31,244,31,79,31,24,31,32,31,32,30,32,29,198,31,198,30,116,31,180,31,27,31,27,30,27,29,59,31,59,30,208,31,219,31,139,31,24,31,104,31,114,31,226,31,226,30,226,29,218,31,230,31,191,31,191,30,196,31,65,31,65,30,164,31,38,31,232,31,51,31,158,31,249,31,96,31,12,31,236,31,236,30,236,29,133,31,69,31,69,30,69,29,108,31,3,31,13,31,72,31,118,31,145,31,169,31,169,30,188,31,109,31,109,30,109,29,109,28,37,31,37,30,69,31,69,30,149,31,8,31,8,30,212,31,212,30,55,31,37,31,111,31,143,31,120,31,120,30,43,31,38,31,38,30,162,31,162,30,168,31,56,31,251,31,251,30,208,31,208,30,32,31,32,30,204,31,106,31,109,31,60,31,62,31,62,30,62,29,180,31,71,31,186,31,28,31,158,31,226,31,226,30,17,31,59,31,32,31,132,31,138,31,175,31,2,31,2,30,2,29,25,31,25,30,10,31,28,31,19,31,152,31,151,31,144,31,144,30,66,31,38,31,70,31,70,30,91,31,82,31,10,31,10,31,109,31,109,30,69,31,15,31,155,31,70,31,71,31,71,30,241,31,34,31,34,30,193,31,124,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
