-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 268;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (167,0,7,0,156,0,129,0,0,0,100,0,0,0,145,0,60,0,233,0,0,0,91,0,74,0,242,0,218,0,147,0,0,0,206,0,208,0,67,0,212,0,9,0,134,0,165,0,151,0,87,0,153,0,0,0,41,0,184,0,236,0,36,0,200,0,0,0,114,0,236,0,26,0,23,0,142,0,209,0,188,0,133,0,0,0,164,0,0,0,159,0,185,0,98,0,0,0,249,0,54,0,142,0,39,0,186,0,0,0,63,0,69,0,0,0,85,0,110,0,101,0,177,0,0,0,197,0,168,0,0,0,74,0,250,0,113,0,0,0,13,0,197,0,185,0,79,0,0,0,172,0,167,0,143,0,32,0,0,0,173,0,40,0,89,0,210,0,7,0,19,0,142,0,104,0,0,0,0,0,193,0,176,0,215,0,0,0,133,0,178,0,5,0,41,0,191,0,234,0,33,0,189,0,189,0,152,0,248,0,17,0,251,0,0,0,136,0,58,0,0,0,220,0,54,0,226,0,96,0,100,0,78,0,247,0,192,0,0,0,253,0,108,0,137,0,21,0,204,0,180,0,0,0,215,0,206,0,0,0,207,0,27,0,192,0,144,0,149,0,159,0,244,0,60,0,128,0,99,0,133,0,123,0,94,0,160,0,141,0,51,0,34,0,46,0,30,0,0,0,54,0,247,0,84,0,209,0,179,0,140,0,157,0,0,0,202,0,49,0,196,0,81,0,155,0,238,0,237,0,131,0,62,0,157,0,0,0,90,0,84,0,0,0,114,0,115,0,0,0,110,0,13,0,55,0,227,0,0,0,16,0,195,0,0,0,78,0,108,0,108,0,63,0,121,0,0,0,35,0,121,0,44,0,0,0,77,0,113,0,93,0,0,0,149,0,97,0,0,0,246,0,124,0,0,0,46,0,36,0,130,0,234,0,161,0,119,0,170,0,181,0,0,0,114,0,218,0,0,0,59,0,108,0,209,0,162,0,11,0,96,0,65,0,75,0,128,0,42,0,0,0,0,0,23,0,138,0,0,0,0,0,189,0,95,0,252,0,249,0,228,0,255,0,194,0,0,0,0,0,176,0,111,0,42,0,251,0,149,0,0,0,2,0,204,0,151,0,208,0,250,0,41,0,0,0,6,0,132,0,219,0,89,0,150,0,229,0,150,0,182,0,57,0,60,0,80,0,0,0,0,0,193,0,129,0);
signal scenario_full  : scenario_type := (167,31,7,31,156,31,129,31,129,30,100,31,100,30,145,31,60,31,233,31,233,30,91,31,74,31,242,31,218,31,147,31,147,30,206,31,208,31,67,31,212,31,9,31,134,31,165,31,151,31,87,31,153,31,153,30,41,31,184,31,236,31,36,31,200,31,200,30,114,31,236,31,26,31,23,31,142,31,209,31,188,31,133,31,133,30,164,31,164,30,159,31,185,31,98,31,98,30,249,31,54,31,142,31,39,31,186,31,186,30,63,31,69,31,69,30,85,31,110,31,101,31,177,31,177,30,197,31,168,31,168,30,74,31,250,31,113,31,113,30,13,31,197,31,185,31,79,31,79,30,172,31,167,31,143,31,32,31,32,30,173,31,40,31,89,31,210,31,7,31,19,31,142,31,104,31,104,30,104,29,193,31,176,31,215,31,215,30,133,31,178,31,5,31,41,31,191,31,234,31,33,31,189,31,189,31,152,31,248,31,17,31,251,31,251,30,136,31,58,31,58,30,220,31,54,31,226,31,96,31,100,31,78,31,247,31,192,31,192,30,253,31,108,31,137,31,21,31,204,31,180,31,180,30,215,31,206,31,206,30,207,31,27,31,192,31,144,31,149,31,159,31,244,31,60,31,128,31,99,31,133,31,123,31,94,31,160,31,141,31,51,31,34,31,46,31,30,31,30,30,54,31,247,31,84,31,209,31,179,31,140,31,157,31,157,30,202,31,49,31,196,31,81,31,155,31,238,31,237,31,131,31,62,31,157,31,157,30,90,31,84,31,84,30,114,31,115,31,115,30,110,31,13,31,55,31,227,31,227,30,16,31,195,31,195,30,78,31,108,31,108,31,63,31,121,31,121,30,35,31,121,31,44,31,44,30,77,31,113,31,93,31,93,30,149,31,97,31,97,30,246,31,124,31,124,30,46,31,36,31,130,31,234,31,161,31,119,31,170,31,181,31,181,30,114,31,218,31,218,30,59,31,108,31,209,31,162,31,11,31,96,31,65,31,75,31,128,31,42,31,42,30,42,29,23,31,138,31,138,30,138,29,189,31,95,31,252,31,249,31,228,31,255,31,194,31,194,30,194,29,176,31,111,31,42,31,251,31,149,31,149,30,2,31,204,31,151,31,208,31,250,31,41,31,41,30,6,31,132,31,219,31,89,31,150,31,229,31,150,31,182,31,57,31,60,31,80,31,80,30,80,29,193,31,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
