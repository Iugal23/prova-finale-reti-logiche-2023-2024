-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 867;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,0,0,0,0,0,0,35,0,218,0,195,0,109,0,93,0,44,0,25,0,107,0,72,0,149,0,233,0,112,0,171,0,40,0,103,0,6,0,0,0,136,0,55,0,78,0,93,0,207,0,207,0,0,0,236,0,10,0,32,0,125,0,113,0,252,0,17,0,192,0,32,0,159,0,77,0,134,0,80,0,20,0,24,0,149,0,172,0,34,0,223,0,209,0,177,0,91,0,116,0,146,0,6,0,181,0,32,0,204,0,225,0,36,0,0,0,148,0,106,0,30,0,229,0,84,0,178,0,200,0,177,0,155,0,0,0,87,0,230,0,96,0,0,0,60,0,25,0,48,0,192,0,144,0,148,0,0,0,0,0,31,0,76,0,144,0,86,0,0,0,145,0,0,0,195,0,73,0,148,0,167,0,112,0,189,0,160,0,130,0,48,0,144,0,0,0,121,0,155,0,0,0,199,0,0,0,150,0,55,0,183,0,0,0,0,0,38,0,0,0,205,0,150,0,128,0,98,0,4,0,33,0,247,0,138,0,193,0,23,0,132,0,0,0,75,0,0,0,237,0,190,0,254,0,236,0,0,0,115,0,13,0,0,0,85,0,0,0,125,0,0,0,91,0,228,0,71,0,162,0,0,0,229,0,10,0,219,0,15,0,170,0,242,0,225,0,0,0,82,0,140,0,0,0,219,0,177,0,249,0,168,0,147,0,84,0,35,0,233,0,142,0,79,0,0,0,132,0,0,0,28,0,0,0,101,0,153,0,194,0,113,0,125,0,194,0,170,0,202,0,203,0,123,0,0,0,225,0,0,0,141,0,0,0,128,0,187,0,0,0,0,0,162,0,196,0,26,0,0,0,209,0,204,0,185,0,32,0,0,0,61,0,156,0,0,0,161,0,213,0,169,0,159,0,134,0,0,0,150,0,0,0,241,0,100,0,236,0,139,0,19,0,0,0,65,0,17,0,165,0,73,0,181,0,0,0,77,0,0,0,0,0,48,0,0,0,218,0,66,0,100,0,177,0,190,0,151,0,142,0,220,0,21,0,79,0,5,0,130,0,91,0,79,0,35,0,94,0,235,0,243,0,0,0,0,0,56,0,252,0,101,0,78,0,0,0,0,0,0,0,76,0,0,0,14,0,7,0,60,0,0,0,63,0,172,0,60,0,149,0,165,0,193,0,0,0,0,0,60,0,0,0,115,0,84,0,171,0,136,0,46,0,0,0,70,0,198,0,163,0,47,0,68,0,86,0,100,0,143,0,0,0,0,0,49,0,95,0,0,0,147,0,19,0,130,0,172,0,19,0,133,0,74,0,64,0,220,0,37,0,94,0,0,0,118,0,227,0,143,0,110,0,0,0,145,0,17,0,44,0,167,0,182,0,95,0,0,0,155,0,48,0,0,0,216,0,191,0,0,0,239,0,105,0,0,0,0,0,40,0,154,0,117,0,52,0,92,0,238,0,165,0,64,0,151,0,124,0,215,0,31,0,0,0,31,0,101,0,204,0,237,0,228,0,41,0,93,0,20,0,33,0,82,0,95,0,124,0,82,0,200,0,200,0,0,0,58,0,220,0,138,0,166,0,0,0,92,0,179,0,146,0,152,0,240,0,228,0,43,0,0,0,223,0,233,0,247,0,0,0,0,0,127,0,67,0,0,0,5,0,139,0,83,0,116,0,28,0,0,0,91,0,123,0,205,0,132,0,213,0,114,0,166,0,108,0,183,0,69,0,218,0,137,0,222,0,11,0,29,0,187,0,229,0,52,0,0,0,208,0,198,0,102,0,44,0,152,0,238,0,188,0,177,0,47,0,11,0,64,0,169,0,64,0,0,0,210,0,76,0,80,0,6,0,98,0,110,0,134,0,127,0,6,0,118,0,87,0,0,0,83,0,103,0,0,0,34,0,40,0,220,0,199,0,121,0,152,0,90,0,0,0,118,0,45,0,126,0,158,0,0,0,159,0,189,0,0,0,0,0,184,0,0,0,35,0,0,0,60,0,41,0,112,0,214,0,104,0,213,0,0,0,0,0,148,0,124,0,115,0,188,0,237,0,53,0,207,0,165,0,0,0,189,0,0,0,0,0,0,0,38,0,41,0,134,0,0,0,0,0,209,0,108,0,146,0,115,0,228,0,0,0,0,0,198,0,15,0,52,0,0,0,106,0,116,0,109,0,195,0,37,0,0,0,96,0,84,0,71,0,0,0,0,0,85,0,72,0,0,0,232,0,100,0,168,0,251,0,184,0,158,0,0,0,119,0,0,0,75,0,204,0,65,0,157,0,184,0,81,0,64,0,0,0,185,0,67,0,178,0,88,0,140,0,186,0,207,0,64,0,188,0,197,0,76,0,27,0,158,0,171,0,15,0,207,0,170,0,214,0,81,0,225,0,25,0,0,0,5,0,75,0,161,0,134,0,0,0,26,0,150,0,0,0,10,0,118,0,204,0,118,0,35,0,89,0,229,0,128,0,13,0,22,0,171,0,92,0,63,0,144,0,6,0,216,0,71,0,0,0,23,0,0,0,197,0,208,0,27,0,145,0,203,0,171,0,93,0,147,0,122,0,0,0,40,0,0,0,155,0,42,0,103,0,94,0,0,0,122,0,39,0,0,0,183,0,219,0,0,0,32,0,74,0,145,0,101,0,132,0,0,0,138,0,0,0,0,0,218,0,200,0,181,0,33,0,38,0,146,0,0,0,154,0,78,0,62,0,253,0,223,0,132,0,13,0,165,0,217,0,0,0,0,0,0,0,126,0,32,0,60,0,205,0,0,0,145,0,0,0,66,0,0,0,53,0,0,0,62,0,198,0,0,0,118,0,195,0,232,0,248,0,182,0,56,0,60,0,119,0,0,0,0,0,140,0,7,0,0,0,13,0,8,0,57,0,167,0,234,0,105,0,52,0,165,0,214,0,136,0,22,0,198,0,220,0,86,0,0,0,36,0,100,0,84,0,228,0,194,0,19,0,247,0,61,0,84,0,186,0,226,0,200,0,0,0,1,0,0,0,0,0,53,0,145,0,53,0,0,0,211,0,252,0,175,0,235,0,236,0,254,0,178,0,150,0,41,0,0,0,112,0,119,0,102,0,227,0,163,0,111,0,226,0,0,0,0,0,255,0,202,0,105,0,186,0,237,0,36,0,127,0,0,0,0,0,222,0,47,0,0,0,167,0,115,0,97,0,146,0,155,0,39,0,248,0,162,0,224,0,92,0,0,0,37,0,0,0,202,0,231,0,55,0,0,0,196,0,246,0,86,0,165,0,199,0,103,0,0,0,0,0,211,0,116,0,254,0,0,0,145,0,0,0,235,0,245,0,0,0,255,0,0,0,11,0,54,0,254,0,192,0,0,0,252,0,62,0,103,0,139,0,0,0,122,0,91,0,113,0,229,0,155,0,42,0,0,0,133,0,255,0,124,0,0,0,56,0,208,0,117,0,181,0,9,0,42,0,252,0,32,0,0,0,177,0,170,0,0,0,61,0,40,0,97,0,0,0,0,0,38,0,31,0,96,0,162,0,28,0,247,0,118,0,162,0,201,0,206,0,54,0,125,0,147,0,252,0,138,0,182,0,0,0,114,0,0,0,121,0,161,0,55,0,37,0,231,0,84,0,69,0,0,0,169,0,70,0,34,0,19,0,183,0,74,0,66,0,0,0,239,0,159,0,191,0,0,0,49,0,233,0,254,0,0,0,225,0,0,0,0,0,196,0,135,0,231,0,74,0,226,0,0,0,177,0,0,0,230,0,0,0,32,0,165,0,145,0,49,0,0,0,243,0,198,0,59,0,162,0,0,0,83,0,147,0,37,0,59,0,242,0,0,0,0,0,0,0,93,0,156,0,80,0,119,0,254,0,82,0,203,0,116,0,108,0,0,0,161,0,41,0);
signal scenario_full  : scenario_type := (24,31,24,30,24,29,24,28,35,31,218,31,195,31,109,31,93,31,44,31,25,31,107,31,72,31,149,31,233,31,112,31,171,31,40,31,103,31,6,31,6,30,136,31,55,31,78,31,93,31,207,31,207,31,207,30,236,31,10,31,32,31,125,31,113,31,252,31,17,31,192,31,32,31,159,31,77,31,134,31,80,31,20,31,24,31,149,31,172,31,34,31,223,31,209,31,177,31,91,31,116,31,146,31,6,31,181,31,32,31,204,31,225,31,36,31,36,30,148,31,106,31,30,31,229,31,84,31,178,31,200,31,177,31,155,31,155,30,87,31,230,31,96,31,96,30,60,31,25,31,48,31,192,31,144,31,148,31,148,30,148,29,31,31,76,31,144,31,86,31,86,30,145,31,145,30,195,31,73,31,148,31,167,31,112,31,189,31,160,31,130,31,48,31,144,31,144,30,121,31,155,31,155,30,199,31,199,30,150,31,55,31,183,31,183,30,183,29,38,31,38,30,205,31,150,31,128,31,98,31,4,31,33,31,247,31,138,31,193,31,23,31,132,31,132,30,75,31,75,30,237,31,190,31,254,31,236,31,236,30,115,31,13,31,13,30,85,31,85,30,125,31,125,30,91,31,228,31,71,31,162,31,162,30,229,31,10,31,219,31,15,31,170,31,242,31,225,31,225,30,82,31,140,31,140,30,219,31,177,31,249,31,168,31,147,31,84,31,35,31,233,31,142,31,79,31,79,30,132,31,132,30,28,31,28,30,101,31,153,31,194,31,113,31,125,31,194,31,170,31,202,31,203,31,123,31,123,30,225,31,225,30,141,31,141,30,128,31,187,31,187,30,187,29,162,31,196,31,26,31,26,30,209,31,204,31,185,31,32,31,32,30,61,31,156,31,156,30,161,31,213,31,169,31,159,31,134,31,134,30,150,31,150,30,241,31,100,31,236,31,139,31,19,31,19,30,65,31,17,31,165,31,73,31,181,31,181,30,77,31,77,30,77,29,48,31,48,30,218,31,66,31,100,31,177,31,190,31,151,31,142,31,220,31,21,31,79,31,5,31,130,31,91,31,79,31,35,31,94,31,235,31,243,31,243,30,243,29,56,31,252,31,101,31,78,31,78,30,78,29,78,28,76,31,76,30,14,31,7,31,60,31,60,30,63,31,172,31,60,31,149,31,165,31,193,31,193,30,193,29,60,31,60,30,115,31,84,31,171,31,136,31,46,31,46,30,70,31,198,31,163,31,47,31,68,31,86,31,100,31,143,31,143,30,143,29,49,31,95,31,95,30,147,31,19,31,130,31,172,31,19,31,133,31,74,31,64,31,220,31,37,31,94,31,94,30,118,31,227,31,143,31,110,31,110,30,145,31,17,31,44,31,167,31,182,31,95,31,95,30,155,31,48,31,48,30,216,31,191,31,191,30,239,31,105,31,105,30,105,29,40,31,154,31,117,31,52,31,92,31,238,31,165,31,64,31,151,31,124,31,215,31,31,31,31,30,31,31,101,31,204,31,237,31,228,31,41,31,93,31,20,31,33,31,82,31,95,31,124,31,82,31,200,31,200,31,200,30,58,31,220,31,138,31,166,31,166,30,92,31,179,31,146,31,152,31,240,31,228,31,43,31,43,30,223,31,233,31,247,31,247,30,247,29,127,31,67,31,67,30,5,31,139,31,83,31,116,31,28,31,28,30,91,31,123,31,205,31,132,31,213,31,114,31,166,31,108,31,183,31,69,31,218,31,137,31,222,31,11,31,29,31,187,31,229,31,52,31,52,30,208,31,198,31,102,31,44,31,152,31,238,31,188,31,177,31,47,31,11,31,64,31,169,31,64,31,64,30,210,31,76,31,80,31,6,31,98,31,110,31,134,31,127,31,6,31,118,31,87,31,87,30,83,31,103,31,103,30,34,31,40,31,220,31,199,31,121,31,152,31,90,31,90,30,118,31,45,31,126,31,158,31,158,30,159,31,189,31,189,30,189,29,184,31,184,30,35,31,35,30,60,31,41,31,112,31,214,31,104,31,213,31,213,30,213,29,148,31,124,31,115,31,188,31,237,31,53,31,207,31,165,31,165,30,189,31,189,30,189,29,189,28,38,31,41,31,134,31,134,30,134,29,209,31,108,31,146,31,115,31,228,31,228,30,228,29,198,31,15,31,52,31,52,30,106,31,116,31,109,31,195,31,37,31,37,30,96,31,84,31,71,31,71,30,71,29,85,31,72,31,72,30,232,31,100,31,168,31,251,31,184,31,158,31,158,30,119,31,119,30,75,31,204,31,65,31,157,31,184,31,81,31,64,31,64,30,185,31,67,31,178,31,88,31,140,31,186,31,207,31,64,31,188,31,197,31,76,31,27,31,158,31,171,31,15,31,207,31,170,31,214,31,81,31,225,31,25,31,25,30,5,31,75,31,161,31,134,31,134,30,26,31,150,31,150,30,10,31,118,31,204,31,118,31,35,31,89,31,229,31,128,31,13,31,22,31,171,31,92,31,63,31,144,31,6,31,216,31,71,31,71,30,23,31,23,30,197,31,208,31,27,31,145,31,203,31,171,31,93,31,147,31,122,31,122,30,40,31,40,30,155,31,42,31,103,31,94,31,94,30,122,31,39,31,39,30,183,31,219,31,219,30,32,31,74,31,145,31,101,31,132,31,132,30,138,31,138,30,138,29,218,31,200,31,181,31,33,31,38,31,146,31,146,30,154,31,78,31,62,31,253,31,223,31,132,31,13,31,165,31,217,31,217,30,217,29,217,28,126,31,32,31,60,31,205,31,205,30,145,31,145,30,66,31,66,30,53,31,53,30,62,31,198,31,198,30,118,31,195,31,232,31,248,31,182,31,56,31,60,31,119,31,119,30,119,29,140,31,7,31,7,30,13,31,8,31,57,31,167,31,234,31,105,31,52,31,165,31,214,31,136,31,22,31,198,31,220,31,86,31,86,30,36,31,100,31,84,31,228,31,194,31,19,31,247,31,61,31,84,31,186,31,226,31,200,31,200,30,1,31,1,30,1,29,53,31,145,31,53,31,53,30,211,31,252,31,175,31,235,31,236,31,254,31,178,31,150,31,41,31,41,30,112,31,119,31,102,31,227,31,163,31,111,31,226,31,226,30,226,29,255,31,202,31,105,31,186,31,237,31,36,31,127,31,127,30,127,29,222,31,47,31,47,30,167,31,115,31,97,31,146,31,155,31,39,31,248,31,162,31,224,31,92,31,92,30,37,31,37,30,202,31,231,31,55,31,55,30,196,31,246,31,86,31,165,31,199,31,103,31,103,30,103,29,211,31,116,31,254,31,254,30,145,31,145,30,235,31,245,31,245,30,255,31,255,30,11,31,54,31,254,31,192,31,192,30,252,31,62,31,103,31,139,31,139,30,122,31,91,31,113,31,229,31,155,31,42,31,42,30,133,31,255,31,124,31,124,30,56,31,208,31,117,31,181,31,9,31,42,31,252,31,32,31,32,30,177,31,170,31,170,30,61,31,40,31,97,31,97,30,97,29,38,31,31,31,96,31,162,31,28,31,247,31,118,31,162,31,201,31,206,31,54,31,125,31,147,31,252,31,138,31,182,31,182,30,114,31,114,30,121,31,161,31,55,31,37,31,231,31,84,31,69,31,69,30,169,31,70,31,34,31,19,31,183,31,74,31,66,31,66,30,239,31,159,31,191,31,191,30,49,31,233,31,254,31,254,30,225,31,225,30,225,29,196,31,135,31,231,31,74,31,226,31,226,30,177,31,177,30,230,31,230,30,32,31,165,31,145,31,49,31,49,30,243,31,198,31,59,31,162,31,162,30,83,31,147,31,37,31,59,31,242,31,242,30,242,29,242,28,93,31,156,31,80,31,119,31,254,31,82,31,203,31,116,31,108,31,108,30,161,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
