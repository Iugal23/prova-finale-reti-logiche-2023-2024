-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 418;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (137,0,128,0,154,0,196,0,0,0,4,0,138,0,140,0,148,0,0,0,106,0,0,0,0,0,206,0,108,0,133,0,109,0,147,0,153,0,132,0,119,0,121,0,212,0,1,0,53,0,196,0,151,0,70,0,3,0,233,0,72,0,0,0,229,0,53,0,165,0,142,0,254,0,163,0,187,0,231,0,218,0,171,0,100,0,0,0,229,0,0,0,20,0,115,0,130,0,20,0,0,0,162,0,77,0,132,0,2,0,0,0,0,0,66,0,104,0,91,0,178,0,0,0,25,0,0,0,79,0,41,0,154,0,29,0,250,0,127,0,39,0,229,0,156,0,50,0,76,0,154,0,90,0,26,0,0,0,39,0,0,0,154,0,254,0,0,0,144,0,161,0,179,0,161,0,161,0,159,0,65,0,218,0,120,0,66,0,200,0,0,0,137,0,61,0,235,0,5,0,31,0,243,0,115,0,0,0,48,0,235,0,249,0,221,0,97,0,52,0,201,0,214,0,0,0,225,0,0,0,28,0,50,0,73,0,0,0,209,0,114,0,232,0,157,0,211,0,241,0,106,0,87,0,185,0,179,0,194,0,171,0,0,0,36,0,0,0,207,0,0,0,61,0,0,0,212,0,0,0,40,0,0,0,122,0,247,0,75,0,19,0,115,0,5,0,0,0,23,0,175,0,142,0,165,0,0,0,123,0,254,0,166,0,0,0,0,0,82,0,21,0,59,0,0,0,0,0,0,0,48,0,214,0,203,0,153,0,250,0,185,0,56,0,137,0,217,0,160,0,216,0,24,0,113,0,118,0,0,0,189,0,148,0,0,0,0,0,0,0,0,0,218,0,249,0,0,0,39,0,127,0,84,0,134,0,30,0,126,0,188,0,0,0,205,0,123,0,0,0,18,0,215,0,140,0,119,0,134,0,93,0,89,0,143,0,219,0,0,0,0,0,248,0,73,0,5,0,163,0,14,0,0,0,0,0,166,0,0,0,196,0,140,0,44,0,188,0,0,0,152,0,95,0,0,0,54,0,20,0,0,0,52,0,168,0,190,0,186,0,65,0,150,0,54,0,88,0,156,0,203,0,0,0,214,0,0,0,158,0,80,0,84,0,231,0,135,0,22,0,236,0,200,0,0,0,153,0,153,0,193,0,248,0,0,0,73,0,239,0,229,0,0,0,0,0,144,0,0,0,63,0,254,0,213,0,165,0,126,0,182,0,103,0,0,0,163,0,1,0,5,0,112,0,211,0,0,0,69,0,131,0,0,0,154,0,217,0,186,0,0,0,233,0,236,0,0,0,219,0,0,0,50,0,115,0,41,0,133,0,255,0,161,0,77,0,79,0,216,0,0,0,129,0,208,0,98,0,0,0,231,0,0,0,154,0,133,0,8,0,183,0,215,0,158,0,181,0,182,0,8,0,0,0,100,0,174,0,0,0,183,0,37,0,201,0,149,0,94,0,0,0,0,0,180,0,204,0,0,0,27,0,248,0,33,0,215,0,107,0,233,0,253,0,183,0,0,0,0,0,8,0,239,0,0,0,157,0,108,0,147,0,73,0,244,0,196,0,151,0,104,0,0,0,175,0,0,0,101,0,117,0,0,0,0,0,177,0,0,0,110,0,190,0,1,0,187,0,23,0,6,0,157,0,0,0,212,0,230,0,54,0,248,0,31,0,0,0,225,0,46,0,97,0,3,0,109,0,188,0,30,0,193,0,132,0,225,0,203,0,26,0,107,0,116,0,123,0,0,0,88,0,0,0,0,0,226,0,180,0,0,0,216,0,184,0,174,0,186,0,170,0,247,0,84,0,40,0,167,0,171,0,120,0,0,0,0,0,207,0,47,0,208,0,240,0,0,0,170,0,0,0,0,0,153,0);
signal scenario_full  : scenario_type := (137,31,128,31,154,31,196,31,196,30,4,31,138,31,140,31,148,31,148,30,106,31,106,30,106,29,206,31,108,31,133,31,109,31,147,31,153,31,132,31,119,31,121,31,212,31,1,31,53,31,196,31,151,31,70,31,3,31,233,31,72,31,72,30,229,31,53,31,165,31,142,31,254,31,163,31,187,31,231,31,218,31,171,31,100,31,100,30,229,31,229,30,20,31,115,31,130,31,20,31,20,30,162,31,77,31,132,31,2,31,2,30,2,29,66,31,104,31,91,31,178,31,178,30,25,31,25,30,79,31,41,31,154,31,29,31,250,31,127,31,39,31,229,31,156,31,50,31,76,31,154,31,90,31,26,31,26,30,39,31,39,30,154,31,254,31,254,30,144,31,161,31,179,31,161,31,161,31,159,31,65,31,218,31,120,31,66,31,200,31,200,30,137,31,61,31,235,31,5,31,31,31,243,31,115,31,115,30,48,31,235,31,249,31,221,31,97,31,52,31,201,31,214,31,214,30,225,31,225,30,28,31,50,31,73,31,73,30,209,31,114,31,232,31,157,31,211,31,241,31,106,31,87,31,185,31,179,31,194,31,171,31,171,30,36,31,36,30,207,31,207,30,61,31,61,30,212,31,212,30,40,31,40,30,122,31,247,31,75,31,19,31,115,31,5,31,5,30,23,31,175,31,142,31,165,31,165,30,123,31,254,31,166,31,166,30,166,29,82,31,21,31,59,31,59,30,59,29,59,28,48,31,214,31,203,31,153,31,250,31,185,31,56,31,137,31,217,31,160,31,216,31,24,31,113,31,118,31,118,30,189,31,148,31,148,30,148,29,148,28,148,27,218,31,249,31,249,30,39,31,127,31,84,31,134,31,30,31,126,31,188,31,188,30,205,31,123,31,123,30,18,31,215,31,140,31,119,31,134,31,93,31,89,31,143,31,219,31,219,30,219,29,248,31,73,31,5,31,163,31,14,31,14,30,14,29,166,31,166,30,196,31,140,31,44,31,188,31,188,30,152,31,95,31,95,30,54,31,20,31,20,30,52,31,168,31,190,31,186,31,65,31,150,31,54,31,88,31,156,31,203,31,203,30,214,31,214,30,158,31,80,31,84,31,231,31,135,31,22,31,236,31,200,31,200,30,153,31,153,31,193,31,248,31,248,30,73,31,239,31,229,31,229,30,229,29,144,31,144,30,63,31,254,31,213,31,165,31,126,31,182,31,103,31,103,30,163,31,1,31,5,31,112,31,211,31,211,30,69,31,131,31,131,30,154,31,217,31,186,31,186,30,233,31,236,31,236,30,219,31,219,30,50,31,115,31,41,31,133,31,255,31,161,31,77,31,79,31,216,31,216,30,129,31,208,31,98,31,98,30,231,31,231,30,154,31,133,31,8,31,183,31,215,31,158,31,181,31,182,31,8,31,8,30,100,31,174,31,174,30,183,31,37,31,201,31,149,31,94,31,94,30,94,29,180,31,204,31,204,30,27,31,248,31,33,31,215,31,107,31,233,31,253,31,183,31,183,30,183,29,8,31,239,31,239,30,157,31,108,31,147,31,73,31,244,31,196,31,151,31,104,31,104,30,175,31,175,30,101,31,117,31,117,30,117,29,177,31,177,30,110,31,190,31,1,31,187,31,23,31,6,31,157,31,157,30,212,31,230,31,54,31,248,31,31,31,31,30,225,31,46,31,97,31,3,31,109,31,188,31,30,31,193,31,132,31,225,31,203,31,26,31,107,31,116,31,123,31,123,30,88,31,88,30,88,29,226,31,180,31,180,30,216,31,184,31,174,31,186,31,170,31,247,31,84,31,40,31,167,31,171,31,120,31,120,30,120,29,207,31,47,31,208,31,240,31,240,30,170,31,170,30,170,29,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
