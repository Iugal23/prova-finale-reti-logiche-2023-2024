-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 255;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (90,0,245,0,0,0,53,0,117,0,173,0,5,0,47,0,251,0,111,0,43,0,109,0,70,0,68,0,25,0,94,0,186,0,187,0,69,0,0,0,202,0,212,0,25,0,228,0,238,0,41,0,142,0,233,0,0,0,157,0,73,0,247,0,0,0,79,0,97,0,33,0,105,0,0,0,83,0,190,0,165,0,0,0,127,0,0,0,0,0,169,0,94,0,0,0,110,0,122,0,0,0,215,0,184,0,161,0,110,0,187,0,16,0,178,0,91,0,0,0,71,0,88,0,46,0,102,0,111,0,212,0,79,0,55,0,182,0,66,0,56,0,156,0,233,0,130,0,11,0,75,0,0,0,206,0,255,0,208,0,0,0,208,0,103,0,0,0,16,0,111,0,165,0,109,0,173,0,173,0,135,0,20,0,217,0,0,0,250,0,0,0,93,0,236,0,214,0,0,0,0,0,149,0,218,0,198,0,0,0,0,0,0,0,218,0,175,0,19,0,91,0,0,0,0,0,8,0,0,0,77,0,57,0,43,0,4,0,134,0,7,0,153,0,140,0,21,0,239,0,86,0,120,0,113,0,0,0,0,0,97,0,46,0,155,0,26,0,43,0,16,0,167,0,106,0,48,0,212,0,0,0,107,0,37,0,176,0,159,0,0,0,53,0,33,0,120,0,239,0,41,0,67,0,220,0,168,0,129,0,76,0,171,0,0,0,70,0,106,0,197,0,103,0,0,0,6,0,79,0,146,0,216,0,197,0,18,0,35,0,91,0,193,0,63,0,239,0,250,0,174,0,238,0,57,0,46,0,7,0,130,0,0,0,0,0,30,0,0,0,219,0,68,0,110,0,57,0,0,0,43,0,49,0,0,0,168,0,0,0,53,0,28,0,0,0,119,0,0,0,56,0,77,0,175,0,70,0,104,0,31,0,28,0,87,0,76,0,127,0,0,0,12,0,98,0,246,0,16,0,164,0,157,0,7,0,255,0,104,0,190,0,7,0,8,0,174,0,23,0,242,0,21,0,34,0,72,0,49,0,230,0,130,0,0,0,0,0,0,0,122,0,0,0,30,0,9,0,239,0,117,0,2,0,235,0,0,0,41,0,0,0,0,0,113,0,251,0,126,0,160,0,53,0,69,0,0,0,236,0);
signal scenario_full  : scenario_type := (90,31,245,31,245,30,53,31,117,31,173,31,5,31,47,31,251,31,111,31,43,31,109,31,70,31,68,31,25,31,94,31,186,31,187,31,69,31,69,30,202,31,212,31,25,31,228,31,238,31,41,31,142,31,233,31,233,30,157,31,73,31,247,31,247,30,79,31,97,31,33,31,105,31,105,30,83,31,190,31,165,31,165,30,127,31,127,30,127,29,169,31,94,31,94,30,110,31,122,31,122,30,215,31,184,31,161,31,110,31,187,31,16,31,178,31,91,31,91,30,71,31,88,31,46,31,102,31,111,31,212,31,79,31,55,31,182,31,66,31,56,31,156,31,233,31,130,31,11,31,75,31,75,30,206,31,255,31,208,31,208,30,208,31,103,31,103,30,16,31,111,31,165,31,109,31,173,31,173,31,135,31,20,31,217,31,217,30,250,31,250,30,93,31,236,31,214,31,214,30,214,29,149,31,218,31,198,31,198,30,198,29,198,28,218,31,175,31,19,31,91,31,91,30,91,29,8,31,8,30,77,31,57,31,43,31,4,31,134,31,7,31,153,31,140,31,21,31,239,31,86,31,120,31,113,31,113,30,113,29,97,31,46,31,155,31,26,31,43,31,16,31,167,31,106,31,48,31,212,31,212,30,107,31,37,31,176,31,159,31,159,30,53,31,33,31,120,31,239,31,41,31,67,31,220,31,168,31,129,31,76,31,171,31,171,30,70,31,106,31,197,31,103,31,103,30,6,31,79,31,146,31,216,31,197,31,18,31,35,31,91,31,193,31,63,31,239,31,250,31,174,31,238,31,57,31,46,31,7,31,130,31,130,30,130,29,30,31,30,30,219,31,68,31,110,31,57,31,57,30,43,31,49,31,49,30,168,31,168,30,53,31,28,31,28,30,119,31,119,30,56,31,77,31,175,31,70,31,104,31,31,31,28,31,87,31,76,31,127,31,127,30,12,31,98,31,246,31,16,31,164,31,157,31,7,31,255,31,104,31,190,31,7,31,8,31,174,31,23,31,242,31,21,31,34,31,72,31,49,31,230,31,130,31,130,30,130,29,130,28,122,31,122,30,30,31,9,31,239,31,117,31,2,31,235,31,235,30,41,31,41,30,41,29,113,31,251,31,126,31,160,31,53,31,69,31,69,30,236,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
