-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 761;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,203,0,147,0,0,0,140,0,75,0,151,0,0,0,14,0,253,0,51,0,147,0,94,0,36,0,123,0,184,0,30,0,201,0,149,0,223,0,0,0,75,0,159,0,248,0,173,0,183,0,182,0,0,0,76,0,29,0,180,0,184,0,0,0,191,0,89,0,78,0,232,0,123,0,133,0,207,0,185,0,83,0,229,0,0,0,196,0,158,0,111,0,164,0,34,0,55,0,0,0,245,0,245,0,0,0,85,0,147,0,69,0,59,0,0,0,23,0,0,0,47,0,92,0,185,0,8,0,236,0,114,0,55,0,125,0,65,0,241,0,243,0,193,0,140,0,0,0,239,0,0,0,143,0,176,0,214,0,132,0,169,0,35,0,37,0,84,0,15,0,162,0,76,0,190,0,152,0,202,0,0,0,0,0,104,0,109,0,169,0,0,0,188,0,179,0,224,0,46,0,93,0,159,0,0,0,0,0,10,0,83,0,63,0,52,0,217,0,131,0,133,0,231,0,74,0,195,0,123,0,64,0,15,0,38,0,219,0,249,0,234,0,153,0,0,0,185,0,69,0,195,0,206,0,178,0,127,0,109,0,115,0,121,0,166,0,169,0,160,0,202,0,163,0,0,0,35,0,183,0,154,0,200,0,200,0,211,0,194,0,97,0,156,0,124,0,140,0,0,0,14,0,84,0,140,0,49,0,0,0,0,0,0,0,0,0,0,0,143,0,214,0,145,0,148,0,118,0,43,0,0,0,138,0,113,0,0,0,188,0,145,0,41,0,18,0,127,0,93,0,90,0,227,0,0,0,209,0,180,0,66,0,88,0,133,0,99,0,192,0,133,0,166,0,205,0,173,0,88,0,59,0,126,0,182,0,238,0,57,0,216,0,160,0,158,0,0,0,48,0,20,0,247,0,12,0,36,0,247,0,125,0,101,0,225,0,132,0,150,0,117,0,86,0,185,0,0,0,33,0,0,0,0,0,29,0,235,0,235,0,150,0,126,0,0,0,202,0,12,0,142,0,150,0,198,0,217,0,103,0,148,0,0,0,212,0,0,0,102,0,100,0,252,0,187,0,219,0,190,0,82,0,0,0,0,0,212,0,0,0,0,0,8,0,141,0,202,0,0,0,238,0,166,0,129,0,53,0,87,0,186,0,0,0,0,0,126,0,243,0,179,0,162,0,0,0,0,0,3,0,188,0,85,0,42,0,0,0,0,0,35,0,59,0,135,0,64,0,0,0,219,0,0,0,0,0,33,0,0,0,0,0,232,0,20,0,191,0,65,0,179,0,87,0,36,0,0,0,0,0,242,0,18,0,5,0,45,0,0,0,118,0,192,0,137,0,93,0,0,0,80,0,8,0,90,0,110,0,23,0,0,0,79,0,238,0,213,0,123,0,107,0,0,0,20,0,0,0,0,0,107,0,11,0,89,0,41,0,53,0,0,0,85,0,236,0,211,0,0,0,226,0,158,0,0,0,0,0,0,0,162,0,178,0,20,0,89,0,55,0,0,0,0,0,86,0,123,0,237,0,56,0,139,0,105,0,23,0,218,0,150,0,45,0,0,0,127,0,0,0,136,0,0,0,61,0,76,0,242,0,68,0,245,0,39,0,122,0,211,0,61,0,215,0,23,0,82,0,168,0,1,0,15,0,99,0,0,0,121,0,151,0,225,0,147,0,245,0,68,0,190,0,181,0,243,0,0,0,192,0,197,0,0,0,188,0,31,0,44,0,3,0,121,0,81,0,113,0,0,0,11,0,138,0,152,0,156,0,67,0,0,0,0,0,12,0,251,0,0,0,14,0,32,0,165,0,81,0,0,0,0,0,79,0,0,0,0,0,113,0,66,0,66,0,0,0,104,0,162,0,19,0,17,0,118,0,108,0,0,0,0,0,174,0,95,0,0,0,63,0,77,0,42,0,140,0,241,0,234,0,0,0,79,0,75,0,254,0,80,0,225,0,62,0,19,0,211,0,46,0,142,0,30,0,88,0,249,0,143,0,229,0,8,0,82,0,0,0,145,0,92,0,4,0,234,0,9,0,17,0,32,0,4,0,52,0,40,0,238,0,0,0,252,0,72,0,226,0,0,0,154,0,31,0,218,0,14,0,105,0,114,0,0,0,11,0,3,0,163,0,115,0,0,0,205,0,0,0,67,0,69,0,0,0,130,0,0,0,242,0,0,0,205,0,0,0,0,0,180,0,205,0,211,0,86,0,113,0,0,0,115,0,46,0,92,0,215,0,16,0,225,0,74,0,0,0,240,0,111,0,197,0,40,0,151,0,135,0,254,0,0,0,161,0,135,0,28,0,109,0,111,0,77,0,253,0,58,0,185,0,81,0,0,0,34,0,229,0,63,0,107,0,47,0,190,0,0,0,92,0,73,0,181,0,105,0,138,0,23,0,197,0,0,0,51,0,0,0,1,0,206,0,0,0,182,0,110,0,204,0,102,0,0,0,80,0,182,0,250,0,233,0,158,0,125,0,0,0,61,0,121,0,149,0,99,0,0,0,129,0,220,0,0,0,0,0,122,0,0,0,139,0,74,0,253,0,219,0,249,0,110,0,195,0,114,0,127,0,174,0,237,0,182,0,7,0,83,0,231,0,0,0,168,0,168,0,62,0,248,0,0,0,162,0,204,0,0,0,248,0,45,0,218,0,102,0,83,0,181,0,110,0,79,0,171,0,207,0,151,0,67,0,112,0,139,0,251,0,0,0,0,0,38,0,60,0,181,0,151,0,198,0,140,0,195,0,33,0,77,0,151,0,63,0,0,0,134,0,14,0,0,0,205,0,0,0,70,0,71,0,69,0,58,0,0,0,71,0,15,0,49,0,69,0,41,0,0,0,159,0,110,0,118,0,208,0,0,0,0,0,152,0,94,0,51,0,170,0,85,0,82,0,176,0,0,0,185,0,72,0,124,0,125,0,9,0,136,0,0,0,63,0,107,0,229,0,0,0,202,0,203,0,242,0,223,0,152,0,0,0,170,0,195,0,18,0,22,0,255,0,235,0,0,0,43,0,46,0,179,0,212,0,26,0,0,0,14,0,228,0,69,0,250,0,246,0,198,0,12,0,28,0,94,0,101,0,0,0,22,0,14,0,52,0,226,0,212,0,5,0,228,0,15,0,0,0,120,0,174,0,135,0,53,0,13,0,162,0,77,0,199,0,231,0,0,0,106,0,157,0,228,0,76,0,25,0,36,0,65,0,0,0,14,0,0,0,207,0,3,0,0,0,32,0,76,0,31,0,139,0,0,0,216,0,128,0,217,0,53,0,204,0,0,0,144,0,0,0,60,0,0,0,207,0,0,0,115,0,77,0,138,0,54,0,0,0,216,0,0,0,129,0,0,0,228,0,41,0,241,0,24,0,152,0,0,0,45,0,0,0,88,0,252,0,18,0,0,0,190,0);
signal scenario_full  : scenario_type := (0,0,203,31,147,31,147,30,140,31,75,31,151,31,151,30,14,31,253,31,51,31,147,31,94,31,36,31,123,31,184,31,30,31,201,31,149,31,223,31,223,30,75,31,159,31,248,31,173,31,183,31,182,31,182,30,76,31,29,31,180,31,184,31,184,30,191,31,89,31,78,31,232,31,123,31,133,31,207,31,185,31,83,31,229,31,229,30,196,31,158,31,111,31,164,31,34,31,55,31,55,30,245,31,245,31,245,30,85,31,147,31,69,31,59,31,59,30,23,31,23,30,47,31,92,31,185,31,8,31,236,31,114,31,55,31,125,31,65,31,241,31,243,31,193,31,140,31,140,30,239,31,239,30,143,31,176,31,214,31,132,31,169,31,35,31,37,31,84,31,15,31,162,31,76,31,190,31,152,31,202,31,202,30,202,29,104,31,109,31,169,31,169,30,188,31,179,31,224,31,46,31,93,31,159,31,159,30,159,29,10,31,83,31,63,31,52,31,217,31,131,31,133,31,231,31,74,31,195,31,123,31,64,31,15,31,38,31,219,31,249,31,234,31,153,31,153,30,185,31,69,31,195,31,206,31,178,31,127,31,109,31,115,31,121,31,166,31,169,31,160,31,202,31,163,31,163,30,35,31,183,31,154,31,200,31,200,31,211,31,194,31,97,31,156,31,124,31,140,31,140,30,14,31,84,31,140,31,49,31,49,30,49,29,49,28,49,27,49,26,143,31,214,31,145,31,148,31,118,31,43,31,43,30,138,31,113,31,113,30,188,31,145,31,41,31,18,31,127,31,93,31,90,31,227,31,227,30,209,31,180,31,66,31,88,31,133,31,99,31,192,31,133,31,166,31,205,31,173,31,88,31,59,31,126,31,182,31,238,31,57,31,216,31,160,31,158,31,158,30,48,31,20,31,247,31,12,31,36,31,247,31,125,31,101,31,225,31,132,31,150,31,117,31,86,31,185,31,185,30,33,31,33,30,33,29,29,31,235,31,235,31,150,31,126,31,126,30,202,31,12,31,142,31,150,31,198,31,217,31,103,31,148,31,148,30,212,31,212,30,102,31,100,31,252,31,187,31,219,31,190,31,82,31,82,30,82,29,212,31,212,30,212,29,8,31,141,31,202,31,202,30,238,31,166,31,129,31,53,31,87,31,186,31,186,30,186,29,126,31,243,31,179,31,162,31,162,30,162,29,3,31,188,31,85,31,42,31,42,30,42,29,35,31,59,31,135,31,64,31,64,30,219,31,219,30,219,29,33,31,33,30,33,29,232,31,20,31,191,31,65,31,179,31,87,31,36,31,36,30,36,29,242,31,18,31,5,31,45,31,45,30,118,31,192,31,137,31,93,31,93,30,80,31,8,31,90,31,110,31,23,31,23,30,79,31,238,31,213,31,123,31,107,31,107,30,20,31,20,30,20,29,107,31,11,31,89,31,41,31,53,31,53,30,85,31,236,31,211,31,211,30,226,31,158,31,158,30,158,29,158,28,162,31,178,31,20,31,89,31,55,31,55,30,55,29,86,31,123,31,237,31,56,31,139,31,105,31,23,31,218,31,150,31,45,31,45,30,127,31,127,30,136,31,136,30,61,31,76,31,242,31,68,31,245,31,39,31,122,31,211,31,61,31,215,31,23,31,82,31,168,31,1,31,15,31,99,31,99,30,121,31,151,31,225,31,147,31,245,31,68,31,190,31,181,31,243,31,243,30,192,31,197,31,197,30,188,31,31,31,44,31,3,31,121,31,81,31,113,31,113,30,11,31,138,31,152,31,156,31,67,31,67,30,67,29,12,31,251,31,251,30,14,31,32,31,165,31,81,31,81,30,81,29,79,31,79,30,79,29,113,31,66,31,66,31,66,30,104,31,162,31,19,31,17,31,118,31,108,31,108,30,108,29,174,31,95,31,95,30,63,31,77,31,42,31,140,31,241,31,234,31,234,30,79,31,75,31,254,31,80,31,225,31,62,31,19,31,211,31,46,31,142,31,30,31,88,31,249,31,143,31,229,31,8,31,82,31,82,30,145,31,92,31,4,31,234,31,9,31,17,31,32,31,4,31,52,31,40,31,238,31,238,30,252,31,72,31,226,31,226,30,154,31,31,31,218,31,14,31,105,31,114,31,114,30,11,31,3,31,163,31,115,31,115,30,205,31,205,30,67,31,69,31,69,30,130,31,130,30,242,31,242,30,205,31,205,30,205,29,180,31,205,31,211,31,86,31,113,31,113,30,115,31,46,31,92,31,215,31,16,31,225,31,74,31,74,30,240,31,111,31,197,31,40,31,151,31,135,31,254,31,254,30,161,31,135,31,28,31,109,31,111,31,77,31,253,31,58,31,185,31,81,31,81,30,34,31,229,31,63,31,107,31,47,31,190,31,190,30,92,31,73,31,181,31,105,31,138,31,23,31,197,31,197,30,51,31,51,30,1,31,206,31,206,30,182,31,110,31,204,31,102,31,102,30,80,31,182,31,250,31,233,31,158,31,125,31,125,30,61,31,121,31,149,31,99,31,99,30,129,31,220,31,220,30,220,29,122,31,122,30,139,31,74,31,253,31,219,31,249,31,110,31,195,31,114,31,127,31,174,31,237,31,182,31,7,31,83,31,231,31,231,30,168,31,168,31,62,31,248,31,248,30,162,31,204,31,204,30,248,31,45,31,218,31,102,31,83,31,181,31,110,31,79,31,171,31,207,31,151,31,67,31,112,31,139,31,251,31,251,30,251,29,38,31,60,31,181,31,151,31,198,31,140,31,195,31,33,31,77,31,151,31,63,31,63,30,134,31,14,31,14,30,205,31,205,30,70,31,71,31,69,31,58,31,58,30,71,31,15,31,49,31,69,31,41,31,41,30,159,31,110,31,118,31,208,31,208,30,208,29,152,31,94,31,51,31,170,31,85,31,82,31,176,31,176,30,185,31,72,31,124,31,125,31,9,31,136,31,136,30,63,31,107,31,229,31,229,30,202,31,203,31,242,31,223,31,152,31,152,30,170,31,195,31,18,31,22,31,255,31,235,31,235,30,43,31,46,31,179,31,212,31,26,31,26,30,14,31,228,31,69,31,250,31,246,31,198,31,12,31,28,31,94,31,101,31,101,30,22,31,14,31,52,31,226,31,212,31,5,31,228,31,15,31,15,30,120,31,174,31,135,31,53,31,13,31,162,31,77,31,199,31,231,31,231,30,106,31,157,31,228,31,76,31,25,31,36,31,65,31,65,30,14,31,14,30,207,31,3,31,3,30,32,31,76,31,31,31,139,31,139,30,216,31,128,31,217,31,53,31,204,31,204,30,144,31,144,30,60,31,60,30,207,31,207,30,115,31,77,31,138,31,54,31,54,30,216,31,216,30,129,31,129,30,228,31,41,31,241,31,24,31,152,31,152,30,45,31,45,30,88,31,252,31,18,31,18,30,190,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
