-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_248 is
end project_tb_248;

architecture project_tb_arch_248 of project_tb_248 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 969;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (172,0,5,0,0,0,107,0,219,0,121,0,19,0,129,0,34,0,64,0,185,0,69,0,198,0,111,0,100,0,0,0,85,0,0,0,0,0,125,0,216,0,0,0,203,0,142,0,142,0,168,0,158,0,112,0,128,0,227,0,127,0,155,0,105,0,68,0,214,0,251,0,232,0,41,0,137,0,4,0,149,0,117,0,136,0,237,0,254,0,192,0,0,0,45,0,114,0,183,0,113,0,0,0,62,0,85,0,137,0,79,0,232,0,136,0,26,0,190,0,92,0,169,0,118,0,135,0,50,0,196,0,186,0,195,0,87,0,0,0,192,0,0,0,0,0,148,0,211,0,238,0,0,0,164,0,69,0,134,0,204,0,0,0,50,0,37,0,80,0,195,0,22,0,118,0,215,0,76,0,0,0,0,0,61,0,0,0,0,0,0,0,230,0,54,0,20,0,243,0,0,0,0,0,211,0,229,0,220,0,13,0,237,0,170,0,61,0,0,0,15,0,169,0,69,0,0,0,101,0,93,0,30,0,22,0,73,0,163,0,146,0,253,0,206,0,0,0,0,0,0,0,200,0,116,0,116,0,0,0,45,0,144,0,144,0,64,0,0,0,56,0,25,0,0,0,121,0,62,0,0,0,119,0,0,0,0,0,31,0,180,0,54,0,193,0,74,0,0,0,139,0,0,0,134,0,106,0,0,0,6,0,64,0,0,0,224,0,206,0,188,0,193,0,174,0,4,0,177,0,121,0,172,0,97,0,0,0,197,0,17,0,144,0,199,0,128,0,87,0,239,0,183,0,113,0,197,0,91,0,248,0,63,0,208,0,38,0,4,0,233,0,153,0,231,0,79,0,206,0,181,0,125,0,95,0,156,0,16,0,190,0,6,0,164,0,119,0,0,0,49,0,0,0,0,0,61,0,58,0,171,0,89,0,74,0,95,0,155,0,84,0,171,0,39,0,102,0,0,0,45,0,100,0,242,0,0,0,213,0,0,0,95,0,162,0,164,0,59,0,222,0,75,0,216,0,23,0,8,0,0,0,226,0,251,0,112,0,188,0,185,0,177,0,0,0,55,0,208,0,30,0,0,0,0,0,10,0,191,0,0,0,176,0,74,0,196,0,216,0,49,0,183,0,110,0,100,0,0,0,7,0,119,0,4,0,241,0,0,0,0,0,91,0,0,0,1,0,179,0,86,0,251,0,102,0,91,0,224,0,64,0,180,0,220,0,57,0,204,0,103,0,108,0,238,0,173,0,93,0,255,0,161,0,16,0,226,0,0,0,137,0,218,0,21,0,151,0,58,0,27,0,208,0,95,0,92,0,142,0,46,0,194,0,0,0,0,0,21,0,0,0,226,0,132,0,32,0,159,0,36,0,9,0,82,0,13,0,13,0,0,0,0,0,80,0,0,0,78,0,143,0,93,0,169,0,159,0,113,0,230,0,168,0,155,0,133,0,44,0,26,0,0,0,190,0,225,0,2,0,72,0,166,0,0,0,41,0,146,0,87,0,38,0,234,0,117,0,0,0,239,0,253,0,4,0,116,0,38,0,160,0,104,0,0,0,239,0,147,0,63,0,108,0,0,0,176,0,161,0,36,0,188,0,113,0,71,0,204,0,192,0,127,0,18,0,140,0,179,0,0,0,214,0,92,0,108,0,0,0,21,0,134,0,136,0,26,0,11,0,85,0,22,0,0,0,244,0,0,0,167,0,112,0,99,0,114,0,0,0,151,0,101,0,233,0,0,0,174,0,12,0,82,0,104,0,0,0,160,0,197,0,91,0,85,0,194,0,206,0,202,0,66,0,166,0,205,0,32,0,50,0,0,0,79,0,168,0,0,0,5,0,173,0,213,0,35,0,0,0,155,0,0,0,215,0,0,0,150,0,17,0,220,0,135,0,143,0,107,0,94,0,183,0,0,0,122,0,119,0,166,0,189,0,62,0,158,0,220,0,24,0,227,0,32,0,50,0,57,0,231,0,126,0,143,0,4,0,46,0,0,0,200,0,0,0,116,0,134,0,230,0,36,0,132,0,223,0,83,0,66,0,204,0,0,0,164,0,61,0,0,0,189,0,181,0,19,0,170,0,201,0,197,0,56,0,99,0,198,0,148,0,14,0,170,0,71,0,194,0,200,0,160,0,191,0,0,0,175,0,20,0,178,0,0,0,0,0,36,0,123,0,114,0,243,0,157,0,54,0,66,0,18,0,228,0,45,0,108,0,0,0,235,0,0,0,166,0,241,0,214,0,0,0,17,0,17,0,6,0,0,0,0,0,251,0,0,0,116,0,18,0,141,0,12,0,183,0,170,0,0,0,0,0,203,0,44,0,226,0,241,0,0,0,0,0,28,0,0,0,41,0,246,0,156,0,78,0,0,0,192,0,178,0,87,0,0,0,0,0,0,0,201,0,0,0,0,0,219,0,31,0,0,0,56,0,69,0,132,0,242,0,27,0,127,0,13,0,0,0,158,0,103,0,23,0,150,0,246,0,227,0,73,0,214,0,166,0,0,0,211,0,209,0,179,0,39,0,0,0,236,0,66,0,169,0,188,0,1,0,30,0,6,0,164,0,138,0,72,0,34,0,49,0,105,0,0,0,214,0,49,0,0,0,221,0,0,0,79,0,64,0,191,0,0,0,0,0,71,0,107,0,239,0,141,0,36,0,147,0,182,0,0,0,254,0,14,0,0,0,220,0,45,0,230,0,0,0,105,0,108,0,117,0,240,0,0,0,0,0,252,0,0,0,19,0,187,0,232,0,0,0,208,0,0,0,176,0,253,0,186,0,128,0,89,0,23,0,217,0,243,0,15,0,78,0,147,0,87,0,47,0,0,0,0,0,118,0,130,0,0,0,0,0,81,0,148,0,230,0,138,0,0,0,141,0,134,0,0,0,210,0,33,0,201,0,180,0,192,0,49,0,0,0,208,0,0,0,0,0,63,0,139,0,16,0,27,0,19,0,199,0,227,0,79,0,197,0,191,0,43,0,156,0,16,0,81,0,130,0,207,0,213,0,184,0,89,0,94,0,179,0,143,0,234,0,159,0,84,0,32,0,214,0,37,0,0,0,237,0,199,0,128,0,138,0,235,0,149,0,121,0,0,0,191,0,0,0,49,0,0,0,25,0,34,0,0,0,168,0,0,0,87,0,241,0,139,0,28,0,108,0,109,0,8,0,0,0,218,0,89,0,63,0,223,0,232,0,253,0,0,0,253,0,2,0,0,0,169,0,48,0,0,0,209,0,248,0,0,0,198,0,100,0,0,0,135,0,152,0,28,0,24,0,178,0,90,0,143,0,123,0,105,0,0,0,153,0,118,0,0,0,108,0,0,0,244,0,141,0,0,0,222,0,250,0,72,0,0,0,90,0,50,0,155,0,126,0,235,0,57,0,0,0,0,0,29,0,0,0,0,0,170,0,13,0,38,0,126,0,219,0,173,0,74,0,197,0,31,0,0,0,212,0,110,0,14,0,90,0,113,0,130,0,197,0,0,0,0,0,143,0,202,0,177,0,104,0,92,0,80,0,0,0,75,0,226,0,0,0,82,0,34,0,205,0,28,0,201,0,0,0,94,0,0,0,208,0,124,0,55,0,0,0,100,0,213,0,237,0,185,0,227,0,0,0,2,0,168,0,34,0,204,0,126,0,124,0,95,0,0,0,5,0,79,0,0,0,0,0,0,0,0,0,85,0,67,0,132,0,245,0,238,0,162,0,24,0,109,0,220,0,197,0,0,0,98,0,0,0,139,0,109,0,40,0,220,0,0,0,246,0,205,0,0,0,106,0,196,0,159,0,92,0,49,0,78,0,190,0,29,0,176,0,0,0,138,0,0,0,16,0,120,0,191,0,189,0,1,0,93,0,0,0,57,0,146,0,0,0,0,0,188,0,154,0,117,0,74,0,227,0,244,0,39,0,136,0,69,0,167,0,5,0,87,0,124,0,160,0,120,0,41,0,124,0,206,0,86,0,128,0,66,0,0,0,65,0,0,0,15,0,166,0,111,0,0,0,0,0,173,0,183,0,204,0,0,0,0,0,192,0,159,0,8,0,121,0,210,0,0,0,218,0,136,0,178,0,64,0,246,0,0,0,122,0,91,0,148,0,175,0,192,0,82,0,220,0,97,0,109,0,0,0,218,0,208,0,39,0,93,0,227,0,1,0,0,0,0,0,136,0,181,0,238,0,157,0,171,0,188,0,31,0,43,0,47,0,1,0,27,0,215,0,194,0,201,0,133,0,11,0,0,0,1,0,199,0,235,0,22,0,0,0,0,0,0,0,213,0,0,0,121,0,233,0,35,0,30,0,0,0,0,0,91,0,106,0,9,0,138,0,165,0,0,0,96,0);
signal scenario_full  : scenario_type := (172,31,5,31,5,30,107,31,219,31,121,31,19,31,129,31,34,31,64,31,185,31,69,31,198,31,111,31,100,31,100,30,85,31,85,30,85,29,125,31,216,31,216,30,203,31,142,31,142,31,168,31,158,31,112,31,128,31,227,31,127,31,155,31,105,31,68,31,214,31,251,31,232,31,41,31,137,31,4,31,149,31,117,31,136,31,237,31,254,31,192,31,192,30,45,31,114,31,183,31,113,31,113,30,62,31,85,31,137,31,79,31,232,31,136,31,26,31,190,31,92,31,169,31,118,31,135,31,50,31,196,31,186,31,195,31,87,31,87,30,192,31,192,30,192,29,148,31,211,31,238,31,238,30,164,31,69,31,134,31,204,31,204,30,50,31,37,31,80,31,195,31,22,31,118,31,215,31,76,31,76,30,76,29,61,31,61,30,61,29,61,28,230,31,54,31,20,31,243,31,243,30,243,29,211,31,229,31,220,31,13,31,237,31,170,31,61,31,61,30,15,31,169,31,69,31,69,30,101,31,93,31,30,31,22,31,73,31,163,31,146,31,253,31,206,31,206,30,206,29,206,28,200,31,116,31,116,31,116,30,45,31,144,31,144,31,64,31,64,30,56,31,25,31,25,30,121,31,62,31,62,30,119,31,119,30,119,29,31,31,180,31,54,31,193,31,74,31,74,30,139,31,139,30,134,31,106,31,106,30,6,31,64,31,64,30,224,31,206,31,188,31,193,31,174,31,4,31,177,31,121,31,172,31,97,31,97,30,197,31,17,31,144,31,199,31,128,31,87,31,239,31,183,31,113,31,197,31,91,31,248,31,63,31,208,31,38,31,4,31,233,31,153,31,231,31,79,31,206,31,181,31,125,31,95,31,156,31,16,31,190,31,6,31,164,31,119,31,119,30,49,31,49,30,49,29,61,31,58,31,171,31,89,31,74,31,95,31,155,31,84,31,171,31,39,31,102,31,102,30,45,31,100,31,242,31,242,30,213,31,213,30,95,31,162,31,164,31,59,31,222,31,75,31,216,31,23,31,8,31,8,30,226,31,251,31,112,31,188,31,185,31,177,31,177,30,55,31,208,31,30,31,30,30,30,29,10,31,191,31,191,30,176,31,74,31,196,31,216,31,49,31,183,31,110,31,100,31,100,30,7,31,119,31,4,31,241,31,241,30,241,29,91,31,91,30,1,31,179,31,86,31,251,31,102,31,91,31,224,31,64,31,180,31,220,31,57,31,204,31,103,31,108,31,238,31,173,31,93,31,255,31,161,31,16,31,226,31,226,30,137,31,218,31,21,31,151,31,58,31,27,31,208,31,95,31,92,31,142,31,46,31,194,31,194,30,194,29,21,31,21,30,226,31,132,31,32,31,159,31,36,31,9,31,82,31,13,31,13,31,13,30,13,29,80,31,80,30,78,31,143,31,93,31,169,31,159,31,113,31,230,31,168,31,155,31,133,31,44,31,26,31,26,30,190,31,225,31,2,31,72,31,166,31,166,30,41,31,146,31,87,31,38,31,234,31,117,31,117,30,239,31,253,31,4,31,116,31,38,31,160,31,104,31,104,30,239,31,147,31,63,31,108,31,108,30,176,31,161,31,36,31,188,31,113,31,71,31,204,31,192,31,127,31,18,31,140,31,179,31,179,30,214,31,92,31,108,31,108,30,21,31,134,31,136,31,26,31,11,31,85,31,22,31,22,30,244,31,244,30,167,31,112,31,99,31,114,31,114,30,151,31,101,31,233,31,233,30,174,31,12,31,82,31,104,31,104,30,160,31,197,31,91,31,85,31,194,31,206,31,202,31,66,31,166,31,205,31,32,31,50,31,50,30,79,31,168,31,168,30,5,31,173,31,213,31,35,31,35,30,155,31,155,30,215,31,215,30,150,31,17,31,220,31,135,31,143,31,107,31,94,31,183,31,183,30,122,31,119,31,166,31,189,31,62,31,158,31,220,31,24,31,227,31,32,31,50,31,57,31,231,31,126,31,143,31,4,31,46,31,46,30,200,31,200,30,116,31,134,31,230,31,36,31,132,31,223,31,83,31,66,31,204,31,204,30,164,31,61,31,61,30,189,31,181,31,19,31,170,31,201,31,197,31,56,31,99,31,198,31,148,31,14,31,170,31,71,31,194,31,200,31,160,31,191,31,191,30,175,31,20,31,178,31,178,30,178,29,36,31,123,31,114,31,243,31,157,31,54,31,66,31,18,31,228,31,45,31,108,31,108,30,235,31,235,30,166,31,241,31,214,31,214,30,17,31,17,31,6,31,6,30,6,29,251,31,251,30,116,31,18,31,141,31,12,31,183,31,170,31,170,30,170,29,203,31,44,31,226,31,241,31,241,30,241,29,28,31,28,30,41,31,246,31,156,31,78,31,78,30,192,31,178,31,87,31,87,30,87,29,87,28,201,31,201,30,201,29,219,31,31,31,31,30,56,31,69,31,132,31,242,31,27,31,127,31,13,31,13,30,158,31,103,31,23,31,150,31,246,31,227,31,73,31,214,31,166,31,166,30,211,31,209,31,179,31,39,31,39,30,236,31,66,31,169,31,188,31,1,31,30,31,6,31,164,31,138,31,72,31,34,31,49,31,105,31,105,30,214,31,49,31,49,30,221,31,221,30,79,31,64,31,191,31,191,30,191,29,71,31,107,31,239,31,141,31,36,31,147,31,182,31,182,30,254,31,14,31,14,30,220,31,45,31,230,31,230,30,105,31,108,31,117,31,240,31,240,30,240,29,252,31,252,30,19,31,187,31,232,31,232,30,208,31,208,30,176,31,253,31,186,31,128,31,89,31,23,31,217,31,243,31,15,31,78,31,147,31,87,31,47,31,47,30,47,29,118,31,130,31,130,30,130,29,81,31,148,31,230,31,138,31,138,30,141,31,134,31,134,30,210,31,33,31,201,31,180,31,192,31,49,31,49,30,208,31,208,30,208,29,63,31,139,31,16,31,27,31,19,31,199,31,227,31,79,31,197,31,191,31,43,31,156,31,16,31,81,31,130,31,207,31,213,31,184,31,89,31,94,31,179,31,143,31,234,31,159,31,84,31,32,31,214,31,37,31,37,30,237,31,199,31,128,31,138,31,235,31,149,31,121,31,121,30,191,31,191,30,49,31,49,30,25,31,34,31,34,30,168,31,168,30,87,31,241,31,139,31,28,31,108,31,109,31,8,31,8,30,218,31,89,31,63,31,223,31,232,31,253,31,253,30,253,31,2,31,2,30,169,31,48,31,48,30,209,31,248,31,248,30,198,31,100,31,100,30,135,31,152,31,28,31,24,31,178,31,90,31,143,31,123,31,105,31,105,30,153,31,118,31,118,30,108,31,108,30,244,31,141,31,141,30,222,31,250,31,72,31,72,30,90,31,50,31,155,31,126,31,235,31,57,31,57,30,57,29,29,31,29,30,29,29,170,31,13,31,38,31,126,31,219,31,173,31,74,31,197,31,31,31,31,30,212,31,110,31,14,31,90,31,113,31,130,31,197,31,197,30,197,29,143,31,202,31,177,31,104,31,92,31,80,31,80,30,75,31,226,31,226,30,82,31,34,31,205,31,28,31,201,31,201,30,94,31,94,30,208,31,124,31,55,31,55,30,100,31,213,31,237,31,185,31,227,31,227,30,2,31,168,31,34,31,204,31,126,31,124,31,95,31,95,30,5,31,79,31,79,30,79,29,79,28,79,27,85,31,67,31,132,31,245,31,238,31,162,31,24,31,109,31,220,31,197,31,197,30,98,31,98,30,139,31,109,31,40,31,220,31,220,30,246,31,205,31,205,30,106,31,196,31,159,31,92,31,49,31,78,31,190,31,29,31,176,31,176,30,138,31,138,30,16,31,120,31,191,31,189,31,1,31,93,31,93,30,57,31,146,31,146,30,146,29,188,31,154,31,117,31,74,31,227,31,244,31,39,31,136,31,69,31,167,31,5,31,87,31,124,31,160,31,120,31,41,31,124,31,206,31,86,31,128,31,66,31,66,30,65,31,65,30,15,31,166,31,111,31,111,30,111,29,173,31,183,31,204,31,204,30,204,29,192,31,159,31,8,31,121,31,210,31,210,30,218,31,136,31,178,31,64,31,246,31,246,30,122,31,91,31,148,31,175,31,192,31,82,31,220,31,97,31,109,31,109,30,218,31,208,31,39,31,93,31,227,31,1,31,1,30,1,29,136,31,181,31,238,31,157,31,171,31,188,31,31,31,43,31,47,31,1,31,27,31,215,31,194,31,201,31,133,31,11,31,11,30,1,31,199,31,235,31,22,31,22,30,22,29,22,28,213,31,213,30,121,31,233,31,35,31,30,31,30,30,30,29,91,31,106,31,9,31,138,31,165,31,165,30,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
