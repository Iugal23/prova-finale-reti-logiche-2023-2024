-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_40 is
end project_tb_40;

architecture project_tb_arch_40 of project_tb_40 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 460;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,5,0,102,0,0,0,220,0,0,0,76,0,115,0,248,0,0,0,237,0,235,0,19,0,19,0,202,0,175,0,239,0,55,0,0,0,117,0,126,0,199,0,16,0,0,0,234,0,0,0,0,0,163,0,43,0,162,0,185,0,0,0,0,0,184,0,248,0,239,0,14,0,150,0,190,0,168,0,0,0,161,0,22,0,32,0,0,0,81,0,194,0,189,0,9,0,0,0,181,0,0,0,0,0,228,0,137,0,38,0,31,0,0,0,18,0,219,0,152,0,0,0,94,0,0,0,149,0,16,0,97,0,211,0,0,0,93,0,179,0,95,0,244,0,49,0,8,0,57,0,98,0,188,0,130,0,221,0,0,0,170,0,0,0,27,0,209,0,75,0,0,0,0,0,46,0,0,0,0,0,40,0,129,0,13,0,4,0,163,0,0,0,232,0,0,0,40,0,0,0,11,0,52,0,74,0,32,0,0,0,87,0,218,0,251,0,0,0,0,0,110,0,48,0,125,0,212,0,2,0,236,0,140,0,0,0,36,0,61,0,209,0,135,0,4,0,13,0,10,0,238,0,0,0,102,0,5,0,0,0,101,0,243,0,17,0,181,0,24,0,233,0,71,0,0,0,117,0,21,0,243,0,103,0,0,0,21,0,220,0,213,0,15,0,47,0,151,0,206,0,212,0,252,0,0,0,98,0,47,0,2,0,97,0,91,0,10,0,19,0,0,0,191,0,0,0,57,0,148,0,124,0,154,0,34,0,222,0,179,0,0,0,0,0,84,0,222,0,26,0,134,0,214,0,205,0,150,0,166,0,0,0,229,0,131,0,7,0,143,0,172,0,0,0,83,0,47,0,241,0,150,0,0,0,42,0,109,0,133,0,139,0,252,0,91,0,116,0,128,0,47,0,62,0,0,0,150,0,212,0,0,0,69,0,169,0,67,0,115,0,221,0,224,0,194,0,144,0,113,0,0,0,38,0,4,0,203,0,182,0,219,0,47,0,194,0,38,0,229,0,142,0,0,0,74,0,55,0,0,0,46,0,127,0,0,0,0,0,0,0,149,0,0,0,0,0,185,0,57,0,147,0,178,0,219,0,179,0,224,0,41,0,184,0,193,0,173,0,119,0,0,0,170,0,183,0,0,0,0,0,45,0,220,0,0,0,0,0,254,0,101,0,54,0,60,0,7,0,98,0,47,0,7,0,0,0,0,0,187,0,45,0,0,0,209,0,0,0,79,0,67,0,43,0,40,0,0,0,211,0,0,0,0,0,0,0,0,0,112,0,115,0,46,0,26,0,0,0,121,0,0,0,0,0,174,0,0,0,212,0,6,0,0,0,238,0,122,0,212,0,0,0,202,0,52,0,207,0,55,0,204,0,5,0,236,0,112,0,156,0,244,0,78,0,47,0,143,0,0,0,0,0,0,0,51,0,105,0,31,0,103,0,250,0,158,0,116,0,77,0,210,0,102,0,38,0,181,0,11,0,82,0,78,0,77,0,191,0,0,0,65,0,195,0,0,0,51,0,132,0,138,0,116,0,185,0,220,0,44,0,63,0,0,0,80,0,243,0,216,0,160,0,141,0,0,0,149,0,252,0,0,0,32,0,125,0,146,0,195,0,129,0,120,0,68,0,0,0,70,0,207,0,0,0,130,0,12,0,0,0,0,0,123,0,147,0,194,0,57,0,39,0,168,0,0,0,151,0,141,0,26,0,86,0,103,0,0,0,0,0,243,0,102,0,0,0,121,0,10,0,173,0,99,0,31,0,107,0,43,0,250,0,25,0,87,0,103,0,176,0,222,0,87,0,240,0,0,0,62,0,121,0,0,0,0,0,236,0,0,0,53,0,127,0,227,0,153,0,84,0,0,0,104,0,218,0,222,0,10,0,118,0,156,0,229,0,152,0,110,0,180,0,0,0,85,0,185,0,120,0,114,0,147,0,87,0,215,0,143,0,50,0,0,0,0,0,192,0,9,0,0,0,38,0,55,0,0,0,93,0,85,0,26,0,238,0,159,0,200,0,217,0,0,0,30,0,164,0,124,0,46,0,0,0,0,0,159,0);
signal scenario_full  : scenario_type := (0,0,5,31,102,31,102,30,220,31,220,30,76,31,115,31,248,31,248,30,237,31,235,31,19,31,19,31,202,31,175,31,239,31,55,31,55,30,117,31,126,31,199,31,16,31,16,30,234,31,234,30,234,29,163,31,43,31,162,31,185,31,185,30,185,29,184,31,248,31,239,31,14,31,150,31,190,31,168,31,168,30,161,31,22,31,32,31,32,30,81,31,194,31,189,31,9,31,9,30,181,31,181,30,181,29,228,31,137,31,38,31,31,31,31,30,18,31,219,31,152,31,152,30,94,31,94,30,149,31,16,31,97,31,211,31,211,30,93,31,179,31,95,31,244,31,49,31,8,31,57,31,98,31,188,31,130,31,221,31,221,30,170,31,170,30,27,31,209,31,75,31,75,30,75,29,46,31,46,30,46,29,40,31,129,31,13,31,4,31,163,31,163,30,232,31,232,30,40,31,40,30,11,31,52,31,74,31,32,31,32,30,87,31,218,31,251,31,251,30,251,29,110,31,48,31,125,31,212,31,2,31,236,31,140,31,140,30,36,31,61,31,209,31,135,31,4,31,13,31,10,31,238,31,238,30,102,31,5,31,5,30,101,31,243,31,17,31,181,31,24,31,233,31,71,31,71,30,117,31,21,31,243,31,103,31,103,30,21,31,220,31,213,31,15,31,47,31,151,31,206,31,212,31,252,31,252,30,98,31,47,31,2,31,97,31,91,31,10,31,19,31,19,30,191,31,191,30,57,31,148,31,124,31,154,31,34,31,222,31,179,31,179,30,179,29,84,31,222,31,26,31,134,31,214,31,205,31,150,31,166,31,166,30,229,31,131,31,7,31,143,31,172,31,172,30,83,31,47,31,241,31,150,31,150,30,42,31,109,31,133,31,139,31,252,31,91,31,116,31,128,31,47,31,62,31,62,30,150,31,212,31,212,30,69,31,169,31,67,31,115,31,221,31,224,31,194,31,144,31,113,31,113,30,38,31,4,31,203,31,182,31,219,31,47,31,194,31,38,31,229,31,142,31,142,30,74,31,55,31,55,30,46,31,127,31,127,30,127,29,127,28,149,31,149,30,149,29,185,31,57,31,147,31,178,31,219,31,179,31,224,31,41,31,184,31,193,31,173,31,119,31,119,30,170,31,183,31,183,30,183,29,45,31,220,31,220,30,220,29,254,31,101,31,54,31,60,31,7,31,98,31,47,31,7,31,7,30,7,29,187,31,45,31,45,30,209,31,209,30,79,31,67,31,43,31,40,31,40,30,211,31,211,30,211,29,211,28,211,27,112,31,115,31,46,31,26,31,26,30,121,31,121,30,121,29,174,31,174,30,212,31,6,31,6,30,238,31,122,31,212,31,212,30,202,31,52,31,207,31,55,31,204,31,5,31,236,31,112,31,156,31,244,31,78,31,47,31,143,31,143,30,143,29,143,28,51,31,105,31,31,31,103,31,250,31,158,31,116,31,77,31,210,31,102,31,38,31,181,31,11,31,82,31,78,31,77,31,191,31,191,30,65,31,195,31,195,30,51,31,132,31,138,31,116,31,185,31,220,31,44,31,63,31,63,30,80,31,243,31,216,31,160,31,141,31,141,30,149,31,252,31,252,30,32,31,125,31,146,31,195,31,129,31,120,31,68,31,68,30,70,31,207,31,207,30,130,31,12,31,12,30,12,29,123,31,147,31,194,31,57,31,39,31,168,31,168,30,151,31,141,31,26,31,86,31,103,31,103,30,103,29,243,31,102,31,102,30,121,31,10,31,173,31,99,31,31,31,107,31,43,31,250,31,25,31,87,31,103,31,176,31,222,31,87,31,240,31,240,30,62,31,121,31,121,30,121,29,236,31,236,30,53,31,127,31,227,31,153,31,84,31,84,30,104,31,218,31,222,31,10,31,118,31,156,31,229,31,152,31,110,31,180,31,180,30,85,31,185,31,120,31,114,31,147,31,87,31,215,31,143,31,50,31,50,30,50,29,192,31,9,31,9,30,38,31,55,31,55,30,93,31,85,31,26,31,238,31,159,31,200,31,217,31,217,30,30,31,164,31,124,31,46,31,46,30,46,29,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
