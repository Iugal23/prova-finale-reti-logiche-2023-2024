-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 615;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (18,0,190,0,0,0,0,0,0,0,26,0,100,0,72,0,0,0,252,0,45,0,139,0,200,0,0,0,0,0,77,0,70,0,45,0,7,0,0,0,117,0,30,0,10,0,8,0,1,0,251,0,144,0,190,0,37,0,14,0,99,0,11,0,132,0,0,0,0,0,251,0,69,0,173,0,101,0,195,0,0,0,65,0,224,0,14,0,167,0,0,0,150,0,218,0,0,0,0,0,83,0,187,0,92,0,0,0,24,0,8,0,180,0,88,0,236,0,223,0,0,0,20,0,121,0,249,0,0,0,222,0,37,0,0,0,66,0,133,0,53,0,19,0,0,0,242,0,17,0,186,0,142,0,55,0,2,0,11,0,124,0,0,0,182,0,159,0,129,0,129,0,184,0,0,0,187,0,155,0,54,0,63,0,190,0,223,0,112,0,31,0,0,0,30,0,27,0,36,0,224,0,226,0,49,0,227,0,169,0,17,0,6,0,1,0,0,0,209,0,0,0,66,0,230,0,229,0,0,0,10,0,174,0,132,0,47,0,90,0,24,0,97,0,66,0,199,0,0,0,65,0,87,0,81,0,152,0,69,0,0,0,219,0,129,0,138,0,0,0,28,0,243,0,35,0,11,0,244,0,251,0,208,0,190,0,44,0,123,0,155,0,88,0,2,0,47,0,195,0,211,0,0,0,0,0,98,0,178,0,0,0,0,0,0,0,1,0,0,0,150,0,2,0,10,0,106,0,198,0,140,0,0,0,0,0,146,0,107,0,15,0,201,0,33,0,155,0,63,0,0,0,20,0,17,0,154,0,16,0,240,0,168,0,48,0,250,0,240,0,171,0,234,0,212,0,99,0,245,0,135,0,180,0,36,0,236,0,0,0,61,0,169,0,132,0,145,0,210,0,219,0,179,0,231,0,125,0,89,0,25,0,0,0,154,0,26,0,76,0,93,0,192,0,44,0,0,0,204,0,119,0,0,0,0,0,90,0,57,0,251,0,127,0,33,0,61,0,0,0,182,0,216,0,238,0,133,0,232,0,143,0,200,0,192,0,226,0,240,0,0,0,252,0,253,0,195,0,209,0,122,0,37,0,0,0,253,0,243,0,15,0,220,0,152,0,0,0,51,0,63,0,14,0,158,0,0,0,101,0,34,0,41,0,200,0,134,0,249,0,37,0,199,0,247,0,123,0,154,0,0,0,170,0,20,0,78,0,0,0,139,0,108,0,0,0,17,0,0,0,154,0,247,0,82,0,106,0,46,0,94,0,114,0,90,0,0,0,64,0,146,0,106,0,239,0,0,0,16,0,0,0,73,0,226,0,37,0,177,0,0,0,0,0,91,0,55,0,133,0,241,0,220,0,163,0,41,0,168,0,1,0,0,0,111,0,70,0,128,0,244,0,142,0,149,0,0,0,54,0,128,0,233,0,26,0,0,0,148,0,202,0,32,0,228,0,242,0,41,0,233,0,245,0,12,0,216,0,192,0,223,0,103,0,0,0,0,0,0,0,18,0,201,0,87,0,83,0,0,0,83,0,189,0,60,0,183,0,135,0,243,0,16,0,57,0,147,0,0,0,47,0,0,0,69,0,113,0,22,0,122,0,99,0,197,0,229,0,124,0,211,0,0,0,59,0,255,0,220,0,231,0,0,0,59,0,80,0,103,0,247,0,0,0,91,0,166,0,0,0,64,0,103,0,193,0,57,0,163,0,186,0,0,0,158,0,115,0,32,0,208,0,57,0,198,0,247,0,76,0,201,0,18,0,109,0,165,0,216,0,115,0,0,0,9,0,199,0,141,0,166,0,0,0,253,0,233,0,5,0,90,0,64,0,6,0,56,0,169,0,34,0,67,0,193,0,228,0,16,0,221,0,98,0,58,0,251,0,14,0,39,0,93,0,219,0,218,0,102,0,167,0,13,0,98,0,183,0,40,0,53,0,223,0,122,0,100,0,7,0,239,0,206,0,254,0,36,0,183,0,168,0,164,0,23,0,103,0,98,0,172,0,38,0,200,0,248,0,0,0,158,0,216,0,254,0,23,0,137,0,228,0,191,0,87,0,128,0,192,0,0,0,171,0,131,0,179,0,140,0,48,0,22,0,191,0,104,0,199,0,104,0,183,0,100,0,0,0,35,0,224,0,172,0,175,0,0,0,0,0,34,0,0,0,114,0,18,0,24,0,22,0,0,0,123,0,8,0,233,0,64,0,0,0,49,0,151,0,0,0,0,0,131,0,196,0,243,0,217,0,0,0,0,0,148,0,157,0,96,0,52,0,222,0,94,0,129,0,128,0,66,0,70,0,45,0,143,0,4,0,98,0,88,0,0,0,168,0,0,0,0,0,148,0,15,0,0,0,201,0,0,0,122,0,248,0,52,0,18,0,11,0,126,0,225,0,66,0,0,0,188,0,0,0,0,0,0,0,0,0,141,0,187,0,0,0,37,0,0,0,124,0,0,0,106,0,130,0,254,0,0,0,162,0,227,0,96,0,12,0,124,0,242,0,92,0,156,0,115,0,40,0,104,0,154,0,144,0,163,0,113,0,215,0,240,0,26,0,56,0,198,0,14,0,0,0,121,0,149,0,0,0,89,0,60,0,106,0,127,0,53,0,121,0,150,0,224,0,156,0,161,0,5,0,6,0,16,0,0,0,1,0,0,0,134,0,0,0,4,0,58,0,91,0,252,0,233,0,113,0,185,0,203,0,179,0,98,0,40,0,0,0,191,0,0,0,0,0,0,0,132,0,193,0,121,0,0,0,72,0);
signal scenario_full  : scenario_type := (18,31,190,31,190,30,190,29,190,28,26,31,100,31,72,31,72,30,252,31,45,31,139,31,200,31,200,30,200,29,77,31,70,31,45,31,7,31,7,30,117,31,30,31,10,31,8,31,1,31,251,31,144,31,190,31,37,31,14,31,99,31,11,31,132,31,132,30,132,29,251,31,69,31,173,31,101,31,195,31,195,30,65,31,224,31,14,31,167,31,167,30,150,31,218,31,218,30,218,29,83,31,187,31,92,31,92,30,24,31,8,31,180,31,88,31,236,31,223,31,223,30,20,31,121,31,249,31,249,30,222,31,37,31,37,30,66,31,133,31,53,31,19,31,19,30,242,31,17,31,186,31,142,31,55,31,2,31,11,31,124,31,124,30,182,31,159,31,129,31,129,31,184,31,184,30,187,31,155,31,54,31,63,31,190,31,223,31,112,31,31,31,31,30,30,31,27,31,36,31,224,31,226,31,49,31,227,31,169,31,17,31,6,31,1,31,1,30,209,31,209,30,66,31,230,31,229,31,229,30,10,31,174,31,132,31,47,31,90,31,24,31,97,31,66,31,199,31,199,30,65,31,87,31,81,31,152,31,69,31,69,30,219,31,129,31,138,31,138,30,28,31,243,31,35,31,11,31,244,31,251,31,208,31,190,31,44,31,123,31,155,31,88,31,2,31,47,31,195,31,211,31,211,30,211,29,98,31,178,31,178,30,178,29,178,28,1,31,1,30,150,31,2,31,10,31,106,31,198,31,140,31,140,30,140,29,146,31,107,31,15,31,201,31,33,31,155,31,63,31,63,30,20,31,17,31,154,31,16,31,240,31,168,31,48,31,250,31,240,31,171,31,234,31,212,31,99,31,245,31,135,31,180,31,36,31,236,31,236,30,61,31,169,31,132,31,145,31,210,31,219,31,179,31,231,31,125,31,89,31,25,31,25,30,154,31,26,31,76,31,93,31,192,31,44,31,44,30,204,31,119,31,119,30,119,29,90,31,57,31,251,31,127,31,33,31,61,31,61,30,182,31,216,31,238,31,133,31,232,31,143,31,200,31,192,31,226,31,240,31,240,30,252,31,253,31,195,31,209,31,122,31,37,31,37,30,253,31,243,31,15,31,220,31,152,31,152,30,51,31,63,31,14,31,158,31,158,30,101,31,34,31,41,31,200,31,134,31,249,31,37,31,199,31,247,31,123,31,154,31,154,30,170,31,20,31,78,31,78,30,139,31,108,31,108,30,17,31,17,30,154,31,247,31,82,31,106,31,46,31,94,31,114,31,90,31,90,30,64,31,146,31,106,31,239,31,239,30,16,31,16,30,73,31,226,31,37,31,177,31,177,30,177,29,91,31,55,31,133,31,241,31,220,31,163,31,41,31,168,31,1,31,1,30,111,31,70,31,128,31,244,31,142,31,149,31,149,30,54,31,128,31,233,31,26,31,26,30,148,31,202,31,32,31,228,31,242,31,41,31,233,31,245,31,12,31,216,31,192,31,223,31,103,31,103,30,103,29,103,28,18,31,201,31,87,31,83,31,83,30,83,31,189,31,60,31,183,31,135,31,243,31,16,31,57,31,147,31,147,30,47,31,47,30,69,31,113,31,22,31,122,31,99,31,197,31,229,31,124,31,211,31,211,30,59,31,255,31,220,31,231,31,231,30,59,31,80,31,103,31,247,31,247,30,91,31,166,31,166,30,64,31,103,31,193,31,57,31,163,31,186,31,186,30,158,31,115,31,32,31,208,31,57,31,198,31,247,31,76,31,201,31,18,31,109,31,165,31,216,31,115,31,115,30,9,31,199,31,141,31,166,31,166,30,253,31,233,31,5,31,90,31,64,31,6,31,56,31,169,31,34,31,67,31,193,31,228,31,16,31,221,31,98,31,58,31,251,31,14,31,39,31,93,31,219,31,218,31,102,31,167,31,13,31,98,31,183,31,40,31,53,31,223,31,122,31,100,31,7,31,239,31,206,31,254,31,36,31,183,31,168,31,164,31,23,31,103,31,98,31,172,31,38,31,200,31,248,31,248,30,158,31,216,31,254,31,23,31,137,31,228,31,191,31,87,31,128,31,192,31,192,30,171,31,131,31,179,31,140,31,48,31,22,31,191,31,104,31,199,31,104,31,183,31,100,31,100,30,35,31,224,31,172,31,175,31,175,30,175,29,34,31,34,30,114,31,18,31,24,31,22,31,22,30,123,31,8,31,233,31,64,31,64,30,49,31,151,31,151,30,151,29,131,31,196,31,243,31,217,31,217,30,217,29,148,31,157,31,96,31,52,31,222,31,94,31,129,31,128,31,66,31,70,31,45,31,143,31,4,31,98,31,88,31,88,30,168,31,168,30,168,29,148,31,15,31,15,30,201,31,201,30,122,31,248,31,52,31,18,31,11,31,126,31,225,31,66,31,66,30,188,31,188,30,188,29,188,28,188,27,141,31,187,31,187,30,37,31,37,30,124,31,124,30,106,31,130,31,254,31,254,30,162,31,227,31,96,31,12,31,124,31,242,31,92,31,156,31,115,31,40,31,104,31,154,31,144,31,163,31,113,31,215,31,240,31,26,31,56,31,198,31,14,31,14,30,121,31,149,31,149,30,89,31,60,31,106,31,127,31,53,31,121,31,150,31,224,31,156,31,161,31,5,31,6,31,16,31,16,30,1,31,1,30,134,31,134,30,4,31,58,31,91,31,252,31,233,31,113,31,185,31,203,31,179,31,98,31,40,31,40,30,191,31,191,30,191,29,191,28,132,31,193,31,121,31,121,30,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
