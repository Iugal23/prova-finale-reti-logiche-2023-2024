-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_258 is
end project_tb_258;

architecture project_tb_arch_258 of project_tb_258 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 933;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (242,0,212,0,0,0,0,0,0,0,33,0,230,0,37,0,111,0,0,0,190,0,44,0,223,0,31,0,34,0,76,0,44,0,30,0,24,0,16,0,191,0,0,0,63,0,193,0,59,0,23,0,225,0,25,0,110,0,218,0,112,0,71,0,240,0,0,0,0,0,4,0,50,0,0,0,0,0,172,0,193,0,18,0,118,0,0,0,227,0,236,0,32,0,26,0,242,0,135,0,170,0,238,0,113,0,253,0,172,0,166,0,253,0,0,0,72,0,200,0,171,0,175,0,213,0,21,0,0,0,100,0,61,0,0,0,238,0,189,0,249,0,157,0,222,0,0,0,67,0,0,0,246,0,0,0,0,0,250,0,236,0,0,0,6,0,114,0,181,0,0,0,100,0,188,0,24,0,36,0,172,0,0,0,196,0,129,0,242,0,68,0,0,0,0,0,61,0,160,0,54,0,126,0,0,0,151,0,165,0,0,0,169,0,131,0,208,0,152,0,72,0,0,0,235,0,0,0,233,0,107,0,0,0,0,0,67,0,0,0,115,0,254,0,181,0,80,0,242,0,129,0,231,0,0,0,0,0,0,0,100,0,134,0,198,0,194,0,121,0,86,0,248,0,99,0,0,0,0,0,170,0,250,0,161,0,231,0,237,0,247,0,0,0,53,0,32,0,236,0,231,0,10,0,165,0,138,0,190,0,111,0,148,0,243,0,238,0,10,0,24,0,153,0,59,0,0,0,195,0,57,0,248,0,246,0,67,0,0,0,124,0,59,0,214,0,0,0,195,0,159,0,161,0,79,0,192,0,0,0,106,0,105,0,213,0,0,0,66,0,76,0,113,0,224,0,80,0,103,0,172,0,0,0,198,0,204,0,203,0,166,0,0,0,138,0,0,0,226,0,189,0,240,0,0,0,59,0,167,0,61,0,153,0,171,0,84,0,78,0,141,0,183,0,156,0,105,0,172,0,58,0,0,0,57,0,165,0,235,0,159,0,201,0,0,0,16,0,76,0,101,0,0,0,155,0,72,0,231,0,129,0,0,0,144,0,136,0,243,0,202,0,126,0,102,0,0,0,0,0,0,0,80,0,0,0,0,0,156,0,226,0,96,0,74,0,245,0,155,0,183,0,99,0,0,0,0,0,42,0,49,0,0,0,79,0,0,0,30,0,243,0,6,0,167,0,20,0,44,0,57,0,0,0,0,0,225,0,145,0,253,0,212,0,56,0,165,0,154,0,209,0,0,0,0,0,0,0,143,0,194,0,0,0,113,0,18,0,248,0,204,0,179,0,243,0,7,0,5,0,164,0,120,0,219,0,130,0,192,0,0,0,228,0,180,0,0,0,239,0,105,0,238,0,251,0,0,0,37,0,0,0,137,0,145,0,187,0,68,0,252,0,98,0,239,0,157,0,3,0,0,0,24,0,251,0,177,0,55,0,0,0,171,0,47,0,162,0,0,0,21,0,0,0,40,0,3,0,65,0,143,0,225,0,232,0,0,0,87,0,74,0,0,0,83,0,0,0,188,0,137,0,0,0,169,0,159,0,127,0,152,0,166,0,76,0,18,0,234,0,56,0,71,0,145,0,234,0,0,0,244,0,31,0,152,0,179,0,0,0,8,0,0,0,73,0,96,0,39,0,182,0,0,0,125,0,208,0,0,0,0,0,0,0,12,0,84,0,166,0,155,0,0,0,201,0,103,0,182,0,0,0,53,0,0,0,42,0,248,0,29,0,11,0,0,0,36,0,167,0,220,0,7,0,0,0,165,0,147,0,120,0,0,0,0,0,109,0,0,0,0,0,207,0,59,0,230,0,102,0,0,0,111,0,137,0,37,0,138,0,80,0,43,0,231,0,18,0,0,0,190,0,87,0,129,0,53,0,56,0,123,0,203,0,204,0,161,0,242,0,201,0,131,0,182,0,79,0,0,0,150,0,52,0,41,0,215,0,39,0,237,0,128,0,80,0,0,0,0,0,82,0,47,0,109,0,0,0,0,0,218,0,89,0,106,0,216,0,52,0,47,0,214,0,118,0,172,0,229,0,240,0,164,0,0,0,0,0,69,0,0,0,81,0,232,0,0,0,33,0,122,0,99,0,252,0,192,0,23,0,55,0,252,0,10,0,0,0,57,0,208,0,0,0,114,0,114,0,51,0,213,0,140,0,35,0,239,0,77,0,208,0,70,0,69,0,0,0,51,0,240,0,131,0,43,0,0,0,45,0,207,0,51,0,111,0,40,0,185,0,229,0,154,0,223,0,0,0,8,0,0,0,152,0,180,0,0,0,167,0,134,0,236,0,146,0,185,0,127,0,36,0,17,0,248,0,166,0,150,0,251,0,249,0,0,0,28,0,0,0,120,0,59,0,212,0,121,0,57,0,98,0,14,0,0,0,0,0,214,0,49,0,0,0,59,0,0,0,1,0,0,0,242,0,191,0,120,0,136,0,59,0,0,0,149,0,33,0,138,0,139,0,0,0,38,0,0,0,0,0,163,0,13,0,0,0,198,0,39,0,0,0,45,0,0,0,220,0,204,0,53,0,231,0,238,0,159,0,0,0,54,0,222,0,92,0,0,0,0,0,235,0,91,0,216,0,190,0,227,0,247,0,0,0,23,0,244,0,0,0,58,0,106,0,252,0,109,0,123,0,13,0,124,0,0,0,55,0,227,0,0,0,43,0,121,0,13,0,16,0,81,0,0,0,183,0,179,0,64,0,225,0,223,0,223,0,125,0,81,0,97,0,125,0,242,0,0,0,0,0,89,0,3,0,0,0,64,0,0,0,0,0,0,0,138,0,199,0,32,0,91,0,21,0,208,0,146,0,155,0,121,0,216,0,184,0,0,0,98,0,181,0,100,0,110,0,247,0,143,0,172,0,174,0,46,0,236,0,50,0,167,0,0,0,24,0,155,0,141,0,0,0,180,0,111,0,45,0,139,0,234,0,181,0,0,0,85,0,0,0,201,0,0,0,0,0,72,0,222,0,0,0,252,0,174,0,169,0,0,0,137,0,62,0,242,0,110,0,74,0,188,0,21,0,187,0,151,0,104,0,0,0,0,0,40,0,136,0,4,0,0,0,0,0,36,0,58,0,140,0,176,0,0,0,96,0,152,0,2,0,7,0,117,0,0,0,0,0,205,0,0,0,158,0,254,0,10,0,179,0,0,0,0,0,0,0,0,0,8,0,0,0,0,0,49,0,49,0,52,0,109,0,252,0,149,0,230,0,32,0,139,0,95,0,0,0,133,0,86,0,220,0,126,0,224,0,15,0,221,0,34,0,45,0,192,0,65,0,32,0,121,0,171,0,225,0,255,0,177,0,178,0,7,0,217,0,156,0,159,0,74,0,81,0,198,0,101,0,39,0,78,0,178,0,157,0,0,0,121,0,1,0,0,0,5,0,137,0,0,0,10,0,162,0,18,0,210,0,244,0,218,0,0,0,179,0,23,0,206,0,19,0,0,0,234,0,139,0,0,0,213,0,7,0,169,0,77,0,172,0,115,0,66,0,213,0,97,0,22,0,157,0,0,0,39,0,0,0,40,0,91,0,137,0,60,0,13,0,35,0,180,0,94,0,170,0,88,0,4,0,75,0,60,0,33,0,143,0,0,0,198,0,0,0,0,0,215,0,234,0,84,0,162,0,34,0,201,0,222,0,240,0,199,0,167,0,0,0,220,0,29,0,28,0,94,0,0,0,27,0,73,0,160,0,0,0,228,0,16,0,107,0,241,0,0,0,41,0,104,0,176,0,31,0,255,0,204,0,0,0,9,0,0,0,0,0,34,0,88,0,0,0,191,0,8,0,184,0,127,0,241,0,171,0,229,0,25,0,179,0,229,0,139,0,245,0,0,0,129,0,0,0,129,0,95,0,38,0,0,0,111,0,0,0,59,0,249,0,210,0,253,0,0,0,14,0,188,0,45,0,217,0,0,0,47,0,0,0,191,0,59,0,8,0,215,0,0,0,176,0,70,0,103,0,142,0,174,0,0,0,247,0,235,0,194,0,249,0,174,0,0,0,195,0,155,0,229,0,227,0,0,0,107,0,64,0,172,0,141,0,218,0,254,0,118,0,36,0,61,0,238,0,156,0,8,0,167,0,63,0,136,0,168,0,116,0,0,0,21,0,188,0,111,0,196,0,245,0,165,0,189,0,23,0,0,0,0,0,160,0,180,0,172,0,229,0);
signal scenario_full  : scenario_type := (242,31,212,31,212,30,212,29,212,28,33,31,230,31,37,31,111,31,111,30,190,31,44,31,223,31,31,31,34,31,76,31,44,31,30,31,24,31,16,31,191,31,191,30,63,31,193,31,59,31,23,31,225,31,25,31,110,31,218,31,112,31,71,31,240,31,240,30,240,29,4,31,50,31,50,30,50,29,172,31,193,31,18,31,118,31,118,30,227,31,236,31,32,31,26,31,242,31,135,31,170,31,238,31,113,31,253,31,172,31,166,31,253,31,253,30,72,31,200,31,171,31,175,31,213,31,21,31,21,30,100,31,61,31,61,30,238,31,189,31,249,31,157,31,222,31,222,30,67,31,67,30,246,31,246,30,246,29,250,31,236,31,236,30,6,31,114,31,181,31,181,30,100,31,188,31,24,31,36,31,172,31,172,30,196,31,129,31,242,31,68,31,68,30,68,29,61,31,160,31,54,31,126,31,126,30,151,31,165,31,165,30,169,31,131,31,208,31,152,31,72,31,72,30,235,31,235,30,233,31,107,31,107,30,107,29,67,31,67,30,115,31,254,31,181,31,80,31,242,31,129,31,231,31,231,30,231,29,231,28,100,31,134,31,198,31,194,31,121,31,86,31,248,31,99,31,99,30,99,29,170,31,250,31,161,31,231,31,237,31,247,31,247,30,53,31,32,31,236,31,231,31,10,31,165,31,138,31,190,31,111,31,148,31,243,31,238,31,10,31,24,31,153,31,59,31,59,30,195,31,57,31,248,31,246,31,67,31,67,30,124,31,59,31,214,31,214,30,195,31,159,31,161,31,79,31,192,31,192,30,106,31,105,31,213,31,213,30,66,31,76,31,113,31,224,31,80,31,103,31,172,31,172,30,198,31,204,31,203,31,166,31,166,30,138,31,138,30,226,31,189,31,240,31,240,30,59,31,167,31,61,31,153,31,171,31,84,31,78,31,141,31,183,31,156,31,105,31,172,31,58,31,58,30,57,31,165,31,235,31,159,31,201,31,201,30,16,31,76,31,101,31,101,30,155,31,72,31,231,31,129,31,129,30,144,31,136,31,243,31,202,31,126,31,102,31,102,30,102,29,102,28,80,31,80,30,80,29,156,31,226,31,96,31,74,31,245,31,155,31,183,31,99,31,99,30,99,29,42,31,49,31,49,30,79,31,79,30,30,31,243,31,6,31,167,31,20,31,44,31,57,31,57,30,57,29,225,31,145,31,253,31,212,31,56,31,165,31,154,31,209,31,209,30,209,29,209,28,143,31,194,31,194,30,113,31,18,31,248,31,204,31,179,31,243,31,7,31,5,31,164,31,120,31,219,31,130,31,192,31,192,30,228,31,180,31,180,30,239,31,105,31,238,31,251,31,251,30,37,31,37,30,137,31,145,31,187,31,68,31,252,31,98,31,239,31,157,31,3,31,3,30,24,31,251,31,177,31,55,31,55,30,171,31,47,31,162,31,162,30,21,31,21,30,40,31,3,31,65,31,143,31,225,31,232,31,232,30,87,31,74,31,74,30,83,31,83,30,188,31,137,31,137,30,169,31,159,31,127,31,152,31,166,31,76,31,18,31,234,31,56,31,71,31,145,31,234,31,234,30,244,31,31,31,152,31,179,31,179,30,8,31,8,30,73,31,96,31,39,31,182,31,182,30,125,31,208,31,208,30,208,29,208,28,12,31,84,31,166,31,155,31,155,30,201,31,103,31,182,31,182,30,53,31,53,30,42,31,248,31,29,31,11,31,11,30,36,31,167,31,220,31,7,31,7,30,165,31,147,31,120,31,120,30,120,29,109,31,109,30,109,29,207,31,59,31,230,31,102,31,102,30,111,31,137,31,37,31,138,31,80,31,43,31,231,31,18,31,18,30,190,31,87,31,129,31,53,31,56,31,123,31,203,31,204,31,161,31,242,31,201,31,131,31,182,31,79,31,79,30,150,31,52,31,41,31,215,31,39,31,237,31,128,31,80,31,80,30,80,29,82,31,47,31,109,31,109,30,109,29,218,31,89,31,106,31,216,31,52,31,47,31,214,31,118,31,172,31,229,31,240,31,164,31,164,30,164,29,69,31,69,30,81,31,232,31,232,30,33,31,122,31,99,31,252,31,192,31,23,31,55,31,252,31,10,31,10,30,57,31,208,31,208,30,114,31,114,31,51,31,213,31,140,31,35,31,239,31,77,31,208,31,70,31,69,31,69,30,51,31,240,31,131,31,43,31,43,30,45,31,207,31,51,31,111,31,40,31,185,31,229,31,154,31,223,31,223,30,8,31,8,30,152,31,180,31,180,30,167,31,134,31,236,31,146,31,185,31,127,31,36,31,17,31,248,31,166,31,150,31,251,31,249,31,249,30,28,31,28,30,120,31,59,31,212,31,121,31,57,31,98,31,14,31,14,30,14,29,214,31,49,31,49,30,59,31,59,30,1,31,1,30,242,31,191,31,120,31,136,31,59,31,59,30,149,31,33,31,138,31,139,31,139,30,38,31,38,30,38,29,163,31,13,31,13,30,198,31,39,31,39,30,45,31,45,30,220,31,204,31,53,31,231,31,238,31,159,31,159,30,54,31,222,31,92,31,92,30,92,29,235,31,91,31,216,31,190,31,227,31,247,31,247,30,23,31,244,31,244,30,58,31,106,31,252,31,109,31,123,31,13,31,124,31,124,30,55,31,227,31,227,30,43,31,121,31,13,31,16,31,81,31,81,30,183,31,179,31,64,31,225,31,223,31,223,31,125,31,81,31,97,31,125,31,242,31,242,30,242,29,89,31,3,31,3,30,64,31,64,30,64,29,64,28,138,31,199,31,32,31,91,31,21,31,208,31,146,31,155,31,121,31,216,31,184,31,184,30,98,31,181,31,100,31,110,31,247,31,143,31,172,31,174,31,46,31,236,31,50,31,167,31,167,30,24,31,155,31,141,31,141,30,180,31,111,31,45,31,139,31,234,31,181,31,181,30,85,31,85,30,201,31,201,30,201,29,72,31,222,31,222,30,252,31,174,31,169,31,169,30,137,31,62,31,242,31,110,31,74,31,188,31,21,31,187,31,151,31,104,31,104,30,104,29,40,31,136,31,4,31,4,30,4,29,36,31,58,31,140,31,176,31,176,30,96,31,152,31,2,31,7,31,117,31,117,30,117,29,205,31,205,30,158,31,254,31,10,31,179,31,179,30,179,29,179,28,179,27,8,31,8,30,8,29,49,31,49,31,52,31,109,31,252,31,149,31,230,31,32,31,139,31,95,31,95,30,133,31,86,31,220,31,126,31,224,31,15,31,221,31,34,31,45,31,192,31,65,31,32,31,121,31,171,31,225,31,255,31,177,31,178,31,7,31,217,31,156,31,159,31,74,31,81,31,198,31,101,31,39,31,78,31,178,31,157,31,157,30,121,31,1,31,1,30,5,31,137,31,137,30,10,31,162,31,18,31,210,31,244,31,218,31,218,30,179,31,23,31,206,31,19,31,19,30,234,31,139,31,139,30,213,31,7,31,169,31,77,31,172,31,115,31,66,31,213,31,97,31,22,31,157,31,157,30,39,31,39,30,40,31,91,31,137,31,60,31,13,31,35,31,180,31,94,31,170,31,88,31,4,31,75,31,60,31,33,31,143,31,143,30,198,31,198,30,198,29,215,31,234,31,84,31,162,31,34,31,201,31,222,31,240,31,199,31,167,31,167,30,220,31,29,31,28,31,94,31,94,30,27,31,73,31,160,31,160,30,228,31,16,31,107,31,241,31,241,30,41,31,104,31,176,31,31,31,255,31,204,31,204,30,9,31,9,30,9,29,34,31,88,31,88,30,191,31,8,31,184,31,127,31,241,31,171,31,229,31,25,31,179,31,229,31,139,31,245,31,245,30,129,31,129,30,129,31,95,31,38,31,38,30,111,31,111,30,59,31,249,31,210,31,253,31,253,30,14,31,188,31,45,31,217,31,217,30,47,31,47,30,191,31,59,31,8,31,215,31,215,30,176,31,70,31,103,31,142,31,174,31,174,30,247,31,235,31,194,31,249,31,174,31,174,30,195,31,155,31,229,31,227,31,227,30,107,31,64,31,172,31,141,31,218,31,254,31,118,31,36,31,61,31,238,31,156,31,8,31,167,31,63,31,136,31,168,31,116,31,116,30,21,31,188,31,111,31,196,31,245,31,165,31,189,31,23,31,23,30,23,29,160,31,180,31,172,31,229,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
