-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_483 is
end project_tb_483;

architecture project_tb_arch_483 of project_tb_483 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 807;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (18,0,216,0,155,0,0,0,130,0,139,0,156,0,0,0,187,0,0,0,1,0,0,0,57,0,14,0,154,0,33,0,0,0,140,0,33,0,52,0,0,0,191,0,155,0,0,0,155,0,0,0,93,0,116,0,0,0,0,0,72,0,31,0,142,0,195,0,10,0,162,0,76,0,100,0,0,0,38,0,127,0,0,0,230,0,238,0,78,0,68,0,63,0,180,0,5,0,150,0,203,0,0,0,0,0,121,0,0,0,0,0,140,0,166,0,246,0,54,0,164,0,0,0,92,0,168,0,119,0,202,0,0,0,113,0,234,0,0,0,213,0,206,0,32,0,166,0,153,0,135,0,187,0,136,0,119,0,0,0,239,0,62,0,87,0,172,0,153,0,232,0,230,0,28,0,51,0,0,0,72,0,0,0,164,0,0,0,148,0,215,0,243,0,114,0,47,0,9,0,180,0,115,0,163,0,136,0,76,0,54,0,0,0,37,0,0,0,213,0,0,0,174,0,117,0,11,0,221,0,29,0,239,0,0,0,42,0,0,0,73,0,0,0,198,0,235,0,22,0,223,0,0,0,197,0,227,0,154,0,0,0,93,0,51,0,81,0,128,0,183,0,145,0,171,0,33,0,0,0,73,0,87,0,12,0,0,0,43,0,42,0,0,0,0,0,68,0,77,0,0,0,0,0,162,0,106,0,55,0,68,0,221,0,153,0,0,0,0,0,203,0,6,0,0,0,0,0,90,0,128,0,0,0,11,0,229,0,233,0,0,0,114,0,146,0,39,0,17,0,205,0,0,0,158,0,43,0,21,0,0,0,255,0,31,0,134,0,111,0,0,0,69,0,171,0,8,0,12,0,132,0,0,0,235,0,39,0,89,0,219,0,139,0,225,0,0,0,86,0,148,0,222,0,187,0,0,0,172,0,0,0,44,0,73,0,0,0,172,0,32,0,218,0,52,0,194,0,32,0,29,0,205,0,103,0,0,0,148,0,84,0,0,0,0,0,46,0,200,0,0,0,55,0,0,0,0,0,13,0,0,0,136,0,244,0,253,0,15,0,26,0,0,0,132,0,61,0,166,0,0,0,72,0,0,0,127,0,0,0,69,0,160,0,0,0,163,0,198,0,145,0,51,0,206,0,167,0,227,0,39,0,88,0,12,0,40,0,188,0,0,0,0,0,96,0,200,0,0,0,20,0,0,0,0,0,139,0,117,0,0,0,198,0,149,0,240,0,92,0,213,0,0,0,71,0,207,0,24,0,49,0,158,0,203,0,0,0,70,0,28,0,160,0,144,0,26,0,144,0,103,0,8,0,93,0,216,0,0,0,0,0,253,0,214,0,143,0,0,0,54,0,0,0,156,0,28,0,85,0,234,0,56,0,36,0,0,0,178,0,50,0,94,0,86,0,211,0,98,0,150,0,183,0,164,0,124,0,0,0,43,0,121,0,254,0,0,0,28,0,211,0,190,0,183,0,68,0,115,0,143,0,173,0,228,0,0,0,0,0,194,0,162,0,127,0,52,0,170,0,75,0,5,0,205,0,80,0,216,0,224,0,254,0,53,0,170,0,0,0,0,0,42,0,0,0,220,0,90,0,129,0,148,0,205,0,191,0,122,0,239,0,254,0,0,0,224,0,133,0,108,0,75,0,212,0,0,0,149,0,0,0,159,0,88,0,0,0,103,0,120,0,167,0,21,0,1,0,73,0,0,0,107,0,0,0,219,0,182,0,104,0,103,0,41,0,0,0,108,0,243,0,221,0,52,0,50,0,222,0,0,0,72,0,103,0,144,0,88,0,147,0,17,0,162,0,0,0,209,0,160,0,0,0,93,0,0,0,108,0,56,0,83,0,239,0,0,0,228,0,20,0,138,0,51,0,219,0,209,0,0,0,0,0,149,0,122,0,138,0,233,0,140,0,69,0,246,0,235,0,230,0,78,0,213,0,39,0,242,0,208,0,235,0,0,0,253,0,16,0,238,0,62,0,108,0,94,0,38,0,206,0,231,0,11,0,74,0,246,0,0,0,158,0,161,0,129,0,185,0,0,0,115,0,45,0,93,0,129,0,31,0,0,0,12,0,56,0,0,0,0,0,26,0,39,0,213,0,218,0,197,0,122,0,0,0,60,0,51,0,227,0,4,0,152,0,252,0,13,0,0,0,199,0,222,0,177,0,0,0,86,0,155,0,12,0,23,0,144,0,0,0,214,0,233,0,63,0,0,0,0,0,247,0,0,0,120,0,154,0,223,0,118,0,0,0,245,0,208,0,67,0,0,0,87,0,145,0,195,0,133,0,2,0,154,0,172,0,189,0,0,0,161,0,174,0,213,0,116,0,83,0,103,0,43,0,0,0,183,0,243,0,99,0,67,0,66,0,0,0,79,0,89,0,151,0,165,0,0,0,197,0,251,0,143,0,34,0,10,0,161,0,167,0,55,0,218,0,185,0,222,0,44,0,132,0,111,0,169,0,26,0,31,0,81,0,5,0,205,0,144,0,181,0,84,0,0,0,0,0,60,0,106,0,150,0,4,0,146,0,44,0,0,0,81,0,146,0,35,0,117,0,13,0,11,0,102,0,220,0,67,0,58,0,0,0,0,0,73,0,30,0,63,0,0,0,0,0,0,0,70,0,133,0,232,0,78,0,0,0,221,0,172,0,33,0,100,0,0,0,90,0,255,0,139,0,14,0,0,0,40,0,21,0,62,0,109,0,62,0,40,0,96,0,0,0,167,0,236,0,31,0,31,0,223,0,0,0,147,0,128,0,4,0,213,0,197,0,112,0,189,0,0,0,93,0,90,0,21,0,169,0,234,0,0,0,123,0,191,0,0,0,113,0,208,0,214,0,0,0,83,0,219,0,111,0,255,0,181,0,64,0,206,0,44,0,0,0,168,0,204,0,20,0,0,0,188,0,34,0,36,0,99,0,36,0,132,0,71,0,0,0,5,0,218,0,77,0,0,0,0,0,21,0,77,0,125,0,123,0,19,0,210,0,151,0,41,0,253,0,140,0,0,0,71,0,65,0,243,0,49,0,173,0,212,0,240,0,168,0,210,0,127,0,109,0,118,0,72,0,238,0,35,0,0,0,0,0,0,0,169,0,253,0,0,0,30,0,37,0,58,0,106,0,114,0,38,0,4,0,29,0,10,0,9,0,0,0,219,0,0,0,123,0,0,0,108,0,148,0,12,0,30,0,0,0,241,0,140,0,223,0,98,0,31,0,0,0,248,0,135,0,0,0,112,0,240,0,177,0,223,0,80,0,9,0,193,0,0,0,36,0,80,0,189,0,0,0,0,0,94,0,154,0,0,0,0,0,90,0,51,0,96,0,159,0,60,0,142,0,50,0,12,0,53,0,21,0,143,0,10,0,251,0,0,0,97,0,61,0,0,0,129,0,0,0,239,0,53,0,0,0,0,0,103,0,12,0,95,0,0,0,113,0,110,0,176,0,0,0,0,0,24,0,39,0,246,0,11,0,0,0,197,0,73,0,19,0,232,0,0,0,117,0,161,0,101,0,0,0,235,0,0,0,0,0,224,0,114,0,203,0,158,0,231,0,0,0,9,0,169,0,93,0,0,0,0,0,208,0,132,0,46,0,124,0,17,0,108,0,41,0,184,0);
signal scenario_full  : scenario_type := (18,31,216,31,155,31,155,30,130,31,139,31,156,31,156,30,187,31,187,30,1,31,1,30,57,31,14,31,154,31,33,31,33,30,140,31,33,31,52,31,52,30,191,31,155,31,155,30,155,31,155,30,93,31,116,31,116,30,116,29,72,31,31,31,142,31,195,31,10,31,162,31,76,31,100,31,100,30,38,31,127,31,127,30,230,31,238,31,78,31,68,31,63,31,180,31,5,31,150,31,203,31,203,30,203,29,121,31,121,30,121,29,140,31,166,31,246,31,54,31,164,31,164,30,92,31,168,31,119,31,202,31,202,30,113,31,234,31,234,30,213,31,206,31,32,31,166,31,153,31,135,31,187,31,136,31,119,31,119,30,239,31,62,31,87,31,172,31,153,31,232,31,230,31,28,31,51,31,51,30,72,31,72,30,164,31,164,30,148,31,215,31,243,31,114,31,47,31,9,31,180,31,115,31,163,31,136,31,76,31,54,31,54,30,37,31,37,30,213,31,213,30,174,31,117,31,11,31,221,31,29,31,239,31,239,30,42,31,42,30,73,31,73,30,198,31,235,31,22,31,223,31,223,30,197,31,227,31,154,31,154,30,93,31,51,31,81,31,128,31,183,31,145,31,171,31,33,31,33,30,73,31,87,31,12,31,12,30,43,31,42,31,42,30,42,29,68,31,77,31,77,30,77,29,162,31,106,31,55,31,68,31,221,31,153,31,153,30,153,29,203,31,6,31,6,30,6,29,90,31,128,31,128,30,11,31,229,31,233,31,233,30,114,31,146,31,39,31,17,31,205,31,205,30,158,31,43,31,21,31,21,30,255,31,31,31,134,31,111,31,111,30,69,31,171,31,8,31,12,31,132,31,132,30,235,31,39,31,89,31,219,31,139,31,225,31,225,30,86,31,148,31,222,31,187,31,187,30,172,31,172,30,44,31,73,31,73,30,172,31,32,31,218,31,52,31,194,31,32,31,29,31,205,31,103,31,103,30,148,31,84,31,84,30,84,29,46,31,200,31,200,30,55,31,55,30,55,29,13,31,13,30,136,31,244,31,253,31,15,31,26,31,26,30,132,31,61,31,166,31,166,30,72,31,72,30,127,31,127,30,69,31,160,31,160,30,163,31,198,31,145,31,51,31,206,31,167,31,227,31,39,31,88,31,12,31,40,31,188,31,188,30,188,29,96,31,200,31,200,30,20,31,20,30,20,29,139,31,117,31,117,30,198,31,149,31,240,31,92,31,213,31,213,30,71,31,207,31,24,31,49,31,158,31,203,31,203,30,70,31,28,31,160,31,144,31,26,31,144,31,103,31,8,31,93,31,216,31,216,30,216,29,253,31,214,31,143,31,143,30,54,31,54,30,156,31,28,31,85,31,234,31,56,31,36,31,36,30,178,31,50,31,94,31,86,31,211,31,98,31,150,31,183,31,164,31,124,31,124,30,43,31,121,31,254,31,254,30,28,31,211,31,190,31,183,31,68,31,115,31,143,31,173,31,228,31,228,30,228,29,194,31,162,31,127,31,52,31,170,31,75,31,5,31,205,31,80,31,216,31,224,31,254,31,53,31,170,31,170,30,170,29,42,31,42,30,220,31,90,31,129,31,148,31,205,31,191,31,122,31,239,31,254,31,254,30,224,31,133,31,108,31,75,31,212,31,212,30,149,31,149,30,159,31,88,31,88,30,103,31,120,31,167,31,21,31,1,31,73,31,73,30,107,31,107,30,219,31,182,31,104,31,103,31,41,31,41,30,108,31,243,31,221,31,52,31,50,31,222,31,222,30,72,31,103,31,144,31,88,31,147,31,17,31,162,31,162,30,209,31,160,31,160,30,93,31,93,30,108,31,56,31,83,31,239,31,239,30,228,31,20,31,138,31,51,31,219,31,209,31,209,30,209,29,149,31,122,31,138,31,233,31,140,31,69,31,246,31,235,31,230,31,78,31,213,31,39,31,242,31,208,31,235,31,235,30,253,31,16,31,238,31,62,31,108,31,94,31,38,31,206,31,231,31,11,31,74,31,246,31,246,30,158,31,161,31,129,31,185,31,185,30,115,31,45,31,93,31,129,31,31,31,31,30,12,31,56,31,56,30,56,29,26,31,39,31,213,31,218,31,197,31,122,31,122,30,60,31,51,31,227,31,4,31,152,31,252,31,13,31,13,30,199,31,222,31,177,31,177,30,86,31,155,31,12,31,23,31,144,31,144,30,214,31,233,31,63,31,63,30,63,29,247,31,247,30,120,31,154,31,223,31,118,31,118,30,245,31,208,31,67,31,67,30,87,31,145,31,195,31,133,31,2,31,154,31,172,31,189,31,189,30,161,31,174,31,213,31,116,31,83,31,103,31,43,31,43,30,183,31,243,31,99,31,67,31,66,31,66,30,79,31,89,31,151,31,165,31,165,30,197,31,251,31,143,31,34,31,10,31,161,31,167,31,55,31,218,31,185,31,222,31,44,31,132,31,111,31,169,31,26,31,31,31,81,31,5,31,205,31,144,31,181,31,84,31,84,30,84,29,60,31,106,31,150,31,4,31,146,31,44,31,44,30,81,31,146,31,35,31,117,31,13,31,11,31,102,31,220,31,67,31,58,31,58,30,58,29,73,31,30,31,63,31,63,30,63,29,63,28,70,31,133,31,232,31,78,31,78,30,221,31,172,31,33,31,100,31,100,30,90,31,255,31,139,31,14,31,14,30,40,31,21,31,62,31,109,31,62,31,40,31,96,31,96,30,167,31,236,31,31,31,31,31,223,31,223,30,147,31,128,31,4,31,213,31,197,31,112,31,189,31,189,30,93,31,90,31,21,31,169,31,234,31,234,30,123,31,191,31,191,30,113,31,208,31,214,31,214,30,83,31,219,31,111,31,255,31,181,31,64,31,206,31,44,31,44,30,168,31,204,31,20,31,20,30,188,31,34,31,36,31,99,31,36,31,132,31,71,31,71,30,5,31,218,31,77,31,77,30,77,29,21,31,77,31,125,31,123,31,19,31,210,31,151,31,41,31,253,31,140,31,140,30,71,31,65,31,243,31,49,31,173,31,212,31,240,31,168,31,210,31,127,31,109,31,118,31,72,31,238,31,35,31,35,30,35,29,35,28,169,31,253,31,253,30,30,31,37,31,58,31,106,31,114,31,38,31,4,31,29,31,10,31,9,31,9,30,219,31,219,30,123,31,123,30,108,31,148,31,12,31,30,31,30,30,241,31,140,31,223,31,98,31,31,31,31,30,248,31,135,31,135,30,112,31,240,31,177,31,223,31,80,31,9,31,193,31,193,30,36,31,80,31,189,31,189,30,189,29,94,31,154,31,154,30,154,29,90,31,51,31,96,31,159,31,60,31,142,31,50,31,12,31,53,31,21,31,143,31,10,31,251,31,251,30,97,31,61,31,61,30,129,31,129,30,239,31,53,31,53,30,53,29,103,31,12,31,95,31,95,30,113,31,110,31,176,31,176,30,176,29,24,31,39,31,246,31,11,31,11,30,197,31,73,31,19,31,232,31,232,30,117,31,161,31,101,31,101,30,235,31,235,30,235,29,224,31,114,31,203,31,158,31,231,31,231,30,9,31,169,31,93,31,93,30,93,29,208,31,132,31,46,31,124,31,17,31,108,31,41,31,184,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
