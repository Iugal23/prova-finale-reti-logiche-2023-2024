-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_369 is
end project_tb_369;

architecture project_tb_arch_369 of project_tb_369 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 601;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,195,0,188,0,190,0,237,0,0,0,125,0,89,0,236,0,0,0,105,0,12,0,184,0,84,0,174,0,28,0,47,0,78,0,0,0,0,0,191,0,99,0,171,0,89,0,236,0,0,0,149,0,218,0,43,0,155,0,0,0,64,0,101,0,204,0,0,0,0,0,90,0,130,0,0,0,239,0,235,0,237,0,87,0,233,0,0,0,89,0,34,0,243,0,0,0,0,0,0,0,20,0,0,0,202,0,0,0,122,0,84,0,10,0,0,0,0,0,151,0,240,0,53,0,131,0,90,0,114,0,225,0,0,0,49,0,31,0,0,0,76,0,79,0,127,0,174,0,53,0,142,0,41,0,44,0,0,0,216,0,0,0,30,0,11,0,254,0,14,0,47,0,6,0,219,0,0,0,167,0,225,0,184,0,191,0,254,0,0,0,64,0,227,0,31,0,212,0,0,0,136,0,36,0,105,0,37,0,0,0,0,0,34,0,229,0,129,0,186,0,250,0,8,0,136,0,67,0,180,0,96,0,221,0,81,0,86,0,68,0,4,0,39,0,58,0,0,0,14,0,121,0,241,0,235,0,35,0,119,0,137,0,0,0,0,0,94,0,22,0,99,0,151,0,207,0,184,0,23,0,186,0,44,0,233,0,73,0,39,0,184,0,247,0,68,0,31,0,195,0,0,0,0,0,0,0,0,0,108,0,189,0,0,0,0,0,219,0,155,0,135,0,195,0,97,0,38,0,91,0,0,0,0,0,213,0,187,0,66,0,232,0,202,0,62,0,227,0,0,0,51,0,0,0,78,0,210,0,0,0,154,0,203,0,0,0,57,0,102,0,141,0,0,0,0,0,184,0,174,0,109,0,0,0,155,0,46,0,39,0,77,0,72,0,139,0,42,0,215,0,119,0,37,0,59,0,188,0,223,0,242,0,0,0,0,0,253,0,109,0,0,0,239,0,193,0,0,0,187,0,212,0,243,0,146,0,216,0,63,0,236,0,0,0,195,0,5,0,0,0,205,0,246,0,0,0,164,0,206,0,0,0,11,0,88,0,6,0,0,0,140,0,141,0,174,0,67,0,56,0,0,0,14,0,77,0,10,0,66,0,21,0,155,0,0,0,16,0,129,0,89,0,0,0,18,0,143,0,47,0,180,0,83,0,27,0,66,0,137,0,198,0,168,0,217,0,29,0,163,0,118,0,252,0,72,0,0,0,95,0,0,0,0,0,211,0,123,0,0,0,133,0,0,0,0,0,244,0,69,0,146,0,0,0,155,0,241,0,64,0,56,0,193,0,14,0,82,0,148,0,0,0,0,0,206,0,255,0,4,0,63,0,213,0,151,0,0,0,194,0,33,0,91,0,69,0,0,0,200,0,0,0,64,0,0,0,0,0,0,0,0,0,0,0,106,0,0,0,165,0,115,0,0,0,174,0,224,0,61,0,173,0,39,0,150,0,173,0,179,0,0,0,146,0,130,0,39,0,0,0,42,0,159,0,231,0,0,0,147,0,58,0,163,0,240,0,66,0,150,0,92,0,68,0,124,0,0,0,204,0,169,0,216,0,169,0,229,0,53,0,193,0,0,0,223,0,0,0,99,0,184,0,219,0,174,0,103,0,0,0,162,0,35,0,0,0,0,0,0,0,214,0,147,0,75,0,156,0,18,0,0,0,58,0,16,0,216,0,0,0,119,0,248,0,52,0,0,0,34,0,117,0,31,0,0,0,119,0,0,0,239,0,0,0,138,0,182,0,0,0,62,0,13,0,33,0,0,0,229,0,0,0,134,0,78,0,35,0,202,0,248,0,0,0,33,0,159,0,0,0,106,0,123,0,94,0,53,0,175,0,126,0,97,0,20,0,54,0,214,0,0,0,218,0,0,0,34,0,136,0,241,0,137,0,216,0,0,0,53,0,196,0,0,0,12,0,241,0,42,0,208,0,95,0,186,0,84,0,63,0,88,0,99,0,242,0,0,0,172,0,136,0,70,0,104,0,5,0,0,0,131,0,0,0,53,0,82,0,83,0,228,0,51,0,117,0,42,0,23,0,243,0,183,0,197,0,30,0,60,0,3,0,28,0,38,0,123,0,129,0,0,0,147,0,92,0,227,0,0,0,26,0,193,0,40,0,0,0,0,0,0,0,68,0,45,0,135,0,60,0,147,0,0,0,33,0,0,0,90,0,118,0,0,0,251,0,0,0,54,0,175,0,49,0,175,0,185,0,155,0,0,0,36,0,129,0,0,0,0,0,155,0,0,0,100,0,143,0,171,0,61,0,51,0,113,0,0,0,246,0,152,0,0,0,0,0,70,0,0,0,77,0,185,0,53,0,212,0,175,0,35,0,25,0,157,0,3,0,48,0,167,0,242,0,235,0,164,0,50,0,145,0,193,0,0,0,204,0,16,0,254,0,215,0,80,0,223,0,60,0,160,0,110,0,26,0,0,0,244,0,146,0,223,0,0,0,163,0,37,0,219,0,97,0,65,0,231,0,227,0,28,0,120,0,53,0,146,0,143,0,29,0,66,0,118,0,182,0,201,0,206,0,227,0,0,0,148,0,11,0,228,0,58,0,203,0,243,0,68,0,217,0,249,0,244,0,237,0,0,0,172,0,218,0,13,0,0,0,166,0,28,0,203,0,0,0,129,0,0,0,87,0,0,0,0,0,0,0,0,0,83,0,192,0,120,0,0,0,16,0);
signal scenario_full  : scenario_type := (105,31,195,31,188,31,190,31,237,31,237,30,125,31,89,31,236,31,236,30,105,31,12,31,184,31,84,31,174,31,28,31,47,31,78,31,78,30,78,29,191,31,99,31,171,31,89,31,236,31,236,30,149,31,218,31,43,31,155,31,155,30,64,31,101,31,204,31,204,30,204,29,90,31,130,31,130,30,239,31,235,31,237,31,87,31,233,31,233,30,89,31,34,31,243,31,243,30,243,29,243,28,20,31,20,30,202,31,202,30,122,31,84,31,10,31,10,30,10,29,151,31,240,31,53,31,131,31,90,31,114,31,225,31,225,30,49,31,31,31,31,30,76,31,79,31,127,31,174,31,53,31,142,31,41,31,44,31,44,30,216,31,216,30,30,31,11,31,254,31,14,31,47,31,6,31,219,31,219,30,167,31,225,31,184,31,191,31,254,31,254,30,64,31,227,31,31,31,212,31,212,30,136,31,36,31,105,31,37,31,37,30,37,29,34,31,229,31,129,31,186,31,250,31,8,31,136,31,67,31,180,31,96,31,221,31,81,31,86,31,68,31,4,31,39,31,58,31,58,30,14,31,121,31,241,31,235,31,35,31,119,31,137,31,137,30,137,29,94,31,22,31,99,31,151,31,207,31,184,31,23,31,186,31,44,31,233,31,73,31,39,31,184,31,247,31,68,31,31,31,195,31,195,30,195,29,195,28,195,27,108,31,189,31,189,30,189,29,219,31,155,31,135,31,195,31,97,31,38,31,91,31,91,30,91,29,213,31,187,31,66,31,232,31,202,31,62,31,227,31,227,30,51,31,51,30,78,31,210,31,210,30,154,31,203,31,203,30,57,31,102,31,141,31,141,30,141,29,184,31,174,31,109,31,109,30,155,31,46,31,39,31,77,31,72,31,139,31,42,31,215,31,119,31,37,31,59,31,188,31,223,31,242,31,242,30,242,29,253,31,109,31,109,30,239,31,193,31,193,30,187,31,212,31,243,31,146,31,216,31,63,31,236,31,236,30,195,31,5,31,5,30,205,31,246,31,246,30,164,31,206,31,206,30,11,31,88,31,6,31,6,30,140,31,141,31,174,31,67,31,56,31,56,30,14,31,77,31,10,31,66,31,21,31,155,31,155,30,16,31,129,31,89,31,89,30,18,31,143,31,47,31,180,31,83,31,27,31,66,31,137,31,198,31,168,31,217,31,29,31,163,31,118,31,252,31,72,31,72,30,95,31,95,30,95,29,211,31,123,31,123,30,133,31,133,30,133,29,244,31,69,31,146,31,146,30,155,31,241,31,64,31,56,31,193,31,14,31,82,31,148,31,148,30,148,29,206,31,255,31,4,31,63,31,213,31,151,31,151,30,194,31,33,31,91,31,69,31,69,30,200,31,200,30,64,31,64,30,64,29,64,28,64,27,64,26,106,31,106,30,165,31,115,31,115,30,174,31,224,31,61,31,173,31,39,31,150,31,173,31,179,31,179,30,146,31,130,31,39,31,39,30,42,31,159,31,231,31,231,30,147,31,58,31,163,31,240,31,66,31,150,31,92,31,68,31,124,31,124,30,204,31,169,31,216,31,169,31,229,31,53,31,193,31,193,30,223,31,223,30,99,31,184,31,219,31,174,31,103,31,103,30,162,31,35,31,35,30,35,29,35,28,214,31,147,31,75,31,156,31,18,31,18,30,58,31,16,31,216,31,216,30,119,31,248,31,52,31,52,30,34,31,117,31,31,31,31,30,119,31,119,30,239,31,239,30,138,31,182,31,182,30,62,31,13,31,33,31,33,30,229,31,229,30,134,31,78,31,35,31,202,31,248,31,248,30,33,31,159,31,159,30,106,31,123,31,94,31,53,31,175,31,126,31,97,31,20,31,54,31,214,31,214,30,218,31,218,30,34,31,136,31,241,31,137,31,216,31,216,30,53,31,196,31,196,30,12,31,241,31,42,31,208,31,95,31,186,31,84,31,63,31,88,31,99,31,242,31,242,30,172,31,136,31,70,31,104,31,5,31,5,30,131,31,131,30,53,31,82,31,83,31,228,31,51,31,117,31,42,31,23,31,243,31,183,31,197,31,30,31,60,31,3,31,28,31,38,31,123,31,129,31,129,30,147,31,92,31,227,31,227,30,26,31,193,31,40,31,40,30,40,29,40,28,68,31,45,31,135,31,60,31,147,31,147,30,33,31,33,30,90,31,118,31,118,30,251,31,251,30,54,31,175,31,49,31,175,31,185,31,155,31,155,30,36,31,129,31,129,30,129,29,155,31,155,30,100,31,143,31,171,31,61,31,51,31,113,31,113,30,246,31,152,31,152,30,152,29,70,31,70,30,77,31,185,31,53,31,212,31,175,31,35,31,25,31,157,31,3,31,48,31,167,31,242,31,235,31,164,31,50,31,145,31,193,31,193,30,204,31,16,31,254,31,215,31,80,31,223,31,60,31,160,31,110,31,26,31,26,30,244,31,146,31,223,31,223,30,163,31,37,31,219,31,97,31,65,31,231,31,227,31,28,31,120,31,53,31,146,31,143,31,29,31,66,31,118,31,182,31,201,31,206,31,227,31,227,30,148,31,11,31,228,31,58,31,203,31,243,31,68,31,217,31,249,31,244,31,237,31,237,30,172,31,218,31,13,31,13,30,166,31,28,31,203,31,203,30,129,31,129,30,87,31,87,30,87,29,87,28,87,27,83,31,192,31,120,31,120,30,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
