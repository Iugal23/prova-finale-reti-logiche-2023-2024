-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_397 is
end project_tb_397;

architecture project_tb_arch_397 of project_tb_397 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 876;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,74,0,204,0,254,0,140,0,168,0,148,0,222,0,0,0,73,0,230,0,189,0,0,0,248,0,134,0,114,0,56,0,183,0,61,0,110,0,108,0,115,0,196,0,14,0,102,0,0,0,81,0,171,0,242,0,236,0,52,0,203,0,159,0,247,0,206,0,132,0,0,0,239,0,183,0,50,0,162,0,0,0,41,0,0,0,42,0,200,0,67,0,0,0,245,0,241,0,33,0,139,0,0,0,54,0,0,0,0,0,145,0,0,0,0,0,108,0,0,0,0,0,27,0,37,0,248,0,32,0,171,0,125,0,55,0,0,0,134,0,134,0,0,0,250,0,25,0,84,0,0,0,0,0,27,0,224,0,31,0,242,0,99,0,168,0,77,0,145,0,23,0,230,0,232,0,212,0,0,0,116,0,142,0,224,0,203,0,20,0,0,0,0,0,0,0,0,0,205,0,209,0,125,0,149,0,152,0,89,0,0,0,115,0,0,0,136,0,122,0,0,0,226,0,85,0,0,0,175,0,192,0,160,0,0,0,166,0,158,0,226,0,141,0,0,0,0,0,108,0,0,0,77,0,226,0,65,0,32,0,217,0,229,0,82,0,11,0,240,0,78,0,91,0,35,0,0,0,5,0,172,0,27,0,116,0,194,0,253,0,216,0,88,0,54,0,242,0,0,0,69,0,27,0,33,0,121,0,0,0,81,0,104,0,0,0,23,0,84,0,99,0,110,0,156,0,192,0,81,0,109,0,149,0,0,0,85,0,118,0,31,0,77,0,78,0,0,0,42,0,0,0,0,0,127,0,0,0,126,0,150,0,195,0,209,0,190,0,76,0,48,0,124,0,136,0,131,0,182,0,0,0,207,0,0,0,117,0,0,0,213,0,112,0,215,0,7,0,34,0,215,0,132,0,201,0,123,0,121,0,223,0,13,0,0,0,124,0,255,0,118,0,0,0,66,0,108,0,167,0,179,0,248,0,0,0,239,0,192,0,42,0,56,0,103,0,52,0,58,0,158,0,160,0,111,0,0,0,158,0,31,0,132,0,216,0,230,0,0,0,113,0,0,0,212,0,94,0,206,0,225,0,177,0,29,0,183,0,228,0,126,0,168,0,128,0,0,0,51,0,1,0,20,0,145,0,74,0,177,0,221,0,26,0,129,0,0,0,0,0,14,0,47,0,237,0,137,0,235,0,50,0,69,0,0,0,104,0,151,0,1,0,0,0,12,0,151,0,58,0,246,0,144,0,0,0,0,0,201,0,242,0,30,0,0,0,101,0,238,0,254,0,29,0,0,0,0,0,126,0,49,0,200,0,65,0,185,0,0,0,49,0,178,0,182,0,187,0,142,0,194,0,209,0,75,0,91,0,0,0,135,0,46,0,17,0,85,0,135,0,103,0,0,0,136,0,85,0,0,0,198,0,155,0,215,0,150,0,0,0,167,0,171,0,119,0,27,0,166,0,82,0,170,0,153,0,0,0,199,0,0,0,188,0,221,0,177,0,186,0,43,0,148,0,231,0,132,0,248,0,0,0,141,0,139,0,161,0,115,0,0,0,253,0,54,0,71,0,208,0,0,0,106,0,175,0,162,0,21,0,178,0,253,0,0,0,207,0,155,0,0,0,200,0,0,0,5,0,0,0,23,0,0,0,152,0,0,0,59,0,0,0,0,0,21,0,0,0,173,0,250,0,26,0,182,0,194,0,97,0,45,0,38,0,85,0,244,0,0,0,58,0,0,0,137,0,206,0,0,0,130,0,160,0,39,0,73,0,108,0,10,0,84,0,225,0,181,0,0,0,46,0,9,0,150,0,74,0,123,0,0,0,26,0,40,0,232,0,23,0,240,0,139,0,188,0,57,0,0,0,219,0,0,0,114,0,141,0,12,0,0,0,0,0,105,0,14,0,0,0,195,0,62,0,109,0,74,0,81,0,146,0,27,0,0,0,203,0,230,0,96,0,240,0,209,0,144,0,212,0,227,0,0,0,28,0,0,0,163,0,0,0,102,0,155,0,142,0,41,0,196,0,0,0,110,0,42,0,0,0,37,0,142,0,0,0,151,0,162,0,227,0,122,0,171,0,0,0,235,0,198,0,0,0,0,0,211,0,72,0,97,0,181,0,194,0,48,0,0,0,0,0,83,0,137,0,1,0,183,0,39,0,85,0,173,0,195,0,232,0,241,0,0,0,0,0,149,0,151,0,0,0,191,0,124,0,157,0,25,0,1,0,37,0,0,0,2,0,87,0,9,0,88,0,156,0,3,0,75,0,4,0,36,0,199,0,107,0,240,0,243,0,0,0,0,0,0,0,0,0,129,0,0,0,183,0,131,0,0,0,21,0,192,0,244,0,197,0,85,0,142,0,24,0,0,0,191,0,241,0,0,0,104,0,165,0,175,0,0,0,149,0,36,0,6,0,80,0,96,0,213,0,129,0,6,0,143,0,0,0,18,0,45,0,0,0,174,0,55,0,98,0,167,0,9,0,80,0,201,0,11,0,109,0,23,0,0,0,78,0,231,0,10,0,132,0,0,0,91,0,119,0,110,0,92,0,130,0,175,0,234,0,22,0,173,0,0,0,252,0,61,0,155,0,80,0,56,0,142,0,244,0,186,0,217,0,0,0,0,0,235,0,17,0,109,0,0,0,255,0,9,0,194,0,61,0,103,0,237,0,0,0,209,0,58,0,236,0,65,0,38,0,213,0,150,0,0,0,130,0,0,0,36,0,145,0,105,0,233,0,88,0,53,0,40,0,248,0,0,0,184,0,0,0,17,0,0,0,161,0,0,0,154,0,115,0,208,0,37,0,169,0,197,0,231,0,90,0,0,0,59,0,98,0,195,0,47,0,0,0,144,0,144,0,191,0,165,0,0,0,0,0,62,0,229,0,225,0,61,0,55,0,24,0,147,0,47,0,228,0,145,0,41,0,0,0,112,0,0,0,249,0,98,0,110,0,0,0,35,0,130,0,156,0,122,0,0,0,222,0,6,0,110,0,133,0,51,0,38,0,230,0,80,0,70,0,193,0,246,0,52,0,254,0,125,0,0,0,118,0,0,0,15,0,238,0,0,0,204,0,175,0,10,0,118,0,39,0,0,0,71,0,0,0,186,0,60,0,236,0,185,0,19,0,162,0,136,0,94,0,0,0,0,0,223,0,0,0,111,0,11,0,0,0,55,0,231,0,72,0,116,0,0,0,138,0,74,0,0,0,52,0,58,0,0,0,54,0,63,0,142,0,247,0,0,0,65,0,217,0,76,0,128,0,64,0,0,0,59,0,120,0,27,0,4,0,1,0,103,0,0,0,0,0,0,0,107,0,114,0,238,0,136,0,29,0,180,0,220,0,231,0,250,0,73,0,0,0,102,0,132,0,0,0,204,0,79,0,54,0,69,0,80,0,72,0,234,0,176,0,50,0,195,0,26,0,60,0,0,0,225,0,7,0,0,0,107,0,24,0,233,0,188,0,76,0,88,0,158,0,6,0,236,0,81,0,0,0,19,0,111,0,0,0,0,0,235,0,239,0,219,0,0,0,246,0,0,0,136,0,194,0,152,0,48,0,111,0,211,0,68,0,38,0,0,0,248,0,91,0,241,0,218,0,240,0,229,0,123,0,26,0,107,0,11,0,0,0,96,0,207,0,64,0,219,0,211,0,158,0,33,0,211,0,179,0,0,0,7,0,0,0,0,0,191,0,0,0,0,0,197,0,250,0,169,0,84,0,199,0,163,0,59,0,12,0,7,0,109,0,233,0,6,0,184,0,67,0,0,0,0,0,96,0,92,0,254,0,147,0,238,0,51,0,0,0,208,0,219,0,106,0,220,0,207,0,108,0,117,0,211,0,83,0,94,0,199,0,119,0,126,0,228,0,4,0,113,0,21,0,0,0,20,0,155,0,154,0,73,0,239,0,194,0,0,0,206,0,0,0);
signal scenario_full  : scenario_type := (0,0,74,31,204,31,254,31,140,31,168,31,148,31,222,31,222,30,73,31,230,31,189,31,189,30,248,31,134,31,114,31,56,31,183,31,61,31,110,31,108,31,115,31,196,31,14,31,102,31,102,30,81,31,171,31,242,31,236,31,52,31,203,31,159,31,247,31,206,31,132,31,132,30,239,31,183,31,50,31,162,31,162,30,41,31,41,30,42,31,200,31,67,31,67,30,245,31,241,31,33,31,139,31,139,30,54,31,54,30,54,29,145,31,145,30,145,29,108,31,108,30,108,29,27,31,37,31,248,31,32,31,171,31,125,31,55,31,55,30,134,31,134,31,134,30,250,31,25,31,84,31,84,30,84,29,27,31,224,31,31,31,242,31,99,31,168,31,77,31,145,31,23,31,230,31,232,31,212,31,212,30,116,31,142,31,224,31,203,31,20,31,20,30,20,29,20,28,20,27,205,31,209,31,125,31,149,31,152,31,89,31,89,30,115,31,115,30,136,31,122,31,122,30,226,31,85,31,85,30,175,31,192,31,160,31,160,30,166,31,158,31,226,31,141,31,141,30,141,29,108,31,108,30,77,31,226,31,65,31,32,31,217,31,229,31,82,31,11,31,240,31,78,31,91,31,35,31,35,30,5,31,172,31,27,31,116,31,194,31,253,31,216,31,88,31,54,31,242,31,242,30,69,31,27,31,33,31,121,31,121,30,81,31,104,31,104,30,23,31,84,31,99,31,110,31,156,31,192,31,81,31,109,31,149,31,149,30,85,31,118,31,31,31,77,31,78,31,78,30,42,31,42,30,42,29,127,31,127,30,126,31,150,31,195,31,209,31,190,31,76,31,48,31,124,31,136,31,131,31,182,31,182,30,207,31,207,30,117,31,117,30,213,31,112,31,215,31,7,31,34,31,215,31,132,31,201,31,123,31,121,31,223,31,13,31,13,30,124,31,255,31,118,31,118,30,66,31,108,31,167,31,179,31,248,31,248,30,239,31,192,31,42,31,56,31,103,31,52,31,58,31,158,31,160,31,111,31,111,30,158,31,31,31,132,31,216,31,230,31,230,30,113,31,113,30,212,31,94,31,206,31,225,31,177,31,29,31,183,31,228,31,126,31,168,31,128,31,128,30,51,31,1,31,20,31,145,31,74,31,177,31,221,31,26,31,129,31,129,30,129,29,14,31,47,31,237,31,137,31,235,31,50,31,69,31,69,30,104,31,151,31,1,31,1,30,12,31,151,31,58,31,246,31,144,31,144,30,144,29,201,31,242,31,30,31,30,30,101,31,238,31,254,31,29,31,29,30,29,29,126,31,49,31,200,31,65,31,185,31,185,30,49,31,178,31,182,31,187,31,142,31,194,31,209,31,75,31,91,31,91,30,135,31,46,31,17,31,85,31,135,31,103,31,103,30,136,31,85,31,85,30,198,31,155,31,215,31,150,31,150,30,167,31,171,31,119,31,27,31,166,31,82,31,170,31,153,31,153,30,199,31,199,30,188,31,221,31,177,31,186,31,43,31,148,31,231,31,132,31,248,31,248,30,141,31,139,31,161,31,115,31,115,30,253,31,54,31,71,31,208,31,208,30,106,31,175,31,162,31,21,31,178,31,253,31,253,30,207,31,155,31,155,30,200,31,200,30,5,31,5,30,23,31,23,30,152,31,152,30,59,31,59,30,59,29,21,31,21,30,173,31,250,31,26,31,182,31,194,31,97,31,45,31,38,31,85,31,244,31,244,30,58,31,58,30,137,31,206,31,206,30,130,31,160,31,39,31,73,31,108,31,10,31,84,31,225,31,181,31,181,30,46,31,9,31,150,31,74,31,123,31,123,30,26,31,40,31,232,31,23,31,240,31,139,31,188,31,57,31,57,30,219,31,219,30,114,31,141,31,12,31,12,30,12,29,105,31,14,31,14,30,195,31,62,31,109,31,74,31,81,31,146,31,27,31,27,30,203,31,230,31,96,31,240,31,209,31,144,31,212,31,227,31,227,30,28,31,28,30,163,31,163,30,102,31,155,31,142,31,41,31,196,31,196,30,110,31,42,31,42,30,37,31,142,31,142,30,151,31,162,31,227,31,122,31,171,31,171,30,235,31,198,31,198,30,198,29,211,31,72,31,97,31,181,31,194,31,48,31,48,30,48,29,83,31,137,31,1,31,183,31,39,31,85,31,173,31,195,31,232,31,241,31,241,30,241,29,149,31,151,31,151,30,191,31,124,31,157,31,25,31,1,31,37,31,37,30,2,31,87,31,9,31,88,31,156,31,3,31,75,31,4,31,36,31,199,31,107,31,240,31,243,31,243,30,243,29,243,28,243,27,129,31,129,30,183,31,131,31,131,30,21,31,192,31,244,31,197,31,85,31,142,31,24,31,24,30,191,31,241,31,241,30,104,31,165,31,175,31,175,30,149,31,36,31,6,31,80,31,96,31,213,31,129,31,6,31,143,31,143,30,18,31,45,31,45,30,174,31,55,31,98,31,167,31,9,31,80,31,201,31,11,31,109,31,23,31,23,30,78,31,231,31,10,31,132,31,132,30,91,31,119,31,110,31,92,31,130,31,175,31,234,31,22,31,173,31,173,30,252,31,61,31,155,31,80,31,56,31,142,31,244,31,186,31,217,31,217,30,217,29,235,31,17,31,109,31,109,30,255,31,9,31,194,31,61,31,103,31,237,31,237,30,209,31,58,31,236,31,65,31,38,31,213,31,150,31,150,30,130,31,130,30,36,31,145,31,105,31,233,31,88,31,53,31,40,31,248,31,248,30,184,31,184,30,17,31,17,30,161,31,161,30,154,31,115,31,208,31,37,31,169,31,197,31,231,31,90,31,90,30,59,31,98,31,195,31,47,31,47,30,144,31,144,31,191,31,165,31,165,30,165,29,62,31,229,31,225,31,61,31,55,31,24,31,147,31,47,31,228,31,145,31,41,31,41,30,112,31,112,30,249,31,98,31,110,31,110,30,35,31,130,31,156,31,122,31,122,30,222,31,6,31,110,31,133,31,51,31,38,31,230,31,80,31,70,31,193,31,246,31,52,31,254,31,125,31,125,30,118,31,118,30,15,31,238,31,238,30,204,31,175,31,10,31,118,31,39,31,39,30,71,31,71,30,186,31,60,31,236,31,185,31,19,31,162,31,136,31,94,31,94,30,94,29,223,31,223,30,111,31,11,31,11,30,55,31,231,31,72,31,116,31,116,30,138,31,74,31,74,30,52,31,58,31,58,30,54,31,63,31,142,31,247,31,247,30,65,31,217,31,76,31,128,31,64,31,64,30,59,31,120,31,27,31,4,31,1,31,103,31,103,30,103,29,103,28,107,31,114,31,238,31,136,31,29,31,180,31,220,31,231,31,250,31,73,31,73,30,102,31,132,31,132,30,204,31,79,31,54,31,69,31,80,31,72,31,234,31,176,31,50,31,195,31,26,31,60,31,60,30,225,31,7,31,7,30,107,31,24,31,233,31,188,31,76,31,88,31,158,31,6,31,236,31,81,31,81,30,19,31,111,31,111,30,111,29,235,31,239,31,219,31,219,30,246,31,246,30,136,31,194,31,152,31,48,31,111,31,211,31,68,31,38,31,38,30,248,31,91,31,241,31,218,31,240,31,229,31,123,31,26,31,107,31,11,31,11,30,96,31,207,31,64,31,219,31,211,31,158,31,33,31,211,31,179,31,179,30,7,31,7,30,7,29,191,31,191,30,191,29,197,31,250,31,169,31,84,31,199,31,163,31,59,31,12,31,7,31,109,31,233,31,6,31,184,31,67,31,67,30,67,29,96,31,92,31,254,31,147,31,238,31,51,31,51,30,208,31,219,31,106,31,220,31,207,31,108,31,117,31,211,31,83,31,94,31,199,31,119,31,126,31,228,31,4,31,113,31,21,31,21,30,20,31,155,31,154,31,73,31,239,31,194,31,194,30,206,31,206,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
