-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_144 is
end project_tb_144;

architecture project_tb_arch_144 of project_tb_144 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 173;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (117,0,13,0,144,0,160,0,0,0,231,0,8,0,0,0,36,0,229,0,0,0,99,0,61,0,65,0,135,0,164,0,0,0,132,0,68,0,14,0,119,0,200,0,69,0,71,0,240,0,143,0,96,0,3,0,175,0,31,0,85,0,35,0,204,0,79,0,213,0,199,0,1,0,205,0,195,0,33,0,203,0,112,0,119,0,15,0,37,0,155,0,57,0,152,0,212,0,167,0,23,0,0,0,103,0,142,0,162,0,0,0,0,0,27,0,0,0,112,0,105,0,157,0,0,0,57,0,4,0,202,0,0,0,196,0,0,0,0,0,253,0,0,0,224,0,42,0,112,0,67,0,38,0,229,0,67,0,74,0,64,0,115,0,83,0,0,0,247,0,53,0,205,0,18,0,158,0,0,0,140,0,237,0,0,0,0,0,226,0,145,0,113,0,233,0,229,0,17,0,105,0,0,0,129,0,95,0,98,0,0,0,70,0,39,0,228,0,109,0,220,0,78,0,6,0,174,0,170,0,255,0,32,0,0,0,0,0,168,0,0,0,49,0,197,0,191,0,83,0,15,0,222,0,242,0,198,0,147,0,0,0,15,0,36,0,113,0,78,0,125,0,0,0,191,0,109,0,21,0,0,0,216,0,68,0,171,0,168,0,5,0,171,0,205,0,0,0,15,0,109,0,124,0,8,0,225,0,0,0,44,0,175,0,180,0,202,0,40,0,161,0,0,0,251,0,161,0,143,0,225,0,0,0,0,0,0,0,197,0,0,0,200,0,135,0);
signal scenario_full  : scenario_type := (117,31,13,31,144,31,160,31,160,30,231,31,8,31,8,30,36,31,229,31,229,30,99,31,61,31,65,31,135,31,164,31,164,30,132,31,68,31,14,31,119,31,200,31,69,31,71,31,240,31,143,31,96,31,3,31,175,31,31,31,85,31,35,31,204,31,79,31,213,31,199,31,1,31,205,31,195,31,33,31,203,31,112,31,119,31,15,31,37,31,155,31,57,31,152,31,212,31,167,31,23,31,23,30,103,31,142,31,162,31,162,30,162,29,27,31,27,30,112,31,105,31,157,31,157,30,57,31,4,31,202,31,202,30,196,31,196,30,196,29,253,31,253,30,224,31,42,31,112,31,67,31,38,31,229,31,67,31,74,31,64,31,115,31,83,31,83,30,247,31,53,31,205,31,18,31,158,31,158,30,140,31,237,31,237,30,237,29,226,31,145,31,113,31,233,31,229,31,17,31,105,31,105,30,129,31,95,31,98,31,98,30,70,31,39,31,228,31,109,31,220,31,78,31,6,31,174,31,170,31,255,31,32,31,32,30,32,29,168,31,168,30,49,31,197,31,191,31,83,31,15,31,222,31,242,31,198,31,147,31,147,30,15,31,36,31,113,31,78,31,125,31,125,30,191,31,109,31,21,31,21,30,216,31,68,31,171,31,168,31,5,31,171,31,205,31,205,30,15,31,109,31,124,31,8,31,225,31,225,30,44,31,175,31,180,31,202,31,40,31,161,31,161,30,251,31,161,31,143,31,225,31,225,30,225,29,225,28,197,31,197,30,200,31,135,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
