-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 427;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (117,0,0,0,251,0,184,0,221,0,181,0,180,0,245,0,252,0,107,0,0,0,173,0,0,0,197,0,135,0,67,0,213,0,104,0,237,0,0,0,0,0,38,0,144,0,128,0,0,0,108,0,0,0,133,0,181,0,122,0,46,0,176,0,15,0,20,0,141,0,2,0,0,0,160,0,124,0,120,0,0,0,0,0,54,0,0,0,0,0,85,0,0,0,167,0,2,0,0,0,202,0,160,0,255,0,78,0,0,0,0,0,184,0,75,0,43,0,187,0,211,0,220,0,0,0,240,0,25,0,15,0,72,0,168,0,0,0,232,0,0,0,95,0,128,0,0,0,171,0,92,0,17,0,46,0,131,0,95,0,204,0,0,0,109,0,63,0,213,0,173,0,129,0,161,0,5,0,21,0,222,0,169,0,0,0,116,0,17,0,38,0,245,0,176,0,30,0,0,0,0,0,194,0,172,0,186,0,48,0,67,0,88,0,0,0,245,0,235,0,203,0,240,0,15,0,0,0,9,0,215,0,17,0,27,0,0,0,0,0,2,0,86,0,149,0,217,0,159,0,84,0,92,0,15,0,179,0,247,0,127,0,26,0,0,0,0,0,152,0,179,0,122,0,183,0,50,0,233,0,0,0,0,0,204,0,190,0,89,0,0,0,169,0,13,0,234,0,0,0,199,0,124,0,168,0,0,0,135,0,102,0,173,0,85,0,6,0,102,0,33,0,17,0,0,0,221,0,104,0,102,0,78,0,247,0,41,0,5,0,30,0,0,0,67,0,45,0,179,0,0,0,123,0,112,0,30,0,167,0,204,0,0,0,72,0,22,0,107,0,141,0,253,0,83,0,143,0,158,0,146,0,127,0,117,0,204,0,0,0,86,0,185,0,0,0,214,0,119,0,149,0,0,0,0,0,0,0,24,0,0,0,50,0,52,0,91,0,87,0,71,0,212,0,106,0,197,0,204,0,157,0,161,0,229,0,0,0,3,0,114,0,0,0,134,0,0,0,188,0,223,0,50,0,52,0,92,0,229,0,64,0,205,0,160,0,103,0,95,0,54,0,44,0,123,0,67,0,250,0,211,0,96,0,157,0,118,0,10,0,65,0,31,0,0,0,172,0,0,0,76,0,244,0,0,0,119,0,0,0,46,0,113,0,87,0,0,0,43,0,64,0,0,0,33,0,184,0,204,0,165,0,59,0,115,0,161,0,107,0,103,0,0,0,209,0,0,0,0,0,237,0,35,0,171,0,201,0,1,0,32,0,165,0,181,0,86,0,121,0,92,0,88,0,149,0,0,0,132,0,0,0,0,0,117,0,255,0,64,0,192,0,0,0,72,0,128,0,56,0,0,0,219,0,77,0,251,0,52,0,0,0,137,0,0,0,0,0,16,0,98,0,21,0,89,0,94,0,90,0,25,0,213,0,0,0,0,0,0,0,230,0,90,0,149,0,129,0,12,0,224,0,190,0,83,0,26,0,173,0,56,0,0,0,98,0,197,0,150,0,159,0,219,0,42,0,187,0,15,0,0,0,151,0,178,0,8,0,0,0,99,0,151,0,118,0,189,0,107,0,197,0,4,0,116,0,180,0,166,0,71,0,253,0,0,0,26,0,0,0,179,0,106,0,222,0,27,0,208,0,91,0,26,0,181,0,129,0,255,0,0,0,236,0,10,0,176,0,228,0,8,0,18,0,81,0,0,0,70,0,0,0,111,0,102,0,0,0,129,0,234,0,225,0,254,0,0,0,205,0,178,0,56,0,172,0,46,0,0,0,0,0,23,0,142,0,163,0,102,0,0,0,228,0,0,0,214,0,151,0,163,0,199,0,251,0,0,0,190,0,30,0,213,0,131,0,83,0,0,0,0,0,152,0,221,0,49,0,193,0,44,0,0,0,0,0,147,0,78,0,22,0,138,0);
signal scenario_full  : scenario_type := (117,31,117,30,251,31,184,31,221,31,181,31,180,31,245,31,252,31,107,31,107,30,173,31,173,30,197,31,135,31,67,31,213,31,104,31,237,31,237,30,237,29,38,31,144,31,128,31,128,30,108,31,108,30,133,31,181,31,122,31,46,31,176,31,15,31,20,31,141,31,2,31,2,30,160,31,124,31,120,31,120,30,120,29,54,31,54,30,54,29,85,31,85,30,167,31,2,31,2,30,202,31,160,31,255,31,78,31,78,30,78,29,184,31,75,31,43,31,187,31,211,31,220,31,220,30,240,31,25,31,15,31,72,31,168,31,168,30,232,31,232,30,95,31,128,31,128,30,171,31,92,31,17,31,46,31,131,31,95,31,204,31,204,30,109,31,63,31,213,31,173,31,129,31,161,31,5,31,21,31,222,31,169,31,169,30,116,31,17,31,38,31,245,31,176,31,30,31,30,30,30,29,194,31,172,31,186,31,48,31,67,31,88,31,88,30,245,31,235,31,203,31,240,31,15,31,15,30,9,31,215,31,17,31,27,31,27,30,27,29,2,31,86,31,149,31,217,31,159,31,84,31,92,31,15,31,179,31,247,31,127,31,26,31,26,30,26,29,152,31,179,31,122,31,183,31,50,31,233,31,233,30,233,29,204,31,190,31,89,31,89,30,169,31,13,31,234,31,234,30,199,31,124,31,168,31,168,30,135,31,102,31,173,31,85,31,6,31,102,31,33,31,17,31,17,30,221,31,104,31,102,31,78,31,247,31,41,31,5,31,30,31,30,30,67,31,45,31,179,31,179,30,123,31,112,31,30,31,167,31,204,31,204,30,72,31,22,31,107,31,141,31,253,31,83,31,143,31,158,31,146,31,127,31,117,31,204,31,204,30,86,31,185,31,185,30,214,31,119,31,149,31,149,30,149,29,149,28,24,31,24,30,50,31,52,31,91,31,87,31,71,31,212,31,106,31,197,31,204,31,157,31,161,31,229,31,229,30,3,31,114,31,114,30,134,31,134,30,188,31,223,31,50,31,52,31,92,31,229,31,64,31,205,31,160,31,103,31,95,31,54,31,44,31,123,31,67,31,250,31,211,31,96,31,157,31,118,31,10,31,65,31,31,31,31,30,172,31,172,30,76,31,244,31,244,30,119,31,119,30,46,31,113,31,87,31,87,30,43,31,64,31,64,30,33,31,184,31,204,31,165,31,59,31,115,31,161,31,107,31,103,31,103,30,209,31,209,30,209,29,237,31,35,31,171,31,201,31,1,31,32,31,165,31,181,31,86,31,121,31,92,31,88,31,149,31,149,30,132,31,132,30,132,29,117,31,255,31,64,31,192,31,192,30,72,31,128,31,56,31,56,30,219,31,77,31,251,31,52,31,52,30,137,31,137,30,137,29,16,31,98,31,21,31,89,31,94,31,90,31,25,31,213,31,213,30,213,29,213,28,230,31,90,31,149,31,129,31,12,31,224,31,190,31,83,31,26,31,173,31,56,31,56,30,98,31,197,31,150,31,159,31,219,31,42,31,187,31,15,31,15,30,151,31,178,31,8,31,8,30,99,31,151,31,118,31,189,31,107,31,197,31,4,31,116,31,180,31,166,31,71,31,253,31,253,30,26,31,26,30,179,31,106,31,222,31,27,31,208,31,91,31,26,31,181,31,129,31,255,31,255,30,236,31,10,31,176,31,228,31,8,31,18,31,81,31,81,30,70,31,70,30,111,31,102,31,102,30,129,31,234,31,225,31,254,31,254,30,205,31,178,31,56,31,172,31,46,31,46,30,46,29,23,31,142,31,163,31,102,31,102,30,228,31,228,30,214,31,151,31,163,31,199,31,251,31,251,30,190,31,30,31,213,31,131,31,83,31,83,30,83,29,152,31,221,31,49,31,193,31,44,31,44,30,44,29,147,31,78,31,22,31,138,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
